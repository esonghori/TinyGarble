
module matrixMult_N_M_0_N5_M8 ( clk, rst, x, y, o );
  input [199:0] x;
  input [199:0] y;
  output [199:0] o;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320;

  XNOR U1 ( .A(n5704), .B(n5703), .Z(n5759) );
  XNOR U2 ( .A(n5698), .B(n5697), .Z(n5763) );
  XNOR U3 ( .A(n7943), .B(n8003), .Z(n7952) );
  XNOR U4 ( .A(n7901), .B(n7900), .Z(n7958) );
  XNOR U5 ( .A(n12270), .B(n12269), .Z(n12243) );
  XNOR U6 ( .A(n12367), .B(n12296), .Z(n12299) );
  XNOR U7 ( .A(n12995), .B(n12994), .Z(n13038) );
  XNOR U8 ( .A(n15890), .B(n15889), .Z(n15933) );
  XNOR U9 ( .A(n15884), .B(n15883), .Z(n15937) );
  XNOR U10 ( .A(n17407), .B(n17347), .Z(n17356) );
  XNOR U11 ( .A(n17304), .B(n17303), .Z(n17362) );
  NAND U12 ( .A(n7261), .B(n7260), .Z(n1) );
  NAND U13 ( .A(n7259), .B(n7258), .Z(n2) );
  AND U14 ( .A(n1), .B(n2), .Z(n7267) );
  NAND U15 ( .A(n13775), .B(n13774), .Z(n3) );
  NAND U16 ( .A(n13772), .B(n13773), .Z(n4) );
  NAND U17 ( .A(n3), .B(n4), .Z(n13848) );
  NAND U18 ( .A(n15229), .B(n15228), .Z(n5) );
  NAND U19 ( .A(n15227), .B(n15226), .Z(n6) );
  AND U20 ( .A(n5), .B(n6), .Z(n15361) );
  NAND U21 ( .A(n1500), .B(n1499), .Z(n7) );
  NAND U22 ( .A(n1498), .B(n1497), .Z(n8) );
  AND U23 ( .A(n7), .B(n8), .Z(n1778) );
  NAND U24 ( .A(n2913), .B(n2912), .Z(n9) );
  NAND U25 ( .A(n2910), .B(n2911), .Z(n10) );
  AND U26 ( .A(n9), .B(n10), .Z(n3307) );
  NANDN U27 ( .A(n7438), .B(n7437), .Z(n11) );
  NANDN U28 ( .A(n7436), .B(n7476), .Z(n12) );
  AND U29 ( .A(n11), .B(n12), .Z(n13) );
  NAND U30 ( .A(n7442), .B(n7441), .Z(n14) );
  NAND U31 ( .A(n7439), .B(n7440), .Z(n15) );
  AND U32 ( .A(n14), .B(n15), .Z(n16) );
  NANDN U33 ( .A(n7446), .B(n7445), .Z(n17) );
  NANDN U34 ( .A(n7444), .B(n7443), .Z(n18) );
  NAND U35 ( .A(n17), .B(n18), .Z(n19) );
  XNOR U36 ( .A(n13), .B(n16), .Z(n20) );
  XNOR U37 ( .A(n19), .B(n20), .Z(n7447) );
  XOR U38 ( .A(n8878), .B(n8877), .Z(n8876) );
  XNOR U39 ( .A(n9136), .B(n9135), .Z(n9129) );
  NAND U40 ( .A(n10851), .B(n10850), .Z(n21) );
  NAND U41 ( .A(n10848), .B(n10849), .Z(n22) );
  NAND U42 ( .A(n21), .B(n22), .Z(n10991) );
  NAND U43 ( .A(n10881), .B(n10880), .Z(n23) );
  NAND U44 ( .A(n10878), .B(n10879), .Z(n24) );
  NAND U45 ( .A(n23), .B(n24), .Z(n11033) );
  XNOR U46 ( .A(n11753), .B(n11752), .Z(n11751) );
  XNOR U47 ( .A(n12700), .B(n12699), .Z(n12749) );
  NAND U48 ( .A(n16902), .B(n16903), .Z(n25) );
  NAND U49 ( .A(n16904), .B(n16905), .Z(n26) );
  AND U50 ( .A(n25), .B(n26), .Z(n27) );
  NAND U51 ( .A(n16908), .B(n16909), .Z(n28) );
  NAND U52 ( .A(n16906), .B(n16907), .Z(n29) );
  AND U53 ( .A(n28), .B(n29), .Z(n30) );
  NAND U54 ( .A(n16910), .B(n16911), .Z(n31) );
  NAND U55 ( .A(n16912), .B(n16913), .Z(n32) );
  AND U56 ( .A(n31), .B(n32), .Z(n33) );
  XOR U57 ( .A(n16991), .B(n16990), .Z(n34) );
  XNOR U58 ( .A(n16929), .B(n16928), .Z(n35) );
  XNOR U59 ( .A(n34), .B(n35), .Z(n36) );
  XOR U60 ( .A(n33), .B(n36), .Z(n37) );
  XNOR U61 ( .A(n27), .B(n30), .Z(n38) );
  XNOR U62 ( .A(n37), .B(n38), .Z(n39) );
  NAND U63 ( .A(n16898), .B(n16899), .Z(n40) );
  NANDN U64 ( .A(n16901), .B(n16900), .Z(n41) );
  NAND U65 ( .A(n40), .B(n41), .Z(n42) );
  XNOR U66 ( .A(n39), .B(n42), .Z(n17008) );
  NAND U67 ( .A(n2923), .B(n2922), .Z(n43) );
  NAND U68 ( .A(n2920), .B(n2921), .Z(n44) );
  NAND U69 ( .A(n43), .B(n44), .Z(n3034) );
  XNOR U70 ( .A(n3780), .B(n3779), .Z(n3778) );
  XNOR U71 ( .A(n4771), .B(n4770), .Z(n4768) );
  XNOR U72 ( .A(n5217), .B(n5216), .Z(n5215) );
  NAND U73 ( .A(n6594), .B(n6593), .Z(n45) );
  NANDN U74 ( .A(n6592), .B(n6591), .Z(n46) );
  AND U75 ( .A(n45), .B(n46), .Z(n6673) );
  NAND U76 ( .A(n8786), .B(n8785), .Z(n47) );
  NANDN U77 ( .A(n8784), .B(n8783), .Z(n48) );
  AND U78 ( .A(n47), .B(n48), .Z(n8865) );
  XNOR U79 ( .A(n9569), .B(n9568), .Z(n9567) );
  XNOR U80 ( .A(n10288), .B(n10287), .Z(n10286) );
  NAND U81 ( .A(n10995), .B(n10994), .Z(n49) );
  NANDN U82 ( .A(n10997), .B(n10996), .Z(n50) );
  NAND U83 ( .A(n49), .B(n50), .Z(n11288) );
  XNOR U84 ( .A(n14667), .B(n14666), .Z(n14665) );
  NAND U85 ( .A(n15289), .B(n15288), .Z(n51) );
  NANDN U86 ( .A(n15287), .B(n15286), .Z(n52) );
  AND U87 ( .A(n51), .B(n52), .Z(n15375) );
  XNOR U88 ( .A(n17086), .B(n17085), .Z(n17083) );
  XNOR U89 ( .A(n18271), .B(n18270), .Z(n18268) );
  XNOR U90 ( .A(n6523), .B(n6522), .Z(n6524) );
  NAND U91 ( .A(n7071), .B(n7072), .Z(n53) );
  NAND U92 ( .A(n7211), .B(n7208), .Z(n54) );
  NAND U93 ( .A(n53), .B(n54), .Z(n7079) );
  XNOR U94 ( .A(n7907), .B(n7906), .Z(n7954) );
  XOR U95 ( .A(n12292), .B(n12291), .Z(n12242) );
  NAND U96 ( .A(n13627), .B(n13626), .Z(n55) );
  NAND U97 ( .A(n13624), .B(n13625), .Z(n56) );
  NAND U98 ( .A(n55), .B(n56), .Z(n13764) );
  NAND U99 ( .A(n13647), .B(n13646), .Z(n57) );
  NANDN U100 ( .A(n13645), .B(n13644), .Z(n58) );
  NAND U101 ( .A(n57), .B(n58), .Z(n13776) );
  XNOR U102 ( .A(n17310), .B(n17309), .Z(n17358) );
  XOR U103 ( .A(n3273), .B(n3272), .Z(n3271) );
  NAND U104 ( .A(n2881), .B(n2880), .Z(n59) );
  NAND U105 ( .A(n2878), .B(n2879), .Z(n60) );
  NAND U106 ( .A(n59), .B(n60), .Z(n2912) );
  XOR U107 ( .A(n3788), .B(n3789), .Z(n61) );
  XNOR U108 ( .A(n3787), .B(n61), .Z(n3903) );
  NAND U109 ( .A(n4322), .B(n4321), .Z(n62) );
  NAND U110 ( .A(n4319), .B(n4320), .Z(n63) );
  NAND U111 ( .A(n62), .B(n63), .Z(n4412) );
  XNOR U112 ( .A(n5766), .B(n5765), .Z(n5779) );
  XNOR U113 ( .A(n6519), .B(n6518), .Z(n6512) );
  NAND U114 ( .A(n7182), .B(n7181), .Z(n64) );
  NANDN U115 ( .A(n7184), .B(n7183), .Z(n65) );
  NAND U116 ( .A(n64), .B(n65), .Z(n7311) );
  XNOR U117 ( .A(n7961), .B(n7960), .Z(n7968) );
  NAND U118 ( .A(n10126), .B(n10125), .Z(n66) );
  NAND U119 ( .A(n10123), .B(n10124), .Z(n67) );
  NAND U120 ( .A(n66), .B(n67), .Z(n10227) );
  XNOR U121 ( .A(n10523), .B(n10522), .Z(n10520) );
  NAND U122 ( .A(n10831), .B(n10830), .Z(n68) );
  NAND U123 ( .A(n10828), .B(n10829), .Z(n69) );
  NAND U124 ( .A(n68), .B(n69), .Z(n10939) );
  XOR U125 ( .A(n11242), .B(n11243), .Z(n11241) );
  XNOR U126 ( .A(n12308), .B(n12307), .Z(n12321) );
  XNOR U127 ( .A(n12591), .B(n12385), .Z(n12372) );
  XNOR U128 ( .A(n12711), .B(n12712), .Z(n12713) );
  XNOR U129 ( .A(n12411), .B(n12410), .Z(n12412) );
  NAND U130 ( .A(n13771), .B(n13770), .Z(n70) );
  NAND U131 ( .A(n13768), .B(n13769), .Z(n71) );
  NAND U132 ( .A(n70), .B(n71), .Z(n13847) );
  NAND U133 ( .A(n13783), .B(n13782), .Z(n72) );
  NAND U134 ( .A(n13780), .B(n13781), .Z(n73) );
  NAND U135 ( .A(n72), .B(n73), .Z(n13900) );
  XNOR U136 ( .A(n14810), .B(n14809), .Z(n14807) );
  XNOR U137 ( .A(n15940), .B(n15939), .Z(n15953) );
  NAND U138 ( .A(n16673), .B(n16672), .Z(n74) );
  NAND U139 ( .A(n16670), .B(n16671), .Z(n75) );
  NAND U140 ( .A(n74), .B(n75), .Z(n16762) );
  XNOR U141 ( .A(n17365), .B(n17364), .Z(n17372) );
  XNOR U142 ( .A(n18116), .B(n18115), .Z(n18109) );
  NAND U143 ( .A(n1479), .B(n1478), .Z(n76) );
  NAND U144 ( .A(n1476), .B(n1477), .Z(n77) );
  NAND U145 ( .A(n76), .B(n77), .Z(n1546) );
  XNOR U146 ( .A(n2239), .B(n2238), .Z(n2148) );
  XOR U147 ( .A(n2317), .B(n2316), .Z(n2315) );
  XNOR U148 ( .A(n3046), .B(n3045), .Z(n3043) );
  NAND U149 ( .A(n2907), .B(n2906), .Z(n78) );
  NANDN U150 ( .A(n2909), .B(n2908), .Z(n79) );
  AND U151 ( .A(n78), .B(n79), .Z(n3308) );
  NAND U152 ( .A(n4344), .B(n4343), .Z(n80) );
  NANDN U153 ( .A(n4342), .B(n4341), .Z(n81) );
  AND U154 ( .A(n80), .B(n81), .Z(n4759) );
  XNOR U155 ( .A(n5083), .B(n5082), .Z(n5072) );
  XNOR U156 ( .A(n5485), .B(n5484), .Z(n5478) );
  XNOR U157 ( .A(n5844), .B(n5843), .Z(n5845) );
  XNOR U158 ( .A(n5870), .B(n5869), .Z(n5927) );
  NAND U159 ( .A(n7283), .B(n7282), .Z(n82) );
  NAND U160 ( .A(n7280), .B(n7281), .Z(n83) );
  AND U161 ( .A(n82), .B(n83), .Z(n7401) );
  NAND U162 ( .A(n7269), .B(n7268), .Z(n84) );
  NAND U163 ( .A(n7266), .B(n7267), .Z(n85) );
  NAND U164 ( .A(n84), .B(n85), .Z(n7656) );
  XNOR U165 ( .A(n8033), .B(n8032), .Z(n8035) );
  XNOR U166 ( .A(n8735), .B(n8734), .Z(n8724) );
  XOR U167 ( .A(n9117), .B(n9118), .Z(n9111) );
  NAND U168 ( .A(n8794), .B(n8793), .Z(n86) );
  NANDN U169 ( .A(n8796), .B(n8795), .Z(n87) );
  AND U170 ( .A(n86), .B(n87), .Z(n9070) );
  XNOR U171 ( .A(n9444), .B(n9443), .Z(n9433) );
  XNOR U172 ( .A(n10162), .B(n10161), .Z(n10151) );
  XNOR U173 ( .A(n10306), .B(n10305), .Z(n10303) );
  NAND U174 ( .A(n10944), .B(n10943), .Z(n88) );
  NANDN U175 ( .A(n10946), .B(n10945), .Z(n89) );
  NAND U176 ( .A(n88), .B(n89), .Z(n11268) );
  XNOR U177 ( .A(n11025), .B(n11026), .Z(n11028) );
  XOR U178 ( .A(n10756), .B(n10757), .Z(n90) );
  NANDN U179 ( .A(n10758), .B(n90), .Z(n91) );
  NAND U180 ( .A(n10756), .B(n10757), .Z(n92) );
  AND U181 ( .A(n91), .B(n92), .Z(n10865) );
  XNOR U182 ( .A(n11773), .B(n11772), .Z(n11771) );
  XOR U183 ( .A(n12425), .B(n12424), .Z(n12401) );
  XNOR U184 ( .A(n12407), .B(n12406), .Z(n12464) );
  XNOR U185 ( .A(n12516), .B(n12515), .Z(n12513) );
  XNOR U186 ( .A(n12502), .B(n12501), .Z(n12499) );
  XNOR U187 ( .A(n13153), .B(n13152), .Z(n13210) );
  NAND U188 ( .A(n14444), .B(n14443), .Z(n93) );
  NAND U189 ( .A(n14442), .B(n14441), .Z(n94) );
  AND U190 ( .A(n93), .B(n94), .Z(n14515) );
  XNOR U191 ( .A(n14915), .B(n14916), .Z(n14910) );
  XNOR U192 ( .A(n15241), .B(n15240), .Z(n15243) );
  XOR U193 ( .A(n15648), .B(n15649), .Z(n15642) );
  NAND U194 ( .A(n15363), .B(n15362), .Z(n95) );
  NAND U195 ( .A(n15360), .B(n15361), .Z(n96) );
  NAND U196 ( .A(n95), .B(n96), .Z(n15654) );
  XNOR U197 ( .A(n16017), .B(n16016), .Z(n16019) );
  XNOR U198 ( .A(n16043), .B(n16042), .Z(n16100) );
  NAND U199 ( .A(n16882), .B(n16883), .Z(n97) );
  NAND U200 ( .A(n16966), .B(n16884), .Z(n98) );
  AND U201 ( .A(n97), .B(n98), .Z(n99) );
  NAND U202 ( .A(n16885), .B(n16886), .Z(n100) );
  NAND U203 ( .A(n16887), .B(n16888), .Z(n101) );
  NAND U204 ( .A(n100), .B(n101), .Z(n102) );
  XNOR U205 ( .A(n99), .B(n102), .Z(n16889) );
  NAND U206 ( .A(n16695), .B(n16694), .Z(n103) );
  NANDN U207 ( .A(n16693), .B(n16692), .Z(n104) );
  AND U208 ( .A(n103), .B(n104), .Z(n17074) );
  XNOR U209 ( .A(n17438), .B(n17437), .Z(n17440) );
  XNOR U210 ( .A(n19072), .B(n19071), .Z(n19070) );
  XOR U211 ( .A(n3058), .B(n3057), .Z(n3033) );
  NAND U212 ( .A(n3627), .B(n3626), .Z(n105) );
  NANDN U213 ( .A(n3625), .B(n3624), .Z(n106) );
  AND U214 ( .A(n105), .B(n106), .Z(n3774) );
  NAND U215 ( .A(n4364), .B(n4363), .Z(n107) );
  NAND U216 ( .A(n4361), .B(n4362), .Z(n108) );
  AND U217 ( .A(n107), .B(n108), .Z(n4487) );
  NAND U218 ( .A(n5228), .B(n5229), .Z(n109) );
  NANDN U219 ( .A(n5231), .B(n5230), .Z(n110) );
  AND U220 ( .A(n109), .B(n110), .Z(n111) );
  NAND U221 ( .A(n5233), .B(n5232), .Z(n112) );
  NAND U222 ( .A(n5234), .B(n5235), .Z(n113) );
  AND U223 ( .A(n112), .B(n113), .Z(n114) );
  NAND U224 ( .A(n5237), .B(n5236), .Z(n115) );
  NANDN U225 ( .A(n5239), .B(n5238), .Z(n116) );
  AND U226 ( .A(n115), .B(n116), .Z(n117) );
  AND U227 ( .A(n5357), .B(n5356), .Z(n118) );
  XNOR U228 ( .A(n5351), .B(n5350), .Z(n119) );
  XNOR U229 ( .A(n118), .B(n119), .Z(n120) );
  AND U230 ( .A(n5245), .B(n5244), .Z(n121) );
  XNOR U231 ( .A(n5455), .B(n120), .Z(n122) );
  XNOR U232 ( .A(n121), .B(n122), .Z(n123) );
  XOR U233 ( .A(n117), .B(n123), .Z(n124) );
  XNOR U234 ( .A(n111), .B(n114), .Z(n125) );
  XNOR U235 ( .A(n124), .B(n125), .Z(n5456) );
  XNOR U236 ( .A(n6674), .B(n6673), .Z(n6672) );
  XNOR U237 ( .A(n8866), .B(n8865), .Z(n8864) );
  XNOR U238 ( .A(n9852), .B(n9851), .Z(n9850) );
  XNOR U239 ( .A(n10572), .B(n10571), .Z(n10570) );
  NAND U240 ( .A(n10991), .B(n10990), .Z(n126) );
  NANDN U241 ( .A(n10993), .B(n10992), .Z(n127) );
  NAND U242 ( .A(n126), .B(n127), .Z(n11289) );
  XNOR U243 ( .A(n12762), .B(n12761), .Z(n12488) );
  XNOR U244 ( .A(n13227), .B(n13226), .Z(n13225) );
  NAND U245 ( .A(n13830), .B(n13829), .Z(n128) );
  NAND U246 ( .A(n13827), .B(n13828), .Z(n129) );
  AND U247 ( .A(n128), .B(n129), .Z(n13921) );
  NAND U248 ( .A(n14521), .B(n14520), .Z(n130) );
  NANDN U249 ( .A(n14523), .B(n14522), .Z(n131) );
  AND U250 ( .A(n130), .B(n131), .Z(n14671) );
  XNOR U251 ( .A(n15376), .B(n15375), .Z(n15373) );
  NAND U252 ( .A(n16715), .B(n16714), .Z(n132) );
  NAND U253 ( .A(n16712), .B(n16713), .Z(n133) );
  AND U254 ( .A(n132), .B(n133), .Z(n16838) );
  NAND U255 ( .A(n18144), .B(n18143), .Z(n134) );
  NANDN U256 ( .A(n18142), .B(n18141), .Z(n135) );
  AND U257 ( .A(n134), .B(n135), .Z(n18269) );
  NAND U258 ( .A(n18885), .B(n18884), .Z(n136) );
  NANDN U259 ( .A(n18883), .B(n18882), .Z(n137) );
  AND U260 ( .A(n136), .B(n137), .Z(n19033) );
  XNOR U261 ( .A(n4919), .B(n4918), .Z(n4920) );
  XNOR U262 ( .A(n6377), .B(n6376), .Z(n6378) );
  XNOR U263 ( .A(n17957), .B(n17956), .Z(n17958) );
  XNOR U264 ( .A(n3646), .B(n3585), .Z(n3594) );
  XOR U265 ( .A(n3581), .B(n3580), .Z(n3550) );
  NAND U266 ( .A(n4231), .B(n4230), .Z(n138) );
  NANDN U267 ( .A(n4233), .B(n4232), .Z(n139) );
  AND U268 ( .A(n138), .B(n139), .Z(n4321) );
  NAND U269 ( .A(n4864), .B(n4865), .Z(n140) );
  NAND U270 ( .A(n5005), .B(n5002), .Z(n141) );
  NAND U271 ( .A(n140), .B(n141), .Z(n4894) );
  XNOR U272 ( .A(n5758), .B(n5757), .Z(n5760) );
  NAND U273 ( .A(n6322), .B(n6323), .Z(n142) );
  NAND U274 ( .A(n6465), .B(n6461), .Z(n143) );
  NAND U275 ( .A(n142), .B(n143), .Z(n6352) );
  NAND U276 ( .A(n7776), .B(n7777), .Z(n144) );
  NAND U277 ( .A(n7916), .B(n7919), .Z(n145) );
  NAND U278 ( .A(n144), .B(n145), .Z(n7806) );
  XNOR U279 ( .A(n7953), .B(n7952), .Z(n7955) );
  NAND U280 ( .A(n9230), .B(n9231), .Z(n146) );
  NAND U281 ( .A(n9353), .B(n9368), .Z(n147) );
  NAND U282 ( .A(n146), .B(n147), .Z(n9260) );
  XNOR U283 ( .A(n9286), .B(n9285), .Z(n9287) );
  XNOR U284 ( .A(n9305), .B(n9304), .Z(n9291) );
  NAND U285 ( .A(n9950), .B(n9951), .Z(n148) );
  NAND U286 ( .A(n10084), .B(n10087), .Z(n149) );
  NAND U287 ( .A(n148), .B(n149), .Z(n9980) );
  XNOR U288 ( .A(n10006), .B(n10005), .Z(n10007) );
  NAND U289 ( .A(n10645), .B(n10644), .Z(n150) );
  NAND U290 ( .A(n10642), .B(n10643), .Z(n151) );
  NAND U291 ( .A(n150), .B(n151), .Z(n10707) );
  NAND U292 ( .A(n10730), .B(n10729), .Z(n152) );
  NAND U293 ( .A(n10727), .B(n10728), .Z(n153) );
  AND U294 ( .A(n152), .B(n153), .Z(n10796) );
  XNOR U295 ( .A(n12379), .B(n12378), .Z(n12380) );
  XNOR U296 ( .A(n12384), .B(n12383), .Z(n12385) );
  XNOR U297 ( .A(n12312), .B(n12311), .Z(n12313) );
  XNOR U298 ( .A(n12999), .B(n12998), .Z(n13000) );
  XNOR U299 ( .A(n13037), .B(n13036), .Z(n13039) );
  XNOR U300 ( .A(n12989), .B(n12988), .Z(n13042) );
  XNOR U301 ( .A(n15041), .B(n15040), .Z(n15043) );
  NAND U302 ( .A(n15758), .B(n15759), .Z(n154) );
  NAND U303 ( .A(n15902), .B(n15901), .Z(n155) );
  NAND U304 ( .A(n154), .B(n155), .Z(n15788) );
  XNOR U305 ( .A(n15932), .B(n15931), .Z(n15934) );
  NAND U306 ( .A(n16584), .B(n16583), .Z(n156) );
  NANDN U307 ( .A(n16586), .B(n16585), .Z(n157) );
  AND U308 ( .A(n156), .B(n157), .Z(n16672) );
  XNOR U309 ( .A(n17357), .B(n17356), .Z(n17359) );
  NAND U310 ( .A(n17914), .B(n17915), .Z(n158) );
  NAND U311 ( .A(n18055), .B(n18059), .Z(n159) );
  NAND U312 ( .A(n158), .B(n159), .Z(n17944) );
  NAND U313 ( .A(n1389), .B(n1388), .Z(n160) );
  NANDN U314 ( .A(n1391), .B(n1390), .Z(n161) );
  NAND U315 ( .A(n160), .B(n161), .Z(n1485) );
  NAND U316 ( .A(n1458), .B(n1723), .Z(n162) );
  NAND U317 ( .A(n1457), .B(n1456), .Z(n163) );
  AND U318 ( .A(n162), .B(n163), .Z(n1758) );
  NAND U319 ( .A(n1447), .B(n1448), .Z(n164) );
  NAND U320 ( .A(n1511), .B(n1446), .Z(n165) );
  AND U321 ( .A(n164), .B(n165), .Z(n1741) );
  NAND U322 ( .A(n2934), .B(n2933), .Z(n166) );
  NAND U323 ( .A(n2931), .B(n2932), .Z(n167) );
  NAND U324 ( .A(n166), .B(n167), .Z(n3179) );
  NAND U325 ( .A(n2937), .B(n2936), .Z(n168) );
  NANDN U326 ( .A(n2935), .B(n3145), .Z(n169) );
  AND U327 ( .A(n168), .B(n169), .Z(n3264) );
  XNOR U328 ( .A(n3613), .B(n3612), .Z(n3614) );
  XNOR U329 ( .A(n3619), .B(n3618), .Z(n3620) );
  XNOR U330 ( .A(n3643), .B(n3642), .Z(n3723) );
  NAND U331 ( .A(n4318), .B(n4317), .Z(n170) );
  NAND U332 ( .A(n4315), .B(n4316), .Z(n171) );
  NAND U333 ( .A(n170), .B(n171), .Z(n4411) );
  XOR U334 ( .A(n5364), .B(n5365), .Z(n5366) );
  XNOR U335 ( .A(n5796), .B(n5795), .Z(n5798) );
  XNOR U336 ( .A(n5836), .B(n5835), .Z(n5880) );
  XNOR U337 ( .A(n6511), .B(n6510), .Z(n6513) );
  XNOR U338 ( .A(n6539), .B(n6538), .Z(n6540) );
  NAND U339 ( .A(n7297), .B(n7341), .Z(n172) );
  NANDN U340 ( .A(n7215), .B(n7214), .Z(n173) );
  AND U341 ( .A(n172), .B(n173), .Z(n7328) );
  NAND U342 ( .A(n7257), .B(n7256), .Z(n174) );
  NAND U343 ( .A(n7254), .B(n7255), .Z(n175) );
  NAND U344 ( .A(n174), .B(n175), .Z(n7266) );
  XNOR U345 ( .A(n7993), .B(n7992), .Z(n8050) );
  XNOR U346 ( .A(n7985), .B(n7984), .Z(n7987) );
  XNOR U347 ( .A(n9422), .B(n9421), .Z(n9415) );
  NAND U348 ( .A(n9408), .B(n9407), .Z(n176) );
  NAND U349 ( .A(n9405), .B(n9406), .Z(n177) );
  NAND U350 ( .A(n176), .B(n177), .Z(n9508) );
  XNOR U351 ( .A(n9804), .B(n9803), .Z(n9801) );
  XNOR U352 ( .A(n10140), .B(n10139), .Z(n10133) );
  NAND U353 ( .A(n10181), .B(n10180), .Z(n178) );
  AND U354 ( .A(n10179), .B(y[59]), .Z(n179) );
  NAND U355 ( .A(x[91]), .B(n179), .Z(n180) );
  AND U356 ( .A(n178), .B(n180), .Z(n10521) );
  AND U357 ( .A(n10717), .B(n10716), .Z(n181) );
  AND U358 ( .A(n10715), .B(x[99]), .Z(n182) );
  NAND U359 ( .A(y[105]), .B(n182), .Z(n183) );
  NANDN U360 ( .A(n181), .B(n183), .Z(n10848) );
  NAND U361 ( .A(n10841), .B(n10840), .Z(n184) );
  NANDN U362 ( .A(n10843), .B(n10842), .Z(n185) );
  AND U363 ( .A(n184), .B(n185), .Z(n10941) );
  XNOR U364 ( .A(n12332), .B(n12331), .Z(n12334) );
  XNOR U365 ( .A(n12728), .B(n12727), .Z(n12725) );
  XNOR U366 ( .A(n12453), .B(n12452), .Z(n12337) );
  XNOR U367 ( .A(n12405), .B(n12404), .Z(n12406) );
  XOR U368 ( .A(n13029), .B(n13028), .Z(n12983) );
  NAND U369 ( .A(n13107), .B(n13162), .Z(n186) );
  NANDN U370 ( .A(n13014), .B(n13013), .Z(n187) );
  AND U371 ( .A(n186), .B(n187), .Z(n13144) );
  XNOR U372 ( .A(n13093), .B(n13092), .Z(n13132) );
  XOR U373 ( .A(n13380), .B(n13379), .Z(n13378) );
  XNOR U374 ( .A(n13109), .B(n13108), .Z(n13181) );
  NAND U375 ( .A(n13765), .B(n13764), .Z(n188) );
  NANDN U376 ( .A(n13767), .B(n13766), .Z(n189) );
  AND U377 ( .A(n188), .B(n189), .Z(n13850) );
  XNOR U378 ( .A(n14138), .B(n14137), .Z(n14135) );
  XNOR U379 ( .A(n14144), .B(n14143), .Z(n14141) );
  XNOR U380 ( .A(n14895), .B(n14896), .Z(n14897) );
  NAND U381 ( .A(n15225), .B(n15224), .Z(n190) );
  NAND U382 ( .A(n15222), .B(n15223), .Z(n191) );
  NAND U383 ( .A(n190), .B(n191), .Z(n15360) );
  XNOR U384 ( .A(n15970), .B(n15969), .Z(n15972) );
  XNOR U385 ( .A(n16010), .B(n16009), .Z(n16071) );
  NAND U386 ( .A(n16669), .B(n16668), .Z(n192) );
  NAND U387 ( .A(n16666), .B(n16667), .Z(n193) );
  NAND U388 ( .A(n192), .B(n193), .Z(n16761) );
  XNOR U389 ( .A(n17389), .B(n17388), .Z(n17391) );
  XNOR U390 ( .A(n17430), .B(n17429), .Z(n17474) );
  XNOR U391 ( .A(n18108), .B(n18107), .Z(n18110) );
  XNOR U392 ( .A(n18166), .B(n18165), .Z(n18167) );
  XNOR U393 ( .A(n18136), .B(n18135), .Z(n18137) );
  NAND U394 ( .A(n1475), .B(n1474), .Z(n194) );
  NAND U395 ( .A(n1472), .B(n1473), .Z(n195) );
  AND U396 ( .A(n194), .B(n195), .Z(n1545) );
  XOR U397 ( .A(n2148), .B(n2147), .Z(n2150) );
  XNOR U398 ( .A(n2331), .B(n2330), .Z(n2329) );
  NAND U399 ( .A(n2974), .B(n2973), .Z(n196) );
  NAND U400 ( .A(n2971), .B(n2972), .Z(n197) );
  AND U401 ( .A(n196), .B(n197), .Z(n3051) );
  XOR U402 ( .A(n3039), .B(n3038), .Z(n3037) );
  NAND U403 ( .A(n2927), .B(n2926), .Z(n198) );
  NAND U404 ( .A(n2924), .B(n2925), .Z(n199) );
  NAND U405 ( .A(n198), .B(n199), .Z(n3177) );
  NAND U406 ( .A(n2978), .B(n2977), .Z(n200) );
  NAND U407 ( .A(n2976), .B(n2975), .Z(n201) );
  AND U408 ( .A(n200), .B(n201), .Z(n3290) );
  XOR U409 ( .A(n3750), .B(n3749), .Z(n3759) );
  XNOR U410 ( .A(n4466), .B(n4465), .Z(n4343) );
  NAND U411 ( .A(n4268), .B(n4267), .Z(n202) );
  NANDN U412 ( .A(n4266), .B(n4265), .Z(n203) );
  NAND U413 ( .A(n202), .B(n203), .Z(n4346) );
  XNOR U414 ( .A(n4769), .B(n4768), .Z(n4758) );
  XNOR U415 ( .A(n5231), .B(n5230), .Z(n5229) );
  XNOR U416 ( .A(n5481), .B(n5480), .Z(n5479) );
  NAND U417 ( .A(n5073), .B(n5072), .Z(n204) );
  NANDN U418 ( .A(n5071), .B(n5070), .Z(n205) );
  AND U419 ( .A(n204), .B(n205), .Z(n5475) );
  XOR U420 ( .A(n5876), .B(n5875), .Z(n5928) );
  NAND U421 ( .A(n5782), .B(n5781), .Z(n206) );
  NANDN U422 ( .A(n5780), .B(n5779), .Z(n207) );
  AND U423 ( .A(n206), .B(n207), .Z(n5922) );
  XNOR U424 ( .A(n5961), .B(n5962), .Z(n5964) );
  XNOR U425 ( .A(n6945), .B(n6944), .Z(n6943) );
  NAND U426 ( .A(n7308), .B(n7307), .Z(n208) );
  NANDN U427 ( .A(n7436), .B(n7310), .Z(n209) );
  AND U428 ( .A(n208), .B(n209), .Z(n7607) );
  NAND U429 ( .A(n7263), .B(n7262), .Z(n210) );
  NANDN U430 ( .A(n7265), .B(n7264), .Z(n211) );
  AND U431 ( .A(n210), .B(n211), .Z(n7655) );
  XOR U432 ( .A(n8065), .B(n8064), .Z(n8117) );
  NAND U433 ( .A(n7971), .B(n7970), .Z(n212) );
  NANDN U434 ( .A(n7969), .B(n7968), .Z(n213) );
  AND U435 ( .A(n212), .B(n213), .Z(n8111) );
  XOR U436 ( .A(n8141), .B(n8140), .Z(n8139) );
  XNOR U437 ( .A(n8739), .B(n8738), .Z(n8741) );
  NAND U438 ( .A(n9052), .B(n9051), .Z(n214) );
  NAND U439 ( .A(n9053), .B(n9054), .Z(n215) );
  AND U440 ( .A(n214), .B(n215), .Z(n216) );
  NAND U441 ( .A(n9058), .B(n9057), .Z(n217) );
  NAND U442 ( .A(n9055), .B(n9056), .Z(n218) );
  NAND U443 ( .A(n217), .B(n218), .Z(n219) );
  XNOR U444 ( .A(n216), .B(n219), .Z(n9059) );
  XNOR U445 ( .A(n9132), .B(n9131), .Z(n9130) );
  NAND U446 ( .A(n8725), .B(n8724), .Z(n220) );
  NANDN U447 ( .A(n8723), .B(n8722), .Z(n221) );
  AND U448 ( .A(n220), .B(n221), .Z(n9126) );
  XNOR U449 ( .A(n9450), .B(n9449), .Z(n9490) );
  XNOR U450 ( .A(n9821), .B(n9822), .Z(n9816) );
  NAND U451 ( .A(n9460), .B(n9459), .Z(n222) );
  NAND U452 ( .A(n9457), .B(n9458), .Z(n223) );
  NAND U453 ( .A(n222), .B(n223), .Z(n9595) );
  NAND U454 ( .A(n10178), .B(n10177), .Z(n224) );
  NAND U455 ( .A(n10175), .B(n10176), .Z(n225) );
  NAND U456 ( .A(n224), .B(n225), .Z(n10314) );
  XNOR U457 ( .A(n11275), .B(n11274), .Z(n11273) );
  XOR U458 ( .A(n11021), .B(n11022), .Z(n11020) );
  NAND U459 ( .A(n11610), .B(n11609), .Z(n226) );
  NAND U460 ( .A(n11607), .B(n11608), .Z(n227) );
  NAND U461 ( .A(n226), .B(n227), .Z(n11766) );
  NAND U462 ( .A(n12224), .B(n12223), .Z(n228) );
  XOR U463 ( .A(n12224), .B(n12223), .Z(n229) );
  NANDN U464 ( .A(n12225), .B(n229), .Z(n230) );
  NAND U465 ( .A(n228), .B(n230), .Z(n12475) );
  XOR U466 ( .A(n12413), .B(n12412), .Z(n12465) );
  NAND U467 ( .A(n12320), .B(n12319), .Z(n231) );
  NANDN U468 ( .A(n12318), .B(n12317), .Z(n232) );
  AND U469 ( .A(n231), .B(n232), .Z(n12461) );
  XNOR U470 ( .A(n12747), .B(n12748), .Z(n12750) );
  XNOR U471 ( .A(n12770), .B(n12769), .Z(n12495) );
  XNOR U472 ( .A(n13241), .B(n13240), .Z(n13239) );
  XNOR U473 ( .A(n14179), .B(n14180), .Z(n14174) );
  XOR U474 ( .A(n13940), .B(n13939), .Z(n13938) );
  NAND U475 ( .A(n13900), .B(n13899), .Z(n233) );
  NANDN U476 ( .A(n13902), .B(n13901), .Z(n234) );
  NAND U477 ( .A(n233), .B(n234), .Z(n14192) );
  XNOR U478 ( .A(n14582), .B(n14581), .Z(n14516) );
  NAND U479 ( .A(n15249), .B(n15248), .Z(n235) );
  NAND U480 ( .A(n15246), .B(n15247), .Z(n236) );
  NAND U481 ( .A(n235), .B(n236), .Z(n15401) );
  XNOR U482 ( .A(n15231), .B(n15230), .Z(n15233) );
  XOR U483 ( .A(n16049), .B(n16048), .Z(n16101) );
  NAND U484 ( .A(n15956), .B(n15955), .Z(n237) );
  NANDN U485 ( .A(n15954), .B(n15953), .Z(n238) );
  AND U486 ( .A(n237), .B(n238), .Z(n16095) );
  XNOR U487 ( .A(n16131), .B(n16130), .Z(n16129) );
  XNOR U488 ( .A(n16817), .B(n16816), .Z(n16694) );
  NAND U489 ( .A(n16612), .B(n16611), .Z(n239) );
  NANDN U490 ( .A(n16614), .B(n16613), .Z(n240) );
  NAND U491 ( .A(n239), .B(n240), .Z(n16697) );
  NAND U492 ( .A(n16875), .B(n16874), .Z(n241) );
  NAND U493 ( .A(n16876), .B(n16877), .Z(n242) );
  AND U494 ( .A(n241), .B(n242), .Z(n243) );
  NAND U495 ( .A(n16879), .B(n16878), .Z(n244) );
  NAND U496 ( .A(n16880), .B(n16881), .Z(n245) );
  NAND U497 ( .A(n244), .B(n245), .Z(n246) );
  XNOR U498 ( .A(n243), .B(n246), .Z(n16890) );
  XNOR U499 ( .A(n17084), .B(n17083), .Z(n17073) );
  XOR U500 ( .A(n17470), .B(n17469), .Z(n17522) );
  NAND U501 ( .A(n17375), .B(n17374), .Z(n247) );
  NANDN U502 ( .A(n17373), .B(n17372), .Z(n248) );
  AND U503 ( .A(n247), .B(n248), .Z(n17516) );
  XNOR U504 ( .A(n17555), .B(n17556), .Z(n17558) );
  XNOR U505 ( .A(n18180), .B(n18179), .Z(n18145) );
  XNOR U506 ( .A(n18967), .B(n18966), .Z(n19019) );
  XNOR U507 ( .A(n19313), .B(n19312), .Z(n19311) );
  XNOR U508 ( .A(n19065), .B(n19066), .Z(n19064) );
  NAND U509 ( .A(n1523), .B(n1522), .Z(n249) );
  NAND U510 ( .A(n1520), .B(n1521), .Z(n250) );
  AND U511 ( .A(n249), .B(n250), .Z(n1830) );
  NAND U512 ( .A(n2905), .B(n2904), .Z(n251) );
  NANDN U513 ( .A(n2903), .B(n2902), .Z(n252) );
  NAND U514 ( .A(n251), .B(n252), .Z(n3317) );
  NAND U515 ( .A(n3791), .B(n3790), .Z(n253) );
  NANDN U516 ( .A(n3793), .B(n3792), .Z(n254) );
  AND U517 ( .A(n253), .B(n254), .Z(n255) );
  AND U518 ( .A(n3911), .B(n3910), .Z(n256) );
  NAND U519 ( .A(n3905), .B(n3904), .Z(n257) );
  XNOR U520 ( .A(n256), .B(n257), .Z(n258) );
  AND U521 ( .A(n3798), .B(n3797), .Z(n259) );
  XNOR U522 ( .A(n3899), .B(n3898), .Z(n260) );
  XNOR U523 ( .A(n259), .B(n260), .Z(n261) );
  XNOR U524 ( .A(n255), .B(n258), .Z(n262) );
  XNOR U525 ( .A(n261), .B(n262), .Z(n263) );
  NANDN U526 ( .A(n3788), .B(n3789), .Z(n264) );
  XNOR U527 ( .A(n3788), .B(n3789), .Z(n265) );
  NAND U528 ( .A(n3787), .B(n265), .Z(n266) );
  NAND U529 ( .A(n264), .B(n266), .Z(n267) );
  XNOR U530 ( .A(n263), .B(n267), .Z(n268) );
  NAND U531 ( .A(n3784), .B(n3783), .Z(n269) );
  NANDN U532 ( .A(n3786), .B(n3785), .Z(n270) );
  NAND U533 ( .A(n269), .B(n270), .Z(n271) );
  XNOR U534 ( .A(n268), .B(n271), .Z(n4023) );
  NAND U535 ( .A(n4360), .B(n4359), .Z(n272) );
  NAND U536 ( .A(n4357), .B(n4358), .Z(n273) );
  AND U537 ( .A(n272), .B(n273), .Z(n4488) );
  NAND U538 ( .A(n5112), .B(n5111), .Z(n274) );
  NAND U539 ( .A(n5109), .B(n5110), .Z(n275) );
  NAND U540 ( .A(n274), .B(n275), .Z(n5220) );
  XNOR U541 ( .A(n6219), .B(n6220), .Z(n6218) );
  XNOR U542 ( .A(n5944), .B(n5943), .Z(n5942) );
  XNOR U543 ( .A(n6957), .B(n6956), .Z(n6955) );
  XNOR U544 ( .A(n8408), .B(n8407), .Z(n8406) );
  XNOR U545 ( .A(n8133), .B(n8132), .Z(n8131) );
  NAND U546 ( .A(n8872), .B(n8871), .Z(n276) );
  NANDN U547 ( .A(n8874), .B(n8873), .Z(n277) );
  AND U548 ( .A(n276), .B(n277), .Z(n9108) );
  XNOR U549 ( .A(n9834), .B(n9833), .Z(n9832) );
  XNOR U550 ( .A(n10554), .B(n10553), .Z(n10552) );
  XNOR U551 ( .A(n10861), .B(n10860), .Z(n10866) );
  XNOR U552 ( .A(n11287), .B(n11286), .Z(n11004) );
  NAND U553 ( .A(n11650), .B(n11649), .Z(n278) );
  NANDN U554 ( .A(n11648), .B(n11647), .Z(n279) );
  AND U555 ( .A(n278), .B(n279), .Z(n11742) );
  XNOR U556 ( .A(n12488), .B(n12487), .Z(n12486) );
  NAND U557 ( .A(n13211), .B(n13210), .Z(n280) );
  NAND U558 ( .A(n13212), .B(n13213), .Z(n281) );
  NAND U559 ( .A(n280), .B(n281), .Z(n13221) );
  XNOR U560 ( .A(n13922), .B(n13921), .Z(n13920) );
  NAND U561 ( .A(n14923), .B(n14924), .Z(n14928) );
  XNOR U562 ( .A(n15663), .B(n15662), .Z(n15658) );
  XNOR U563 ( .A(n16392), .B(n16393), .Z(n16391) );
  XNOR U564 ( .A(n16117), .B(n16116), .Z(n16115) );
  NAND U565 ( .A(n16711), .B(n16710), .Z(n282) );
  NAND U566 ( .A(n16708), .B(n16709), .Z(n283) );
  AND U567 ( .A(n282), .B(n283), .Z(n16839) );
  XNOR U568 ( .A(n17813), .B(n17814), .Z(n17812) );
  XNOR U569 ( .A(n17538), .B(n17537), .Z(n17536) );
  XNOR U570 ( .A(n18554), .B(n18553), .Z(n18552) );
  XNOR U571 ( .A(n19305), .B(n19304), .Z(n19037) );
  XNOR U572 ( .A(n4939), .B(n4938), .Z(n4924) );
  XNOR U573 ( .A(n8568), .B(n8567), .Z(n8569) );
  XNOR U574 ( .A(n8588), .B(n8587), .Z(n8573) );
  XOR U575 ( .A(n1377), .B(n1376), .Z(n1331) );
  XOR U576 ( .A(n2100), .B(n2099), .Z(n2075) );
  XOR U577 ( .A(n2090), .B(n2089), .Z(n2069) );
  XNOR U578 ( .A(n3471), .B(n3470), .Z(n3472) );
  XNOR U579 ( .A(n3500), .B(n3499), .Z(n3476) );
  NAND U580 ( .A(n3412), .B(n3413), .Z(n284) );
  NAND U581 ( .A(n3546), .B(n3561), .Z(n285) );
  NAND U582 ( .A(n284), .B(n285), .Z(n3444) );
  XNOR U583 ( .A(n3595), .B(n3594), .Z(n3597) );
  NAND U584 ( .A(n4152), .B(n4153), .Z(n286) );
  NAND U585 ( .A(n4282), .B(n4285), .Z(n287) );
  NAND U586 ( .A(n286), .B(n287), .Z(n4182) );
  XNOR U587 ( .A(n4225), .B(n4224), .Z(n4210) );
  XNOR U588 ( .A(n4921), .B(n4920), .Z(n4896) );
  XNOR U589 ( .A(n5710), .B(n5709), .Z(n5764) );
  XOR U590 ( .A(n7227), .B(n7226), .Z(n7186) );
  AND U591 ( .A(n7123), .B(n7122), .Z(n288) );
  AND U592 ( .A(n7121), .B(x[59]), .Z(n289) );
  NAND U593 ( .A(y[105]), .B(n289), .Z(n290) );
  NANDN U594 ( .A(n288), .B(n290), .Z(n7254) );
  NAND U595 ( .A(n8068), .B(n8024), .Z(n291) );
  NANDN U596 ( .A(n7925), .B(n7924), .Z(n292) );
  AND U597 ( .A(n291), .B(n292), .Z(n8044) );
  XNOR U598 ( .A(n7913), .B(n7912), .Z(n7959) );
  NAND U599 ( .A(n8503), .B(n8504), .Z(n293) );
  NAND U600 ( .A(n8658), .B(n8655), .Z(n294) );
  NAND U601 ( .A(n293), .B(n294), .Z(n8541) );
  XNOR U602 ( .A(n9392), .B(n9391), .Z(n9393) );
  XNOR U603 ( .A(n10110), .B(n10109), .Z(n10111) );
  NAND U604 ( .A(n10698), .B(n10697), .Z(n295) );
  NAND U605 ( .A(n10695), .B(n10696), .Z(n296) );
  AND U606 ( .A(n295), .B(n296), .Z(n10792) );
  NAND U607 ( .A(n11376), .B(n11377), .Z(n297) );
  NAND U608 ( .A(n11531), .B(n11530), .Z(n298) );
  NAND U609 ( .A(n297), .B(n298), .Z(n11414) );
  XNOR U610 ( .A(n12290), .B(n12289), .Z(n12291) );
  XOR U611 ( .A(n12281), .B(n12280), .Z(n12237) );
  XNOR U612 ( .A(n12260), .B(n12259), .Z(n12261) );
  XNOR U613 ( .A(n12300), .B(n12299), .Z(n12302) );
  NAND U614 ( .A(n12864), .B(n12865), .Z(n299) );
  NAND U615 ( .A(n13008), .B(n13005), .Z(n300) );
  NAND U616 ( .A(n299), .B(n300), .Z(n12894) );
  XNOR U617 ( .A(n13001), .B(n13000), .Z(n13043) );
  NAND U618 ( .A(n13662), .B(n13661), .Z(n301) );
  NAND U619 ( .A(n13659), .B(n13660), .Z(n302) );
  AND U620 ( .A(n301), .B(n302), .Z(n13774) );
  NAND U621 ( .A(n13821), .B(n13881), .Z(n303) );
  NANDN U622 ( .A(n13744), .B(n13743), .Z(n304) );
  AND U623 ( .A(n303), .B(n304), .Z(n13838) );
  NAND U624 ( .A(n14074), .B(n13762), .Z(n305) );
  NAND U625 ( .A(n13763), .B(n13804), .Z(n306) );
  NAND U626 ( .A(n305), .B(n306), .Z(n13833) );
  NAND U627 ( .A(n13658), .B(n13654), .Z(n307) );
  NAND U628 ( .A(n13655), .B(n13656), .Z(n308) );
  NAND U629 ( .A(n307), .B(n308), .Z(n13780) );
  XNOR U630 ( .A(n15024), .B(n15025), .Z(n14991) );
  NAND U631 ( .A(n15069), .B(n15068), .Z(n309) );
  NAND U632 ( .A(n15066), .B(n15067), .Z(n310) );
  AND U633 ( .A(n309), .B(n310), .Z(n15227) );
  XNOR U634 ( .A(n15896), .B(n15895), .Z(n15938) );
  XNOR U635 ( .A(n16578), .B(n16577), .Z(n16555) );
  NAND U636 ( .A(n17180), .B(n17181), .Z(n311) );
  NAND U637 ( .A(n17320), .B(n17323), .Z(n312) );
  NAND U638 ( .A(n311), .B(n312), .Z(n17210) );
  XNOR U639 ( .A(n17316), .B(n17315), .Z(n17363) );
  XOR U640 ( .A(n18828), .B(n18827), .Z(n18787) );
  XOR U641 ( .A(n18839), .B(n18838), .Z(n18793) );
  NAND U642 ( .A(n1455), .B(n1685), .Z(n313) );
  NAND U643 ( .A(n1453), .B(n1454), .Z(n314) );
  AND U644 ( .A(n313), .B(n314), .Z(n1759) );
  NAND U645 ( .A(n1445), .B(n1444), .Z(n315) );
  NAND U646 ( .A(n1443), .B(n1442), .Z(n316) );
  AND U647 ( .A(n315), .B(n316), .Z(n1753) );
  NAND U648 ( .A(n1515), .B(n1514), .Z(n317) );
  NAND U649 ( .A(n1513), .B(n1512), .Z(n318) );
  AND U650 ( .A(n317), .B(n318), .Z(n1613) );
  NAND U651 ( .A(n1342), .B(n1341), .Z(n319) );
  NAND U652 ( .A(n1339), .B(n1340), .Z(n320) );
  NAND U653 ( .A(n319), .B(n320), .Z(n1451) );
  NAND U654 ( .A(n1346), .B(n1345), .Z(n321) );
  NAND U655 ( .A(n1343), .B(n1344), .Z(n322) );
  NAND U656 ( .A(n321), .B(n322), .Z(n1508) );
  NAND U657 ( .A(n1338), .B(n1337), .Z(n323) );
  NANDN U658 ( .A(n1461), .B(n1336), .Z(n324) );
  NAND U659 ( .A(n323), .B(n324), .Z(n1432) );
  XOR U660 ( .A(n3267), .B(n3266), .Z(n3265) );
  XNOR U661 ( .A(n3748), .B(n3747), .Z(n3749) );
  XNOR U662 ( .A(n3921), .B(n3920), .Z(n3918) );
  NAND U663 ( .A(n3729), .B(n3667), .Z(n325) );
  NANDN U664 ( .A(n3567), .B(n3566), .Z(n326) );
  AND U665 ( .A(n325), .B(n326), .Z(n3687) );
  XNOR U666 ( .A(n3676), .B(n3675), .Z(n3677) );
  NAND U667 ( .A(n4201), .B(n4200), .Z(n327) );
  NANDN U668 ( .A(n4203), .B(n4202), .Z(n328) );
  AND U669 ( .A(n327), .B(n328), .Z(n4261) );
  XNOR U670 ( .A(n4637), .B(n4636), .Z(n4634) );
  XNOR U671 ( .A(n5360), .B(n5361), .Z(n5358) );
  XNOR U672 ( .A(n5081), .B(n5080), .Z(n5082) );
  XNOR U673 ( .A(n5075), .B(n5074), .Z(n5076) );
  XOR U674 ( .A(n5750), .B(n5749), .Z(n5723) );
  XNOR U675 ( .A(n5772), .B(n5771), .Z(n5786) );
  XOR U676 ( .A(n6182), .B(n6183), .Z(n6184) );
  NAND U677 ( .A(n5834), .B(n5908), .Z(n329) );
  NANDN U678 ( .A(n5735), .B(n5734), .Z(n330) );
  AND U679 ( .A(n329), .B(n330), .Z(n5855) );
  XNOR U680 ( .A(n5815), .B(n5814), .Z(n5862) );
  XNOR U681 ( .A(n5802), .B(n5801), .Z(n5803) );
  XNOR U682 ( .A(n6097), .B(n6096), .Z(n6094) );
  NAND U683 ( .A(n6355), .B(n6354), .Z(n331) );
  NANDN U684 ( .A(n6353), .B(n6352), .Z(n332) );
  AND U685 ( .A(n331), .B(n332), .Z(n6427) );
  XOR U686 ( .A(n6846), .B(n6845), .Z(n6844) );
  XOR U687 ( .A(n6835), .B(n6836), .Z(n6837) );
  XNOR U688 ( .A(n6533), .B(n6532), .Z(n6534) );
  NAND U689 ( .A(n7299), .B(n7298), .Z(n333) );
  NANDN U690 ( .A(n7297), .B(n7440), .Z(n334) );
  AND U691 ( .A(n333), .B(n334), .Z(n7457) );
  NAND U692 ( .A(n7211), .B(n7417), .Z(n335) );
  NAND U693 ( .A(n7212), .B(n7213), .Z(n336) );
  NAND U694 ( .A(n335), .B(n336), .Z(n7327) );
  NAND U695 ( .A(n7219), .B(n7218), .Z(n337) );
  NANDN U696 ( .A(n7221), .B(n7220), .Z(n338) );
  AND U697 ( .A(n337), .B(n338), .Z(n7317) );
  XOR U698 ( .A(n7939), .B(n7938), .Z(n7893) );
  XNOR U699 ( .A(n8005), .B(n8004), .Z(n8051) );
  XNOR U700 ( .A(n7949), .B(n7948), .Z(n7975) );
  XNOR U701 ( .A(n7991), .B(n7990), .Z(n7992) );
  XNOR U702 ( .A(n8363), .B(n8362), .Z(n8360) );
  XNOR U703 ( .A(n8026), .B(n8025), .Z(n8105) );
  XNOR U704 ( .A(n8713), .B(n8712), .Z(n8706) );
  XNOR U705 ( .A(n9082), .B(n9081), .Z(n9079) );
  XNOR U706 ( .A(n8733), .B(n8732), .Z(n8734) );
  XNOR U707 ( .A(n8727), .B(n8726), .Z(n8728) );
  NAND U708 ( .A(n9263), .B(n9262), .Z(n339) );
  NANDN U709 ( .A(n9261), .B(n9260), .Z(n340) );
  AND U710 ( .A(n339), .B(n340), .Z(n9336) );
  XNOR U711 ( .A(n9370), .B(n9369), .Z(n9362) );
  XOR U712 ( .A(n9382), .B(n9381), .Z(n9357) );
  XNOR U713 ( .A(n9414), .B(n9413), .Z(n9416) );
  NAND U714 ( .A(n9410), .B(n9409), .Z(n341) );
  NANDN U715 ( .A(n9412), .B(n9411), .Z(n342) );
  NAND U716 ( .A(n341), .B(n342), .Z(n9509) );
  NAND U717 ( .A(n9753), .B(n9397), .Z(n343) );
  NAND U718 ( .A(n9398), .B(n9461), .Z(n344) );
  NAND U719 ( .A(n343), .B(n344), .Z(n9496) );
  NAND U720 ( .A(n9983), .B(n9982), .Z(n345) );
  NANDN U721 ( .A(n9981), .B(n9980), .Z(n346) );
  AND U722 ( .A(n345), .B(n346), .Z(n10056) );
  XNOR U723 ( .A(n10089), .B(n10088), .Z(n10067) );
  XOR U724 ( .A(n10101), .B(n10100), .Z(n10062) );
  XNOR U725 ( .A(n10132), .B(n10131), .Z(n10134) );
  NAND U726 ( .A(n10128), .B(n10127), .Z(n347) );
  NANDN U727 ( .A(n10130), .B(n10129), .Z(n348) );
  NAND U728 ( .A(n347), .B(n348), .Z(n10228) );
  NAND U729 ( .A(n10472), .B(n10115), .Z(n349) );
  NAND U730 ( .A(n10116), .B(n10179), .Z(n350) );
  NAND U731 ( .A(n349), .B(n350), .Z(n10215) );
  NAND U732 ( .A(n10797), .B(n10796), .Z(n351) );
  NAND U733 ( .A(n10794), .B(n10795), .Z(n352) );
  NAND U734 ( .A(n351), .B(n352), .Z(n10917) );
  XNOR U735 ( .A(n11042), .B(n11041), .Z(n11039) );
  XOR U736 ( .A(n11161), .B(n11160), .Z(n11159) );
  NAND U737 ( .A(n10779), .B(n10778), .Z(n353) );
  NAND U738 ( .A(n10776), .B(n10777), .Z(n354) );
  NAND U739 ( .A(n353), .B(n354), .Z(n10893) );
  XOR U740 ( .A(n11988), .B(n11987), .Z(n11986) );
  XNOR U741 ( .A(n12549), .B(n12440), .Z(n12441) );
  XNOR U742 ( .A(n12707), .B(n12708), .Z(n12705) );
  XNOR U743 ( .A(n13051), .B(n13050), .Z(n13069) );
  XNOR U744 ( .A(n13462), .B(n13461), .Z(n13459) );
  XNOR U745 ( .A(n13098), .B(n13097), .Z(n13133) );
  XNOR U746 ( .A(n13091), .B(n13090), .Z(n13092) );
  XNOR U747 ( .A(n13079), .B(n13078), .Z(n13081) );
  NAND U748 ( .A(n13532), .B(n13531), .Z(n355) );
  NAND U749 ( .A(n13530), .B(n13738), .Z(n356) );
  NAND U750 ( .A(n355), .B(n356), .Z(n13594) );
  NAND U751 ( .A(n13669), .B(n13668), .Z(n357) );
  NAND U752 ( .A(n13666), .B(n13667), .Z(n358) );
  AND U753 ( .A(n357), .B(n358), .Z(n13717) );
  NAND U754 ( .A(n13637), .B(n13636), .Z(n359) );
  NAND U755 ( .A(n13634), .B(n13635), .Z(n360) );
  AND U756 ( .A(n359), .B(n360), .Z(n13713) );
  XNOR U757 ( .A(n13999), .B(n13998), .Z(n13996) );
  NAND U758 ( .A(n13803), .B(n13802), .Z(n361) );
  NAND U759 ( .A(n13800), .B(n13801), .Z(n362) );
  NAND U760 ( .A(n361), .B(n362), .Z(n14158) );
  XNOR U761 ( .A(n15617), .B(n15616), .Z(n15614) );
  XNOR U762 ( .A(n15479), .B(n15480), .Z(n15477) );
  NAND U763 ( .A(n15221), .B(n15220), .Z(n363) );
  NAND U764 ( .A(n15218), .B(n15219), .Z(n364) );
  NAND U765 ( .A(n363), .B(n364), .Z(n15362) );
  XOR U766 ( .A(n15924), .B(n15923), .Z(n15876) );
  XNOR U767 ( .A(n15946), .B(n15945), .Z(n15959) );
  XNOR U768 ( .A(n16352), .B(n16351), .Z(n16349) );
  NAND U769 ( .A(n16008), .B(n16057), .Z(n365) );
  NANDN U770 ( .A(n15908), .B(n15907), .Z(n366) );
  AND U771 ( .A(n365), .B(n366), .Z(n16034) );
  XNOR U772 ( .A(n15995), .B(n15994), .Z(n16023) );
  XNOR U773 ( .A(n15982), .B(n15981), .Z(n15983) );
  XNOR U774 ( .A(n16271), .B(n16270), .Z(n16268) );
  NAND U775 ( .A(n16546), .B(n16545), .Z(n367) );
  NANDN U776 ( .A(n16548), .B(n16547), .Z(n368) );
  AND U777 ( .A(n367), .B(n368), .Z(n16607) );
  XNOR U778 ( .A(n17030), .B(n17029), .Z(n17027) );
  XOR U779 ( .A(n17343), .B(n17342), .Z(n17296) );
  XNOR U780 ( .A(n17353), .B(n17352), .Z(n17379) );
  XOR U781 ( .A(n17776), .B(n17777), .Z(n17778) );
  NAND U782 ( .A(n17428), .B(n17502), .Z(n369) );
  NANDN U783 ( .A(n17329), .B(n17328), .Z(n370) );
  AND U784 ( .A(n369), .B(n370), .Z(n17449) );
  XNOR U785 ( .A(n17409), .B(n17408), .Z(n17456) );
  XNOR U786 ( .A(n17395), .B(n17394), .Z(n17396) );
  XNOR U787 ( .A(n17691), .B(n17690), .Z(n17688) );
  NAND U788 ( .A(n17947), .B(n17946), .Z(n371) );
  NANDN U789 ( .A(n17945), .B(n17944), .Z(n372) );
  AND U790 ( .A(n371), .B(n372), .Z(n18021) );
  XNOR U791 ( .A(n18239), .B(n18238), .Z(n18241) );
  XNOR U792 ( .A(n18510), .B(n18509), .Z(n18507) );
  XNOR U793 ( .A(n18130), .B(n18129), .Z(n18131) );
  NAND U794 ( .A(n18916), .B(n18999), .Z(n373) );
  NANDN U795 ( .A(n18824), .B(n18823), .Z(n374) );
  AND U796 ( .A(n373), .B(n374), .Z(n18946) );
  NAND U797 ( .A(n1310), .B(n1311), .Z(n375) );
  XOR U798 ( .A(n1310), .B(n1311), .Z(n376) );
  NANDN U799 ( .A(n1309), .B(n376), .Z(n377) );
  NAND U800 ( .A(n375), .B(n377), .Z(n1417) );
  NAND U801 ( .A(n1483), .B(n1482), .Z(n378) );
  NAND U802 ( .A(n1480), .B(n1481), .Z(n379) );
  NAND U803 ( .A(n378), .B(n379), .Z(n1544) );
  NAND U804 ( .A(n1505), .B(n1504), .Z(n380) );
  NANDN U805 ( .A(n1503), .B(n1596), .Z(n381) );
  NAND U806 ( .A(n380), .B(n381), .Z(n1537) );
  XNOR U807 ( .A(n2573), .B(n2572), .Z(n2571) );
  XNOR U808 ( .A(n2537), .B(n2536), .Z(n2535) );
  XNOR U809 ( .A(n2305), .B(n2304), .Z(n2303) );
  NAND U810 ( .A(n2964), .B(n2963), .Z(n382) );
  NAND U811 ( .A(n2962), .B(n2961), .Z(n383) );
  AND U812 ( .A(n382), .B(n383), .Z(n3050) );
  XNOR U813 ( .A(n3180), .B(n3179), .Z(n3178) );
  XOR U814 ( .A(n3297), .B(n3296), .Z(n3293) );
  NAND U815 ( .A(n2786), .B(n2787), .Z(n384) );
  XOR U816 ( .A(n2786), .B(n2787), .Z(n385) );
  NANDN U817 ( .A(n2785), .B(n385), .Z(n386) );
  NAND U818 ( .A(n384), .B(n386), .Z(n2897) );
  XNOR U819 ( .A(n3629), .B(n3628), .Z(n3631) );
  XNOR U820 ( .A(n3756), .B(n3755), .Z(n3626) );
  XNOR U821 ( .A(n4034), .B(n4035), .Z(n4028) );
  XNOR U822 ( .A(n3793), .B(n3792), .Z(n3790) );
  NAND U823 ( .A(n4246), .B(n4245), .Z(n387) );
  NAND U824 ( .A(n4244), .B(n4243), .Z(n388) );
  AND U825 ( .A(n387), .B(n388), .Z(n4475) );
  XNOR U826 ( .A(n4464), .B(n4463), .Z(n4465) );
  NAND U827 ( .A(n4412), .B(n4411), .Z(n389) );
  NANDN U828 ( .A(n4414), .B(n4413), .Z(n390) );
  AND U829 ( .A(n389), .B(n390), .Z(n4742) );
  XNOR U830 ( .A(n4518), .B(n4517), .Z(n4515) );
  NAND U831 ( .A(n4397), .B(n4445), .Z(n391) );
  NANDN U832 ( .A(n4291), .B(n4290), .Z(n392) );
  AND U833 ( .A(n391), .B(n392), .Z(n4362) );
  NAND U834 ( .A(n4674), .B(n4309), .Z(n393) );
  NAND U835 ( .A(n4310), .B(n4376), .Z(n394) );
  NAND U836 ( .A(n393), .B(n394), .Z(n4359) );
  XNOR U837 ( .A(n4765), .B(n4764), .Z(n4763) );
  NAND U838 ( .A(n4962), .B(n4961), .Z(n395) );
  NAND U839 ( .A(n4960), .B(n4959), .Z(n396) );
  AND U840 ( .A(n395), .B(n396), .Z(n5208) );
  NAND U841 ( .A(n4982), .B(n4981), .Z(n397) );
  NAND U842 ( .A(n4983), .B(n4984), .Z(n398) );
  NAND U843 ( .A(n397), .B(n398), .Z(n5131) );
  XNOR U844 ( .A(n5087), .B(n5086), .Z(n5089) );
  XOR U845 ( .A(n5466), .B(n5467), .Z(n5460) );
  NAND U846 ( .A(n5139), .B(n5138), .Z(n399) );
  NANDN U847 ( .A(n5141), .B(n5140), .Z(n400) );
  AND U848 ( .A(n399), .B(n400), .Z(n5225) );
  XNOR U849 ( .A(n5239), .B(n5238), .Z(n5237) );
  NAND U850 ( .A(n5778), .B(n5777), .Z(n401) );
  NANDN U851 ( .A(n5776), .B(n5775), .Z(n402) );
  AND U852 ( .A(n401), .B(n402), .Z(n5924) );
  XNOR U853 ( .A(n6210), .B(n6211), .Z(n6205) );
  NAND U854 ( .A(n6333), .B(n6332), .Z(n403) );
  NAND U855 ( .A(n6331), .B(n6330), .Z(n404) );
  AND U856 ( .A(n403), .B(n404), .Z(n6417) );
  XNOR U857 ( .A(n6541), .B(n6540), .Z(n6530) );
  XNOR U858 ( .A(n6547), .B(n6546), .Z(n6593) );
  XNOR U859 ( .A(n6692), .B(n6691), .Z(n6689) );
  NAND U860 ( .A(n7167), .B(n7168), .Z(n405) );
  XOR U861 ( .A(n7167), .B(n7168), .Z(n406) );
  NANDN U862 ( .A(n7166), .B(n406), .Z(n407) );
  NAND U863 ( .A(n405), .B(n407), .Z(n7380) );
  NAND U864 ( .A(n7374), .B(n7373), .Z(n408) );
  NAND U865 ( .A(n7371), .B(n7372), .Z(n409) );
  AND U866 ( .A(n408), .B(n409), .Z(n7626) );
  NAND U867 ( .A(n7306), .B(n7538), .Z(n410) );
  NAND U868 ( .A(n7305), .B(n7304), .Z(n411) );
  AND U869 ( .A(n410), .B(n411), .Z(n7608) );
  NAND U870 ( .A(n7874), .B(n7873), .Z(n412) );
  NAND U871 ( .A(n7872), .B(n7871), .Z(n413) );
  AND U872 ( .A(n412), .B(n413), .Z(n8121) );
  NAND U873 ( .A(n7967), .B(n7966), .Z(n414) );
  NANDN U874 ( .A(n7965), .B(n7964), .Z(n415) );
  AND U875 ( .A(n414), .B(n415), .Z(n8113) );
  XNOR U876 ( .A(n8147), .B(n8146), .Z(n8144) );
  XNOR U877 ( .A(n8399), .B(n8398), .Z(n8397) );
  NAND U878 ( .A(n8923), .B(n8922), .Z(n416) );
  NAND U879 ( .A(n8924), .B(n8925), .Z(n417) );
  AND U880 ( .A(n416), .B(n417), .Z(n418) );
  NAND U881 ( .A(n8927), .B(n8926), .Z(n419) );
  NAND U882 ( .A(n8928), .B(n8929), .Z(n420) );
  NAND U883 ( .A(n419), .B(n420), .Z(n421) );
  XNOR U884 ( .A(n418), .B(n421), .Z(n8930) );
  XNOR U885 ( .A(n8874), .B(n8873), .Z(n8872) );
  NAND U886 ( .A(n9241), .B(n9240), .Z(n422) );
  NAND U887 ( .A(n9239), .B(n9238), .Z(n423) );
  AND U888 ( .A(n422), .B(n423), .Z(n9326) );
  XNOR U889 ( .A(n9442), .B(n9441), .Z(n9443) );
  NAND U890 ( .A(n9501), .B(n9500), .Z(n424) );
  NAND U891 ( .A(n9498), .B(n9499), .Z(n425) );
  AND U892 ( .A(n424), .B(n425), .Z(n9580) );
  NAND U893 ( .A(n9347), .B(n9346), .Z(n426) );
  NAND U894 ( .A(n9344), .B(n9345), .Z(n427) );
  NAND U895 ( .A(n426), .B(n427), .Z(n9466) );
  NAND U896 ( .A(n9961), .B(n9960), .Z(n428) );
  NAND U897 ( .A(n9959), .B(n9958), .Z(n429) );
  AND U898 ( .A(n428), .B(n429), .Z(n10046) );
  XNOR U899 ( .A(n10160), .B(n10159), .Z(n10161) );
  NAND U900 ( .A(n10220), .B(n10219), .Z(n430) );
  NAND U901 ( .A(n10217), .B(n10218), .Z(n431) );
  AND U902 ( .A(n430), .B(n431), .Z(n10299) );
  NAND U903 ( .A(n10078), .B(n10077), .Z(n432) );
  NAND U904 ( .A(n10075), .B(n10076), .Z(n433) );
  NAND U905 ( .A(n432), .B(n433), .Z(n10184) );
  NAND U906 ( .A(n10847), .B(n10846), .Z(n434) );
  NAND U907 ( .A(n10844), .B(n10845), .Z(n435) );
  NAND U908 ( .A(n434), .B(n435), .Z(n10992) );
  NAND U909 ( .A(n10942), .B(n10941), .Z(n436) );
  NAND U910 ( .A(n10940), .B(n10939), .Z(n437) );
  AND U911 ( .A(n436), .B(n437), .Z(n11267) );
  NAND U912 ( .A(n10932), .B(n10931), .Z(n438) );
  NAND U913 ( .A(n10929), .B(n10930), .Z(n439) );
  AND U914 ( .A(n438), .B(n439), .Z(n11015) );
  NAND U915 ( .A(n11652), .B(n11651), .Z(n440) );
  NANDN U916 ( .A(n11654), .B(n11653), .Z(n441) );
  AND U917 ( .A(n440), .B(n441), .Z(n11759) );
  XOR U918 ( .A(n11747), .B(n11746), .Z(n11745) );
  XNOR U919 ( .A(n11602), .B(n11601), .Z(n11604) );
  XNOR U920 ( .A(n12375), .B(n12374), .Z(n12399) );
  NAND U921 ( .A(n12324), .B(n12323), .Z(n442) );
  NANDN U922 ( .A(n12322), .B(n12321), .Z(n443) );
  AND U923 ( .A(n442), .B(n443), .Z(n12459) );
  XNOR U924 ( .A(n12514), .B(n12513), .Z(n12748) );
  XNOR U925 ( .A(n12505), .B(n12506), .Z(n12508) );
  XNOR U926 ( .A(n12496), .B(n12495), .Z(n12493) );
  NAND U927 ( .A(n12235), .B(n12234), .Z(n444) );
  NANDN U928 ( .A(n12233), .B(n12232), .Z(n445) );
  AND U929 ( .A(n444), .B(n445), .Z(n12469) );
  NAND U930 ( .A(n12962), .B(n12961), .Z(n446) );
  NAND U931 ( .A(n12960), .B(n12959), .Z(n447) );
  AND U932 ( .A(n446), .B(n447), .Z(n13215) );
  XNOR U933 ( .A(n13127), .B(n13126), .Z(n13129) );
  XOR U934 ( .A(n13159), .B(n13158), .Z(n13211) );
  XNOR U935 ( .A(n13374), .B(n13373), .Z(n13372) );
  XNOR U936 ( .A(n13493), .B(n13494), .Z(n13488) );
  NAND U937 ( .A(n14114), .B(n14113), .Z(n448) );
  NAND U938 ( .A(n14115), .B(n14116), .Z(n449) );
  AND U939 ( .A(n448), .B(n449), .Z(n450) );
  NAND U940 ( .A(n14120), .B(n14119), .Z(n451) );
  NAND U941 ( .A(n14117), .B(n14118), .Z(n452) );
  NAND U942 ( .A(n451), .B(n452), .Z(n453) );
  XNOR U943 ( .A(n450), .B(n453), .Z(n14121) );
  NAND U944 ( .A(n13904), .B(n13903), .Z(n454) );
  NANDN U945 ( .A(n13906), .B(n13905), .Z(n455) );
  NAND U946 ( .A(n454), .B(n455), .Z(n14191) );
  NAND U947 ( .A(n14626), .B(n14570), .Z(n456) );
  NANDN U948 ( .A(n14457), .B(n14456), .Z(n457) );
  AND U949 ( .A(n456), .B(n457), .Z(n14524) );
  NAND U950 ( .A(n14407), .B(n14408), .Z(n458) );
  XOR U951 ( .A(n14407), .B(n14408), .Z(n459) );
  NANDN U952 ( .A(n14406), .B(n459), .Z(n460) );
  NAND U953 ( .A(n458), .B(n460), .Z(n14658) );
  XNOR U954 ( .A(n14926), .B(n14925), .Z(n14924) );
  XOR U955 ( .A(n15037), .B(n15036), .Z(n14979) );
  XNOR U956 ( .A(n15113), .B(n15112), .Z(n15115) );
  NAND U957 ( .A(n15297), .B(n15296), .Z(n461) );
  NANDN U958 ( .A(n15299), .B(n15298), .Z(n462) );
  AND U959 ( .A(n461), .B(n462), .Z(n15394) );
  XNOR U960 ( .A(n15381), .B(n15380), .Z(n15378) );
  XOR U961 ( .A(n15125), .B(n15126), .Z(n463) );
  NANDN U962 ( .A(n15127), .B(n463), .Z(n464) );
  NAND U963 ( .A(n15125), .B(n15126), .Z(n465) );
  AND U964 ( .A(n464), .B(n465), .Z(n15366) );
  NAND U965 ( .A(n15857), .B(n15856), .Z(n466) );
  NAND U966 ( .A(n15855), .B(n15854), .Z(n467) );
  AND U967 ( .A(n466), .B(n467), .Z(n16105) );
  NAND U968 ( .A(n15952), .B(n15951), .Z(n468) );
  NANDN U969 ( .A(n15950), .B(n15949), .Z(n469) );
  AND U970 ( .A(n468), .B(n469), .Z(n16097) );
  XNOR U971 ( .A(n16383), .B(n16384), .Z(n16378) );
  XNOR U972 ( .A(n16815), .B(n16814), .Z(n16816) );
  XNOR U973 ( .A(n17063), .B(n17064), .Z(n17066) );
  NAND U974 ( .A(n16762), .B(n16761), .Z(n470) );
  NANDN U975 ( .A(n16764), .B(n16763), .Z(n471) );
  AND U976 ( .A(n470), .B(n471), .Z(n17057) );
  NAND U977 ( .A(n16866), .B(n16865), .Z(n472) );
  NAND U978 ( .A(n16967), .B(n16867), .Z(n473) );
  AND U979 ( .A(n472), .B(n473), .Z(n474) );
  NAND U980 ( .A(n16869), .B(n16868), .Z(n475) );
  NAND U981 ( .A(n16870), .B(n16871), .Z(n476) );
  NAND U982 ( .A(n475), .B(n476), .Z(n477) );
  XNOR U983 ( .A(n474), .B(n477), .Z(n16872) );
  NAND U984 ( .A(n16782), .B(n16748), .Z(n478) );
  NANDN U985 ( .A(n16638), .B(n16637), .Z(n479) );
  AND U986 ( .A(n478), .B(n479), .Z(n16713) );
  XNOR U987 ( .A(n17080), .B(n17079), .Z(n17078) );
  NAND U988 ( .A(n17277), .B(n17276), .Z(n480) );
  NAND U989 ( .A(n17275), .B(n17274), .Z(n481) );
  AND U990 ( .A(n480), .B(n481), .Z(n17526) );
  NAND U991 ( .A(n17371), .B(n17370), .Z(n482) );
  NANDN U992 ( .A(n17369), .B(n17368), .Z(n483) );
  AND U993 ( .A(n482), .B(n483), .Z(n17518) );
  XNOR U994 ( .A(n17804), .B(n17805), .Z(n17799) );
  NAND U995 ( .A(n17925), .B(n17924), .Z(n484) );
  NAND U996 ( .A(n17923), .B(n17922), .Z(n485) );
  AND U997 ( .A(n484), .B(n485), .Z(n18011) );
  XNOR U998 ( .A(n18138), .B(n18137), .Z(n18127) );
  XNOR U999 ( .A(n18205), .B(n18204), .Z(n18143) );
  XNOR U1000 ( .A(n18536), .B(n18535), .Z(n18533) );
  XNOR U1001 ( .A(n18289), .B(n18288), .Z(n18286) );
  XNOR U1002 ( .A(n18168), .B(n18167), .Z(n18146) );
  XNOR U1003 ( .A(n18887), .B(n18886), .Z(n18889) );
  XOR U1004 ( .A(n19019), .B(n19018), .Z(n19021) );
  XOR U1005 ( .A(n19172), .B(n19171), .Z(n19044) );
  XNOR U1006 ( .A(n18918), .B(n18917), .Z(n18971) );
  XOR U1007 ( .A(n19052), .B(n19051), .Z(n19050) );
  NAND U1008 ( .A(n1425), .B(n1424), .Z(n486) );
  NAND U1009 ( .A(n1422), .B(n1423), .Z(n487) );
  AND U1010 ( .A(n486), .B(n487), .Z(n1825) );
  NAND U1011 ( .A(n2146), .B(n2145), .Z(n488) );
  NANDN U1012 ( .A(n2144), .B(n2143), .Z(n489) );
  AND U1013 ( .A(n488), .B(n489), .Z(n2293) );
  NAND U1014 ( .A(n3305), .B(n3306), .Z(n3310) );
  XNOR U1015 ( .A(n4053), .B(n4052), .Z(n3773) );
  XNOR U1016 ( .A(n4759), .B(n4758), .Z(n4757) );
  NAND U1017 ( .A(n4356), .B(n4355), .Z(n490) );
  NAND U1018 ( .A(n4354), .B(n4353), .Z(n491) );
  AND U1019 ( .A(n490), .B(n491), .Z(n4486) );
  XNOR U1020 ( .A(n5475), .B(n5474), .Z(n5473) );
  XOR U1021 ( .A(n5353), .B(n5352), .Z(n5219) );
  NAND U1022 ( .A(n5928), .B(n5927), .Z(n492) );
  NAND U1023 ( .A(n5929), .B(n5930), .Z(n493) );
  NAND U1024 ( .A(n492), .B(n493), .Z(n5938) );
  NAND U1025 ( .A(n6571), .B(n6570), .Z(n494) );
  NAND U1026 ( .A(n6568), .B(n6569), .Z(n495) );
  NAND U1027 ( .A(n494), .B(n495), .Z(n6679) );
  NAND U1028 ( .A(n7378), .B(n7377), .Z(n496) );
  NANDN U1029 ( .A(n7376), .B(n7375), .Z(n497) );
  AND U1030 ( .A(n496), .B(n497), .Z(n7661) );
  NAND U1031 ( .A(n7334), .B(n7333), .Z(n498) );
  NAND U1032 ( .A(n7332), .B(n7331), .Z(n499) );
  AND U1033 ( .A(n498), .B(n499), .Z(n7675) );
  NAND U1034 ( .A(n8117), .B(n8116), .Z(n500) );
  NAND U1035 ( .A(n8118), .B(n8119), .Z(n501) );
  NAND U1036 ( .A(n500), .B(n501), .Z(n8127) );
  XNOR U1037 ( .A(n9126), .B(n9125), .Z(n9124) );
  NAND U1038 ( .A(n8747), .B(n8746), .Z(n502) );
  NAND U1039 ( .A(n8744), .B(n8745), .Z(n503) );
  NAND U1040 ( .A(n502), .B(n503), .Z(n8869) );
  NAND U1041 ( .A(n9585), .B(n9584), .Z(n504) );
  NAND U1042 ( .A(n9586), .B(n9587), .Z(n505) );
  AND U1043 ( .A(n504), .B(n505), .Z(n506) );
  NAND U1044 ( .A(n9591), .B(n9590), .Z(n507) );
  NANDN U1045 ( .A(n9588), .B(n9589), .Z(n508) );
  AND U1046 ( .A(n507), .B(n508), .Z(n509) );
  NAND U1047 ( .A(n9593), .B(n9592), .Z(n510) );
  NAND U1048 ( .A(n9594), .B(n9595), .Z(n511) );
  AND U1049 ( .A(n510), .B(n511), .Z(n512) );
  AND U1050 ( .A(n9712), .B(n9711), .Z(n513) );
  XNOR U1051 ( .A(n9810), .B(n9809), .Z(n514) );
  XNOR U1052 ( .A(n513), .B(n514), .Z(n515) );
  AND U1053 ( .A(n9601), .B(n9600), .Z(n516) );
  XNOR U1054 ( .A(n9706), .B(n9705), .Z(n517) );
  XNOR U1055 ( .A(n516), .B(n517), .Z(n518) );
  XOR U1056 ( .A(n515), .B(n518), .Z(n519) );
  XNOR U1057 ( .A(n509), .B(n512), .Z(n520) );
  XNOR U1058 ( .A(n519), .B(n520), .Z(n521) );
  XNOR U1059 ( .A(n506), .B(n521), .Z(n9811) );
  NAND U1060 ( .A(n10304), .B(n10303), .Z(n522) );
  NANDN U1061 ( .A(n10306), .B(n10305), .Z(n523) );
  AND U1062 ( .A(n522), .B(n523), .Z(n524) );
  NAND U1063 ( .A(n10310), .B(n10309), .Z(n525) );
  NAND U1064 ( .A(n10308), .B(n10307), .Z(n526) );
  AND U1065 ( .A(n525), .B(n526), .Z(n527) );
  NAND U1066 ( .A(n10312), .B(n10311), .Z(n528) );
  NAND U1067 ( .A(n10313), .B(n10314), .Z(n529) );
  AND U1068 ( .A(n528), .B(n529), .Z(n530) );
  AND U1069 ( .A(n10431), .B(n10430), .Z(n531) );
  XNOR U1070 ( .A(n10425), .B(n10424), .Z(n532) );
  XNOR U1071 ( .A(n531), .B(n532), .Z(n533) );
  AND U1072 ( .A(n10320), .B(n10319), .Z(n534) );
  XNOR U1073 ( .A(n10530), .B(n533), .Z(n535) );
  XNOR U1074 ( .A(n534), .B(n535), .Z(n536) );
  XOR U1075 ( .A(n530), .B(n536), .Z(n537) );
  XNOR U1076 ( .A(n524), .B(n527), .Z(n538) );
  XNOR U1077 ( .A(n537), .B(n538), .Z(n10531) );
  NOR U1078 ( .A(n11003), .B(n11004), .Z(n11006) );
  XNOR U1079 ( .A(n11743), .B(n11742), .Z(n11741) );
  NAND U1080 ( .A(n12465), .B(n12464), .Z(n539) );
  NAND U1081 ( .A(n12466), .B(n12467), .Z(n540) );
  NAND U1082 ( .A(n539), .B(n540), .Z(n12483) );
  XNOR U1083 ( .A(n13502), .B(n13503), .Z(n13501) );
  XOR U1084 ( .A(n13253), .B(n13252), .Z(n13229) );
  XNOR U1085 ( .A(n13916), .B(n13915), .Z(n13909) );
  NAND U1086 ( .A(n13810), .B(n13809), .Z(n541) );
  NAND U1087 ( .A(n13807), .B(n13808), .Z(n542) );
  NAND U1088 ( .A(n541), .B(n542), .Z(n13927) );
  NAND U1089 ( .A(n14677), .B(n14676), .Z(n543) );
  NAND U1090 ( .A(n14678), .B(n14679), .Z(n544) );
  AND U1091 ( .A(n543), .B(n544), .Z(n545) );
  NAND U1092 ( .A(n14683), .B(n14682), .Z(n546) );
  NANDN U1093 ( .A(n14680), .B(n14681), .Z(n547) );
  AND U1094 ( .A(n546), .B(n547), .Z(n548) );
  NAND U1095 ( .A(n14684), .B(n14685), .Z(n549) );
  NAND U1096 ( .A(n14686), .B(n14687), .Z(n550) );
  AND U1097 ( .A(n549), .B(n550), .Z(n551) );
  XOR U1098 ( .A(n14906), .B(n14905), .Z(n552) );
  XNOR U1099 ( .A(n14800), .B(n14799), .Z(n553) );
  XNOR U1100 ( .A(n552), .B(n553), .Z(n554) );
  XOR U1101 ( .A(n551), .B(n554), .Z(n555) );
  XNOR U1102 ( .A(n545), .B(n548), .Z(n556) );
  XNOR U1103 ( .A(n555), .B(n556), .Z(n557) );
  NAND U1104 ( .A(n14673), .B(n14672), .Z(n558) );
  NAND U1105 ( .A(n14674), .B(n14675), .Z(n559) );
  NAND U1106 ( .A(n558), .B(n559), .Z(n560) );
  XNOR U1107 ( .A(n557), .B(n560), .Z(n14922) );
  NAND U1108 ( .A(n15237), .B(n15236), .Z(n561) );
  NANDN U1109 ( .A(n15239), .B(n15238), .Z(n562) );
  NAND U1110 ( .A(n561), .B(n562), .Z(n15655) );
  NAND U1111 ( .A(n16101), .B(n16100), .Z(n563) );
  NAND U1112 ( .A(n16102), .B(n16103), .Z(n564) );
  NAND U1113 ( .A(n563), .B(n564), .Z(n16111) );
  XNOR U1114 ( .A(n17074), .B(n17073), .Z(n17072) );
  NAND U1115 ( .A(n16707), .B(n16706), .Z(n565) );
  NAND U1116 ( .A(n16705), .B(n16704), .Z(n566) );
  AND U1117 ( .A(n565), .B(n566), .Z(n16837) );
  NAND U1118 ( .A(n17522), .B(n17521), .Z(n567) );
  NAND U1119 ( .A(n17523), .B(n17524), .Z(n568) );
  NAND U1120 ( .A(n567), .B(n568), .Z(n17532) );
  NAND U1121 ( .A(n18150), .B(n18149), .Z(n569) );
  NANDN U1122 ( .A(n18152), .B(n18151), .Z(n570) );
  AND U1123 ( .A(n569), .B(n570), .Z(n18277) );
  XNOR U1124 ( .A(n19033), .B(n19034), .Z(n19032) );
  XNOR U1125 ( .A(n6396), .B(n6395), .Z(n6382) );
  XNOR U1126 ( .A(n17990), .B(n17989), .Z(n17975) );
  XNOR U1127 ( .A(n1178), .B(n1177), .Z(n1211) );
  NAND U1128 ( .A(n1208), .B(n1209), .Z(n571) );
  NAND U1129 ( .A(n1347), .B(n1350), .Z(n572) );
  NAND U1130 ( .A(n571), .B(n572), .Z(n1216) );
  XNOR U1131 ( .A(n1901), .B(n1900), .Z(n1928) );
  NAND U1132 ( .A(n1925), .B(n1926), .Z(n573) );
  NAND U1133 ( .A(n2059), .B(n2080), .Z(n574) );
  NAND U1134 ( .A(n573), .B(n574), .Z(n1963) );
  XNOR U1135 ( .A(n2660), .B(n2659), .Z(n2693) );
  NAND U1136 ( .A(n2690), .B(n2691), .Z(n575) );
  NAND U1137 ( .A(n2832), .B(n2829), .Z(n576) );
  NAND U1138 ( .A(n575), .B(n576), .Z(n2698) );
  NAND U1139 ( .A(n2727), .B(n2726), .Z(n577) );
  NAND U1140 ( .A(n2724), .B(n2725), .Z(n578) );
  AND U1141 ( .A(n577), .B(n578), .Z(n2890) );
  AND U1142 ( .A(n2742), .B(n2741), .Z(n579) );
  AND U1143 ( .A(n2740), .B(y[97]), .Z(n580) );
  NAND U1144 ( .A(x[19]), .B(n580), .Z(n581) );
  NANDN U1145 ( .A(n579), .B(n581), .Z(n2882) );
  XNOR U1146 ( .A(n3382), .B(n3381), .Z(n3414) );
  XNOR U1147 ( .A(n3473), .B(n3472), .Z(n3446) );
  XNOR U1148 ( .A(n3641), .B(n3640), .Z(n3642) );
  XNOR U1149 ( .A(n3635), .B(n3634), .Z(n3636) );
  XOR U1150 ( .A(n3571), .B(n3570), .Z(n3556) );
  XNOR U1151 ( .A(n5059), .B(n5058), .Z(n5061) );
  XNOR U1152 ( .A(n5065), .B(n5064), .Z(n5066) );
  XNOR U1153 ( .A(n5549), .B(n5548), .Z(n5576) );
  NAND U1154 ( .A(n5573), .B(n5574), .Z(n582) );
  NAND U1155 ( .A(n5713), .B(n5729), .Z(n583) );
  NAND U1156 ( .A(n582), .B(n583), .Z(n5611) );
  XNOR U1157 ( .A(n5708), .B(n5707), .Z(n5709) );
  XNOR U1158 ( .A(n5808), .B(n5807), .Z(n5810) );
  XNOR U1159 ( .A(n5770), .B(n5769), .Z(n5771) );
  XNOR U1160 ( .A(n6379), .B(n6378), .Z(n6354) );
  XNOR U1161 ( .A(n6517), .B(n6516), .Z(n6518) );
  XNOR U1162 ( .A(n7041), .B(n7040), .Z(n7074) );
  NAND U1163 ( .A(n7108), .B(n7107), .Z(n584) );
  NAND U1164 ( .A(n7105), .B(n7106), .Z(n585) );
  AND U1165 ( .A(n584), .B(n585), .Z(n7259) );
  XNOR U1166 ( .A(n7911), .B(n7910), .Z(n7912) );
  XNOR U1167 ( .A(n8045), .B(n8044), .Z(n8047) );
  XNOR U1168 ( .A(n7947), .B(n7946), .Z(n7948) );
  XNOR U1169 ( .A(n8478), .B(n8477), .Z(n8505) );
  XNOR U1170 ( .A(n8570), .B(n8569), .Z(n8543) );
  XNOR U1171 ( .A(n8711), .B(n8710), .Z(n8712) );
  XNOR U1172 ( .A(n8717), .B(n8716), .Z(n8718) );
  XNOR U1173 ( .A(n9288), .B(n9287), .Z(n9262) );
  XNOR U1174 ( .A(n9380), .B(n9379), .Z(n9381) );
  XNOR U1175 ( .A(n10008), .B(n10007), .Z(n9982) );
  XNOR U1176 ( .A(n10025), .B(n10024), .Z(n10011) );
  XNOR U1177 ( .A(n10099), .B(n10098), .Z(n10100) );
  NAND U1178 ( .A(n10723), .B(n10722), .Z(n586) );
  NAND U1179 ( .A(n10720), .B(n10721), .Z(n587) );
  AND U1180 ( .A(n586), .B(n587), .Z(n10835) );
  NAND U1181 ( .A(n10688), .B(n10687), .Z(n588) );
  NAND U1182 ( .A(n10685), .B(n10686), .Z(n589) );
  NAND U1183 ( .A(n588), .B(n589), .Z(n10840) );
  XNOR U1184 ( .A(n11351), .B(n11350), .Z(n11379) );
  XNOR U1185 ( .A(n12091), .B(n12090), .Z(n12124) );
  XNOR U1186 ( .A(n12617), .B(n12616), .Z(n12614) );
  XOR U1187 ( .A(n12445), .B(n12388), .Z(n12274) );
  XNOR U1188 ( .A(n12451), .B(n12450), .Z(n12452) );
  XNOR U1189 ( .A(n12279), .B(n12278), .Z(n12280) );
  XNOR U1190 ( .A(n12262), .B(n12261), .Z(n12306) );
  NAND U1191 ( .A(n12122), .B(n12123), .Z(n590) );
  NAND U1192 ( .A(n12265), .B(n12268), .Z(n591) );
  NAND U1193 ( .A(n590), .B(n591), .Z(n12130) );
  XNOR U1194 ( .A(n13102), .B(n13101), .Z(n13104) );
  XNOR U1195 ( .A(n13049), .B(n13048), .Z(n13050) );
  XNOR U1196 ( .A(n14276), .B(n14275), .Z(n14309) );
  NAND U1197 ( .A(n14306), .B(n14307), .Z(n592) );
  NAND U1198 ( .A(n14438), .B(n14451), .Z(n593) );
  NAND U1199 ( .A(n592), .B(n593), .Z(n14314) );
  XNOR U1200 ( .A(n15019), .B(n15018), .Z(n15021) );
  AND U1201 ( .A(n15084), .B(n15083), .Z(n594) );
  AND U1202 ( .A(n15082), .B(x[139]), .Z(n595) );
  NAND U1203 ( .A(y[113]), .B(n595), .Z(n596) );
  NANDN U1204 ( .A(n594), .B(n596), .Z(n15222) );
  XNOR U1205 ( .A(n15894), .B(n15893), .Z(n15895) );
  XNOR U1206 ( .A(n15988), .B(n15987), .Z(n15990) );
  XNOR U1207 ( .A(n15944), .B(n15943), .Z(n15945) );
  XNOR U1208 ( .A(n16463), .B(n16462), .Z(n16490) );
  NAND U1209 ( .A(n16487), .B(n16488), .Z(n597) );
  NAND U1210 ( .A(n16628), .B(n16632), .Z(n598) );
  NAND U1211 ( .A(n597), .B(n598), .Z(n16525) );
  XNOR U1212 ( .A(n17314), .B(n17313), .Z(n17315) );
  XNOR U1213 ( .A(n17351), .B(n17350), .Z(n17352) );
  XNOR U1214 ( .A(n17959), .B(n17958), .Z(n17946) );
  XNOR U1215 ( .A(n18114), .B(n18113), .Z(n18115) );
  XNOR U1216 ( .A(n18120), .B(n18119), .Z(n18122) );
  XNOR U1217 ( .A(n18638), .B(n18637), .Z(n18666) );
  NAND U1218 ( .A(n18663), .B(n18664), .Z(n599) );
  NAND U1219 ( .A(n18815), .B(n18818), .Z(n600) );
  NAND U1220 ( .A(n599), .B(n600), .Z(n18701) );
  XNOR U1221 ( .A(n18899), .B(n18843), .Z(n18846) );
  XOR U1222 ( .A(n19281), .B(n19280), .Z(n19283) );
  NAND U1223 ( .A(n1680), .B(n1380), .Z(n601) );
  NAND U1224 ( .A(n1381), .B(n1446), .Z(n602) );
  NAND U1225 ( .A(n601), .B(n602), .Z(n1474) );
  NAND U1226 ( .A(n1441), .B(n1440), .Z(n603) );
  NAND U1227 ( .A(n1439), .B(n1438), .Z(n604) );
  AND U1228 ( .A(n603), .B(n604), .Z(n1755) );
  XNOR U1229 ( .A(n1375), .B(n1374), .Z(n1376) );
  NAND U1230 ( .A(n2255), .B(n2188), .Z(n605) );
  NANDN U1231 ( .A(n2086), .B(n2085), .Z(n606) );
  AND U1232 ( .A(n605), .B(n606), .Z(n2225) );
  XOR U1233 ( .A(n2354), .B(n2353), .Z(n2352) );
  XOR U1234 ( .A(n2421), .B(n2420), .Z(n2419) );
  XNOR U1235 ( .A(n2237), .B(n2236), .Z(n2238) );
  XOR U1236 ( .A(n2853), .B(n2852), .Z(n2807) );
  XOR U1237 ( .A(n2842), .B(n2841), .Z(n2801) );
  NAND U1238 ( .A(n2935), .B(n2998), .Z(n607) );
  NANDN U1239 ( .A(n2838), .B(n2837), .Z(n608) );
  AND U1240 ( .A(n607), .B(n608), .Z(n2972) );
  NAND U1241 ( .A(n2930), .B(n2929), .Z(n609) );
  AND U1242 ( .A(n2928), .B(x[11]), .Z(n610) );
  NAND U1243 ( .A(y[59]), .B(n610), .Z(n611) );
  AND U1244 ( .A(n609), .B(n611), .Z(n3270) );
  XOR U1245 ( .A(n3186), .B(n3185), .Z(n3184) );
  XNOR U1246 ( .A(n3139), .B(n3138), .Z(n3136) );
  XNOR U1247 ( .A(n3607), .B(n3606), .Z(n3609) );
  XNOR U1248 ( .A(n3669), .B(n3668), .Z(n3724) );
  XNOR U1249 ( .A(n3700), .B(n3699), .Z(n3701) );
  XNOR U1250 ( .A(n3688), .B(n3687), .Z(n3690) );
  XNOR U1251 ( .A(n3648), .B(n3647), .Z(n3694) );
  XNOR U1252 ( .A(n3965), .B(n3964), .Z(n3962) );
  XOR U1253 ( .A(n3903), .B(n3902), .Z(n3901) );
  NAND U1254 ( .A(n4185), .B(n4184), .Z(n612) );
  NANDN U1255 ( .A(n4183), .B(n4182), .Z(n613) );
  AND U1256 ( .A(n612), .B(n613), .Z(n4254) );
  XNOR U1257 ( .A(n4330), .B(n4329), .Z(n4332) );
  XNOR U1258 ( .A(n4336), .B(n4335), .Z(n4337) );
  XNOR U1259 ( .A(n4324), .B(n4323), .Z(n4326) );
  NAND U1260 ( .A(n4312), .B(n4311), .Z(n614) );
  NANDN U1261 ( .A(n4314), .B(n4313), .Z(n615) );
  AND U1262 ( .A(n614), .B(n615), .Z(n4413) );
  NAND U1263 ( .A(n4281), .B(n4280), .Z(n616) );
  NAND U1264 ( .A(n4278), .B(n4279), .Z(n617) );
  NAND U1265 ( .A(n616), .B(n617), .Z(n4441) );
  XNOR U1266 ( .A(n4725), .B(n4724), .Z(n4722) );
  NAND U1267 ( .A(n4399), .B(n4398), .Z(n618) );
  NANDN U1268 ( .A(n4397), .B(n4661), .Z(n619) );
  AND U1269 ( .A(n618), .B(n619), .Z(n4635) );
  NAND U1270 ( .A(n4374), .B(n4373), .Z(n620) );
  NAND U1271 ( .A(n4371), .B(n4372), .Z(n621) );
  NAND U1272 ( .A(n620), .B(n621), .Z(n4631) );
  XOR U1273 ( .A(n4589), .B(n4588), .Z(n4587) );
  NAND U1274 ( .A(n4277), .B(n4276), .Z(n622) );
  NAND U1275 ( .A(n4275), .B(n4274), .Z(n623) );
  AND U1276 ( .A(n622), .B(n623), .Z(n4384) );
  XNOR U1277 ( .A(n5053), .B(n5052), .Z(n5055) );
  NAND U1278 ( .A(n4897), .B(n4896), .Z(n624) );
  NANDN U1279 ( .A(n4895), .B(n4894), .Z(n625) );
  AND U1280 ( .A(n624), .B(n625), .Z(n4970) );
  XOR U1281 ( .A(n5027), .B(n5026), .Z(n4982) );
  XOR U1282 ( .A(n5243), .B(n5242), .Z(n5241) );
  XOR U1283 ( .A(n5375), .B(n5374), .Z(n5373) );
  NAND U1284 ( .A(n5113), .B(n5171), .Z(n626) );
  NANDN U1285 ( .A(n5011), .B(n5010), .Z(n627) );
  AND U1286 ( .A(n626), .B(n627), .Z(n5142) );
  XOR U1287 ( .A(n5739), .B(n5738), .Z(n5718) );
  XNOR U1288 ( .A(n5726), .B(n5725), .Z(n5781) );
  XNOR U1289 ( .A(n6178), .B(n6179), .Z(n6176) );
  XNOR U1290 ( .A(n6049), .B(n6048), .Z(n6046) );
  XNOR U1291 ( .A(n5856), .B(n5855), .Z(n5858) );
  XNOR U1292 ( .A(n5702), .B(n5701), .Z(n5703) );
  XNOR U1293 ( .A(n5874), .B(n5873), .Z(n5875) );
  XNOR U1294 ( .A(n5868), .B(n5867), .Z(n5869) );
  XOR U1295 ( .A(n6485), .B(n6484), .Z(n6439) );
  XOR U1296 ( .A(n6475), .B(n6474), .Z(n6433) );
  NAND U1297 ( .A(n6582), .B(n6623), .Z(n628) );
  NANDN U1298 ( .A(n6471), .B(n6470), .Z(n629) );
  AND U1299 ( .A(n628), .B(n629), .Z(n6599) );
  XNOR U1300 ( .A(n6831), .B(n6832), .Z(n6829) );
  XNOR U1301 ( .A(n6784), .B(n6783), .Z(n6781) );
  NAND U1302 ( .A(n7366), .B(n7365), .Z(n630) );
  NAND U1303 ( .A(n7364), .B(n7363), .Z(n631) );
  AND U1304 ( .A(n630), .B(n631), .Z(n7463) );
  NAND U1305 ( .A(n7253), .B(n7252), .Z(n632) );
  NAND U1306 ( .A(n7250), .B(n7251), .Z(n633) );
  NAND U1307 ( .A(n632), .B(n633), .Z(n7268) );
  NAND U1308 ( .A(n7809), .B(n7808), .Z(n634) );
  NANDN U1309 ( .A(n7807), .B(n7806), .Z(n635) );
  AND U1310 ( .A(n634), .B(n635), .Z(n7882) );
  XOR U1311 ( .A(n7929), .B(n7928), .Z(n7888) );
  XNOR U1312 ( .A(n7896), .B(n7895), .Z(n7970) );
  XNOR U1313 ( .A(n8357), .B(n8356), .Z(n8354) );
  XNOR U1314 ( .A(n7997), .B(n7996), .Z(n7999) );
  XNOR U1315 ( .A(n8218), .B(n8217), .Z(n8215) );
  XNOR U1316 ( .A(n7905), .B(n7904), .Z(n7906) );
  XNOR U1317 ( .A(n8063), .B(n8062), .Z(n8064) );
  XNOR U1318 ( .A(n8057), .B(n8056), .Z(n8058) );
  XNOR U1319 ( .A(n8705), .B(n8704), .Z(n8707) );
  XOR U1320 ( .A(n8679), .B(n8678), .Z(n8633) );
  NAND U1321 ( .A(n8775), .B(n8815), .Z(n636) );
  NANDN U1322 ( .A(n8664), .B(n8663), .Z(n637) );
  AND U1323 ( .A(n636), .B(n637), .Z(n8797) );
  XNOR U1324 ( .A(n9076), .B(n9075), .Z(n9073) );
  XNOR U1325 ( .A(n8937), .B(n8936), .Z(n8934) );
  XOR U1326 ( .A(n9394), .B(n9393), .Z(n9363) );
  XNOR U1327 ( .A(n9420), .B(n9419), .Z(n9421) );
  XNOR U1328 ( .A(n9426), .B(n9425), .Z(n9427) );
  NAND U1329 ( .A(n9351), .B(n9350), .Z(n638) );
  NAND U1330 ( .A(n9348), .B(n9349), .Z(n639) );
  NAND U1331 ( .A(n638), .B(n639), .Z(n9538) );
  XNOR U1332 ( .A(n9669), .B(n9670), .Z(n9667) );
  XOR U1333 ( .A(n9599), .B(n9598), .Z(n9597) );
  NAND U1334 ( .A(n9462), .B(n9463), .Z(n640) );
  NAND U1335 ( .A(n9525), .B(n9461), .Z(n641) );
  AND U1336 ( .A(n640), .B(n641), .Z(n9802) );
  XNOR U1337 ( .A(n9716), .B(n9715), .Z(n9713) );
  NAND U1338 ( .A(n9343), .B(n9342), .Z(n642) );
  NANDN U1339 ( .A(n9480), .B(n9341), .Z(n643) );
  NAND U1340 ( .A(n642), .B(n643), .Z(n9447) );
  XOR U1341 ( .A(n10112), .B(n10111), .Z(n10068) );
  XNOR U1342 ( .A(n10138), .B(n10137), .Z(n10139) );
  XNOR U1343 ( .A(n10144), .B(n10143), .Z(n10145) );
  NAND U1344 ( .A(n10082), .B(n10081), .Z(n644) );
  NAND U1345 ( .A(n10079), .B(n10080), .Z(n645) );
  NAND U1346 ( .A(n644), .B(n645), .Z(n10263) );
  XOR U1347 ( .A(n10389), .B(n10388), .Z(n10387) );
  XNOR U1348 ( .A(n10318), .B(n10317), .Z(n10315) );
  XNOR U1349 ( .A(n10517), .B(n10516), .Z(n10514) );
  AND U1350 ( .A(n10074), .B(n10073), .Z(n646) );
  ANDN U1351 ( .B(y[97]), .A(n10198), .Z(n647) );
  NAND U1352 ( .A(x[98]), .B(n647), .Z(n648) );
  NANDN U1353 ( .A(n646), .B(n648), .Z(n10165) );
  XNOR U1354 ( .A(n10752), .B(n10751), .Z(n10738) );
  NAND U1355 ( .A(n10708), .B(n10707), .Z(n649) );
  NANDN U1356 ( .A(n10706), .B(n10705), .Z(n650) );
  NAND U1357 ( .A(n649), .B(n650), .Z(n10844) );
  NAND U1358 ( .A(n10793), .B(n10792), .Z(n651) );
  NANDN U1359 ( .A(n10791), .B(n10790), .Z(n652) );
  NAND U1360 ( .A(n651), .B(n652), .Z(n10916) );
  NAND U1361 ( .A(n10890), .B(n10889), .Z(n653) );
  ANDN U1362 ( .B(y[67]), .A(n10888), .Z(n654) );
  NAND U1363 ( .A(x[91]), .B(n654), .Z(n655) );
  AND U1364 ( .A(n653), .B(n655), .Z(n11040) );
  XNOR U1365 ( .A(n11246), .B(n11247), .Z(n11248) );
  XNOR U1366 ( .A(n11863), .B(n11862), .Z(n11860) );
  XOR U1367 ( .A(n11779), .B(n11778), .Z(n11777) );
  NAND U1368 ( .A(n11639), .B(n11716), .Z(n656) );
  NANDN U1369 ( .A(n11537), .B(n11536), .Z(n657) );
  AND U1370 ( .A(n656), .B(n657), .Z(n11655) );
  XOR U1371 ( .A(n11950), .B(n11949), .Z(n11948) );
  XOR U1372 ( .A(n11552), .B(n11551), .Z(n11506) );
  XOR U1373 ( .A(n11541), .B(n11540), .Z(n11500) );
  XNOR U1374 ( .A(n12314), .B(n12313), .Z(n12328) );
  XNOR U1375 ( .A(n12245), .B(n12244), .Z(n12323) );
  XNOR U1376 ( .A(n12566), .B(n12380), .Z(n12373) );
  XNOR U1377 ( .A(n12702), .B(n12701), .Z(n12699) );
  XOR U1378 ( .A(n12722), .B(n12721), .Z(n12720) );
  XNOR U1379 ( .A(n12442), .B(n12441), .Z(n12338) );
  NAND U1380 ( .A(n12897), .B(n12896), .Z(n658) );
  NANDN U1381 ( .A(n12895), .B(n12894), .Z(n659) );
  AND U1382 ( .A(n658), .B(n659), .Z(n12970) );
  XOR U1383 ( .A(n13018), .B(n13017), .Z(n12976) );
  XNOR U1384 ( .A(n12982), .B(n12981), .Z(n12984) );
  XNOR U1385 ( .A(n13045), .B(n13044), .Z(n13060) );
  XOR U1386 ( .A(n13468), .B(n13467), .Z(n13466) );
  XOR U1387 ( .A(n13332), .B(n13331), .Z(n13330) );
  XNOR U1388 ( .A(n13145), .B(n13144), .Z(n13147) );
  XNOR U1389 ( .A(n12993), .B(n12992), .Z(n12994) );
  XNOR U1390 ( .A(n13157), .B(n13156), .Z(n13158) );
  XNOR U1391 ( .A(n13151), .B(n13150), .Z(n13152) );
  NAND U1392 ( .A(n13806), .B(n13805), .Z(n660) );
  AND U1393 ( .A(n13804), .B(y[59]), .Z(n661) );
  NAND U1394 ( .A(x[131]), .B(n661), .Z(n662) );
  AND U1395 ( .A(n660), .B(n662), .Z(n13997) );
  NAND U1396 ( .A(n13840), .B(n13839), .Z(n663) );
  NAND U1397 ( .A(n13837), .B(n13838), .Z(n664) );
  AND U1398 ( .A(n663), .B(n664), .Z(n14151) );
  NAND U1399 ( .A(n13733), .B(n13732), .Z(n665) );
  NAND U1400 ( .A(n13730), .B(n13731), .Z(n666) );
  NAND U1401 ( .A(n665), .B(n666), .Z(n13865) );
  NAND U1402 ( .A(n13823), .B(n13822), .Z(n667) );
  NANDN U1403 ( .A(n13821), .B(n13964), .Z(n668) );
  AND U1404 ( .A(n667), .B(n668), .Z(n14142) );
  NAND U1405 ( .A(n13779), .B(n13778), .Z(n669) );
  NAND U1406 ( .A(n13776), .B(n13777), .Z(n670) );
  NAND U1407 ( .A(n669), .B(n670), .Z(n13901) );
  XOR U1408 ( .A(n14471), .B(n14470), .Z(n14446) );
  XOR U1409 ( .A(n14762), .B(n14761), .Z(n14760) );
  XNOR U1410 ( .A(n14891), .B(n14892), .Z(n14889) );
  XNOR U1411 ( .A(n15623), .B(n15622), .Z(n15620) );
  NAND U1412 ( .A(n15278), .B(n15318), .Z(n671) );
  NANDN U1413 ( .A(n15178), .B(n15177), .Z(n672) );
  AND U1414 ( .A(n671), .B(n672), .Z(n15300) );
  XOR U1415 ( .A(n15517), .B(n15516), .Z(n15515) );
  XOR U1416 ( .A(n15193), .B(n15192), .Z(n15147) );
  NAND U1417 ( .A(n15791), .B(n15790), .Z(n673) );
  NANDN U1418 ( .A(n15789), .B(n15788), .Z(n674) );
  AND U1419 ( .A(n673), .B(n674), .Z(n15865) );
  XOR U1420 ( .A(n15912), .B(n15911), .Z(n15871) );
  XNOR U1421 ( .A(n15879), .B(n15878), .Z(n15955) );
  XNOR U1422 ( .A(n16358), .B(n16357), .Z(n16355) );
  XOR U1423 ( .A(n16224), .B(n16223), .Z(n16222) );
  XNOR U1424 ( .A(n16035), .B(n16034), .Z(n16037) );
  XNOR U1425 ( .A(n15888), .B(n15887), .Z(n15889) );
  XNOR U1426 ( .A(n16047), .B(n16046), .Z(n16048) );
  XNOR U1427 ( .A(n16041), .B(n16040), .Z(n16042) );
  XNOR U1428 ( .A(n16681), .B(n16680), .Z(n16682) );
  XNOR U1429 ( .A(n16687), .B(n16686), .Z(n16688) );
  XNOR U1430 ( .A(n16675), .B(n16674), .Z(n16677) );
  NAND U1431 ( .A(n16663), .B(n16662), .Z(n675) );
  NANDN U1432 ( .A(n16665), .B(n16664), .Z(n676) );
  AND U1433 ( .A(n675), .B(n676), .Z(n16763) );
  NAND U1434 ( .A(n16627), .B(n16626), .Z(n677) );
  NAND U1435 ( .A(n16624), .B(n16625), .Z(n678) );
  NAND U1436 ( .A(n677), .B(n678), .Z(n16797) );
  XNOR U1437 ( .A(n17024), .B(n17023), .Z(n17021) );
  XNOR U1438 ( .A(n16901), .B(n16900), .Z(n16898) );
  NAND U1439 ( .A(n16731), .B(n16730), .Z(n679) );
  NAND U1440 ( .A(n16728), .B(n16729), .Z(n680) );
  NAND U1441 ( .A(n679), .B(n680), .Z(n17044) );
  NAND U1442 ( .A(n16750), .B(n16749), .Z(n681) );
  NANDN U1443 ( .A(n16748), .B(n16871), .Z(n682) );
  AND U1444 ( .A(n681), .B(n682), .Z(n17028) );
  NAND U1445 ( .A(n16623), .B(n16622), .Z(n683) );
  NAND U1446 ( .A(n16621), .B(n16620), .Z(n684) );
  AND U1447 ( .A(n683), .B(n684), .Z(n16719) );
  NAND U1448 ( .A(n17213), .B(n17212), .Z(n685) );
  NANDN U1449 ( .A(n17211), .B(n17210), .Z(n686) );
  AND U1450 ( .A(n685), .B(n686), .Z(n17285) );
  XOR U1451 ( .A(n17333), .B(n17332), .Z(n17291) );
  XNOR U1452 ( .A(n17299), .B(n17298), .Z(n17374) );
  XNOR U1453 ( .A(n17772), .B(n17773), .Z(n17770) );
  XNOR U1454 ( .A(n17643), .B(n17642), .Z(n17640) );
  XNOR U1455 ( .A(n17401), .B(n17400), .Z(n17403) );
  XNOR U1456 ( .A(n17450), .B(n17449), .Z(n17452) );
  XNOR U1457 ( .A(n17308), .B(n17307), .Z(n17309) );
  XNOR U1458 ( .A(n17468), .B(n17467), .Z(n17469) );
  XNOR U1459 ( .A(n17462), .B(n17461), .Z(n17463) );
  XOR U1460 ( .A(n18082), .B(n18081), .Z(n18033) );
  XNOR U1461 ( .A(n18516), .B(n18515), .Z(n18513) );
  XNOR U1462 ( .A(n18428), .B(n18427), .Z(n18425) );
  XOR U1463 ( .A(n18380), .B(n18379), .Z(n18378) );
  XNOR U1464 ( .A(n18935), .B(n18934), .Z(n18937) );
  XNOR U1465 ( .A(n18965), .B(n18964), .Z(n18966) );
  XNOR U1466 ( .A(n18893), .B(n18892), .Z(n18894) );
  XOR U1467 ( .A(n19274), .B(n19275), .Z(n19276) );
  XOR U1468 ( .A(n19078), .B(n19077), .Z(n19076) );
  XOR U1469 ( .A(n19156), .B(n19155), .Z(n19154) );
  XNOR U1470 ( .A(n18947), .B(n18946), .Z(n18949) );
  XNOR U1471 ( .A(n18901), .B(n18900), .Z(n18953) );
  XNOR U1472 ( .A(n18905), .B(n18904), .Z(n18907) );
  NAND U1473 ( .A(n1121), .B(n1120), .Z(n687) );
  NAND U1474 ( .A(n1119), .B(n1230), .Z(n688) );
  AND U1475 ( .A(n687), .B(n688), .Z(n1138) );
  NAND U1476 ( .A(n1487), .B(n1486), .Z(n689) );
  NAND U1477 ( .A(n1484), .B(n1485), .Z(n690) );
  AND U1478 ( .A(n689), .B(n690), .Z(n1800) );
  NAND U1479 ( .A(n1471), .B(n1470), .Z(n691) );
  NAND U1480 ( .A(n1468), .B(n1469), .Z(n692) );
  AND U1481 ( .A(n691), .B(n692), .Z(n1794) );
  NAND U1482 ( .A(n1452), .B(n1451), .Z(n693) );
  NAND U1483 ( .A(n1449), .B(n1450), .Z(n694) );
  AND U1484 ( .A(n693), .B(n694), .Z(n1534) );
  NAND U1485 ( .A(n1509), .B(n1508), .Z(n695) );
  NAND U1486 ( .A(n1506), .B(n1507), .Z(n696) );
  AND U1487 ( .A(n695), .B(n696), .Z(n1772) );
  NAND U1488 ( .A(n1494), .B(n1495), .Z(n697) );
  NAND U1489 ( .A(n1496), .B(n1701), .Z(n698) );
  AND U1490 ( .A(n697), .B(n698), .Z(n1540) );
  NAND U1491 ( .A(n1843), .B(n1842), .Z(n699) );
  NAND U1492 ( .A(n1841), .B(n1977), .Z(n700) );
  AND U1493 ( .A(n699), .B(n700), .Z(n1860) );
  XNOR U1494 ( .A(n2209), .B(n2208), .Z(n2149) );
  XOR U1495 ( .A(n2341), .B(n2340), .Z(n2549) );
  XOR U1496 ( .A(n2311), .B(n2310), .Z(n2309) );
  XNOR U1497 ( .A(n2565), .B(n2564), .Z(n2299) );
  NAND U1498 ( .A(n2602), .B(n2601), .Z(n701) );
  NAND U1499 ( .A(n2600), .B(n2712), .Z(n702) );
  AND U1500 ( .A(n701), .B(n702), .Z(n2619) );
  NAND U1501 ( .A(n3324), .B(n3323), .Z(n703) );
  NAND U1502 ( .A(n3322), .B(n3458), .Z(n704) );
  AND U1503 ( .A(n703), .B(n704), .Z(n3341) );
  XOR U1504 ( .A(n3678), .B(n3677), .Z(n3761) );
  XNOR U1505 ( .A(n3754), .B(n3753), .Z(n3755) );
  XNOR U1506 ( .A(n4028), .B(n4029), .Z(n4026) );
  XNOR U1507 ( .A(n3786), .B(n3785), .Z(n3783) );
  NAND U1508 ( .A(n4064), .B(n4063), .Z(n705) );
  NAND U1509 ( .A(n4062), .B(n4194), .Z(n706) );
  AND U1510 ( .A(n705), .B(n706), .Z(n4081) );
  NAND U1511 ( .A(n4163), .B(n4162), .Z(n707) );
  NAND U1512 ( .A(n4161), .B(n4160), .Z(n708) );
  AND U1513 ( .A(n707), .B(n708), .Z(n4244) );
  NAND U1514 ( .A(n4776), .B(n4775), .Z(n709) );
  NAND U1515 ( .A(n4774), .B(n4906), .Z(n710) );
  AND U1516 ( .A(n709), .B(n710), .Z(n4793) );
  NAND U1517 ( .A(n4875), .B(n4874), .Z(n711) );
  NAND U1518 ( .A(n4873), .B(n4872), .Z(n712) );
  AND U1519 ( .A(n711), .B(n712), .Z(n4960) );
  NAND U1520 ( .A(n5492), .B(n5491), .Z(n713) );
  NAND U1521 ( .A(n5490), .B(n5626), .Z(n714) );
  AND U1522 ( .A(n713), .B(n714), .Z(n5509) );
  NAND U1523 ( .A(n6233), .B(n6232), .Z(n715) );
  NAND U1524 ( .A(n6231), .B(n6364), .Z(n716) );
  AND U1525 ( .A(n715), .B(n716), .Z(n6250) );
  NAND U1526 ( .A(n6419), .B(n6418), .Z(n717) );
  NAND U1527 ( .A(n6417), .B(n6416), .Z(n718) );
  AND U1528 ( .A(n717), .B(n718), .Z(n6665) );
  XNOR U1529 ( .A(n6939), .B(n6938), .Z(n6936) );
  NAND U1530 ( .A(n6596), .B(n6595), .Z(n719) );
  NANDN U1531 ( .A(n6598), .B(n6597), .Z(n720) );
  AND U1532 ( .A(n719), .B(n720), .Z(n6698) );
  XNOR U1533 ( .A(n6686), .B(n6685), .Z(n6683) );
  XNOR U1534 ( .A(n6963), .B(n6962), .Z(n6961) );
  NAND U1535 ( .A(n6531), .B(n6530), .Z(n721) );
  NANDN U1536 ( .A(n6529), .B(n6528), .Z(n722) );
  AND U1537 ( .A(n721), .B(n722), .Z(n6957) );
  NAND U1538 ( .A(n6984), .B(n6983), .Z(n723) );
  NAND U1539 ( .A(n6982), .B(n7093), .Z(n724) );
  AND U1540 ( .A(n723), .B(n724), .Z(n7001) );
  NAND U1541 ( .A(n7360), .B(n7359), .Z(n725) );
  NAND U1542 ( .A(n7357), .B(n7358), .Z(n726) );
  AND U1543 ( .A(n725), .B(n726), .Z(n7643) );
  NAND U1544 ( .A(n7314), .B(n7313), .Z(n727) );
  NAND U1545 ( .A(n7311), .B(n7312), .Z(n728) );
  AND U1546 ( .A(n727), .B(n728), .Z(n7639) );
  NAND U1547 ( .A(n7343), .B(n7342), .Z(n729) );
  NANDN U1548 ( .A(n7341), .B(n7527), .Z(n730) );
  AND U1549 ( .A(n729), .B(n730), .Z(n7620) );
  NAND U1550 ( .A(n7330), .B(n7329), .Z(n731) );
  NAND U1551 ( .A(n7327), .B(n7328), .Z(n732) );
  AND U1552 ( .A(n731), .B(n732), .Z(n7393) );
  NAND U1553 ( .A(n7279), .B(n7278), .Z(n733) );
  NAND U1554 ( .A(n7276), .B(n7277), .Z(n734) );
  AND U1555 ( .A(n733), .B(n734), .Z(n7389) );
  NAND U1556 ( .A(n7243), .B(n7242), .Z(n735) );
  NAND U1557 ( .A(n7240), .B(n7241), .Z(n736) );
  NAND U1558 ( .A(n735), .B(n736), .Z(n7331) );
  NAND U1559 ( .A(n7688), .B(n7687), .Z(n737) );
  NAND U1560 ( .A(n7686), .B(n7818), .Z(n738) );
  AND U1561 ( .A(n737), .B(n738), .Z(n7705) );
  NAND U1562 ( .A(n7787), .B(n7786), .Z(n739) );
  NAND U1563 ( .A(n7785), .B(n7784), .Z(n740) );
  AND U1564 ( .A(n739), .B(n740), .Z(n7872) );
  NAND U1565 ( .A(n8421), .B(n8420), .Z(n741) );
  NAND U1566 ( .A(n8419), .B(n8555), .Z(n742) );
  AND U1567 ( .A(n741), .B(n742), .Z(n8438) );
  NAND U1568 ( .A(n9143), .B(n9142), .Z(n743) );
  NAND U1569 ( .A(n9141), .B(n9272), .Z(n744) );
  AND U1570 ( .A(n743), .B(n744), .Z(n9160) );
  NAND U1571 ( .A(n9328), .B(n9327), .Z(n745) );
  NAND U1572 ( .A(n9326), .B(n9325), .Z(n746) );
  AND U1573 ( .A(n745), .B(n746), .Z(n9560) );
  NAND U1574 ( .A(n9509), .B(n9508), .Z(n747) );
  NANDN U1575 ( .A(n9511), .B(n9510), .Z(n748) );
  AND U1576 ( .A(n747), .B(n748), .Z(n9814) );
  NAND U1577 ( .A(n9497), .B(n9496), .Z(n749) );
  NAND U1578 ( .A(n9494), .B(n9495), .Z(n750) );
  AND U1579 ( .A(n749), .B(n750), .Z(n9581) );
  NAND U1580 ( .A(n9456), .B(n9455), .Z(n751) );
  NAND U1581 ( .A(n9453), .B(n9454), .Z(n752) );
  NAND U1582 ( .A(n751), .B(n752), .Z(n9592) );
  NAND U1583 ( .A(n9434), .B(n9433), .Z(n753) );
  NANDN U1584 ( .A(n9432), .B(n9431), .Z(n754) );
  AND U1585 ( .A(n753), .B(n754), .Z(n9834) );
  NAND U1586 ( .A(n9861), .B(n9860), .Z(n755) );
  NAND U1587 ( .A(n9859), .B(n9992), .Z(n756) );
  AND U1588 ( .A(n755), .B(n756), .Z(n9878) );
  NAND U1589 ( .A(n10048), .B(n10047), .Z(n757) );
  NAND U1590 ( .A(n10046), .B(n10045), .Z(n758) );
  AND U1591 ( .A(n757), .B(n758), .Z(n10279) );
  XNOR U1592 ( .A(n10539), .B(n10540), .Z(n10542) );
  NAND U1593 ( .A(n10228), .B(n10227), .Z(n759) );
  NANDN U1594 ( .A(n10230), .B(n10229), .Z(n760) );
  AND U1595 ( .A(n759), .B(n760), .Z(n10534) );
  NAND U1596 ( .A(n10216), .B(n10215), .Z(n761) );
  NAND U1597 ( .A(n10213), .B(n10214), .Z(n762) );
  AND U1598 ( .A(n761), .B(n762), .Z(n10300) );
  NAND U1599 ( .A(n10174), .B(n10173), .Z(n763) );
  NAND U1600 ( .A(n10171), .B(n10172), .Z(n764) );
  NAND U1601 ( .A(n763), .B(n764), .Z(n10311) );
  NAND U1602 ( .A(n10152), .B(n10151), .Z(n765) );
  NANDN U1603 ( .A(n10150), .B(n10149), .Z(n766) );
  AND U1604 ( .A(n765), .B(n766), .Z(n10554) );
  XNOR U1605 ( .A(n10744), .B(n10743), .Z(n10746) );
  NAND U1606 ( .A(n10623), .B(n10622), .Z(n767) );
  NAND U1607 ( .A(n10621), .B(n10620), .Z(n768) );
  AND U1608 ( .A(n767), .B(n768), .Z(n10732) );
  NAND U1609 ( .A(n11294), .B(n11293), .Z(n769) );
  NAND U1610 ( .A(n11292), .B(n11428), .Z(n770) );
  AND U1611 ( .A(n769), .B(n770), .Z(n11311) );
  NAND U1612 ( .A(n12034), .B(n12033), .Z(n771) );
  NAND U1613 ( .A(n12032), .B(n12144), .Z(n772) );
  AND U1614 ( .A(n771), .B(n772), .Z(n12051) );
  NAND U1615 ( .A(n12777), .B(n12776), .Z(n773) );
  NAND U1616 ( .A(n12775), .B(n12907), .Z(n774) );
  AND U1617 ( .A(n773), .B(n774), .Z(n12794) );
  NAND U1618 ( .A(n12875), .B(n12874), .Z(n775) );
  NAND U1619 ( .A(n12873), .B(n12872), .Z(n776) );
  AND U1620 ( .A(n775), .B(n776), .Z(n12960) );
  NAND U1621 ( .A(n13714), .B(n13713), .Z(n777) );
  NANDN U1622 ( .A(n13712), .B(n13711), .Z(n778) );
  NAND U1623 ( .A(n777), .B(n778), .Z(n13827) );
  NAND U1624 ( .A(n13850), .B(n13849), .Z(n779) );
  NAND U1625 ( .A(n13848), .B(n13847), .Z(n780) );
  AND U1626 ( .A(n779), .B(n780), .Z(n14172) );
  NAND U1627 ( .A(n13985), .B(n13984), .Z(n781) );
  NAND U1628 ( .A(n13986), .B(n13987), .Z(n782) );
  AND U1629 ( .A(n781), .B(n782), .Z(n783) );
  NAND U1630 ( .A(n13989), .B(n13988), .Z(n784) );
  NAND U1631 ( .A(n13990), .B(n13991), .Z(n785) );
  NAND U1632 ( .A(n784), .B(n785), .Z(n786) );
  XNOR U1633 ( .A(n783), .B(n786), .Z(n13992) );
  XNOR U1634 ( .A(n13934), .B(n13933), .Z(n13931) );
  NAND U1635 ( .A(n13729), .B(n13728), .Z(n787) );
  NAND U1636 ( .A(n13726), .B(n13727), .Z(n788) );
  NAND U1637 ( .A(n787), .B(n788), .Z(n13809) );
  NAND U1638 ( .A(n13799), .B(n13798), .Z(n789) );
  NAND U1639 ( .A(n13796), .B(n13797), .Z(n790) );
  NAND U1640 ( .A(n789), .B(n790), .Z(n14155) );
  NAND U1641 ( .A(n14219), .B(n14218), .Z(n791) );
  NAND U1642 ( .A(n14217), .B(n14328), .Z(n792) );
  AND U1643 ( .A(n791), .B(n792), .Z(n14236) );
  NAND U1644 ( .A(n14942), .B(n14941), .Z(n793) );
  NAND U1645 ( .A(n14940), .B(n15054), .Z(n794) );
  AND U1646 ( .A(n793), .B(n794), .Z(n14959) );
  XNOR U1647 ( .A(n15135), .B(n15134), .Z(n15137) );
  NAND U1648 ( .A(n15670), .B(n15669), .Z(n795) );
  NAND U1649 ( .A(n15668), .B(n15814), .Z(n796) );
  AND U1650 ( .A(n795), .B(n796), .Z(n15687) );
  NAND U1651 ( .A(n15769), .B(n15768), .Z(n797) );
  NAND U1652 ( .A(n15767), .B(n15766), .Z(n798) );
  AND U1653 ( .A(n797), .B(n798), .Z(n15855) );
  NAND U1654 ( .A(n16406), .B(n16405), .Z(n799) );
  NAND U1655 ( .A(n16404), .B(n16539), .Z(n800) );
  AND U1656 ( .A(n799), .B(n800), .Z(n16423) );
  NAND U1657 ( .A(n17091), .B(n17090), .Z(n801) );
  NAND U1658 ( .A(n17089), .B(n17222), .Z(n802) );
  AND U1659 ( .A(n801), .B(n802), .Z(n17108) );
  NAND U1660 ( .A(n17191), .B(n17190), .Z(n803) );
  NAND U1661 ( .A(n17189), .B(n17188), .Z(n804) );
  AND U1662 ( .A(n803), .B(n804), .Z(n17275) );
  NAND U1663 ( .A(n17827), .B(n17826), .Z(n805) );
  NAND U1664 ( .A(n17825), .B(n17970), .Z(n806) );
  AND U1665 ( .A(n805), .B(n806), .Z(n17844) );
  NAND U1666 ( .A(n18013), .B(n18012), .Z(n807) );
  NAND U1667 ( .A(n18011), .B(n18010), .Z(n808) );
  AND U1668 ( .A(n807), .B(n808), .Z(n18262) );
  XNOR U1669 ( .A(n18542), .B(n18541), .Z(n18540) );
  XNOR U1670 ( .A(n18295), .B(n18294), .Z(n18292) );
  XNOR U1671 ( .A(n18560), .B(n18559), .Z(n18558) );
  NAND U1672 ( .A(n18128), .B(n18127), .Z(n809) );
  NANDN U1673 ( .A(n18126), .B(n18125), .Z(n810) );
  AND U1674 ( .A(n809), .B(n810), .Z(n18554) );
  NAND U1675 ( .A(n18581), .B(n18580), .Z(n811) );
  NAND U1676 ( .A(n18579), .B(n18715), .Z(n812) );
  AND U1677 ( .A(n811), .B(n812), .Z(n18598) );
  XNOR U1678 ( .A(n1315), .B(n1314), .Z(n1310) );
  XOR U1679 ( .A(n1815), .B(n1816), .Z(n813) );
  NAND U1680 ( .A(n1814), .B(n813), .Z(n1817) );
  XNOR U1681 ( .A(n2293), .B(n2292), .Z(n2291) );
  XNOR U1682 ( .A(n2791), .B(n2790), .Z(n2786) );
  XNOR U1683 ( .A(n3774), .B(n3773), .Z(n3772) );
  XNOR U1684 ( .A(n6824), .B(n6823), .Z(n6677) );
  XNOR U1685 ( .A(n7172), .B(n7171), .Z(n7167) );
  XOR U1686 ( .A(n7660), .B(n7661), .Z(n814) );
  NAND U1687 ( .A(n7659), .B(n814), .Z(n7662) );
  NAND U1688 ( .A(n9467), .B(n9466), .Z(n815) );
  NAND U1689 ( .A(n9464), .B(n9465), .Z(n816) );
  NAND U1690 ( .A(n815), .B(n816), .Z(n9574) );
  NAND U1691 ( .A(n10185), .B(n10184), .Z(n817) );
  NAND U1692 ( .A(n10182), .B(n10183), .Z(n818) );
  NAND U1693 ( .A(n817), .B(n818), .Z(n10293) );
  NAND U1694 ( .A(n13671), .B(n13672), .Z(n819) );
  XOR U1695 ( .A(n13671), .B(n13672), .Z(n820) );
  NANDN U1696 ( .A(n13670), .B(n820), .Z(n821) );
  NAND U1697 ( .A(n819), .B(n821), .Z(n13693) );
  XNOR U1698 ( .A(n14210), .B(n14209), .Z(n14208) );
  XNOR U1699 ( .A(n14412), .B(n14411), .Z(n14407) );
  NAND U1700 ( .A(n15105), .B(n15104), .Z(n822) );
  NAND U1701 ( .A(n15102), .B(n15103), .Z(n823) );
  NAND U1702 ( .A(n822), .B(n823), .Z(n15125) );
  NAND U1703 ( .A(n18146), .B(n18145), .Z(n824) );
  NANDN U1704 ( .A(n18148), .B(n18147), .Z(n825) );
  AND U1705 ( .A(n824), .B(n825), .Z(n18275) );
  NAND U1706 ( .A(n3028), .B(n3029), .Z(n826) );
  NANDN U1707 ( .A(n3031), .B(n3030), .Z(n827) );
  AND U1708 ( .A(n826), .B(n827), .Z(n828) );
  NAND U1709 ( .A(n3034), .B(n3035), .Z(n829) );
  NANDN U1710 ( .A(n3033), .B(n3032), .Z(n830) );
  AND U1711 ( .A(n829), .B(n830), .Z(n831) );
  AND U1712 ( .A(n3316), .B(n3315), .Z(n832) );
  NAND U1713 ( .A(n3310), .B(n3309), .Z(n833) );
  XNOR U1714 ( .A(n832), .B(n833), .Z(n834) );
  XOR U1715 ( .A(n3304), .B(n834), .Z(n835) );
  XNOR U1716 ( .A(n3289), .B(n3288), .Z(n836) );
  XNOR U1717 ( .A(n835), .B(n836), .Z(n837) );
  XNOR U1718 ( .A(n828), .B(n831), .Z(n838) );
  XNOR U1719 ( .A(n837), .B(n838), .Z(n839) );
  XOR U1720 ( .A(n3317), .B(n3318), .Z(n840) );
  NANDN U1721 ( .A(n3319), .B(n840), .Z(n841) );
  NAND U1722 ( .A(n3317), .B(n3318), .Z(n842) );
  AND U1723 ( .A(n841), .B(n842), .Z(n843) );
  XNOR U1724 ( .A(n839), .B(n843), .Z(o[23]) );
  XOR U1725 ( .A(n4755), .B(n4754), .Z(n844) );
  XNOR U1726 ( .A(n4741), .B(n4740), .Z(n845) );
  XNOR U1727 ( .A(n844), .B(n845), .Z(n846) );
  AND U1728 ( .A(n4767), .B(n4766), .Z(n847) );
  NAND U1729 ( .A(n4761), .B(n4760), .Z(n848) );
  XNOR U1730 ( .A(n847), .B(n848), .Z(n849) );
  XOR U1731 ( .A(n846), .B(n849), .Z(n850) );
  NAND U1732 ( .A(n4482), .B(n4481), .Z(n851) );
  NANDN U1733 ( .A(n4484), .B(n4483), .Z(n852) );
  AND U1734 ( .A(n851), .B(n852), .Z(n853) );
  NAND U1735 ( .A(n4485), .B(n4486), .Z(n854) );
  NAND U1736 ( .A(n4487), .B(n4488), .Z(n855) );
  AND U1737 ( .A(n854), .B(n855), .Z(n856) );
  XNOR U1738 ( .A(n853), .B(n856), .Z(n857) );
  XNOR U1739 ( .A(n850), .B(n857), .Z(n858) );
  NANDN U1740 ( .A(n4771), .B(n4770), .Z(n859) );
  NANDN U1741 ( .A(n4769), .B(n4768), .Z(n860) );
  NAND U1742 ( .A(n859), .B(n860), .Z(n861) );
  XNOR U1743 ( .A(n858), .B(n861), .Z(o[39]) );
  NAND U1744 ( .A(n5214), .B(n5215), .Z(n862) );
  NANDN U1745 ( .A(n5217), .B(n5216), .Z(n863) );
  AND U1746 ( .A(n862), .B(n863), .Z(n864) );
  NAND U1747 ( .A(n5221), .B(n5220), .Z(n865) );
  NANDN U1748 ( .A(n5219), .B(n5218), .Z(n866) );
  AND U1749 ( .A(n865), .B(n866), .Z(n867) );
  XOR U1750 ( .A(n5471), .B(n5470), .Z(n868) );
  XNOR U1751 ( .A(n5457), .B(n5456), .Z(n869) );
  XNOR U1752 ( .A(n868), .B(n869), .Z(n870) );
  AND U1753 ( .A(n5483), .B(n5482), .Z(n871) );
  NAND U1754 ( .A(n5477), .B(n5476), .Z(n872) );
  XNOR U1755 ( .A(n871), .B(n872), .Z(n873) );
  XOR U1756 ( .A(n870), .B(n873), .Z(n874) );
  XNOR U1757 ( .A(n864), .B(n867), .Z(n875) );
  XNOR U1758 ( .A(n874), .B(n875), .Z(n876) );
  NAND U1759 ( .A(n5487), .B(n5486), .Z(n877) );
  NANDN U1760 ( .A(n5485), .B(n5484), .Z(n878) );
  NAND U1761 ( .A(n877), .B(n878), .Z(n879) );
  XNOR U1762 ( .A(n876), .B(n879), .Z(o[47]) );
  ANDN U1763 ( .B(n6222), .A(n6221), .Z(n880) );
  OR U1764 ( .A(n6227), .B(n6228), .Z(n881) );
  XNOR U1765 ( .A(n880), .B(n881), .Z(n882) );
  XOR U1766 ( .A(n6216), .B(n882), .Z(n883) );
  XNOR U1767 ( .A(n6201), .B(n6200), .Z(n884) );
  XNOR U1768 ( .A(n883), .B(n884), .Z(n885) );
  NAND U1769 ( .A(n5942), .B(n5941), .Z(n886) );
  NANDN U1770 ( .A(n5944), .B(n5943), .Z(n887) );
  AND U1771 ( .A(n886), .B(n887), .Z(n888) );
  NAND U1772 ( .A(n5945), .B(n5946), .Z(n889) );
  NAND U1773 ( .A(n5947), .B(n5948), .Z(n890) );
  AND U1774 ( .A(n889), .B(n890), .Z(n891) );
  XNOR U1775 ( .A(n888), .B(n891), .Z(n892) );
  XNOR U1776 ( .A(n885), .B(n892), .Z(n893) );
  NANDN U1777 ( .A(n5938), .B(n5939), .Z(n894) );
  XNOR U1778 ( .A(n5938), .B(n5939), .Z(n895) );
  NAND U1779 ( .A(n5940), .B(n895), .Z(n896) );
  AND U1780 ( .A(n894), .B(n896), .Z(n897) );
  XNOR U1781 ( .A(n893), .B(n897), .Z(o[55]) );
  NAND U1782 ( .A(n8131), .B(n8130), .Z(n898) );
  NANDN U1783 ( .A(n8133), .B(n8132), .Z(n899) );
  AND U1784 ( .A(n898), .B(n899), .Z(n900) );
  NAND U1785 ( .A(n8134), .B(n8135), .Z(n901) );
  NAND U1786 ( .A(n8136), .B(n8137), .Z(n902) );
  AND U1787 ( .A(n901), .B(n902), .Z(n903) );
  AND U1788 ( .A(n8409), .B(n8410), .Z(n904) );
  OR U1789 ( .A(n8415), .B(n8416), .Z(n905) );
  XNOR U1790 ( .A(n904), .B(n905), .Z(n906) );
  XOR U1791 ( .A(n8404), .B(n906), .Z(n907) );
  XNOR U1792 ( .A(n8389), .B(n8388), .Z(n908) );
  XNOR U1793 ( .A(n907), .B(n908), .Z(n909) );
  XNOR U1794 ( .A(n900), .B(n903), .Z(n910) );
  XNOR U1795 ( .A(n909), .B(n910), .Z(n911) );
  NANDN U1796 ( .A(n8127), .B(n8128), .Z(n912) );
  XNOR U1797 ( .A(n8127), .B(n8128), .Z(n913) );
  NAND U1798 ( .A(n8129), .B(n913), .Z(n914) );
  AND U1799 ( .A(n912), .B(n914), .Z(n915) );
  XNOR U1800 ( .A(n911), .B(n915), .Z(o[79]) );
  NAND U1801 ( .A(n8863), .B(n8864), .Z(n916) );
  NANDN U1802 ( .A(n8866), .B(n8865), .Z(n917) );
  AND U1803 ( .A(n916), .B(n917), .Z(n918) );
  NAND U1804 ( .A(n8867), .B(n8868), .Z(n919) );
  NAND U1805 ( .A(n8870), .B(n8869), .Z(n920) );
  AND U1806 ( .A(n919), .B(n920), .Z(n921) );
  XOR U1807 ( .A(n9122), .B(n9121), .Z(n922) );
  XNOR U1808 ( .A(n9108), .B(n9107), .Z(n923) );
  XNOR U1809 ( .A(n922), .B(n923), .Z(n924) );
  AND U1810 ( .A(n9134), .B(n9133), .Z(n925) );
  NAND U1811 ( .A(n9128), .B(n9127), .Z(n926) );
  XNOR U1812 ( .A(n925), .B(n926), .Z(n927) );
  XOR U1813 ( .A(n924), .B(n927), .Z(n928) );
  XNOR U1814 ( .A(n918), .B(n921), .Z(n929) );
  XNOR U1815 ( .A(n928), .B(n929), .Z(n930) );
  NAND U1816 ( .A(n9138), .B(n9137), .Z(n931) );
  NANDN U1817 ( .A(n9136), .B(n9135), .Z(n932) );
  NAND U1818 ( .A(n931), .B(n932), .Z(n933) );
  XNOR U1819 ( .A(n930), .B(n933), .Z(o[87]) );
  NAND U1820 ( .A(n10999), .B(n11000), .Z(n934) );
  NAND U1821 ( .A(n11001), .B(n11002), .Z(n935) );
  AND U1822 ( .A(n934), .B(n935), .Z(n936) );
  OR U1823 ( .A(n11005), .B(n11006), .Z(n937) );
  NAND U1824 ( .A(n11003), .B(n11004), .Z(n938) );
  AND U1825 ( .A(n937), .B(n938), .Z(n939) );
  AND U1826 ( .A(n11012), .B(n11011), .Z(n940) );
  XNOR U1827 ( .A(n11281), .B(n11280), .Z(n941) );
  XNOR U1828 ( .A(n940), .B(n941), .Z(n942) );
  NAND U1829 ( .A(n11284), .B(n11285), .Z(n943) );
  NAND U1830 ( .A(n11282), .B(n11283), .Z(n944) );
  AND U1831 ( .A(n943), .B(n944), .Z(n945) );
  NAND U1832 ( .A(n11288), .B(n11289), .Z(n946) );
  NANDN U1833 ( .A(n11287), .B(n11286), .Z(n947) );
  AND U1834 ( .A(n946), .B(n947), .Z(n948) );
  XOR U1835 ( .A(n945), .B(n948), .Z(n949) );
  XNOR U1836 ( .A(n939), .B(n942), .Z(n950) );
  XNOR U1837 ( .A(n949), .B(n950), .Z(n951) );
  XNOR U1838 ( .A(n936), .B(n951), .Z(o[111]) );
  NAND U1839 ( .A(n11740), .B(n11741), .Z(n952) );
  NANDN U1840 ( .A(n11743), .B(n11742), .Z(n953) );
  AND U1841 ( .A(n952), .B(n953), .Z(n954) );
  XOR U1842 ( .A(n12018), .B(n12017), .Z(n955) );
  XNOR U1843 ( .A(n12004), .B(n12003), .Z(n956) );
  XNOR U1844 ( .A(n955), .B(n956), .Z(n957) );
  NAND U1845 ( .A(n12025), .B(n12024), .Z(n958) );
  NANDN U1846 ( .A(n12022), .B(n12023), .Z(n959) );
  AND U1847 ( .A(n958), .B(n959), .Z(n960) );
  NAND U1848 ( .A(n12028), .B(n12029), .Z(n961) );
  NAND U1849 ( .A(n12026), .B(n12027), .Z(n962) );
  AND U1850 ( .A(n961), .B(n962), .Z(n963) );
  NANDN U1851 ( .A(n12019), .B(n12020), .Z(n964) );
  XNOR U1852 ( .A(n12019), .B(n12020), .Z(n965) );
  NAND U1853 ( .A(n12021), .B(n965), .Z(n966) );
  AND U1854 ( .A(n964), .B(n966), .Z(n967) );
  XNOR U1855 ( .A(n963), .B(n967), .Z(n968) );
  XOR U1856 ( .A(n960), .B(n968), .Z(n969) );
  XNOR U1857 ( .A(n954), .B(n957), .Z(n970) );
  XNOR U1858 ( .A(n969), .B(n970), .Z(o[119]) );
  NAND U1859 ( .A(n12492), .B(n12491), .Z(n971) );
  XOR U1860 ( .A(n12492), .B(n12491), .Z(n972) );
  NANDN U1861 ( .A(n12490), .B(n972), .Z(n973) );
  NAND U1862 ( .A(n971), .B(n973), .Z(n974) );
  OR U1863 ( .A(n12481), .B(n12482), .Z(n975) );
  NAND U1864 ( .A(n12483), .B(n12484), .Z(n976) );
  AND U1865 ( .A(n975), .B(n976), .Z(n977) );
  NAND U1866 ( .A(n12485), .B(n12486), .Z(n978) );
  NANDN U1867 ( .A(n12488), .B(n12487), .Z(n979) );
  AND U1868 ( .A(n978), .B(n979), .Z(n980) );
  AND U1869 ( .A(n12498), .B(n12497), .Z(n981) );
  XNOR U1870 ( .A(n12760), .B(n12759), .Z(n982) );
  XNOR U1871 ( .A(n981), .B(n982), .Z(n983) );
  AND U1872 ( .A(n12772), .B(n12771), .Z(n984) );
  NAND U1873 ( .A(n12766), .B(n12765), .Z(n985) );
  XNOR U1874 ( .A(n984), .B(n985), .Z(n986) );
  XOR U1875 ( .A(n983), .B(n986), .Z(n987) );
  XNOR U1876 ( .A(n977), .B(n980), .Z(n988) );
  XNOR U1877 ( .A(n987), .B(n988), .Z(n989) );
  XNOR U1878 ( .A(n974), .B(n989), .Z(o[127]) );
  NAND U1879 ( .A(n13225), .B(n13224), .Z(n990) );
  NANDN U1880 ( .A(n13227), .B(n13226), .Z(n991) );
  AND U1881 ( .A(n990), .B(n991), .Z(n992) );
  NAND U1882 ( .A(n13230), .B(n13231), .Z(n993) );
  NANDN U1883 ( .A(n13229), .B(n13228), .Z(n994) );
  AND U1884 ( .A(n993), .B(n994), .Z(n995) );
  ANDN U1885 ( .B(n13505), .A(n13504), .Z(n996) );
  OR U1886 ( .A(n13510), .B(n13511), .Z(n997) );
  XNOR U1887 ( .A(n996), .B(n997), .Z(n998) );
  XOR U1888 ( .A(n13499), .B(n998), .Z(n999) );
  XNOR U1889 ( .A(n13484), .B(n13483), .Z(n1000) );
  XNOR U1890 ( .A(n999), .B(n1000), .Z(n1001) );
  XNOR U1891 ( .A(n992), .B(n995), .Z(n1002) );
  XNOR U1892 ( .A(n1001), .B(n1002), .Z(n1003) );
  NANDN U1893 ( .A(n13221), .B(n13222), .Z(n1004) );
  XNOR U1894 ( .A(n13221), .B(n13222), .Z(n1005) );
  NAND U1895 ( .A(n13223), .B(n1005), .Z(n1006) );
  AND U1896 ( .A(n1004), .B(n1006), .Z(n1007) );
  XNOR U1897 ( .A(n1003), .B(n1007), .Z(o[135]) );
  NAND U1898 ( .A(n14665), .B(n14664), .Z(n1008) );
  NANDN U1899 ( .A(n14667), .B(n14666), .Z(n1009) );
  AND U1900 ( .A(n1008), .B(n1009), .Z(n1010) );
  NAND U1901 ( .A(n14668), .B(n14669), .Z(n1011) );
  NAND U1902 ( .A(n14670), .B(n14671), .Z(n1012) );
  AND U1903 ( .A(n1011), .B(n1012), .Z(n1013) );
  AND U1904 ( .A(n14934), .B(n14933), .Z(n1014) );
  NAND U1905 ( .A(n14928), .B(n14927), .Z(n1015) );
  XNOR U1906 ( .A(n1014), .B(n1015), .Z(n1016) );
  XOR U1907 ( .A(n14921), .B(n1016), .Z(n1017) );
  XNOR U1908 ( .A(n1013), .B(n14922), .Z(n1018) );
  XNOR U1909 ( .A(n1017), .B(n1018), .Z(n1019) );
  NAND U1910 ( .A(n14936), .B(n14935), .Z(n1020) );
  XOR U1911 ( .A(n14936), .B(n14935), .Z(n1021) );
  NAND U1912 ( .A(n1021), .B(n14937), .Z(n1022) );
  NAND U1913 ( .A(n1020), .B(n1022), .Z(n1023) );
  XNOR U1914 ( .A(n1010), .B(n1019), .Z(n1024) );
  XNOR U1915 ( .A(n1023), .B(n1024), .Z(o[151]) );
  NANDN U1916 ( .A(n15374), .B(n15373), .Z(n1025) );
  NANDN U1917 ( .A(n15376), .B(n15375), .Z(n1026) );
  AND U1918 ( .A(n1025), .B(n1026), .Z(n1027) );
  XOR U1919 ( .A(n15653), .B(n15652), .Z(n1028) );
  XNOR U1920 ( .A(n15639), .B(n15638), .Z(n1029) );
  XNOR U1921 ( .A(n1028), .B(n1029), .Z(n1030) );
  OR U1922 ( .A(n15658), .B(n15657), .Z(n1031) );
  NANDN U1923 ( .A(n15656), .B(n15655), .Z(n1032) );
  AND U1924 ( .A(n1031), .B(n1032), .Z(n1033) );
  XNOR U1925 ( .A(n1027), .B(n1030), .Z(n1034) );
  XNOR U1926 ( .A(n1033), .B(n1034), .Z(n1035) );
  NANDN U1927 ( .A(n15659), .B(n15660), .Z(n1036) );
  XNOR U1928 ( .A(n15659), .B(n15660), .Z(n1037) );
  NAND U1929 ( .A(n15661), .B(n1037), .Z(n1038) );
  AND U1930 ( .A(n1036), .B(n1038), .Z(n1039) );
  XNOR U1931 ( .A(n1035), .B(n1039), .Z(n1040) );
  NAND U1932 ( .A(n15665), .B(n15664), .Z(n1041) );
  NANDN U1933 ( .A(n15663), .B(n15662), .Z(n1042) );
  NAND U1934 ( .A(n1041), .B(n1042), .Z(n1043) );
  XNOR U1935 ( .A(n1040), .B(n1043), .Z(o[159]) );
  ANDN U1936 ( .B(n16395), .A(n16394), .Z(n1044) );
  OR U1937 ( .A(n16400), .B(n16401), .Z(n1045) );
  XNOR U1938 ( .A(n1044), .B(n1045), .Z(n1046) );
  XOR U1939 ( .A(n16389), .B(n1046), .Z(n1047) );
  XNOR U1940 ( .A(n16374), .B(n16373), .Z(n1048) );
  XNOR U1941 ( .A(n1047), .B(n1048), .Z(n1049) );
  NAND U1942 ( .A(n16115), .B(n16114), .Z(n1050) );
  NANDN U1943 ( .A(n16117), .B(n16116), .Z(n1051) );
  AND U1944 ( .A(n1050), .B(n1051), .Z(n1052) );
  NAND U1945 ( .A(n16118), .B(n16119), .Z(n1053) );
  NAND U1946 ( .A(n16120), .B(n16121), .Z(n1054) );
  AND U1947 ( .A(n1053), .B(n1054), .Z(n1055) );
  XNOR U1948 ( .A(n1052), .B(n1055), .Z(n1056) );
  XNOR U1949 ( .A(n1049), .B(n1056), .Z(n1057) );
  NANDN U1950 ( .A(n16111), .B(n16112), .Z(n1058) );
  XNOR U1951 ( .A(n16111), .B(n16112), .Z(n1059) );
  NAND U1952 ( .A(n16113), .B(n1059), .Z(n1060) );
  AND U1953 ( .A(n1058), .B(n1060), .Z(n1061) );
  XNOR U1954 ( .A(n1057), .B(n1061), .Z(o[167]) );
  NAND U1955 ( .A(n16833), .B(n16832), .Z(n1062) );
  NANDN U1956 ( .A(n16835), .B(n16834), .Z(n1063) );
  AND U1957 ( .A(n1062), .B(n1063), .Z(n1064) );
  NAND U1958 ( .A(n16836), .B(n16837), .Z(n1065) );
  NAND U1959 ( .A(n16838), .B(n16839), .Z(n1066) );
  AND U1960 ( .A(n1065), .B(n1066), .Z(n1067) );
  XOR U1961 ( .A(n17070), .B(n17069), .Z(n1068) );
  XNOR U1962 ( .A(n17056), .B(n17055), .Z(n1069) );
  XNOR U1963 ( .A(n1068), .B(n1069), .Z(n1070) );
  AND U1964 ( .A(n17082), .B(n17081), .Z(n1071) );
  NAND U1965 ( .A(n17076), .B(n17075), .Z(n1072) );
  XNOR U1966 ( .A(n1071), .B(n1072), .Z(n1073) );
  XOR U1967 ( .A(n1070), .B(n1073), .Z(n1074) );
  XNOR U1968 ( .A(n1064), .B(n1067), .Z(n1075) );
  XNOR U1969 ( .A(n1074), .B(n1075), .Z(n1076) );
  NANDN U1970 ( .A(n17086), .B(n17085), .Z(n1077) );
  NANDN U1971 ( .A(n17084), .B(n17083), .Z(n1078) );
  NAND U1972 ( .A(n1077), .B(n1078), .Z(n1079) );
  XNOR U1973 ( .A(n1076), .B(n1079), .Z(o[175]) );
  NAND U1974 ( .A(n17536), .B(n17535), .Z(n1080) );
  NANDN U1975 ( .A(n17538), .B(n17537), .Z(n1081) );
  AND U1976 ( .A(n1080), .B(n1081), .Z(n1082) );
  NAND U1977 ( .A(n17539), .B(n17540), .Z(n1083) );
  NAND U1978 ( .A(n17541), .B(n17542), .Z(n1084) );
  AND U1979 ( .A(n1083), .B(n1084), .Z(n1085) );
  ANDN U1980 ( .B(n17816), .A(n17815), .Z(n1086) );
  OR U1981 ( .A(n17821), .B(n17822), .Z(n1087) );
  XNOR U1982 ( .A(n1086), .B(n1087), .Z(n1088) );
  XOR U1983 ( .A(n17810), .B(n1088), .Z(n1089) );
  XNOR U1984 ( .A(n17795), .B(n17794), .Z(n1090) );
  XNOR U1985 ( .A(n1089), .B(n1090), .Z(n1091) );
  XNOR U1986 ( .A(n1082), .B(n1085), .Z(n1092) );
  XNOR U1987 ( .A(n1091), .B(n1092), .Z(n1093) );
  NANDN U1988 ( .A(n17532), .B(n17533), .Z(n1094) );
  XNOR U1989 ( .A(n17532), .B(n17533), .Z(n1095) );
  NAND U1990 ( .A(n17534), .B(n1095), .Z(n1096) );
  AND U1991 ( .A(n1094), .B(n1096), .Z(n1097) );
  XNOR U1992 ( .A(n1093), .B(n1097), .Z(o[183]) );
  NAND U1993 ( .A(n19031), .B(n19032), .Z(n1098) );
  NANDN U1994 ( .A(n19033), .B(n19034), .Z(n1099) );
  AND U1995 ( .A(n1098), .B(n1099), .Z(n1100) );
  NAND U1996 ( .A(n19040), .B(n19039), .Z(n1101) );
  NAND U1997 ( .A(n19041), .B(n19042), .Z(n1102) );
  AND U1998 ( .A(n1101), .B(n1102), .Z(n1103) );
  XOR U1999 ( .A(n19317), .B(n19316), .Z(n1104) );
  XNOR U2000 ( .A(n19303), .B(n19302), .Z(n1105) );
  XNOR U2001 ( .A(n1104), .B(n1105), .Z(n1106) );
  NAND U2002 ( .A(n19035), .B(n19036), .Z(n1107) );
  NAND U2003 ( .A(n19037), .B(n19038), .Z(n1108) );
  AND U2004 ( .A(n1107), .B(n1108), .Z(n1109) );
  NAND U2005 ( .A(n19320), .B(n19319), .Z(n1110) );
  XOR U2006 ( .A(n19320), .B(n19319), .Z(n1111) );
  NAND U2007 ( .A(n19318), .B(n1111), .Z(n1112) );
  AND U2008 ( .A(n1110), .B(n1112), .Z(n1113) );
  XNOR U2009 ( .A(n1109), .B(n1113), .Z(n1114) );
  XNOR U2010 ( .A(n1103), .B(n1106), .Z(n1115) );
  XNOR U2011 ( .A(n1114), .B(n1115), .Z(n1116) );
  XNOR U2012 ( .A(n1100), .B(n1116), .Z(o[199]) );
  NAND U2013 ( .A(y[160]), .B(x[32]), .Z(n1230) );
  NAND U2014 ( .A(x[8]), .B(y[40]), .Z(n1119) );
  XOR U2015 ( .A(n1230), .B(n1119), .Z(n1120) );
  AND U2016 ( .A(y[0]), .B(x[0]), .Z(n1127) );
  AND U2017 ( .A(y[80]), .B(x[16]), .Z(n1124) );
  XOR U2018 ( .A(n1127), .B(n1124), .Z(n1123) );
  AND U2019 ( .A(y[120]), .B(x[24]), .Z(n1122) );
  XNOR U2020 ( .A(n1123), .B(n1122), .Z(n1121) );
  XNOR U2021 ( .A(n1120), .B(n1121), .Z(o[0]) );
  AND U2022 ( .A(x[0]), .B(y[1]), .Z(n1118) );
  NAND U2023 ( .A(x[1]), .B(y[0]), .Z(n1117) );
  XNOR U2024 ( .A(n1118), .B(n1117), .Z(n1129) );
  AND U2025 ( .A(x[9]), .B(y[40]), .Z(n1128) );
  XOR U2026 ( .A(n1129), .B(n1128), .Z(n1146) );
  AND U2027 ( .A(y[160]), .B(x[33]), .Z(n1350) );
  AND U2028 ( .A(x[16]), .B(y[81]), .Z(n1132) );
  XOR U2029 ( .A(n1350), .B(n1132), .Z(n1134) );
  AND U2030 ( .A(y[161]), .B(x[32]), .Z(n1156) );
  NAND U2031 ( .A(y[80]), .B(x[17]), .Z(n1155) );
  XNOR U2032 ( .A(n1156), .B(n1155), .Z(n1133) );
  XOR U2033 ( .A(n1134), .B(n1133), .Z(n1144) );
  AND U2034 ( .A(y[41]), .B(x[8]), .Z(n1380) );
  AND U2035 ( .A(y[121]), .B(x[24]), .Z(n1149) );
  XOR U2036 ( .A(n1380), .B(n1149), .Z(n1151) );
  AND U2037 ( .A(y[120]), .B(x[25]), .Z(n1150) );
  XNOR U2038 ( .A(n1151), .B(n1150), .Z(n1143) );
  XNOR U2039 ( .A(n1144), .B(n1143), .Z(n1145) );
  XNOR U2040 ( .A(n1146), .B(n1145), .Z(n1140) );
  NAND U2041 ( .A(n1123), .B(n1122), .Z(n1126) );
  AND U2042 ( .A(n1127), .B(n1124), .Z(n1125) );
  ANDN U2043 ( .B(n1126), .A(n1125), .Z(n1137) );
  XNOR U2044 ( .A(n1138), .B(n1137), .Z(n1139) );
  XNOR U2045 ( .A(n1140), .B(n1139), .Z(o[1]) );
  NAND U2046 ( .A(y[1]), .B(x[1]), .Z(n1178) );
  NANDN U2047 ( .A(n1178), .B(n1127), .Z(n1131) );
  NAND U2048 ( .A(n1129), .B(n1128), .Z(n1130) );
  AND U2049 ( .A(n1131), .B(n1130), .Z(n1198) );
  NAND U2050 ( .A(n1350), .B(n1132), .Z(n1136) );
  NAND U2051 ( .A(n1134), .B(n1133), .Z(n1135) );
  AND U2052 ( .A(n1136), .B(n1135), .Z(n1197) );
  AND U2053 ( .A(y[122]), .B(x[24]), .Z(n1202) );
  NAND U2054 ( .A(y[2]), .B(x[0]), .Z(n1203) );
  XNOR U2055 ( .A(n1202), .B(n1203), .Z(n1204) );
  NAND U2056 ( .A(x[10]), .B(y[40]), .Z(n1205) );
  XNOR U2057 ( .A(n1204), .B(n1205), .Z(n1196) );
  XOR U2058 ( .A(n1197), .B(n1196), .Z(n1199) );
  XOR U2059 ( .A(n1198), .B(n1199), .Z(n1158) );
  NANDN U2060 ( .A(n1138), .B(n1137), .Z(n1142) );
  NAND U2061 ( .A(n1140), .B(n1139), .Z(n1141) );
  NAND U2062 ( .A(n1142), .B(n1141), .Z(n1157) );
  XNOR U2063 ( .A(n1158), .B(n1157), .Z(n1160) );
  NANDN U2064 ( .A(n1144), .B(n1143), .Z(n1148) );
  NANDN U2065 ( .A(n1146), .B(n1145), .Z(n1147) );
  AND U2066 ( .A(n1148), .B(n1147), .Z(n1166) );
  AND U2067 ( .A(y[0]), .B(x[2]), .Z(n1175) );
  NAND U2068 ( .A(x[16]), .B(y[82]), .Z(n1176) );
  XNOR U2069 ( .A(n1175), .B(n1176), .Z(n1177) );
  AND U2070 ( .A(x[26]), .B(y[120]), .Z(n1210) );
  XOR U2071 ( .A(n1211), .B(n1210), .Z(n1213) );
  AND U2072 ( .A(y[80]), .B(x[18]), .Z(n1260) );
  AND U2073 ( .A(y[162]), .B(x[32]), .Z(n1188) );
  XOR U2074 ( .A(n1260), .B(n1188), .Z(n1190) );
  AND U2075 ( .A(y[81]), .B(x[17]), .Z(n1189) );
  XOR U2076 ( .A(n1190), .B(n1189), .Z(n1212) );
  XOR U2077 ( .A(n1213), .B(n1212), .Z(n1163) );
  NAND U2078 ( .A(n1380), .B(n1149), .Z(n1153) );
  AND U2079 ( .A(n1151), .B(n1150), .Z(n1152) );
  ANDN U2080 ( .B(n1153), .A(n1152), .Z(n1172) );
  AND U2081 ( .A(y[161]), .B(x[33]), .Z(n1235) );
  NAND U2082 ( .A(x[34]), .B(y[160]), .Z(n1154) );
  XNOR U2083 ( .A(n1235), .B(n1154), .Z(n1209) );
  ANDN U2084 ( .B(n1156), .A(n1155), .Z(n1208) );
  XOR U2085 ( .A(n1209), .B(n1208), .Z(n1169) );
  AND U2086 ( .A(y[121]), .B(x[25]), .Z(n1181) );
  NAND U2087 ( .A(x[9]), .B(y[41]), .Z(n1182) );
  XNOR U2088 ( .A(n1181), .B(n1182), .Z(n1183) );
  NAND U2089 ( .A(y[42]), .B(x[8]), .Z(n1184) );
  XOR U2090 ( .A(n1183), .B(n1184), .Z(n1170) );
  XNOR U2091 ( .A(n1169), .B(n1170), .Z(n1171) );
  XOR U2092 ( .A(n1172), .B(n1171), .Z(n1164) );
  XNOR U2093 ( .A(n1163), .B(n1164), .Z(n1165) );
  XNOR U2094 ( .A(n1166), .B(n1165), .Z(n1159) );
  XNOR U2095 ( .A(n1160), .B(n1159), .Z(o[2]) );
  NANDN U2096 ( .A(n1158), .B(n1157), .Z(n1162) );
  NAND U2097 ( .A(n1160), .B(n1159), .Z(n1161) );
  AND U2098 ( .A(n1162), .B(n1161), .Z(n1302) );
  NANDN U2099 ( .A(n1164), .B(n1163), .Z(n1168) );
  NAND U2100 ( .A(n1166), .B(n1165), .Z(n1167) );
  AND U2101 ( .A(n1168), .B(n1167), .Z(n1287) );
  NANDN U2102 ( .A(n1170), .B(n1169), .Z(n1174) );
  NANDN U2103 ( .A(n1172), .B(n1171), .Z(n1173) );
  AND U2104 ( .A(n1174), .B(n1173), .Z(n1285) );
  NANDN U2105 ( .A(n1176), .B(n1175), .Z(n1180) );
  NANDN U2106 ( .A(n1178), .B(n1177), .Z(n1179) );
  NAND U2107 ( .A(n1180), .B(n1179), .Z(n1296) );
  NANDN U2108 ( .A(n1182), .B(n1181), .Z(n1186) );
  NANDN U2109 ( .A(n1184), .B(n1183), .Z(n1185) );
  AND U2110 ( .A(n1186), .B(n1185), .Z(n1251) );
  AND U2111 ( .A(y[123]), .B(x[24]), .Z(n1280) );
  AND U2112 ( .A(x[16]), .B(y[83]), .Z(n1279) );
  NAND U2113 ( .A(y[0]), .B(x[3]), .Z(n1278) );
  XOR U2114 ( .A(n1279), .B(n1278), .Z(n1281) );
  XOR U2115 ( .A(n1280), .B(n1281), .Z(n1249) );
  AND U2116 ( .A(x[18]), .B(y[81]), .Z(n1336) );
  NAND U2117 ( .A(x[19]), .B(y[80]), .Z(n1187) );
  XNOR U2118 ( .A(n1336), .B(n1187), .Z(n1262) );
  NAND U2119 ( .A(y[82]), .B(x[17]), .Z(n1263) );
  XNOR U2120 ( .A(n1262), .B(n1263), .Z(n1248) );
  XNOR U2121 ( .A(n1249), .B(n1248), .Z(n1250) );
  XNOR U2122 ( .A(n1251), .B(n1250), .Z(n1297) );
  XOR U2123 ( .A(n1296), .B(n1297), .Z(n1299) );
  NAND U2124 ( .A(n1260), .B(n1188), .Z(n1192) );
  AND U2125 ( .A(n1190), .B(n1189), .Z(n1191) );
  ANDN U2126 ( .B(n1192), .A(n1191), .Z(n1256) );
  AND U2127 ( .A(y[2]), .B(x[1]), .Z(n1226) );
  AND U2128 ( .A(x[2]), .B(y[1]), .Z(n1225) );
  NAND U2129 ( .A(y[122]), .B(x[25]), .Z(n1224) );
  XOR U2130 ( .A(n1225), .B(n1224), .Z(n1227) );
  XOR U2131 ( .A(n1226), .B(n1227), .Z(n1255) );
  AND U2132 ( .A(x[35]), .B(y[160]), .Z(n1194) );
  NAND U2133 ( .A(x[32]), .B(y[163]), .Z(n1193) );
  XNOR U2134 ( .A(n1194), .B(n1193), .Z(n1231) );
  AND U2135 ( .A(x[34]), .B(y[161]), .Z(n1347) );
  NAND U2136 ( .A(y[162]), .B(x[33]), .Z(n1195) );
  XOR U2137 ( .A(n1347), .B(n1195), .Z(n1232) );
  XNOR U2138 ( .A(n1231), .B(n1232), .Z(n1254) );
  XOR U2139 ( .A(n1255), .B(n1254), .Z(n1257) );
  XOR U2140 ( .A(n1256), .B(n1257), .Z(n1298) );
  XOR U2141 ( .A(n1299), .B(n1298), .Z(n1284) );
  XNOR U2142 ( .A(n1285), .B(n1284), .Z(n1286) );
  XOR U2143 ( .A(n1287), .B(n1286), .Z(n1303) );
  XNOR U2144 ( .A(n1302), .B(n1303), .Z(n1305) );
  NANDN U2145 ( .A(n1197), .B(n1196), .Z(n1201) );
  OR U2146 ( .A(n1199), .B(n1198), .Z(n1200) );
  AND U2147 ( .A(n1201), .B(n1200), .Z(n1293) );
  NANDN U2148 ( .A(n1203), .B(n1202), .Z(n1207) );
  NANDN U2149 ( .A(n1205), .B(n1204), .Z(n1206) );
  AND U2150 ( .A(n1207), .B(n1206), .Z(n1217) );
  XNOR U2151 ( .A(n1217), .B(n1216), .Z(n1219) );
  AND U2152 ( .A(x[11]), .B(y[40]), .Z(n1270) );
  AND U2153 ( .A(y[3]), .B(x[0]), .Z(n1269) );
  NAND U2154 ( .A(x[26]), .B(y[121]), .Z(n1268) );
  XOR U2155 ( .A(n1269), .B(n1268), .Z(n1271) );
  XOR U2156 ( .A(n1270), .B(n1271), .Z(n1245) );
  AND U2157 ( .A(y[43]), .B(x[8]), .Z(n1238) );
  AND U2158 ( .A(x[10]), .B(y[41]), .Z(n1237) );
  NAND U2159 ( .A(y[120]), .B(x[27]), .Z(n1236) );
  XOR U2160 ( .A(n1237), .B(n1236), .Z(n1239) );
  XOR U2161 ( .A(n1238), .B(n1239), .Z(n1243) );
  AND U2162 ( .A(y[42]), .B(x[9]), .Z(n1242) );
  XNOR U2163 ( .A(n1243), .B(n1242), .Z(n1244) );
  XNOR U2164 ( .A(n1245), .B(n1244), .Z(n1218) );
  XOR U2165 ( .A(n1219), .B(n1218), .Z(n1291) );
  NAND U2166 ( .A(n1211), .B(n1210), .Z(n1215) );
  NAND U2167 ( .A(n1213), .B(n1212), .Z(n1214) );
  AND U2168 ( .A(n1215), .B(n1214), .Z(n1290) );
  XNOR U2169 ( .A(n1291), .B(n1290), .Z(n1292) );
  XNOR U2170 ( .A(n1293), .B(n1292), .Z(n1304) );
  XOR U2171 ( .A(n1305), .B(n1304), .Z(o[3]) );
  NANDN U2172 ( .A(n1217), .B(n1216), .Z(n1221) );
  NAND U2173 ( .A(n1219), .B(n1218), .Z(n1220) );
  AND U2174 ( .A(n1221), .B(n1220), .Z(n1319) );
  AND U2175 ( .A(y[42]), .B(x[10]), .Z(n1446) );
  AND U2176 ( .A(x[8]), .B(y[44]), .Z(n1223) );
  AND U2177 ( .A(y[41]), .B(x[11]), .Z(n1222) );
  XOR U2178 ( .A(n1223), .B(n1222), .Z(n1381) );
  XOR U2179 ( .A(n1446), .B(n1381), .Z(n1382) );
  NAND U2180 ( .A(y[43]), .B(x[9]), .Z(n1383) );
  XNOR U2181 ( .A(n1382), .B(n1383), .Z(n1385) );
  AND U2182 ( .A(y[120]), .B(x[28]), .Z(n1340) );
  AND U2183 ( .A(y[3]), .B(x[1]), .Z(n1339) );
  XOR U2184 ( .A(n1340), .B(n1339), .Z(n1342) );
  AND U2185 ( .A(x[0]), .B(y[4]), .Z(n1341) );
  XOR U2186 ( .A(n1342), .B(n1341), .Z(n1384) );
  XOR U2187 ( .A(n1385), .B(n1384), .Z(n1395) );
  NANDN U2188 ( .A(n1225), .B(n1224), .Z(n1229) );
  OR U2189 ( .A(n1227), .B(n1226), .Z(n1228) );
  AND U2190 ( .A(n1229), .B(n1228), .Z(n1393) );
  AND U2191 ( .A(y[163]), .B(x[35]), .Z(n1632) );
  NANDN U2192 ( .A(n1230), .B(n1632), .Z(n1234) );
  NANDN U2193 ( .A(n1232), .B(n1231), .Z(n1233) );
  AND U2194 ( .A(n1234), .B(n1233), .Z(n1392) );
  XNOR U2195 ( .A(n1393), .B(n1392), .Z(n1394) );
  XNOR U2196 ( .A(n1395), .B(n1394), .Z(n1413) );
  AND U2197 ( .A(y[0]), .B(x[4]), .Z(n1363) );
  AND U2198 ( .A(y[122]), .B(x[26]), .Z(n1362) );
  NAND U2199 ( .A(y[84]), .B(x[16]), .Z(n1361) );
  XOR U2200 ( .A(n1362), .B(n1361), .Z(n1364) );
  XOR U2201 ( .A(n1363), .B(n1364), .Z(n1325) );
  AND U2202 ( .A(x[34]), .B(y[162]), .Z(n1277) );
  AND U2203 ( .A(n1277), .B(n1235), .Z(n1358) );
  AND U2204 ( .A(y[164]), .B(x[32]), .Z(n1356) );
  IV U2205 ( .A(n1356), .Z(n1503) );
  AND U2206 ( .A(y[80]), .B(x[20]), .Z(n1355) );
  XNOR U2207 ( .A(n1503), .B(n1355), .Z(n1357) );
  XOR U2208 ( .A(n1358), .B(n1357), .Z(n1324) );
  XNOR U2209 ( .A(n1325), .B(n1324), .Z(n1327) );
  NANDN U2210 ( .A(n1237), .B(n1236), .Z(n1241) );
  OR U2211 ( .A(n1239), .B(n1238), .Z(n1240) );
  AND U2212 ( .A(n1241), .B(n1240), .Z(n1326) );
  XOR U2213 ( .A(n1327), .B(n1326), .Z(n1411) );
  NANDN U2214 ( .A(n1243), .B(n1242), .Z(n1247) );
  NANDN U2215 ( .A(n1245), .B(n1244), .Z(n1246) );
  AND U2216 ( .A(n1247), .B(n1246), .Z(n1410) );
  XNOR U2217 ( .A(n1411), .B(n1410), .Z(n1412) );
  XNOR U2218 ( .A(n1413), .B(n1412), .Z(n1318) );
  XNOR U2219 ( .A(n1319), .B(n1318), .Z(n1321) );
  NANDN U2220 ( .A(n1249), .B(n1248), .Z(n1253) );
  NANDN U2221 ( .A(n1251), .B(n1250), .Z(n1252) );
  AND U2222 ( .A(n1253), .B(n1252), .Z(n1399) );
  NANDN U2223 ( .A(n1255), .B(n1254), .Z(n1259) );
  OR U2224 ( .A(n1257), .B(n1256), .Z(n1258) );
  NAND U2225 ( .A(n1259), .B(n1258), .Z(n1398) );
  XNOR U2226 ( .A(n1399), .B(n1398), .Z(n1400) );
  AND U2227 ( .A(y[81]), .B(x[19]), .Z(n1261) );
  NAND U2228 ( .A(n1261), .B(n1260), .Z(n1265) );
  NANDN U2229 ( .A(n1263), .B(n1262), .Z(n1264) );
  AND U2230 ( .A(n1265), .B(n1264), .Z(n1405) );
  AND U2231 ( .A(y[40]), .B(x[12]), .Z(n1344) );
  AND U2232 ( .A(y[124]), .B(x[24]), .Z(n1343) );
  XOR U2233 ( .A(n1344), .B(n1343), .Z(n1346) );
  AND U2234 ( .A(x[25]), .B(y[123]), .Z(n1345) );
  XOR U2235 ( .A(n1346), .B(n1345), .Z(n1389) );
  AND U2236 ( .A(x[18]), .B(y[82]), .Z(n1267) );
  NAND U2237 ( .A(x[19]), .B(y[81]), .Z(n1266) );
  XNOR U2238 ( .A(n1267), .B(n1266), .Z(n1338) );
  AND U2239 ( .A(x[17]), .B(y[83]), .Z(n1337) );
  XOR U2240 ( .A(n1338), .B(n1337), .Z(n1388) );
  XOR U2241 ( .A(n1389), .B(n1388), .Z(n1390) );
  NANDN U2242 ( .A(n1269), .B(n1268), .Z(n1273) );
  OR U2243 ( .A(n1271), .B(n1270), .Z(n1272) );
  NAND U2244 ( .A(n1273), .B(n1272), .Z(n1391) );
  XNOR U2245 ( .A(n1390), .B(n1391), .Z(n1404) );
  XNOR U2246 ( .A(n1405), .B(n1404), .Z(n1406) );
  AND U2247 ( .A(y[2]), .B(x[2]), .Z(n1377) );
  AND U2248 ( .A(y[121]), .B(x[27]), .Z(n1375) );
  NAND U2249 ( .A(x[3]), .B(y[1]), .Z(n1374) );
  AND U2250 ( .A(y[160]), .B(x[36]), .Z(n1275) );
  NAND U2251 ( .A(x[33]), .B(y[163]), .Z(n1274) );
  XNOR U2252 ( .A(n1275), .B(n1274), .Z(n1351) );
  NAND U2253 ( .A(x[35]), .B(y[161]), .Z(n1276) );
  XOR U2254 ( .A(n1277), .B(n1276), .Z(n1352) );
  XNOR U2255 ( .A(n1351), .B(n1352), .Z(n1330) );
  XOR U2256 ( .A(n1331), .B(n1330), .Z(n1332) );
  NANDN U2257 ( .A(n1279), .B(n1278), .Z(n1283) );
  OR U2258 ( .A(n1281), .B(n1280), .Z(n1282) );
  NAND U2259 ( .A(n1283), .B(n1282), .Z(n1333) );
  XOR U2260 ( .A(n1332), .B(n1333), .Z(n1407) );
  XOR U2261 ( .A(n1406), .B(n1407), .Z(n1401) );
  XNOR U2262 ( .A(n1400), .B(n1401), .Z(n1320) );
  XNOR U2263 ( .A(n1321), .B(n1320), .Z(n1311) );
  NANDN U2264 ( .A(n1285), .B(n1284), .Z(n1289) );
  NANDN U2265 ( .A(n1287), .B(n1286), .Z(n1288) );
  AND U2266 ( .A(n1289), .B(n1288), .Z(n1314) );
  NANDN U2267 ( .A(n1291), .B(n1290), .Z(n1295) );
  NAND U2268 ( .A(n1293), .B(n1292), .Z(n1294) );
  NAND U2269 ( .A(n1295), .B(n1294), .Z(n1312) );
  NAND U2270 ( .A(n1297), .B(n1296), .Z(n1301) );
  NAND U2271 ( .A(n1299), .B(n1298), .Z(n1300) );
  AND U2272 ( .A(n1301), .B(n1300), .Z(n1313) );
  XNOR U2273 ( .A(n1312), .B(n1313), .Z(n1315) );
  NANDN U2274 ( .A(n1303), .B(n1302), .Z(n1307) );
  NAND U2275 ( .A(n1305), .B(n1304), .Z(n1306) );
  NAND U2276 ( .A(n1307), .B(n1306), .Z(n1309) );
  XNOR U2277 ( .A(n1310), .B(n1309), .Z(n1308) );
  XNOR U2278 ( .A(n1311), .B(n1308), .Z(o[4]) );
  NAND U2279 ( .A(n1313), .B(n1312), .Z(n1317) );
  NANDN U2280 ( .A(n1315), .B(n1314), .Z(n1316) );
  AND U2281 ( .A(n1317), .B(n1316), .Z(n1416) );
  XNOR U2282 ( .A(n1417), .B(n1416), .Z(n1419) );
  NANDN U2283 ( .A(n1319), .B(n1318), .Z(n1323) );
  NAND U2284 ( .A(n1321), .B(n1320), .Z(n1322) );
  AND U2285 ( .A(n1323), .B(n1322), .Z(n1525) );
  NANDN U2286 ( .A(n1325), .B(n1324), .Z(n1329) );
  NAND U2287 ( .A(n1327), .B(n1326), .Z(n1328) );
  NAND U2288 ( .A(n1329), .B(n1328), .Z(n1468) );
  NAND U2289 ( .A(n1331), .B(n1330), .Z(n1335) );
  NANDN U2290 ( .A(n1333), .B(n1332), .Z(n1334) );
  NAND U2291 ( .A(n1335), .B(n1334), .Z(n1469) );
  XOR U2292 ( .A(n1468), .B(n1469), .Z(n1471) );
  AND U2293 ( .A(y[82]), .B(x[19]), .Z(n1373) );
  IV U2294 ( .A(n1373), .Z(n1461) );
  AND U2295 ( .A(x[24]), .B(y[125]), .Z(n1685) );
  AND U2296 ( .A(y[40]), .B(x[13]), .Z(n1454) );
  AND U2297 ( .A(x[18]), .B(y[83]), .Z(n1453) );
  XOR U2298 ( .A(n1454), .B(n1453), .Z(n1455) );
  XOR U2299 ( .A(n1685), .B(n1455), .Z(n1450) );
  AND U2300 ( .A(y[121]), .B(x[28]), .Z(n1457) );
  AND U2301 ( .A(y[0]), .B(x[5]), .Z(n1456) );
  XOR U2302 ( .A(n1457), .B(n1456), .Z(n1458) );
  AND U2303 ( .A(x[4]), .B(y[1]), .Z(n1723) );
  XOR U2304 ( .A(n1458), .B(n1723), .Z(n1449) );
  XOR U2305 ( .A(n1450), .B(n1449), .Z(n1452) );
  XOR U2306 ( .A(n1451), .B(n1452), .Z(n1433) );
  XOR U2307 ( .A(n1432), .B(n1433), .Z(n1435) );
  AND U2308 ( .A(y[162]), .B(x[35]), .Z(n1370) );
  AND U2309 ( .A(n1347), .B(n1370), .Z(n1505) );
  AND U2310 ( .A(y[165]), .B(x[32]), .Z(n1349) );
  AND U2311 ( .A(y[164]), .B(x[33]), .Z(n1348) );
  XOR U2312 ( .A(n1349), .B(n1348), .Z(n1504) );
  XOR U2313 ( .A(n1505), .B(n1504), .Z(n1507) );
  AND U2314 ( .A(x[8]), .B(y[45]), .Z(n1513) );
  AND U2315 ( .A(x[1]), .B(y[4]), .Z(n1512) );
  XOR U2316 ( .A(n1513), .B(n1512), .Z(n1515) );
  AND U2317 ( .A(y[41]), .B(x[12]), .Z(n1514) );
  XOR U2318 ( .A(n1515), .B(n1514), .Z(n1506) );
  XOR U2319 ( .A(n1507), .B(n1506), .Z(n1509) );
  XOR U2320 ( .A(n1508), .B(n1509), .Z(n1434) );
  XOR U2321 ( .A(n1435), .B(n1434), .Z(n1470) );
  XOR U2322 ( .A(n1471), .B(n1470), .Z(n1425) );
  AND U2323 ( .A(y[163]), .B(x[36]), .Z(n1681) );
  NAND U2324 ( .A(n1681), .B(n1350), .Z(n1354) );
  NANDN U2325 ( .A(n1352), .B(n1351), .Z(n1353) );
  NAND U2326 ( .A(n1354), .B(n1353), .Z(n1476) );
  IV U2327 ( .A(n1355), .Z(n1459) );
  NANDN U2328 ( .A(n1356), .B(n1459), .Z(n1360) );
  NANDN U2329 ( .A(n1358), .B(n1357), .Z(n1359) );
  AND U2330 ( .A(n1360), .B(n1359), .Z(n1477) );
  XOR U2331 ( .A(n1476), .B(n1477), .Z(n1479) );
  NANDN U2332 ( .A(n1362), .B(n1361), .Z(n1366) );
  OR U2333 ( .A(n1364), .B(n1363), .Z(n1365) );
  AND U2334 ( .A(n1366), .B(n1365), .Z(n1483) );
  AND U2335 ( .A(y[43]), .B(x[10]), .Z(n1368) );
  NAND U2336 ( .A(x[11]), .B(y[42]), .Z(n1367) );
  XNOR U2337 ( .A(n1368), .B(n1367), .Z(n1448) );
  AND U2338 ( .A(y[44]), .B(x[9]), .Z(n1447) );
  XOR U2339 ( .A(n1448), .B(n1447), .Z(n1481) );
  AND U2340 ( .A(y[163]), .B(x[34]), .Z(n1439) );
  AND U2341 ( .A(y[160]), .B(x[37]), .Z(n1438) );
  XOR U2342 ( .A(n1439), .B(n1438), .Z(n1441) );
  NAND U2343 ( .A(y[161]), .B(x[36]), .Z(n1369) );
  XNOR U2344 ( .A(n1370), .B(n1369), .Z(n1440) );
  XOR U2345 ( .A(n1441), .B(n1440), .Z(n1480) );
  XOR U2346 ( .A(n1481), .B(n1480), .Z(n1482) );
  XOR U2347 ( .A(n1483), .B(n1482), .Z(n1478) );
  XOR U2348 ( .A(n1479), .B(n1478), .Z(n1491) );
  AND U2349 ( .A(y[81]), .B(x[20]), .Z(n1372) );
  NAND U2350 ( .A(x[21]), .B(y[80]), .Z(n1371) );
  XNOR U2351 ( .A(n1372), .B(n1371), .Z(n1460) );
  XOR U2352 ( .A(n1460), .B(n1373), .Z(n1521) );
  AND U2353 ( .A(y[120]), .B(x[29]), .Z(n1443) );
  AND U2354 ( .A(y[2]), .B(x[3]), .Z(n1442) );
  XOR U2355 ( .A(n1443), .B(n1442), .Z(n1445) );
  AND U2356 ( .A(y[3]), .B(x[2]), .Z(n1444) );
  XOR U2357 ( .A(n1445), .B(n1444), .Z(n1520) );
  XOR U2358 ( .A(n1521), .B(n1520), .Z(n1523) );
  NANDN U2359 ( .A(n1375), .B(n1374), .Z(n1379) );
  NANDN U2360 ( .A(n1377), .B(n1376), .Z(n1378) );
  AND U2361 ( .A(n1379), .B(n1378), .Z(n1522) );
  XOR U2362 ( .A(n1523), .B(n1522), .Z(n1489) );
  AND U2363 ( .A(x[11]), .B(y[44]), .Z(n1680) );
  AND U2364 ( .A(y[84]), .B(x[17]), .Z(n1701) );
  AND U2365 ( .A(y[122]), .B(x[27]), .Z(n1496) );
  XOR U2366 ( .A(n1701), .B(n1496), .Z(n1495) );
  AND U2367 ( .A(x[16]), .B(y[85]), .Z(n1494) );
  XOR U2368 ( .A(n1495), .B(n1494), .Z(n1473) );
  AND U2369 ( .A(y[5]), .B(x[0]), .Z(n1498) );
  AND U2370 ( .A(y[124]), .B(x[25]), .Z(n1497) );
  XOR U2371 ( .A(n1498), .B(n1497), .Z(n1500) );
  AND U2372 ( .A(x[26]), .B(y[123]), .Z(n1499) );
  XOR U2373 ( .A(n1500), .B(n1499), .Z(n1472) );
  XOR U2374 ( .A(n1473), .B(n1472), .Z(n1475) );
  XOR U2375 ( .A(n1474), .B(n1475), .Z(n1488) );
  XOR U2376 ( .A(n1489), .B(n1488), .Z(n1490) );
  XOR U2377 ( .A(n1491), .B(n1490), .Z(n1422) );
  NANDN U2378 ( .A(n1383), .B(n1382), .Z(n1387) );
  NAND U2379 ( .A(n1385), .B(n1384), .Z(n1386) );
  NAND U2380 ( .A(n1387), .B(n1386), .Z(n1484) );
  XOR U2381 ( .A(n1484), .B(n1485), .Z(n1487) );
  NANDN U2382 ( .A(n1393), .B(n1392), .Z(n1397) );
  NANDN U2383 ( .A(n1395), .B(n1394), .Z(n1396) );
  AND U2384 ( .A(n1397), .B(n1396), .Z(n1486) );
  XOR U2385 ( .A(n1487), .B(n1486), .Z(n1423) );
  XOR U2386 ( .A(n1422), .B(n1423), .Z(n1424) );
  XOR U2387 ( .A(n1425), .B(n1424), .Z(n1524) );
  XNOR U2388 ( .A(n1525), .B(n1524), .Z(n1526) );
  NANDN U2389 ( .A(n1399), .B(n1398), .Z(n1403) );
  NANDN U2390 ( .A(n1401), .B(n1400), .Z(n1402) );
  AND U2391 ( .A(n1403), .B(n1402), .Z(n1429) );
  NANDN U2392 ( .A(n1405), .B(n1404), .Z(n1409) );
  NANDN U2393 ( .A(n1407), .B(n1406), .Z(n1408) );
  AND U2394 ( .A(n1409), .B(n1408), .Z(n1427) );
  NANDN U2395 ( .A(n1411), .B(n1410), .Z(n1415) );
  NAND U2396 ( .A(n1413), .B(n1412), .Z(n1414) );
  AND U2397 ( .A(n1415), .B(n1414), .Z(n1426) );
  XNOR U2398 ( .A(n1427), .B(n1426), .Z(n1428) );
  XOR U2399 ( .A(n1429), .B(n1428), .Z(n1527) );
  XNOR U2400 ( .A(n1526), .B(n1527), .Z(n1418) );
  XOR U2401 ( .A(n1419), .B(n1418), .Z(o[5]) );
  NANDN U2402 ( .A(n1417), .B(n1416), .Z(n1421) );
  NAND U2403 ( .A(n1419), .B(n1418), .Z(n1420) );
  AND U2404 ( .A(n1421), .B(n1420), .Z(n1814) );
  NANDN U2405 ( .A(n1427), .B(n1426), .Z(n1431) );
  NANDN U2406 ( .A(n1429), .B(n1428), .Z(n1430) );
  NAND U2407 ( .A(n1431), .B(n1430), .Z(n1826) );
  XNOR U2408 ( .A(n1825), .B(n1826), .Z(n1823) );
  NAND U2409 ( .A(n1433), .B(n1432), .Z(n1437) );
  NAND U2410 ( .A(n1435), .B(n1434), .Z(n1436) );
  AND U2411 ( .A(n1437), .B(n1436), .Z(n1810) );
  AND U2412 ( .A(x[11]), .B(y[43]), .Z(n1511) );
  AND U2413 ( .A(x[27]), .B(y[123]), .Z(n1620) );
  NAND U2414 ( .A(x[19]), .B(y[83]), .Z(n1621) );
  XNOR U2415 ( .A(n1620), .B(n1621), .Z(n1618) );
  NAND U2416 ( .A(x[3]), .B(y[3]), .Z(n1619) );
  XNOR U2417 ( .A(n1618), .B(n1619), .Z(n1743) );
  AND U2418 ( .A(x[26]), .B(y[124]), .Z(n1732) );
  NAND U2419 ( .A(x[20]), .B(y[82]), .Z(n1733) );
  XNOR U2420 ( .A(n1732), .B(n1733), .Z(n1730) );
  AND U2421 ( .A(x[2]), .B(y[4]), .Z(n1731) );
  XNOR U2422 ( .A(n1730), .B(n1731), .Z(n1742) );
  XNOR U2423 ( .A(n1743), .B(n1742), .Z(n1740) );
  XNOR U2424 ( .A(n1741), .B(n1740), .Z(n1752) );
  XNOR U2425 ( .A(n1753), .B(n1752), .Z(n1754) );
  XNOR U2426 ( .A(n1755), .B(n1754), .Z(n1533) );
  XNOR U2427 ( .A(n1533), .B(n1534), .Z(n1531) );
  XOR U2428 ( .A(n1759), .B(n1758), .Z(n1761) );
  AND U2429 ( .A(y[81]), .B(x[21]), .Z(n1717) );
  NANDN U2430 ( .A(n1459), .B(n1717), .Z(n1463) );
  NANDN U2431 ( .A(n1461), .B(n1460), .Z(n1462) );
  AND U2432 ( .A(n1463), .B(n1462), .Z(n1661) );
  AND U2433 ( .A(x[5]), .B(y[1]), .Z(n1465) );
  NAND U2434 ( .A(y[2]), .B(x[4]), .Z(n1464) );
  XNOR U2435 ( .A(n1465), .B(n1464), .Z(n1724) );
  NAND U2436 ( .A(y[120]), .B(x[30]), .Z(n1725) );
  XNOR U2437 ( .A(n1724), .B(n1725), .Z(n1663) );
  AND U2438 ( .A(x[33]), .B(y[165]), .Z(n1596) );
  AND U2439 ( .A(y[161]), .B(x[35]), .Z(n1467) );
  AND U2440 ( .A(x[36]), .B(y[162]), .Z(n1466) );
  AND U2441 ( .A(n1467), .B(n1466), .Z(n1598) );
  NAND U2442 ( .A(x[34]), .B(y[164]), .Z(n1599) );
  XNOR U2443 ( .A(n1598), .B(n1599), .Z(n1597) );
  XNOR U2444 ( .A(n1596), .B(n1597), .Z(n1662) );
  XNOR U2445 ( .A(n1663), .B(n1662), .Z(n1660) );
  XNOR U2446 ( .A(n1661), .B(n1660), .Z(n1760) );
  XNOR U2447 ( .A(n1761), .B(n1760), .Z(n1532) );
  XNOR U2448 ( .A(n1531), .B(n1532), .Z(n1795) );
  XNOR U2449 ( .A(n1795), .B(n1794), .Z(n1792) );
  XNOR U2450 ( .A(n1545), .B(n1546), .Z(n1543) );
  XNOR U2451 ( .A(n1543), .B(n1544), .Z(n1793) );
  XNOR U2452 ( .A(n1792), .B(n1793), .Z(n1811) );
  XNOR U2453 ( .A(n1810), .B(n1811), .Z(n1808) );
  OR U2454 ( .A(n1489), .B(n1488), .Z(n1493) );
  NANDN U2455 ( .A(n1491), .B(n1490), .Z(n1492) );
  AND U2456 ( .A(n1493), .B(n1492), .Z(n1798) );
  AND U2457 ( .A(y[5]), .B(x[1]), .Z(n1696) );
  NAND U2458 ( .A(y[40]), .B(x[14]), .Z(n1697) );
  XNOR U2459 ( .A(n1696), .B(n1697), .Z(n1694) );
  NAND U2460 ( .A(x[8]), .B(y[46]), .Z(n1695) );
  XNOR U2461 ( .A(n1694), .B(n1695), .Z(n1777) );
  AND U2462 ( .A(x[37]), .B(y[161]), .Z(n1502) );
  NAND U2463 ( .A(y[162]), .B(x[36]), .Z(n1501) );
  XNOR U2464 ( .A(n1502), .B(n1501), .Z(n1630) );
  AND U2465 ( .A(y[160]), .B(x[38]), .Z(n1631) );
  XNOR U2466 ( .A(n1630), .B(n1631), .Z(n1633) );
  XNOR U2467 ( .A(n1632), .B(n1633), .Z(n1776) );
  XNOR U2468 ( .A(n1777), .B(n1776), .Z(n1779) );
  XNOR U2469 ( .A(n1778), .B(n1779), .Z(n1538) );
  XNOR U2470 ( .A(n1538), .B(n1537), .Z(n1539) );
  XNOR U2471 ( .A(n1540), .B(n1539), .Z(n1832) );
  AND U2472 ( .A(x[16]), .B(y[86]), .Z(n1592) );
  NAND U2473 ( .A(y[0]), .B(x[6]), .Z(n1593) );
  XNOR U2474 ( .A(n1592), .B(n1593), .Z(n1590) );
  NAND U2475 ( .A(x[29]), .B(y[121]), .Z(n1591) );
  XNOR U2476 ( .A(n1590), .B(n1591), .Z(n1656) );
  AND U2477 ( .A(y[41]), .B(x[13]), .Z(n1668) );
  NAND U2478 ( .A(x[10]), .B(y[44]), .Z(n1669) );
  XNOR U2479 ( .A(n1668), .B(n1669), .Z(n1666) );
  NAND U2480 ( .A(x[9]), .B(y[45]), .Z(n1667) );
  XNOR U2481 ( .A(n1666), .B(n1667), .Z(n1604) );
  NAND U2482 ( .A(x[12]), .B(y[42]), .Z(n1510) );
  XNOR U2483 ( .A(n1511), .B(n1510), .Z(n1605) );
  XNOR U2484 ( .A(n1604), .B(n1605), .Z(n1657) );
  XNOR U2485 ( .A(n1656), .B(n1657), .Z(n1654) );
  AND U2486 ( .A(x[32]), .B(y[166]), .Z(n1716) );
  XOR U2487 ( .A(n1717), .B(n1716), .Z(n1718) );
  AND U2488 ( .A(y[80]), .B(x[22]), .Z(n1719) );
  XNOR U2489 ( .A(n1718), .B(n1719), .Z(n1655) );
  XNOR U2490 ( .A(n1654), .B(n1655), .Z(n1770) );
  AND U2491 ( .A(y[85]), .B(x[17]), .Z(n1517) );
  NAND U2492 ( .A(x[18]), .B(y[84]), .Z(n1516) );
  XNOR U2493 ( .A(n1517), .B(n1516), .Z(n1702) );
  NAND U2494 ( .A(y[122]), .B(x[28]), .Z(n1703) );
  XNOR U2495 ( .A(n1702), .B(n1703), .Z(n1615) );
  AND U2496 ( .A(y[126]), .B(x[24]), .Z(n1519) );
  NAND U2497 ( .A(y[125]), .B(x[25]), .Z(n1518) );
  XNOR U2498 ( .A(n1519), .B(n1518), .Z(n1686) );
  AND U2499 ( .A(x[0]), .B(y[6]), .Z(n1687) );
  XNOR U2500 ( .A(n1686), .B(n1687), .Z(n1614) );
  XNOR U2501 ( .A(n1615), .B(n1614), .Z(n1612) );
  XNOR U2502 ( .A(n1613), .B(n1612), .Z(n1771) );
  XNOR U2503 ( .A(n1770), .B(n1771), .Z(n1773) );
  XNOR U2504 ( .A(n1772), .B(n1773), .Z(n1831) );
  XNOR U2505 ( .A(n1832), .B(n1831), .Z(n1829) );
  XNOR U2506 ( .A(n1829), .B(n1830), .Z(n1799) );
  XNOR U2507 ( .A(n1798), .B(n1799), .Z(n1801) );
  XNOR U2508 ( .A(n1800), .B(n1801), .Z(n1809) );
  XNOR U2509 ( .A(n1808), .B(n1809), .Z(n1824) );
  XNOR U2510 ( .A(n1823), .B(n1824), .Z(n1816) );
  NANDN U2511 ( .A(n1525), .B(n1524), .Z(n1529) );
  NANDN U2512 ( .A(n1527), .B(n1526), .Z(n1528) );
  AND U2513 ( .A(n1529), .B(n1528), .Z(n1815) );
  XNOR U2514 ( .A(n1816), .B(n1815), .Z(n1530) );
  XOR U2515 ( .A(n1814), .B(n1530), .Z(o[6]) );
  NANDN U2516 ( .A(n1532), .B(n1531), .Z(n1536) );
  NANDN U2517 ( .A(n1534), .B(n1533), .Z(n1535) );
  AND U2518 ( .A(n1536), .B(n1535), .Z(n1791) );
  NANDN U2519 ( .A(n1538), .B(n1537), .Z(n1542) );
  NANDN U2520 ( .A(n1540), .B(n1539), .Z(n1541) );
  NAND U2521 ( .A(n1542), .B(n1541), .Z(n1789) );
  NANDN U2522 ( .A(n1544), .B(n1543), .Z(n1548) );
  NANDN U2523 ( .A(n1546), .B(n1545), .Z(n1547) );
  AND U2524 ( .A(n1548), .B(n1547), .Z(n1787) );
  AND U2525 ( .A(y[87]), .B(x[16]), .Z(n1553) );
  AND U2526 ( .A(x[25]), .B(y[126]), .Z(n1684) );
  AND U2527 ( .A(y[7]), .B(x[0]), .Z(n1550) );
  NAND U2528 ( .A(y[124]), .B(x[27]), .Z(n1549) );
  XNOR U2529 ( .A(n1550), .B(n1549), .Z(n1551) );
  XNOR U2530 ( .A(n1684), .B(n1551), .Z(n1552) );
  XNOR U2531 ( .A(n1553), .B(n1552), .Z(n1569) );
  AND U2532 ( .A(y[47]), .B(x[8]), .Z(n1555) );
  NAND U2533 ( .A(x[22]), .B(y[81]), .Z(n1554) );
  XNOR U2534 ( .A(n1555), .B(n1554), .Z(n1559) );
  AND U2535 ( .A(x[6]), .B(y[1]), .Z(n1557) );
  NAND U2536 ( .A(x[7]), .B(y[0]), .Z(n1556) );
  XNOR U2537 ( .A(n1557), .B(n1556), .Z(n1558) );
  XOR U2538 ( .A(n1559), .B(n1558), .Z(n1567) );
  AND U2539 ( .A(x[28]), .B(y[123]), .Z(n1561) );
  NAND U2540 ( .A(x[23]), .B(y[80]), .Z(n1560) );
  XNOR U2541 ( .A(n1561), .B(n1560), .Z(n1565) );
  AND U2542 ( .A(y[167]), .B(x[32]), .Z(n1563) );
  NAND U2543 ( .A(y[166]), .B(x[33]), .Z(n1562) );
  XNOR U2544 ( .A(n1563), .B(n1562), .Z(n1564) );
  XNOR U2545 ( .A(n1565), .B(n1564), .Z(n1566) );
  XNOR U2546 ( .A(n1567), .B(n1566), .Z(n1568) );
  XOR U2547 ( .A(n1569), .B(n1568), .Z(n1589) );
  AND U2548 ( .A(y[86]), .B(x[17]), .Z(n1571) );
  NAND U2549 ( .A(y[3]), .B(x[4]), .Z(n1570) );
  XNOR U2550 ( .A(n1571), .B(n1570), .Z(n1575) );
  AND U2551 ( .A(y[6]), .B(x[1]), .Z(n1573) );
  NAND U2552 ( .A(y[83]), .B(x[20]), .Z(n1572) );
  XNOR U2553 ( .A(n1573), .B(n1572), .Z(n1574) );
  XOR U2554 ( .A(n1575), .B(n1574), .Z(n1583) );
  AND U2555 ( .A(x[14]), .B(y[41]), .Z(n1577) );
  NAND U2556 ( .A(x[39]), .B(y[160]), .Z(n1576) );
  XNOR U2557 ( .A(n1577), .B(n1576), .Z(n1581) );
  AND U2558 ( .A(y[82]), .B(x[21]), .Z(n1579) );
  NAND U2559 ( .A(x[38]), .B(y[161]), .Z(n1578) );
  XNOR U2560 ( .A(n1579), .B(n1578), .Z(n1580) );
  XNOR U2561 ( .A(n1581), .B(n1580), .Z(n1582) );
  XNOR U2562 ( .A(n1583), .B(n1582), .Z(n1587) );
  AND U2563 ( .A(y[43]), .B(x[12]), .Z(n1602) );
  AND U2564 ( .A(y[85]), .B(x[18]), .Z(n1700) );
  XOR U2565 ( .A(n1602), .B(n1700), .Z(n1585) );
  AND U2566 ( .A(y[2]), .B(x[5]), .Z(n1722) );
  AND U2567 ( .A(y[162]), .B(x[37]), .Z(n1674) );
  XNOR U2568 ( .A(n1722), .B(n1674), .Z(n1584) );
  XNOR U2569 ( .A(n1585), .B(n1584), .Z(n1586) );
  XNOR U2570 ( .A(n1587), .B(n1586), .Z(n1588) );
  XNOR U2571 ( .A(n1589), .B(n1588), .Z(n1629) );
  NANDN U2572 ( .A(n1591), .B(n1590), .Z(n1595) );
  NANDN U2573 ( .A(n1593), .B(n1592), .Z(n1594) );
  AND U2574 ( .A(n1595), .B(n1594), .Z(n1611) );
  NAND U2575 ( .A(n1597), .B(n1596), .Z(n1601) );
  NANDN U2576 ( .A(n1599), .B(n1598), .Z(n1600) );
  AND U2577 ( .A(n1601), .B(n1600), .Z(n1609) );
  AND U2578 ( .A(y[42]), .B(x[11]), .Z(n1603) );
  NAND U2579 ( .A(n1603), .B(n1602), .Z(n1607) );
  NAND U2580 ( .A(n1605), .B(n1604), .Z(n1606) );
  NAND U2581 ( .A(n1607), .B(n1606), .Z(n1608) );
  XNOR U2582 ( .A(n1609), .B(n1608), .Z(n1610) );
  XOR U2583 ( .A(n1611), .B(n1610), .Z(n1627) );
  NAND U2584 ( .A(n1613), .B(n1612), .Z(n1617) );
  NANDN U2585 ( .A(n1615), .B(n1614), .Z(n1616) );
  NAND U2586 ( .A(n1617), .B(n1616), .Z(n1625) );
  NANDN U2587 ( .A(n1619), .B(n1618), .Z(n1623) );
  NANDN U2588 ( .A(n1621), .B(n1620), .Z(n1622) );
  AND U2589 ( .A(n1623), .B(n1622), .Z(n1624) );
  XOR U2590 ( .A(n1625), .B(n1624), .Z(n1626) );
  XNOR U2591 ( .A(n1627), .B(n1626), .Z(n1628) );
  XOR U2592 ( .A(n1629), .B(n1628), .Z(n1653) );
  NAND U2593 ( .A(n1631), .B(n1630), .Z(n1635) );
  NANDN U2594 ( .A(n1633), .B(n1632), .Z(n1634) );
  AND U2595 ( .A(n1635), .B(n1634), .Z(n1651) );
  AND U2596 ( .A(y[5]), .B(x[2]), .Z(n1637) );
  NAND U2597 ( .A(y[164]), .B(x[35]), .Z(n1636) );
  XNOR U2598 ( .A(n1637), .B(n1636), .Z(n1641) );
  AND U2599 ( .A(x[30]), .B(y[121]), .Z(n1639) );
  NAND U2600 ( .A(y[4]), .B(x[3]), .Z(n1638) );
  XNOR U2601 ( .A(n1639), .B(n1638), .Z(n1640) );
  XOR U2602 ( .A(n1641), .B(n1640), .Z(n1649) );
  AND U2603 ( .A(x[31]), .B(y[120]), .Z(n1643) );
  NAND U2604 ( .A(x[19]), .B(y[84]), .Z(n1642) );
  XNOR U2605 ( .A(n1643), .B(n1642), .Z(n1647) );
  AND U2606 ( .A(x[29]), .B(y[122]), .Z(n1645) );
  NAND U2607 ( .A(y[165]), .B(x[34]), .Z(n1644) );
  XNOR U2608 ( .A(n1645), .B(n1644), .Z(n1646) );
  XNOR U2609 ( .A(n1647), .B(n1646), .Z(n1648) );
  XNOR U2610 ( .A(n1649), .B(n1648), .Z(n1650) );
  XNOR U2611 ( .A(n1651), .B(n1650), .Z(n1652) );
  XNOR U2612 ( .A(n1653), .B(n1652), .Z(n1769) );
  NANDN U2613 ( .A(n1655), .B(n1654), .Z(n1659) );
  NANDN U2614 ( .A(n1657), .B(n1656), .Z(n1658) );
  AND U2615 ( .A(n1659), .B(n1658), .Z(n1751) );
  NAND U2616 ( .A(n1661), .B(n1660), .Z(n1665) );
  NANDN U2617 ( .A(n1663), .B(n1662), .Z(n1664) );
  NAND U2618 ( .A(n1665), .B(n1664), .Z(n1749) );
  NANDN U2619 ( .A(n1667), .B(n1666), .Z(n1671) );
  NANDN U2620 ( .A(n1669), .B(n1668), .Z(n1670) );
  AND U2621 ( .A(n1671), .B(n1670), .Z(n1715) );
  AND U2622 ( .A(y[127]), .B(x[24]), .Z(n1673) );
  NAND U2623 ( .A(y[46]), .B(x[9]), .Z(n1672) );
  XNOR U2624 ( .A(n1673), .B(n1672), .Z(n1693) );
  AND U2625 ( .A(x[36]), .B(y[161]), .Z(n1675) );
  AND U2626 ( .A(n1675), .B(n1674), .Z(n1679) );
  AND U2627 ( .A(y[45]), .B(x[10]), .Z(n1677) );
  NAND U2628 ( .A(x[13]), .B(y[42]), .Z(n1676) );
  XNOR U2629 ( .A(n1677), .B(n1676), .Z(n1678) );
  XOR U2630 ( .A(n1679), .B(n1678), .Z(n1683) );
  XNOR U2631 ( .A(n1681), .B(n1680), .Z(n1682) );
  XNOR U2632 ( .A(n1683), .B(n1682), .Z(n1691) );
  NAND U2633 ( .A(n1685), .B(n1684), .Z(n1689) );
  NAND U2634 ( .A(n1687), .B(n1686), .Z(n1688) );
  NAND U2635 ( .A(n1689), .B(n1688), .Z(n1690) );
  XNOR U2636 ( .A(n1691), .B(n1690), .Z(n1692) );
  XOR U2637 ( .A(n1693), .B(n1692), .Z(n1713) );
  NANDN U2638 ( .A(n1695), .B(n1694), .Z(n1699) );
  NANDN U2639 ( .A(n1697), .B(n1696), .Z(n1698) );
  AND U2640 ( .A(n1699), .B(n1698), .Z(n1707) );
  NAND U2641 ( .A(n1701), .B(n1700), .Z(n1705) );
  NANDN U2642 ( .A(n1703), .B(n1702), .Z(n1704) );
  NAND U2643 ( .A(n1705), .B(n1704), .Z(n1706) );
  XNOR U2644 ( .A(n1707), .B(n1706), .Z(n1711) );
  AND U2645 ( .A(x[15]), .B(y[40]), .Z(n1709) );
  NAND U2646 ( .A(y[125]), .B(x[26]), .Z(n1708) );
  XNOR U2647 ( .A(n1709), .B(n1708), .Z(n1710) );
  XNOR U2648 ( .A(n1711), .B(n1710), .Z(n1712) );
  XNOR U2649 ( .A(n1713), .B(n1712), .Z(n1714) );
  XOR U2650 ( .A(n1715), .B(n1714), .Z(n1739) );
  NAND U2651 ( .A(n1717), .B(n1716), .Z(n1721) );
  NAND U2652 ( .A(n1719), .B(n1718), .Z(n1720) );
  AND U2653 ( .A(n1721), .B(n1720), .Z(n1729) );
  NAND U2654 ( .A(n1723), .B(n1722), .Z(n1727) );
  NANDN U2655 ( .A(n1725), .B(n1724), .Z(n1726) );
  NAND U2656 ( .A(n1727), .B(n1726), .Z(n1728) );
  XNOR U2657 ( .A(n1729), .B(n1728), .Z(n1737) );
  NAND U2658 ( .A(n1731), .B(n1730), .Z(n1735) );
  NANDN U2659 ( .A(n1733), .B(n1732), .Z(n1734) );
  AND U2660 ( .A(n1735), .B(n1734), .Z(n1736) );
  XNOR U2661 ( .A(n1737), .B(n1736), .Z(n1738) );
  XNOR U2662 ( .A(n1739), .B(n1738), .Z(n1747) );
  NAND U2663 ( .A(n1741), .B(n1740), .Z(n1745) );
  NANDN U2664 ( .A(n1743), .B(n1742), .Z(n1744) );
  NAND U2665 ( .A(n1745), .B(n1744), .Z(n1746) );
  XNOR U2666 ( .A(n1747), .B(n1746), .Z(n1748) );
  XNOR U2667 ( .A(n1749), .B(n1748), .Z(n1750) );
  XOR U2668 ( .A(n1751), .B(n1750), .Z(n1767) );
  NANDN U2669 ( .A(n1753), .B(n1752), .Z(n1757) );
  NANDN U2670 ( .A(n1755), .B(n1754), .Z(n1756) );
  NAND U2671 ( .A(n1757), .B(n1756), .Z(n1765) );
  OR U2672 ( .A(n1759), .B(n1758), .Z(n1763) );
  NAND U2673 ( .A(n1761), .B(n1760), .Z(n1762) );
  AND U2674 ( .A(n1763), .B(n1762), .Z(n1764) );
  XOR U2675 ( .A(n1765), .B(n1764), .Z(n1766) );
  XNOR U2676 ( .A(n1767), .B(n1766), .Z(n1768) );
  XOR U2677 ( .A(n1769), .B(n1768), .Z(n1785) );
  OR U2678 ( .A(n1771), .B(n1770), .Z(n1775) );
  NANDN U2679 ( .A(n1773), .B(n1772), .Z(n1774) );
  AND U2680 ( .A(n1775), .B(n1774), .Z(n1783) );
  OR U2681 ( .A(n1777), .B(n1776), .Z(n1781) );
  NANDN U2682 ( .A(n1779), .B(n1778), .Z(n1780) );
  AND U2683 ( .A(n1781), .B(n1780), .Z(n1782) );
  XNOR U2684 ( .A(n1783), .B(n1782), .Z(n1784) );
  XNOR U2685 ( .A(n1785), .B(n1784), .Z(n1786) );
  XOR U2686 ( .A(n1787), .B(n1786), .Z(n1788) );
  XNOR U2687 ( .A(n1789), .B(n1788), .Z(n1790) );
  XOR U2688 ( .A(n1791), .B(n1790), .Z(n1807) );
  NAND U2689 ( .A(n1793), .B(n1792), .Z(n1797) );
  NANDN U2690 ( .A(n1795), .B(n1794), .Z(n1796) );
  AND U2691 ( .A(n1797), .B(n1796), .Z(n1805) );
  OR U2692 ( .A(n1799), .B(n1798), .Z(n1803) );
  NANDN U2693 ( .A(n1801), .B(n1800), .Z(n1802) );
  AND U2694 ( .A(n1803), .B(n1802), .Z(n1804) );
  XNOR U2695 ( .A(n1805), .B(n1804), .Z(n1806) );
  XNOR U2696 ( .A(n1807), .B(n1806), .Z(n1822) );
  NAND U2697 ( .A(n1809), .B(n1808), .Z(n1813) );
  NANDN U2698 ( .A(n1811), .B(n1810), .Z(n1812) );
  AND U2699 ( .A(n1813), .B(n1812), .Z(n1820) );
  NAND U2700 ( .A(n1816), .B(n1815), .Z(n1818) );
  AND U2701 ( .A(n1818), .B(n1817), .Z(n1819) );
  XNOR U2702 ( .A(n1820), .B(n1819), .Z(n1821) );
  XOR U2703 ( .A(n1822), .B(n1821), .Z(n1838) );
  NANDN U2704 ( .A(n1824), .B(n1823), .Z(n1828) );
  NANDN U2705 ( .A(n1826), .B(n1825), .Z(n1827) );
  AND U2706 ( .A(n1828), .B(n1827), .Z(n1836) );
  NAND U2707 ( .A(n1830), .B(n1829), .Z(n1834) );
  NANDN U2708 ( .A(n1832), .B(n1831), .Z(n1833) );
  AND U2709 ( .A(n1834), .B(n1833), .Z(n1835) );
  XNOR U2710 ( .A(n1836), .B(n1835), .Z(n1837) );
  XNOR U2711 ( .A(n1838), .B(n1837), .Z(o[7]) );
  NAND U2712 ( .A(x[32]), .B(y[168]), .Z(n1977) );
  NAND U2713 ( .A(x[8]), .B(y[48]), .Z(n1841) );
  XOR U2714 ( .A(n1977), .B(n1841), .Z(n1842) );
  AND U2715 ( .A(x[0]), .B(y[8]), .Z(n1849) );
  AND U2716 ( .A(x[16]), .B(y[88]), .Z(n1846) );
  XOR U2717 ( .A(n1849), .B(n1846), .Z(n1845) );
  AND U2718 ( .A(x[24]), .B(y[128]), .Z(n1844) );
  XNOR U2719 ( .A(n1845), .B(n1844), .Z(n1843) );
  XNOR U2720 ( .A(n1842), .B(n1843), .Z(o[8]) );
  AND U2721 ( .A(y[8]), .B(x[1]), .Z(n1840) );
  NAND U2722 ( .A(y[9]), .B(x[0]), .Z(n1839) );
  XNOR U2723 ( .A(n1840), .B(n1839), .Z(n1851) );
  AND U2724 ( .A(x[9]), .B(y[48]), .Z(n1850) );
  XOR U2725 ( .A(n1851), .B(n1850), .Z(n1868) );
  AND U2726 ( .A(x[33]), .B(y[168]), .Z(n2080) );
  AND U2727 ( .A(x[16]), .B(y[89]), .Z(n1854) );
  XOR U2728 ( .A(n2080), .B(n1854), .Z(n1856) );
  AND U2729 ( .A(x[32]), .B(y[169]), .Z(n1879) );
  NAND U2730 ( .A(x[17]), .B(y[88]), .Z(n1878) );
  XNOR U2731 ( .A(n1879), .B(n1878), .Z(n1855) );
  XOR U2732 ( .A(n1856), .B(n1855), .Z(n1866) );
  AND U2733 ( .A(x[8]), .B(y[49]), .Z(n2103) );
  AND U2734 ( .A(x[24]), .B(y[129]), .Z(n1871) );
  XOR U2735 ( .A(n2103), .B(n1871), .Z(n1873) );
  AND U2736 ( .A(x[25]), .B(y[128]), .Z(n1872) );
  XNOR U2737 ( .A(n1873), .B(n1872), .Z(n1865) );
  XNOR U2738 ( .A(n1866), .B(n1865), .Z(n1867) );
  XNOR U2739 ( .A(n1868), .B(n1867), .Z(n1862) );
  NAND U2740 ( .A(n1845), .B(n1844), .Z(n1848) );
  AND U2741 ( .A(n1849), .B(n1846), .Z(n1847) );
  ANDN U2742 ( .B(n1848), .A(n1847), .Z(n1859) );
  XNOR U2743 ( .A(n1860), .B(n1859), .Z(n1861) );
  XNOR U2744 ( .A(n1862), .B(n1861), .Z(o[9]) );
  NAND U2745 ( .A(x[1]), .B(y[9]), .Z(n1901) );
  NANDN U2746 ( .A(n1901), .B(n1849), .Z(n1853) );
  NAND U2747 ( .A(n1851), .B(n1850), .Z(n1852) );
  AND U2748 ( .A(n1853), .B(n1852), .Z(n1935) );
  NAND U2749 ( .A(n2080), .B(n1854), .Z(n1858) );
  NAND U2750 ( .A(n1856), .B(n1855), .Z(n1857) );
  AND U2751 ( .A(n1858), .B(n1857), .Z(n1934) );
  AND U2752 ( .A(x[24]), .B(y[130]), .Z(n1919) );
  NAND U2753 ( .A(x[0]), .B(y[10]), .Z(n1920) );
  XNOR U2754 ( .A(n1919), .B(n1920), .Z(n1921) );
  NAND U2755 ( .A(x[10]), .B(y[48]), .Z(n1922) );
  XNOR U2756 ( .A(n1921), .B(n1922), .Z(n1933) );
  XOR U2757 ( .A(n1934), .B(n1933), .Z(n1936) );
  XOR U2758 ( .A(n1935), .B(n1936), .Z(n1881) );
  NANDN U2759 ( .A(n1860), .B(n1859), .Z(n1864) );
  NAND U2760 ( .A(n1862), .B(n1861), .Z(n1863) );
  NAND U2761 ( .A(n1864), .B(n1863), .Z(n1880) );
  XNOR U2762 ( .A(n1881), .B(n1880), .Z(n1883) );
  NANDN U2763 ( .A(n1866), .B(n1865), .Z(n1870) );
  NANDN U2764 ( .A(n1868), .B(n1867), .Z(n1869) );
  AND U2765 ( .A(n1870), .B(n1869), .Z(n1889) );
  AND U2766 ( .A(x[2]), .B(y[8]), .Z(n1898) );
  NAND U2767 ( .A(x[16]), .B(y[90]), .Z(n1899) );
  XNOR U2768 ( .A(n1898), .B(n1899), .Z(n1900) );
  AND U2769 ( .A(x[26]), .B(y[128]), .Z(n1927) );
  XOR U2770 ( .A(n1928), .B(n1927), .Z(n1930) );
  AND U2771 ( .A(x[18]), .B(y[88]), .Z(n2007) );
  AND U2772 ( .A(x[32]), .B(y[170]), .Z(n1911) );
  XOR U2773 ( .A(n2007), .B(n1911), .Z(n1913) );
  AND U2774 ( .A(x[17]), .B(y[89]), .Z(n1912) );
  XOR U2775 ( .A(n1913), .B(n1912), .Z(n1929) );
  XOR U2776 ( .A(n1930), .B(n1929), .Z(n1886) );
  NAND U2777 ( .A(n2103), .B(n1871), .Z(n1875) );
  AND U2778 ( .A(n1873), .B(n1872), .Z(n1874) );
  ANDN U2779 ( .B(n1875), .A(n1874), .Z(n1895) );
  AND U2780 ( .A(y[168]), .B(x[34]), .Z(n1877) );
  NAND U2781 ( .A(y[169]), .B(x[33]), .Z(n1876) );
  XNOR U2782 ( .A(n1877), .B(n1876), .Z(n1926) );
  ANDN U2783 ( .B(n1879), .A(n1878), .Z(n1925) );
  XOR U2784 ( .A(n1926), .B(n1925), .Z(n1892) );
  AND U2785 ( .A(x[25]), .B(y[129]), .Z(n1904) );
  NAND U2786 ( .A(x[9]), .B(y[49]), .Z(n1905) );
  XNOR U2787 ( .A(n1904), .B(n1905), .Z(n1906) );
  NAND U2788 ( .A(x[8]), .B(y[50]), .Z(n1907) );
  XOR U2789 ( .A(n1906), .B(n1907), .Z(n1893) );
  XNOR U2790 ( .A(n1892), .B(n1893), .Z(n1894) );
  XOR U2791 ( .A(n1895), .B(n1894), .Z(n1887) );
  XNOR U2792 ( .A(n1886), .B(n1887), .Z(n1888) );
  XNOR U2793 ( .A(n1889), .B(n1888), .Z(n1882) );
  XNOR U2794 ( .A(n1883), .B(n1882), .Z(o[10]) );
  NANDN U2795 ( .A(n1881), .B(n1880), .Z(n1885) );
  NAND U2796 ( .A(n1883), .B(n1882), .Z(n1884) );
  AND U2797 ( .A(n1885), .B(n1884), .Z(n1957) );
  NANDN U2798 ( .A(n1887), .B(n1886), .Z(n1891) );
  NAND U2799 ( .A(n1889), .B(n1888), .Z(n1890) );
  AND U2800 ( .A(n1891), .B(n1890), .Z(n1942) );
  NANDN U2801 ( .A(n1893), .B(n1892), .Z(n1897) );
  NANDN U2802 ( .A(n1895), .B(n1894), .Z(n1896) );
  AND U2803 ( .A(n1897), .B(n1896), .Z(n1940) );
  NANDN U2804 ( .A(n1899), .B(n1898), .Z(n1903) );
  NANDN U2805 ( .A(n1901), .B(n1900), .Z(n1902) );
  NAND U2806 ( .A(n1903), .B(n1902), .Z(n1951) );
  NANDN U2807 ( .A(n1905), .B(n1904), .Z(n1909) );
  NANDN U2808 ( .A(n1907), .B(n1906), .Z(n1908) );
  AND U2809 ( .A(n1909), .B(n1908), .Z(n1998) );
  AND U2810 ( .A(x[24]), .B(y[131]), .Z(n2026) );
  AND U2811 ( .A(x[16]), .B(y[91]), .Z(n2025) );
  NAND U2812 ( .A(x[3]), .B(y[8]), .Z(n2024) );
  XOR U2813 ( .A(n2025), .B(n2024), .Z(n2027) );
  XOR U2814 ( .A(n2026), .B(n2027), .Z(n1996) );
  AND U2815 ( .A(x[18]), .B(y[89]), .Z(n2048) );
  NAND U2816 ( .A(y[88]), .B(x[19]), .Z(n1910) );
  XNOR U2817 ( .A(n2048), .B(n1910), .Z(n2010) );
  AND U2818 ( .A(x[17]), .B(y[90]), .Z(n2009) );
  XOR U2819 ( .A(n2010), .B(n2009), .Z(n1995) );
  XNOR U2820 ( .A(n1996), .B(n1995), .Z(n1997) );
  XNOR U2821 ( .A(n1998), .B(n1997), .Z(n1952) );
  XOR U2822 ( .A(n1951), .B(n1952), .Z(n1954) );
  NAND U2823 ( .A(n2007), .B(n1911), .Z(n1915) );
  AND U2824 ( .A(n1913), .B(n1912), .Z(n1914) );
  ANDN U2825 ( .B(n1915), .A(n1914), .Z(n2003) );
  AND U2826 ( .A(x[1]), .B(y[10]), .Z(n1973) );
  AND U2827 ( .A(x[2]), .B(y[9]), .Z(n1972) );
  NAND U2828 ( .A(x[25]), .B(y[130]), .Z(n1971) );
  XOR U2829 ( .A(n1972), .B(n1971), .Z(n1974) );
  XOR U2830 ( .A(n1973), .B(n1974), .Z(n2002) );
  AND U2831 ( .A(y[171]), .B(x[32]), .Z(n1917) );
  NAND U2832 ( .A(y[168]), .B(x[35]), .Z(n1916) );
  XNOR U2833 ( .A(n1917), .B(n1916), .Z(n1978) );
  AND U2834 ( .A(y[169]), .B(x[34]), .Z(n2059) );
  NAND U2835 ( .A(y[170]), .B(x[33]), .Z(n1918) );
  XOR U2836 ( .A(n2059), .B(n1918), .Z(n1979) );
  XNOR U2837 ( .A(n1978), .B(n1979), .Z(n2001) );
  XOR U2838 ( .A(n2002), .B(n2001), .Z(n2004) );
  XOR U2839 ( .A(n2003), .B(n2004), .Z(n1953) );
  XOR U2840 ( .A(n1954), .B(n1953), .Z(n1939) );
  XNOR U2841 ( .A(n1940), .B(n1939), .Z(n1941) );
  XOR U2842 ( .A(n1942), .B(n1941), .Z(n1958) );
  XNOR U2843 ( .A(n1957), .B(n1958), .Z(n1960) );
  NANDN U2844 ( .A(n1920), .B(n1919), .Z(n1924) );
  NANDN U2845 ( .A(n1922), .B(n1921), .Z(n1923) );
  AND U2846 ( .A(n1924), .B(n1923), .Z(n1964) );
  XNOR U2847 ( .A(n1964), .B(n1963), .Z(n1966) );
  AND U2848 ( .A(x[11]), .B(y[48]), .Z(n2018) );
  AND U2849 ( .A(x[0]), .B(y[11]), .Z(n2016) );
  NAND U2850 ( .A(x[26]), .B(y[129]), .Z(n2015) );
  XNOR U2851 ( .A(n2016), .B(n2015), .Z(n2017) );
  XOR U2852 ( .A(n2018), .B(n2017), .Z(n1991) );
  AND U2853 ( .A(x[8]), .B(y[51]), .Z(n1986) );
  AND U2854 ( .A(x[10]), .B(y[49]), .Z(n1984) );
  NAND U2855 ( .A(x[27]), .B(y[128]), .Z(n1983) );
  XNOR U2856 ( .A(n1984), .B(n1983), .Z(n1985) );
  XOR U2857 ( .A(n1986), .B(n1985), .Z(n1989) );
  AND U2858 ( .A(x[9]), .B(y[50]), .Z(n1990) );
  XOR U2859 ( .A(n1989), .B(n1990), .Z(n1992) );
  XOR U2860 ( .A(n1991), .B(n1992), .Z(n1965) );
  XOR U2861 ( .A(n1966), .B(n1965), .Z(n1946) );
  NAND U2862 ( .A(n1928), .B(n1927), .Z(n1932) );
  NAND U2863 ( .A(n1930), .B(n1929), .Z(n1931) );
  AND U2864 ( .A(n1932), .B(n1931), .Z(n1945) );
  XNOR U2865 ( .A(n1946), .B(n1945), .Z(n1948) );
  NANDN U2866 ( .A(n1934), .B(n1933), .Z(n1938) );
  OR U2867 ( .A(n1936), .B(n1935), .Z(n1937) );
  AND U2868 ( .A(n1938), .B(n1937), .Z(n1947) );
  XNOR U2869 ( .A(n1948), .B(n1947), .Z(n1959) );
  XOR U2870 ( .A(n1960), .B(n1959), .Z(o[11]) );
  NANDN U2871 ( .A(n1940), .B(n1939), .Z(n1944) );
  NANDN U2872 ( .A(n1942), .B(n1941), .Z(n1943) );
  AND U2873 ( .A(n1944), .B(n1943), .Z(n2038) );
  NANDN U2874 ( .A(n1946), .B(n1945), .Z(n1950) );
  NAND U2875 ( .A(n1948), .B(n1947), .Z(n1949) );
  NAND U2876 ( .A(n1950), .B(n1949), .Z(n2036) );
  NAND U2877 ( .A(n1952), .B(n1951), .Z(n1956) );
  NAND U2878 ( .A(n1954), .B(n1953), .Z(n1955) );
  AND U2879 ( .A(n1956), .B(n1955), .Z(n2037) );
  XOR U2880 ( .A(n2036), .B(n2037), .Z(n2039) );
  XOR U2881 ( .A(n2038), .B(n2039), .Z(n2030) );
  NANDN U2882 ( .A(n1958), .B(n1957), .Z(n1962) );
  NAND U2883 ( .A(n1960), .B(n1959), .Z(n1961) );
  NAND U2884 ( .A(n1962), .B(n1961), .Z(n2031) );
  XNOR U2885 ( .A(n2030), .B(n2031), .Z(n2033) );
  NANDN U2886 ( .A(n1964), .B(n1963), .Z(n1968) );
  NAND U2887 ( .A(n1966), .B(n1965), .Z(n1967) );
  AND U2888 ( .A(n1968), .B(n1967), .Z(n2043) );
  AND U2889 ( .A(x[10]), .B(y[50]), .Z(n2177) );
  AND U2890 ( .A(y[52]), .B(x[8]), .Z(n1970) );
  NAND U2891 ( .A(y[49]), .B(x[11]), .Z(n1969) );
  XOR U2892 ( .A(n1970), .B(n1969), .Z(n2104) );
  XNOR U2893 ( .A(n2177), .B(n2104), .Z(n2107) );
  NAND U2894 ( .A(x[9]), .B(y[51]), .Z(n2108) );
  XNOR U2895 ( .A(n2107), .B(n2108), .Z(n2110) );
  AND U2896 ( .A(x[28]), .B(y[128]), .Z(n2053) );
  NAND U2897 ( .A(x[1]), .B(y[11]), .Z(n2054) );
  XNOR U2898 ( .A(n2053), .B(n2054), .Z(n2055) );
  NAND U2899 ( .A(x[0]), .B(y[12]), .Z(n2056) );
  XNOR U2900 ( .A(n2055), .B(n2056), .Z(n2109) );
  XOR U2901 ( .A(n2110), .B(n2109), .Z(n2122) );
  NANDN U2902 ( .A(n1972), .B(n1971), .Z(n1976) );
  OR U2903 ( .A(n1974), .B(n1973), .Z(n1975) );
  AND U2904 ( .A(n1976), .B(n1975), .Z(n2120) );
  AND U2905 ( .A(x[35]), .B(y[171]), .Z(n2425) );
  NANDN U2906 ( .A(n1977), .B(n2425), .Z(n1981) );
  NANDN U2907 ( .A(n1979), .B(n1978), .Z(n1980) );
  AND U2908 ( .A(n1981), .B(n1980), .Z(n2119) );
  XNOR U2909 ( .A(n2120), .B(n2119), .Z(n2121) );
  XNOR U2910 ( .A(n2122), .B(n2121), .Z(n2140) );
  NAND U2911 ( .A(x[4]), .B(y[8]), .Z(n2089) );
  NAND U2912 ( .A(x[26]), .B(y[130]), .Z(n2088) );
  NAND U2913 ( .A(x[16]), .B(y[92]), .Z(n2087) );
  XNOR U2914 ( .A(n2088), .B(n2087), .Z(n2090) );
  AND U2915 ( .A(y[170]), .B(x[34]), .Z(n2023) );
  AND U2916 ( .A(x[33]), .B(y[169]), .Z(n1982) );
  NAND U2917 ( .A(n2023), .B(n1982), .Z(n2085) );
  NAND U2918 ( .A(x[20]), .B(y[88]), .Z(n2188) );
  NAND U2919 ( .A(x[32]), .B(y[172]), .Z(n2255) );
  XNOR U2920 ( .A(n2188), .B(n2255), .Z(n2086) );
  XOR U2921 ( .A(n2085), .B(n2086), .Z(n2068) );
  XOR U2922 ( .A(n2069), .B(n2068), .Z(n2070) );
  NANDN U2923 ( .A(n1984), .B(n1983), .Z(n1988) );
  NANDN U2924 ( .A(n1986), .B(n1985), .Z(n1987) );
  NAND U2925 ( .A(n1988), .B(n1987), .Z(n2071) );
  XOR U2926 ( .A(n2070), .B(n2071), .Z(n2137) );
  NAND U2927 ( .A(n1990), .B(n1989), .Z(n1994) );
  NAND U2928 ( .A(n1992), .B(n1991), .Z(n1993) );
  AND U2929 ( .A(n1994), .B(n1993), .Z(n2138) );
  XOR U2930 ( .A(n2137), .B(n2138), .Z(n2139) );
  XNOR U2931 ( .A(n2140), .B(n2139), .Z(n2042) );
  XNOR U2932 ( .A(n2043), .B(n2042), .Z(n2045) );
  NANDN U2933 ( .A(n1996), .B(n1995), .Z(n2000) );
  NANDN U2934 ( .A(n1998), .B(n1997), .Z(n1999) );
  NAND U2935 ( .A(n2000), .B(n1999), .Z(n2126) );
  NANDN U2936 ( .A(n2002), .B(n2001), .Z(n2006) );
  OR U2937 ( .A(n2004), .B(n2003), .Z(n2005) );
  NAND U2938 ( .A(n2006), .B(n2005), .Z(n2125) );
  XOR U2939 ( .A(n2126), .B(n2125), .Z(n2128) );
  AND U2940 ( .A(x[19]), .B(y[89]), .Z(n2008) );
  NAND U2941 ( .A(n2008), .B(n2007), .Z(n2012) );
  NAND U2942 ( .A(n2010), .B(n2009), .Z(n2011) );
  NAND U2943 ( .A(n2012), .B(n2011), .Z(n2131) );
  AND U2944 ( .A(x[12]), .B(y[48]), .Z(n2062) );
  NAND U2945 ( .A(x[24]), .B(y[132]), .Z(n2063) );
  XNOR U2946 ( .A(n2062), .B(n2063), .Z(n2064) );
  NAND U2947 ( .A(x[25]), .B(y[131]), .Z(n2065) );
  XNOR U2948 ( .A(n2064), .B(n2065), .Z(n2113) );
  AND U2949 ( .A(y[90]), .B(x[18]), .Z(n2014) );
  NAND U2950 ( .A(y[89]), .B(x[19]), .Z(n2013) );
  XNOR U2951 ( .A(n2014), .B(n2013), .Z(n2049) );
  NAND U2952 ( .A(x[17]), .B(y[91]), .Z(n2050) );
  XOR U2953 ( .A(n2049), .B(n2050), .Z(n2114) );
  XNOR U2954 ( .A(n2113), .B(n2114), .Z(n2115) );
  NANDN U2955 ( .A(n2016), .B(n2015), .Z(n2020) );
  NANDN U2956 ( .A(n2018), .B(n2017), .Z(n2019) );
  NAND U2957 ( .A(n2020), .B(n2019), .Z(n2116) );
  XNOR U2958 ( .A(n2115), .B(n2116), .Z(n2132) );
  XOR U2959 ( .A(n2131), .B(n2132), .Z(n2134) );
  NAND U2960 ( .A(x[2]), .B(y[10]), .Z(n2099) );
  NAND U2961 ( .A(x[27]), .B(y[129]), .Z(n2098) );
  NAND U2962 ( .A(x[3]), .B(y[9]), .Z(n2097) );
  XNOR U2963 ( .A(n2098), .B(n2097), .Z(n2100) );
  AND U2964 ( .A(y[171]), .B(x[33]), .Z(n2022) );
  NAND U2965 ( .A(y[168]), .B(x[36]), .Z(n2021) );
  XNOR U2966 ( .A(n2022), .B(n2021), .Z(n2082) );
  AND U2967 ( .A(x[35]), .B(y[169]), .Z(n2195) );
  XOR U2968 ( .A(n2195), .B(n2023), .Z(n2081) );
  XOR U2969 ( .A(n2082), .B(n2081), .Z(n2074) );
  XOR U2970 ( .A(n2075), .B(n2074), .Z(n2076) );
  NANDN U2971 ( .A(n2025), .B(n2024), .Z(n2029) );
  OR U2972 ( .A(n2027), .B(n2026), .Z(n2028) );
  NAND U2973 ( .A(n2029), .B(n2028), .Z(n2077) );
  XNOR U2974 ( .A(n2076), .B(n2077), .Z(n2133) );
  XOR U2975 ( .A(n2134), .B(n2133), .Z(n2127) );
  XOR U2976 ( .A(n2128), .B(n2127), .Z(n2044) );
  XNOR U2977 ( .A(n2045), .B(n2044), .Z(n2032) );
  XNOR U2978 ( .A(n2033), .B(n2032), .Z(o[12]) );
  NANDN U2979 ( .A(n2031), .B(n2030), .Z(n2035) );
  NAND U2980 ( .A(n2033), .B(n2032), .Z(n2034) );
  AND U2981 ( .A(n2035), .B(n2034), .Z(n2284) );
  NAND U2982 ( .A(n2037), .B(n2036), .Z(n2041) );
  NAND U2983 ( .A(n2039), .B(n2038), .Z(n2040) );
  NAND U2984 ( .A(n2041), .B(n2040), .Z(n2285) );
  XNOR U2985 ( .A(n2284), .B(n2285), .Z(n2287) );
  NANDN U2986 ( .A(n2043), .B(n2042), .Z(n2047) );
  NAND U2987 ( .A(n2045), .B(n2044), .Z(n2046) );
  AND U2988 ( .A(n2047), .B(n2046), .Z(n2144) );
  AND U2989 ( .A(x[19]), .B(y[90]), .Z(n2190) );
  NAND U2990 ( .A(n2190), .B(n2048), .Z(n2052) );
  NANDN U2991 ( .A(n2050), .B(n2049), .Z(n2051) );
  NAND U2992 ( .A(n2052), .B(n2051), .Z(n2159) );
  NANDN U2993 ( .A(n2054), .B(n2053), .Z(n2058) );
  NANDN U2994 ( .A(n2056), .B(n2055), .Z(n2057) );
  NAND U2995 ( .A(n2058), .B(n2057), .Z(n2167) );
  AND U2996 ( .A(x[13]), .B(y[48]), .Z(n2202) );
  AND U2997 ( .A(x[18]), .B(y[91]), .Z(n2201) );
  XOR U2998 ( .A(n2202), .B(n2201), .Z(n2203) );
  AND U2999 ( .A(x[24]), .B(y[133]), .Z(n2403) );
  XOR U3000 ( .A(n2203), .B(n2403), .Z(n2166) );
  AND U3001 ( .A(x[28]), .B(y[129]), .Z(n2197) );
  AND U3002 ( .A(x[5]), .B(y[8]), .Z(n2196) );
  XOR U3003 ( .A(n2197), .B(n2196), .Z(n2198) );
  AND U3004 ( .A(x[4]), .B(y[9]), .Z(n2379) );
  XOR U3005 ( .A(n2198), .B(n2379), .Z(n2165) );
  XOR U3006 ( .A(n2166), .B(n2165), .Z(n2168) );
  XOR U3007 ( .A(n2167), .B(n2168), .Z(n2160) );
  XOR U3008 ( .A(n2159), .B(n2160), .Z(n2162) );
  AND U3009 ( .A(y[170]), .B(x[35]), .Z(n2094) );
  AND U3010 ( .A(n2094), .B(n2059), .Z(n2257) );
  AND U3011 ( .A(y[173]), .B(x[32]), .Z(n2061) );
  AND U3012 ( .A(y[172]), .B(x[33]), .Z(n2060) );
  XOR U3013 ( .A(n2061), .B(n2060), .Z(n2256) );
  XOR U3014 ( .A(n2257), .B(n2256), .Z(n2279) );
  AND U3015 ( .A(x[8]), .B(y[53]), .Z(n2269) );
  AND U3016 ( .A(x[1]), .B(y[12]), .Z(n2268) );
  XOR U3017 ( .A(n2269), .B(n2268), .Z(n2271) );
  AND U3018 ( .A(x[12]), .B(y[49]), .Z(n2270) );
  XOR U3019 ( .A(n2271), .B(n2270), .Z(n2278) );
  XOR U3020 ( .A(n2279), .B(n2278), .Z(n2281) );
  NANDN U3021 ( .A(n2063), .B(n2062), .Z(n2067) );
  NANDN U3022 ( .A(n2065), .B(n2064), .Z(n2066) );
  NAND U3023 ( .A(n2067), .B(n2066), .Z(n2280) );
  XOR U3024 ( .A(n2281), .B(n2280), .Z(n2161) );
  XOR U3025 ( .A(n2162), .B(n2161), .Z(n2208) );
  NAND U3026 ( .A(n2069), .B(n2068), .Z(n2073) );
  NANDN U3027 ( .A(n2071), .B(n2070), .Z(n2072) );
  NAND U3028 ( .A(n2073), .B(n2072), .Z(n2207) );
  NAND U3029 ( .A(n2075), .B(n2074), .Z(n2079) );
  NANDN U3030 ( .A(n2077), .B(n2076), .Z(n2078) );
  NAND U3031 ( .A(n2079), .B(n2078), .Z(n2206) );
  XNOR U3032 ( .A(n2207), .B(n2206), .Z(n2209) );
  AND U3033 ( .A(x[36]), .B(y[171]), .Z(n2493) );
  NAND U3034 ( .A(n2493), .B(n2080), .Z(n2084) );
  NAND U3035 ( .A(n2082), .B(n2081), .Z(n2083) );
  NAND U3036 ( .A(n2084), .B(n2083), .Z(n2224) );
  XOR U3037 ( .A(n2224), .B(n2225), .Z(n2227) );
  NAND U3038 ( .A(n2088), .B(n2087), .Z(n2092) );
  NANDN U3039 ( .A(n2090), .B(n2089), .Z(n2091) );
  AND U3040 ( .A(n2092), .B(n2091), .Z(n2215) );
  AND U3041 ( .A(x[11]), .B(y[50]), .Z(n2348) );
  NAND U3042 ( .A(y[51]), .B(x[10]), .Z(n2093) );
  XNOR U3043 ( .A(n2348), .B(n2093), .Z(n2179) );
  AND U3044 ( .A(x[9]), .B(y[52]), .Z(n2178) );
  XOR U3045 ( .A(n2179), .B(n2178), .Z(n2213) );
  AND U3046 ( .A(x[34]), .B(y[171]), .Z(n2172) );
  AND U3047 ( .A(x[37]), .B(y[168]), .Z(n2171) );
  XOR U3048 ( .A(n2172), .B(n2171), .Z(n2174) );
  NAND U3049 ( .A(x[36]), .B(y[169]), .Z(n2446) );
  XNOR U3050 ( .A(n2094), .B(n2446), .Z(n2173) );
  XOR U3051 ( .A(n2174), .B(n2173), .Z(n2212) );
  XOR U3052 ( .A(n2213), .B(n2212), .Z(n2214) );
  XOR U3053 ( .A(n2215), .B(n2214), .Z(n2226) );
  XOR U3054 ( .A(n2227), .B(n2226), .Z(n2239) );
  AND U3055 ( .A(x[21]), .B(y[88]), .Z(n2096) );
  AND U3056 ( .A(y[89]), .B(x[20]), .Z(n2095) );
  XOR U3057 ( .A(n2096), .B(n2095), .Z(n2189) );
  XOR U3058 ( .A(n2190), .B(n2189), .Z(n2261) );
  AND U3059 ( .A(x[29]), .B(y[128]), .Z(n2183) );
  AND U3060 ( .A(x[3]), .B(y[10]), .Z(n2182) );
  XOR U3061 ( .A(n2183), .B(n2182), .Z(n2185) );
  AND U3062 ( .A(x[2]), .B(y[11]), .Z(n2184) );
  XOR U3063 ( .A(n2185), .B(n2184), .Z(n2260) );
  XOR U3064 ( .A(n2261), .B(n2260), .Z(n2263) );
  NAND U3065 ( .A(n2098), .B(n2097), .Z(n2102) );
  NANDN U3066 ( .A(n2100), .B(n2099), .Z(n2101) );
  AND U3067 ( .A(n2102), .B(n2101), .Z(n2262) );
  XOR U3068 ( .A(n2263), .B(n2262), .Z(n2237) );
  AND U3069 ( .A(x[11]), .B(y[52]), .Z(n2492) );
  NAND U3070 ( .A(n2492), .B(n2103), .Z(n2106) );
  NANDN U3071 ( .A(n2104), .B(n2177), .Z(n2105) );
  NAND U3072 ( .A(n2106), .B(n2105), .Z(n2220) );
  AND U3073 ( .A(x[27]), .B(y[130]), .Z(n2242) );
  AND U3074 ( .A(x[17]), .B(y[92]), .Z(n2390) );
  XOR U3075 ( .A(n2242), .B(n2390), .Z(n2244) );
  AND U3076 ( .A(x[16]), .B(y[93]), .Z(n2243) );
  XOR U3077 ( .A(n2244), .B(n2243), .Z(n2219) );
  AND U3078 ( .A(x[0]), .B(y[13]), .Z(n2248) );
  AND U3079 ( .A(x[25]), .B(y[132]), .Z(n2247) );
  XOR U3080 ( .A(n2248), .B(n2247), .Z(n2250) );
  AND U3081 ( .A(x[26]), .B(y[131]), .Z(n2249) );
  XOR U3082 ( .A(n2250), .B(n2249), .Z(n2218) );
  XOR U3083 ( .A(n2219), .B(n2218), .Z(n2221) );
  XNOR U3084 ( .A(n2220), .B(n2221), .Z(n2236) );
  NANDN U3085 ( .A(n2108), .B(n2107), .Z(n2112) );
  NAND U3086 ( .A(n2110), .B(n2109), .Z(n2111) );
  NAND U3087 ( .A(n2112), .B(n2111), .Z(n2231) );
  NANDN U3088 ( .A(n2114), .B(n2113), .Z(n2118) );
  NANDN U3089 ( .A(n2116), .B(n2115), .Z(n2117) );
  NAND U3090 ( .A(n2118), .B(n2117), .Z(n2230) );
  XOR U3091 ( .A(n2231), .B(n2230), .Z(n2233) );
  NANDN U3092 ( .A(n2120), .B(n2119), .Z(n2124) );
  NANDN U3093 ( .A(n2122), .B(n2121), .Z(n2123) );
  AND U3094 ( .A(n2124), .B(n2123), .Z(n2232) );
  XOR U3095 ( .A(n2233), .B(n2232), .Z(n2147) );
  XNOR U3096 ( .A(n2149), .B(n2150), .Z(n2143) );
  XNOR U3097 ( .A(n2144), .B(n2143), .Z(n2146) );
  NAND U3098 ( .A(n2126), .B(n2125), .Z(n2130) );
  NAND U3099 ( .A(n2128), .B(n2127), .Z(n2129) );
  NAND U3100 ( .A(n2130), .B(n2129), .Z(n2155) );
  NAND U3101 ( .A(n2132), .B(n2131), .Z(n2136) );
  NAND U3102 ( .A(n2134), .B(n2133), .Z(n2135) );
  NAND U3103 ( .A(n2136), .B(n2135), .Z(n2153) );
  NAND U3104 ( .A(n2138), .B(n2137), .Z(n2142) );
  NAND U3105 ( .A(n2140), .B(n2139), .Z(n2141) );
  AND U3106 ( .A(n2142), .B(n2141), .Z(n2154) );
  XOR U3107 ( .A(n2153), .B(n2154), .Z(n2156) );
  XOR U3108 ( .A(n2155), .B(n2156), .Z(n2145) );
  XOR U3109 ( .A(n2146), .B(n2145), .Z(n2286) );
  XOR U3110 ( .A(n2287), .B(n2286), .Z(o[13]) );
  NANDN U3111 ( .A(n2148), .B(n2147), .Z(n2152) );
  NANDN U3112 ( .A(n2150), .B(n2149), .Z(n2151) );
  AND U3113 ( .A(n2152), .B(n2151), .Z(n2589) );
  NAND U3114 ( .A(n2154), .B(n2153), .Z(n2158) );
  NAND U3115 ( .A(n2156), .B(n2155), .Z(n2157) );
  AND U3116 ( .A(n2158), .B(n2157), .Z(n2588) );
  XOR U3117 ( .A(n2589), .B(n2588), .Z(n2591) );
  NAND U3118 ( .A(n2160), .B(n2159), .Z(n2164) );
  NAND U3119 ( .A(n2162), .B(n2161), .Z(n2163) );
  AND U3120 ( .A(n2164), .B(n2163), .Z(n2583) );
  NAND U3121 ( .A(n2166), .B(n2165), .Z(n2170) );
  NAND U3122 ( .A(n2168), .B(n2167), .Z(n2169) );
  NAND U3123 ( .A(n2170), .B(n2169), .Z(n2550) );
  NAND U3124 ( .A(n2172), .B(n2171), .Z(n2176) );
  NAND U3125 ( .A(n2174), .B(n2173), .Z(n2175) );
  NAND U3126 ( .A(n2176), .B(n2175), .Z(n2328) );
  AND U3127 ( .A(y[51]), .B(x[11]), .Z(n2266) );
  NAND U3128 ( .A(n2177), .B(n2266), .Z(n2181) );
  NAND U3129 ( .A(n2179), .B(n2178), .Z(n2180) );
  AND U3130 ( .A(n2181), .B(n2180), .Z(n2351) );
  AND U3131 ( .A(x[27]), .B(y[131]), .Z(n2441) );
  AND U3132 ( .A(x[19]), .B(y[91]), .Z(n2440) );
  XOR U3133 ( .A(n2441), .B(n2440), .Z(n2439) );
  AND U3134 ( .A(x[3]), .B(y[11]), .Z(n2438) );
  XOR U3135 ( .A(n2439), .B(n2438), .Z(n2354) );
  AND U3136 ( .A(x[26]), .B(y[132]), .Z(n2366) );
  AND U3137 ( .A(x[20]), .B(y[90]), .Z(n2365) );
  XOR U3138 ( .A(n2366), .B(n2365), .Z(n2364) );
  AND U3139 ( .A(x[2]), .B(y[12]), .Z(n2363) );
  XNOR U3140 ( .A(n2364), .B(n2363), .Z(n2353) );
  XNOR U3141 ( .A(n2351), .B(n2352), .Z(n2331) );
  NAND U3142 ( .A(n2183), .B(n2182), .Z(n2187) );
  NAND U3143 ( .A(n2185), .B(n2184), .Z(n2186) );
  NAND U3144 ( .A(n2187), .B(n2186), .Z(n2330) );
  XOR U3145 ( .A(n2328), .B(n2329), .Z(n2551) );
  XOR U3146 ( .A(n2550), .B(n2551), .Z(n2548) );
  AND U3147 ( .A(x[21]), .B(y[89]), .Z(n2360) );
  NANDN U3148 ( .A(n2188), .B(n2360), .Z(n2192) );
  NAND U3149 ( .A(n2190), .B(n2189), .Z(n2191) );
  AND U3150 ( .A(n2192), .B(n2191), .Z(n2314) );
  AND U3151 ( .A(y[9]), .B(x[5]), .Z(n2194) );
  NAND U3152 ( .A(y[10]), .B(x[4]), .Z(n2193) );
  XNOR U3153 ( .A(n2194), .B(n2193), .Z(n2378) );
  AND U3154 ( .A(x[30]), .B(y[128]), .Z(n2377) );
  XOR U3155 ( .A(n2378), .B(n2377), .Z(n2317) );
  AND U3156 ( .A(x[33]), .B(y[173]), .Z(n2433) );
  AND U3157 ( .A(x[36]), .B(y[170]), .Z(n2254) );
  AND U3158 ( .A(n2195), .B(n2254), .Z(n2431) );
  AND U3159 ( .A(x[34]), .B(y[172]), .Z(n2430) );
  XOR U3160 ( .A(n2431), .B(n2430), .Z(n2432) );
  XNOR U3161 ( .A(n2433), .B(n2432), .Z(n2316) );
  XOR U3162 ( .A(n2314), .B(n2315), .Z(n2340) );
  NAND U3163 ( .A(n2197), .B(n2196), .Z(n2200) );
  NAND U3164 ( .A(n2198), .B(n2379), .Z(n2199) );
  NAND U3165 ( .A(n2200), .B(n2199), .Z(n2343) );
  NAND U3166 ( .A(n2202), .B(n2201), .Z(n2205) );
  NAND U3167 ( .A(n2203), .B(n2403), .Z(n2204) );
  NAND U3168 ( .A(n2205), .B(n2204), .Z(n2342) );
  XNOR U3169 ( .A(n2343), .B(n2342), .Z(n2341) );
  XNOR U3170 ( .A(n2548), .B(n2549), .Z(n2573) );
  NAND U3171 ( .A(n2207), .B(n2206), .Z(n2211) );
  NANDN U3172 ( .A(n2209), .B(n2208), .Z(n2210) );
  AND U3173 ( .A(n2211), .B(n2210), .Z(n2572) );
  NAND U3174 ( .A(n2213), .B(n2212), .Z(n2217) );
  NAND U3175 ( .A(n2215), .B(n2214), .Z(n2216) );
  AND U3176 ( .A(n2217), .B(n2216), .Z(n2543) );
  NAND U3177 ( .A(n2219), .B(n2218), .Z(n2223) );
  NAND U3178 ( .A(n2221), .B(n2220), .Z(n2222) );
  AND U3179 ( .A(n2223), .B(n2222), .Z(n2545) );
  NAND U3180 ( .A(n2225), .B(n2224), .Z(n2229) );
  NAND U3181 ( .A(n2227), .B(n2226), .Z(n2228) );
  AND U3182 ( .A(n2229), .B(n2228), .Z(n2544) );
  XOR U3183 ( .A(n2545), .B(n2544), .Z(n2542) );
  XOR U3184 ( .A(n2543), .B(n2542), .Z(n2570) );
  XOR U3185 ( .A(n2571), .B(n2570), .Z(n2582) );
  XOR U3186 ( .A(n2583), .B(n2582), .Z(n2585) );
  NAND U3187 ( .A(n2231), .B(n2230), .Z(n2235) );
  NAND U3188 ( .A(n2233), .B(n2232), .Z(n2234) );
  AND U3189 ( .A(n2235), .B(n2234), .Z(n2297) );
  NANDN U3190 ( .A(n2237), .B(n2236), .Z(n2241) );
  NANDN U3191 ( .A(n2239), .B(n2238), .Z(n2240) );
  NAND U3192 ( .A(n2241), .B(n2240), .Z(n2298) );
  NAND U3193 ( .A(n2242), .B(n2390), .Z(n2246) );
  NAND U3194 ( .A(n2244), .B(n2243), .Z(n2245) );
  NAND U3195 ( .A(n2246), .B(n2245), .Z(n2534) );
  NAND U3196 ( .A(n2248), .B(n2247), .Z(n2252) );
  NAND U3197 ( .A(n2250), .B(n2249), .Z(n2251) );
  AND U3198 ( .A(n2252), .B(n2251), .Z(n2308) );
  AND U3199 ( .A(x[1]), .B(y[13]), .Z(n2374) );
  AND U3200 ( .A(x[14]), .B(y[48]), .Z(n2373) );
  XOR U3201 ( .A(n2374), .B(n2373), .Z(n2372) );
  AND U3202 ( .A(x[8]), .B(y[54]), .Z(n2371) );
  XOR U3203 ( .A(n2372), .B(n2371), .Z(n2311) );
  NAND U3204 ( .A(y[169]), .B(x[37]), .Z(n2253) );
  XNOR U3205 ( .A(n2254), .B(n2253), .Z(n2427) );
  AND U3206 ( .A(x[38]), .B(y[168]), .Z(n2426) );
  XOR U3207 ( .A(n2427), .B(n2426), .Z(n2424) );
  XNOR U3208 ( .A(n2425), .B(n2424), .Z(n2310) );
  XNOR U3209 ( .A(n2308), .B(n2309), .Z(n2537) );
  NANDN U3210 ( .A(n2255), .B(n2433), .Z(n2259) );
  NAND U3211 ( .A(n2257), .B(n2256), .Z(n2258) );
  NAND U3212 ( .A(n2259), .B(n2258), .Z(n2536) );
  XOR U3213 ( .A(n2534), .B(n2535), .Z(n2565) );
  NAND U3214 ( .A(n2261), .B(n2260), .Z(n2265) );
  NAND U3215 ( .A(n2263), .B(n2262), .Z(n2264) );
  AND U3216 ( .A(n2265), .B(n2264), .Z(n2567) );
  AND U3217 ( .A(x[32]), .B(y[174]), .Z(n2359) );
  XOR U3218 ( .A(n2360), .B(n2359), .Z(n2358) );
  AND U3219 ( .A(x[22]), .B(y[88]), .Z(n2357) );
  XOR U3220 ( .A(n2358), .B(n2357), .Z(n2323) );
  AND U3221 ( .A(x[16]), .B(y[94]), .Z(n2409) );
  AND U3222 ( .A(x[6]), .B(y[8]), .Z(n2408) );
  XOR U3223 ( .A(n2409), .B(n2408), .Z(n2407) );
  AND U3224 ( .A(x[29]), .B(y[129]), .Z(n2406) );
  XOR U3225 ( .A(n2407), .B(n2406), .Z(n2325) );
  AND U3226 ( .A(x[13]), .B(y[49]), .Z(n2396) );
  AND U3227 ( .A(x[10]), .B(y[52]), .Z(n2395) );
  XOR U3228 ( .A(n2396), .B(n2395), .Z(n2394) );
  AND U3229 ( .A(x[9]), .B(y[53]), .Z(n2393) );
  XOR U3230 ( .A(n2394), .B(n2393), .Z(n2347) );
  AND U3231 ( .A(x[12]), .B(y[50]), .Z(n2267) );
  XOR U3232 ( .A(n2267), .B(n2266), .Z(n2346) );
  XOR U3233 ( .A(n2347), .B(n2346), .Z(n2324) );
  XOR U3234 ( .A(n2325), .B(n2324), .Z(n2322) );
  XOR U3235 ( .A(n2323), .B(n2322), .Z(n2305) );
  NAND U3236 ( .A(n2269), .B(n2268), .Z(n2273) );
  NAND U3237 ( .A(n2271), .B(n2270), .Z(n2272) );
  AND U3238 ( .A(n2273), .B(n2272), .Z(n2418) );
  AND U3239 ( .A(x[28]), .B(y[130]), .Z(n2389) );
  AND U3240 ( .A(x[18]), .B(y[92]), .Z(n2275) );
  AND U3241 ( .A(y[93]), .B(x[17]), .Z(n2274) );
  XOR U3242 ( .A(n2275), .B(n2274), .Z(n2388) );
  XOR U3243 ( .A(n2389), .B(n2388), .Z(n2421) );
  AND U3244 ( .A(x[0]), .B(y[14]), .Z(n2402) );
  AND U3245 ( .A(y[134]), .B(x[24]), .Z(n2277) );
  AND U3246 ( .A(y[133]), .B(x[25]), .Z(n2276) );
  XOR U3247 ( .A(n2277), .B(n2276), .Z(n2401) );
  XNOR U3248 ( .A(n2402), .B(n2401), .Z(n2420) );
  XNOR U3249 ( .A(n2418), .B(n2419), .Z(n2304) );
  NAND U3250 ( .A(n2279), .B(n2278), .Z(n2283) );
  NAND U3251 ( .A(n2281), .B(n2280), .Z(n2282) );
  AND U3252 ( .A(n2283), .B(n2282), .Z(n2302) );
  XOR U3253 ( .A(n2303), .B(n2302), .Z(n2566) );
  XOR U3254 ( .A(n2567), .B(n2566), .Z(n2564) );
  XOR U3255 ( .A(n2298), .B(n2299), .Z(n2296) );
  XOR U3256 ( .A(n2297), .B(n2296), .Z(n2584) );
  XOR U3257 ( .A(n2585), .B(n2584), .Z(n2590) );
  XNOR U3258 ( .A(n2591), .B(n2590), .Z(n2292) );
  NANDN U3259 ( .A(n2285), .B(n2284), .Z(n2289) );
  NAND U3260 ( .A(n2287), .B(n2286), .Z(n2288) );
  NAND U3261 ( .A(n2289), .B(n2288), .Z(n2290) );
  XOR U3262 ( .A(n2291), .B(n2290), .Z(o[14]) );
  NAND U3263 ( .A(n2291), .B(n2290), .Z(n2295) );
  NANDN U3264 ( .A(n2293), .B(n2292), .Z(n2294) );
  AND U3265 ( .A(n2295), .B(n2294), .Z(n2581) );
  NAND U3266 ( .A(n2297), .B(n2296), .Z(n2301) );
  NAND U3267 ( .A(n2299), .B(n2298), .Z(n2300) );
  AND U3268 ( .A(n2301), .B(n2300), .Z(n2563) );
  NAND U3269 ( .A(n2303), .B(n2302), .Z(n2307) );
  NANDN U3270 ( .A(n2305), .B(n2304), .Z(n2306) );
  AND U3271 ( .A(n2307), .B(n2306), .Z(n2339) );
  NANDN U3272 ( .A(n2309), .B(n2308), .Z(n2313) );
  NANDN U3273 ( .A(n2311), .B(n2310), .Z(n2312) );
  AND U3274 ( .A(n2313), .B(n2312), .Z(n2321) );
  NANDN U3275 ( .A(n2315), .B(n2314), .Z(n2319) );
  NANDN U3276 ( .A(n2317), .B(n2316), .Z(n2318) );
  NAND U3277 ( .A(n2319), .B(n2318), .Z(n2320) );
  XNOR U3278 ( .A(n2321), .B(n2320), .Z(n2337) );
  NAND U3279 ( .A(n2323), .B(n2322), .Z(n2327) );
  NAND U3280 ( .A(n2325), .B(n2324), .Z(n2326) );
  AND U3281 ( .A(n2327), .B(n2326), .Z(n2335) );
  NAND U3282 ( .A(n2329), .B(n2328), .Z(n2333) );
  NANDN U3283 ( .A(n2331), .B(n2330), .Z(n2332) );
  NAND U3284 ( .A(n2333), .B(n2332), .Z(n2334) );
  XNOR U3285 ( .A(n2335), .B(n2334), .Z(n2336) );
  XNOR U3286 ( .A(n2337), .B(n2336), .Z(n2338) );
  XNOR U3287 ( .A(n2339), .B(n2338), .Z(n2561) );
  NANDN U3288 ( .A(n2341), .B(n2340), .Z(n2345) );
  NAND U3289 ( .A(n2343), .B(n2342), .Z(n2344) );
  AND U3290 ( .A(n2345), .B(n2344), .Z(n2559) );
  NAND U3291 ( .A(n2347), .B(n2346), .Z(n2350) );
  AND U3292 ( .A(x[12]), .B(y[51]), .Z(n2490) );
  NAND U3293 ( .A(n2348), .B(n2490), .Z(n2349) );
  AND U3294 ( .A(n2350), .B(n2349), .Z(n2533) );
  NANDN U3295 ( .A(n2352), .B(n2351), .Z(n2356) );
  NANDN U3296 ( .A(n2354), .B(n2353), .Z(n2355) );
  AND U3297 ( .A(n2356), .B(n2355), .Z(n2387) );
  NAND U3298 ( .A(n2358), .B(n2357), .Z(n2362) );
  NAND U3299 ( .A(n2360), .B(n2359), .Z(n2361) );
  AND U3300 ( .A(n2362), .B(n2361), .Z(n2370) );
  NAND U3301 ( .A(n2364), .B(n2363), .Z(n2368) );
  NAND U3302 ( .A(n2366), .B(n2365), .Z(n2367) );
  NAND U3303 ( .A(n2368), .B(n2367), .Z(n2369) );
  XNOR U3304 ( .A(n2370), .B(n2369), .Z(n2385) );
  NAND U3305 ( .A(n2372), .B(n2371), .Z(n2376) );
  NAND U3306 ( .A(n2374), .B(n2373), .Z(n2375) );
  AND U3307 ( .A(n2376), .B(n2375), .Z(n2383) );
  NAND U3308 ( .A(n2378), .B(n2377), .Z(n2381) );
  AND U3309 ( .A(x[5]), .B(y[10]), .Z(n2491) );
  NAND U3310 ( .A(n2379), .B(n2491), .Z(n2380) );
  NAND U3311 ( .A(n2381), .B(n2380), .Z(n2382) );
  XNOR U3312 ( .A(n2383), .B(n2382), .Z(n2384) );
  XNOR U3313 ( .A(n2385), .B(n2384), .Z(n2386) );
  XNOR U3314 ( .A(n2387), .B(n2386), .Z(n2417) );
  NAND U3315 ( .A(n2389), .B(n2388), .Z(n2392) );
  AND U3316 ( .A(x[18]), .B(y[93]), .Z(n2497) );
  NAND U3317 ( .A(n2390), .B(n2497), .Z(n2391) );
  AND U3318 ( .A(n2392), .B(n2391), .Z(n2400) );
  NAND U3319 ( .A(n2394), .B(n2393), .Z(n2398) );
  NAND U3320 ( .A(n2396), .B(n2395), .Z(n2397) );
  NAND U3321 ( .A(n2398), .B(n2397), .Z(n2399) );
  XNOR U3322 ( .A(n2400), .B(n2399), .Z(n2415) );
  NAND U3323 ( .A(n2402), .B(n2401), .Z(n2405) );
  AND U3324 ( .A(x[25]), .B(y[134]), .Z(n2496) );
  NAND U3325 ( .A(n2403), .B(n2496), .Z(n2404) );
  AND U3326 ( .A(n2405), .B(n2404), .Z(n2413) );
  NAND U3327 ( .A(n2407), .B(n2406), .Z(n2411) );
  NAND U3328 ( .A(n2409), .B(n2408), .Z(n2410) );
  NAND U3329 ( .A(n2411), .B(n2410), .Z(n2412) );
  XNOR U3330 ( .A(n2413), .B(n2412), .Z(n2414) );
  XNOR U3331 ( .A(n2415), .B(n2414), .Z(n2416) );
  XNOR U3332 ( .A(n2417), .B(n2416), .Z(n2531) );
  NANDN U3333 ( .A(n2419), .B(n2418), .Z(n2423) );
  NANDN U3334 ( .A(n2421), .B(n2420), .Z(n2422) );
  AND U3335 ( .A(n2423), .B(n2422), .Z(n2529) );
  NAND U3336 ( .A(n2425), .B(n2424), .Z(n2429) );
  AND U3337 ( .A(n2427), .B(n2426), .Z(n2428) );
  ANDN U3338 ( .B(n2429), .A(n2428), .Z(n2437) );
  AND U3339 ( .A(n2431), .B(n2430), .Z(n2435) );
  AND U3340 ( .A(n2433), .B(n2432), .Z(n2434) );
  OR U3341 ( .A(n2435), .B(n2434), .Z(n2436) );
  XNOR U3342 ( .A(n2437), .B(n2436), .Z(n2527) );
  NAND U3343 ( .A(n2439), .B(n2438), .Z(n2443) );
  NAND U3344 ( .A(n2441), .B(n2440), .Z(n2442) );
  AND U3345 ( .A(n2443), .B(n2442), .Z(n2525) );
  AND U3346 ( .A(y[54]), .B(x[9]), .Z(n2445) );
  NAND U3347 ( .A(y[53]), .B(x[10]), .Z(n2444) );
  XNOR U3348 ( .A(n2445), .B(n2444), .Z(n2451) );
  AND U3349 ( .A(y[135]), .B(x[24]), .Z(n2449) );
  AND U3350 ( .A(y[170]), .B(n2446), .Z(n2447) );
  NAND U3351 ( .A(n2447), .B(x[37]), .Z(n2448) );
  XNOR U3352 ( .A(n2449), .B(n2448), .Z(n2450) );
  XOR U3353 ( .A(n2451), .B(n2450), .Z(n2459) );
  AND U3354 ( .A(y[92]), .B(x[19]), .Z(n2453) );
  NAND U3355 ( .A(y[133]), .B(x[26]), .Z(n2452) );
  XNOR U3356 ( .A(n2453), .B(n2452), .Z(n2457) );
  AND U3357 ( .A(y[48]), .B(x[15]), .Z(n2455) );
  NAND U3358 ( .A(y[50]), .B(x[13]), .Z(n2454) );
  XNOR U3359 ( .A(n2455), .B(n2454), .Z(n2456) );
  XNOR U3360 ( .A(n2457), .B(n2456), .Z(n2458) );
  XNOR U3361 ( .A(n2459), .B(n2458), .Z(n2523) );
  AND U3362 ( .A(y[94]), .B(x[17]), .Z(n2461) );
  NAND U3363 ( .A(y[91]), .B(x[20]), .Z(n2460) );
  XNOR U3364 ( .A(n2461), .B(n2460), .Z(n2465) );
  AND U3365 ( .A(y[169]), .B(x[38]), .Z(n2463) );
  NAND U3366 ( .A(y[174]), .B(x[33]), .Z(n2462) );
  XNOR U3367 ( .A(n2463), .B(n2462), .Z(n2464) );
  XOR U3368 ( .A(n2465), .B(n2464), .Z(n2473) );
  AND U3369 ( .A(y[88]), .B(x[23]), .Z(n2467) );
  NAND U3370 ( .A(y[15]), .B(x[0]), .Z(n2466) );
  XNOR U3371 ( .A(n2467), .B(n2466), .Z(n2471) );
  AND U3372 ( .A(y[8]), .B(x[7]), .Z(n2469) );
  NAND U3373 ( .A(y[175]), .B(x[32]), .Z(n2468) );
  XNOR U3374 ( .A(n2469), .B(n2468), .Z(n2470) );
  XNOR U3375 ( .A(n2471), .B(n2470), .Z(n2472) );
  XNOR U3376 ( .A(n2473), .B(n2472), .Z(n2489) );
  AND U3377 ( .A(y[89]), .B(x[22]), .Z(n2475) );
  NAND U3378 ( .A(y[131]), .B(x[28]), .Z(n2474) );
  XNOR U3379 ( .A(n2475), .B(n2474), .Z(n2479) );
  AND U3380 ( .A(y[9]), .B(x[6]), .Z(n2477) );
  NAND U3381 ( .A(y[49]), .B(x[14]), .Z(n2476) );
  XNOR U3382 ( .A(n2477), .B(n2476), .Z(n2478) );
  XOR U3383 ( .A(n2479), .B(n2478), .Z(n2487) );
  AND U3384 ( .A(y[129]), .B(x[30]), .Z(n2481) );
  NAND U3385 ( .A(y[12]), .B(x[3]), .Z(n2480) );
  XNOR U3386 ( .A(n2481), .B(n2480), .Z(n2485) );
  AND U3387 ( .A(y[55]), .B(x[8]), .Z(n2483) );
  NAND U3388 ( .A(y[13]), .B(x[2]), .Z(n2482) );
  XNOR U3389 ( .A(n2483), .B(n2482), .Z(n2484) );
  XNOR U3390 ( .A(n2485), .B(n2484), .Z(n2486) );
  XNOR U3391 ( .A(n2487), .B(n2486), .Z(n2488) );
  XOR U3392 ( .A(n2489), .B(n2488), .Z(n2521) );
  XOR U3393 ( .A(n2491), .B(n2490), .Z(n2495) );
  XNOR U3394 ( .A(n2493), .B(n2492), .Z(n2494) );
  XNOR U3395 ( .A(n2495), .B(n2494), .Z(n2519) );
  AND U3396 ( .A(y[95]), .B(x[16]), .Z(n2517) );
  AND U3397 ( .A(y[132]), .B(x[27]), .Z(n2499) );
  XNOR U3398 ( .A(n2497), .B(n2496), .Z(n2498) );
  XNOR U3399 ( .A(n2499), .B(n2498), .Z(n2515) );
  AND U3400 ( .A(y[168]), .B(x[39]), .Z(n2501) );
  NAND U3401 ( .A(y[128]), .B(x[31]), .Z(n2500) );
  XNOR U3402 ( .A(n2501), .B(n2500), .Z(n2505) );
  AND U3403 ( .A(y[14]), .B(x[1]), .Z(n2503) );
  NAND U3404 ( .A(y[90]), .B(x[21]), .Z(n2502) );
  XNOR U3405 ( .A(n2503), .B(n2502), .Z(n2504) );
  XOR U3406 ( .A(n2505), .B(n2504), .Z(n2513) );
  AND U3407 ( .A(y[130]), .B(x[29]), .Z(n2507) );
  NAND U3408 ( .A(y[172]), .B(x[35]), .Z(n2506) );
  XNOR U3409 ( .A(n2507), .B(n2506), .Z(n2511) );
  AND U3410 ( .A(y[11]), .B(x[4]), .Z(n2509) );
  NAND U3411 ( .A(y[173]), .B(x[34]), .Z(n2508) );
  XNOR U3412 ( .A(n2509), .B(n2508), .Z(n2510) );
  XNOR U3413 ( .A(n2511), .B(n2510), .Z(n2512) );
  XNOR U3414 ( .A(n2513), .B(n2512), .Z(n2514) );
  XNOR U3415 ( .A(n2515), .B(n2514), .Z(n2516) );
  XNOR U3416 ( .A(n2517), .B(n2516), .Z(n2518) );
  XNOR U3417 ( .A(n2519), .B(n2518), .Z(n2520) );
  XNOR U3418 ( .A(n2521), .B(n2520), .Z(n2522) );
  XNOR U3419 ( .A(n2523), .B(n2522), .Z(n2524) );
  XNOR U3420 ( .A(n2525), .B(n2524), .Z(n2526) );
  XNOR U3421 ( .A(n2527), .B(n2526), .Z(n2528) );
  XNOR U3422 ( .A(n2529), .B(n2528), .Z(n2530) );
  XNOR U3423 ( .A(n2531), .B(n2530), .Z(n2532) );
  XNOR U3424 ( .A(n2533), .B(n2532), .Z(n2541) );
  NAND U3425 ( .A(n2535), .B(n2534), .Z(n2539) );
  NANDN U3426 ( .A(n2537), .B(n2536), .Z(n2538) );
  NAND U3427 ( .A(n2539), .B(n2538), .Z(n2540) );
  XNOR U3428 ( .A(n2541), .B(n2540), .Z(n2557) );
  NAND U3429 ( .A(n2543), .B(n2542), .Z(n2547) );
  NAND U3430 ( .A(n2545), .B(n2544), .Z(n2546) );
  AND U3431 ( .A(n2547), .B(n2546), .Z(n2555) );
  NANDN U3432 ( .A(n2549), .B(n2548), .Z(n2553) );
  NAND U3433 ( .A(n2551), .B(n2550), .Z(n2552) );
  NAND U3434 ( .A(n2553), .B(n2552), .Z(n2554) );
  XNOR U3435 ( .A(n2555), .B(n2554), .Z(n2556) );
  XNOR U3436 ( .A(n2557), .B(n2556), .Z(n2558) );
  XNOR U3437 ( .A(n2559), .B(n2558), .Z(n2560) );
  XNOR U3438 ( .A(n2561), .B(n2560), .Z(n2562) );
  XNOR U3439 ( .A(n2563), .B(n2562), .Z(n2579) );
  NANDN U3440 ( .A(n2565), .B(n2564), .Z(n2569) );
  NAND U3441 ( .A(n2567), .B(n2566), .Z(n2568) );
  AND U3442 ( .A(n2569), .B(n2568), .Z(n2577) );
  NAND U3443 ( .A(n2571), .B(n2570), .Z(n2575) );
  NANDN U3444 ( .A(n2573), .B(n2572), .Z(n2574) );
  NAND U3445 ( .A(n2575), .B(n2574), .Z(n2576) );
  XNOR U3446 ( .A(n2577), .B(n2576), .Z(n2578) );
  XNOR U3447 ( .A(n2579), .B(n2578), .Z(n2580) );
  XNOR U3448 ( .A(n2581), .B(n2580), .Z(n2597) );
  AND U3449 ( .A(n2583), .B(n2582), .Z(n2587) );
  AND U3450 ( .A(n2585), .B(n2584), .Z(n2586) );
  NOR U3451 ( .A(n2587), .B(n2586), .Z(n2595) );
  NAND U3452 ( .A(n2589), .B(n2588), .Z(n2593) );
  NAND U3453 ( .A(n2591), .B(n2590), .Z(n2592) );
  AND U3454 ( .A(n2593), .B(n2592), .Z(n2594) );
  XNOR U3455 ( .A(n2595), .B(n2594), .Z(n2596) );
  XNOR U3456 ( .A(n2597), .B(n2596), .Z(o[15]) );
  NAND U3457 ( .A(x[32]), .B(y[176]), .Z(n2712) );
  NAND U3458 ( .A(x[8]), .B(y[56]), .Z(n2600) );
  XOR U3459 ( .A(n2712), .B(n2600), .Z(n2601) );
  AND U3460 ( .A(x[0]), .B(y[16]), .Z(n2608) );
  AND U3461 ( .A(x[16]), .B(y[96]), .Z(n2605) );
  XOR U3462 ( .A(n2608), .B(n2605), .Z(n2604) );
  AND U3463 ( .A(x[24]), .B(y[136]), .Z(n2603) );
  XNOR U3464 ( .A(n2604), .B(n2603), .Z(n2602) );
  XNOR U3465 ( .A(n2601), .B(n2602), .Z(o[16]) );
  AND U3466 ( .A(y[16]), .B(x[1]), .Z(n2599) );
  NAND U3467 ( .A(y[17]), .B(x[0]), .Z(n2598) );
  XNOR U3468 ( .A(n2599), .B(n2598), .Z(n2610) );
  AND U3469 ( .A(x[9]), .B(y[56]), .Z(n2609) );
  XOR U3470 ( .A(n2610), .B(n2609), .Z(n2627) );
  AND U3471 ( .A(x[33]), .B(y[176]), .Z(n2832) );
  AND U3472 ( .A(x[16]), .B(y[97]), .Z(n2613) );
  XOR U3473 ( .A(n2832), .B(n2613), .Z(n2615) );
  AND U3474 ( .A(x[32]), .B(y[177]), .Z(n2638) );
  NAND U3475 ( .A(x[17]), .B(y[96]), .Z(n2637) );
  XNOR U3476 ( .A(n2638), .B(n2637), .Z(n2614) );
  XOR U3477 ( .A(n2615), .B(n2614), .Z(n2625) );
  AND U3478 ( .A(x[8]), .B(y[57]), .Z(n2856) );
  AND U3479 ( .A(x[24]), .B(y[137]), .Z(n2630) );
  XOR U3480 ( .A(n2856), .B(n2630), .Z(n2632) );
  AND U3481 ( .A(x[25]), .B(y[136]), .Z(n2631) );
  XNOR U3482 ( .A(n2632), .B(n2631), .Z(n2624) );
  XNOR U3483 ( .A(n2625), .B(n2624), .Z(n2626) );
  XNOR U3484 ( .A(n2627), .B(n2626), .Z(n2621) );
  NAND U3485 ( .A(n2604), .B(n2603), .Z(n2607) );
  AND U3486 ( .A(n2608), .B(n2605), .Z(n2606) );
  ANDN U3487 ( .B(n2607), .A(n2606), .Z(n2618) );
  XNOR U3488 ( .A(n2619), .B(n2618), .Z(n2620) );
  XNOR U3489 ( .A(n2621), .B(n2620), .Z(o[17]) );
  NAND U3490 ( .A(x[1]), .B(y[17]), .Z(n2660) );
  NANDN U3491 ( .A(n2660), .B(n2608), .Z(n2612) );
  NAND U3492 ( .A(n2610), .B(n2609), .Z(n2611) );
  AND U3493 ( .A(n2612), .B(n2611), .Z(n2680) );
  NAND U3494 ( .A(n2832), .B(n2613), .Z(n2617) );
  NAND U3495 ( .A(n2615), .B(n2614), .Z(n2616) );
  AND U3496 ( .A(n2617), .B(n2616), .Z(n2679) );
  AND U3497 ( .A(x[24]), .B(y[138]), .Z(n2684) );
  NAND U3498 ( .A(x[0]), .B(y[18]), .Z(n2685) );
  XNOR U3499 ( .A(n2684), .B(n2685), .Z(n2686) );
  NAND U3500 ( .A(x[10]), .B(y[56]), .Z(n2687) );
  XNOR U3501 ( .A(n2686), .B(n2687), .Z(n2678) );
  XOR U3502 ( .A(n2679), .B(n2678), .Z(n2681) );
  XOR U3503 ( .A(n2680), .B(n2681), .Z(n2640) );
  NANDN U3504 ( .A(n2619), .B(n2618), .Z(n2623) );
  NAND U3505 ( .A(n2621), .B(n2620), .Z(n2622) );
  NAND U3506 ( .A(n2623), .B(n2622), .Z(n2639) );
  XNOR U3507 ( .A(n2640), .B(n2639), .Z(n2642) );
  NANDN U3508 ( .A(n2625), .B(n2624), .Z(n2629) );
  NANDN U3509 ( .A(n2627), .B(n2626), .Z(n2628) );
  AND U3510 ( .A(n2629), .B(n2628), .Z(n2648) );
  AND U3511 ( .A(x[2]), .B(y[16]), .Z(n2657) );
  NAND U3512 ( .A(x[16]), .B(y[98]), .Z(n2658) );
  XNOR U3513 ( .A(n2657), .B(n2658), .Z(n2659) );
  AND U3514 ( .A(x[26]), .B(y[136]), .Z(n2692) );
  XOR U3515 ( .A(n2693), .B(n2692), .Z(n2695) );
  AND U3516 ( .A(x[18]), .B(y[96]), .Z(n2740) );
  AND U3517 ( .A(x[32]), .B(y[178]), .Z(n2670) );
  XOR U3518 ( .A(n2740), .B(n2670), .Z(n2672) );
  AND U3519 ( .A(x[17]), .B(y[97]), .Z(n2671) );
  XOR U3520 ( .A(n2672), .B(n2671), .Z(n2694) );
  XOR U3521 ( .A(n2695), .B(n2694), .Z(n2645) );
  NAND U3522 ( .A(n2856), .B(n2630), .Z(n2634) );
  AND U3523 ( .A(n2632), .B(n2631), .Z(n2633) );
  ANDN U3524 ( .B(n2634), .A(n2633), .Z(n2654) );
  AND U3525 ( .A(y[176]), .B(x[34]), .Z(n2636) );
  NAND U3526 ( .A(y[177]), .B(x[33]), .Z(n2635) );
  XNOR U3527 ( .A(n2636), .B(n2635), .Z(n2691) );
  ANDN U3528 ( .B(n2638), .A(n2637), .Z(n2690) );
  XOR U3529 ( .A(n2691), .B(n2690), .Z(n2651) );
  AND U3530 ( .A(x[25]), .B(y[137]), .Z(n2663) );
  NAND U3531 ( .A(x[9]), .B(y[57]), .Z(n2664) );
  XNOR U3532 ( .A(n2663), .B(n2664), .Z(n2665) );
  NAND U3533 ( .A(x[8]), .B(y[58]), .Z(n2666) );
  XOR U3534 ( .A(n2665), .B(n2666), .Z(n2652) );
  XNOR U3535 ( .A(n2651), .B(n2652), .Z(n2653) );
  XOR U3536 ( .A(n2654), .B(n2653), .Z(n2646) );
  XNOR U3537 ( .A(n2645), .B(n2646), .Z(n2647) );
  XNOR U3538 ( .A(n2648), .B(n2647), .Z(n2641) );
  XNOR U3539 ( .A(n2642), .B(n2641), .Z(o[18]) );
  NANDN U3540 ( .A(n2640), .B(n2639), .Z(n2644) );
  NAND U3541 ( .A(n2642), .B(n2641), .Z(n2643) );
  AND U3542 ( .A(n2644), .B(n2643), .Z(n2778) );
  NANDN U3543 ( .A(n2646), .B(n2645), .Z(n2650) );
  NAND U3544 ( .A(n2648), .B(n2647), .Z(n2649) );
  AND U3545 ( .A(n2650), .B(n2649), .Z(n2763) );
  NANDN U3546 ( .A(n2652), .B(n2651), .Z(n2656) );
  NANDN U3547 ( .A(n2654), .B(n2653), .Z(n2655) );
  AND U3548 ( .A(n2656), .B(n2655), .Z(n2761) );
  NANDN U3549 ( .A(n2658), .B(n2657), .Z(n2662) );
  NANDN U3550 ( .A(n2660), .B(n2659), .Z(n2661) );
  NAND U3551 ( .A(n2662), .B(n2661), .Z(n2772) );
  NANDN U3552 ( .A(n2664), .B(n2663), .Z(n2668) );
  NANDN U3553 ( .A(n2666), .B(n2665), .Z(n2667) );
  AND U3554 ( .A(n2668), .B(n2667), .Z(n2731) );
  AND U3555 ( .A(x[24]), .B(y[139]), .Z(n2756) );
  AND U3556 ( .A(x[16]), .B(y[99]), .Z(n2755) );
  NAND U3557 ( .A(x[3]), .B(y[16]), .Z(n2754) );
  XOR U3558 ( .A(n2755), .B(n2754), .Z(n2757) );
  XOR U3559 ( .A(n2756), .B(n2757), .Z(n2729) );
  AND U3560 ( .A(y[97]), .B(x[18]), .Z(n2812) );
  NAND U3561 ( .A(y[96]), .B(x[19]), .Z(n2669) );
  XNOR U3562 ( .A(n2812), .B(n2669), .Z(n2742) );
  AND U3563 ( .A(x[17]), .B(y[98]), .Z(n2741) );
  XOR U3564 ( .A(n2742), .B(n2741), .Z(n2728) );
  XNOR U3565 ( .A(n2729), .B(n2728), .Z(n2730) );
  XNOR U3566 ( .A(n2731), .B(n2730), .Z(n2773) );
  XOR U3567 ( .A(n2772), .B(n2773), .Z(n2775) );
  NAND U3568 ( .A(n2740), .B(n2670), .Z(n2674) );
  AND U3569 ( .A(n2672), .B(n2671), .Z(n2673) );
  ANDN U3570 ( .B(n2674), .A(n2673), .Z(n2736) );
  AND U3571 ( .A(x[1]), .B(y[18]), .Z(n2708) );
  AND U3572 ( .A(x[2]), .B(y[17]), .Z(n2707) );
  NAND U3573 ( .A(x[25]), .B(y[138]), .Z(n2706) );
  XOR U3574 ( .A(n2707), .B(n2706), .Z(n2709) );
  XOR U3575 ( .A(n2708), .B(n2709), .Z(n2735) );
  AND U3576 ( .A(y[179]), .B(x[32]), .Z(n2676) );
  NAND U3577 ( .A(y[176]), .B(x[35]), .Z(n2675) );
  XNOR U3578 ( .A(n2676), .B(n2675), .Z(n2713) );
  AND U3579 ( .A(y[177]), .B(x[34]), .Z(n2829) );
  NAND U3580 ( .A(y[178]), .B(x[33]), .Z(n2677) );
  XOR U3581 ( .A(n2829), .B(n2677), .Z(n2714) );
  XNOR U3582 ( .A(n2713), .B(n2714), .Z(n2734) );
  XOR U3583 ( .A(n2735), .B(n2734), .Z(n2737) );
  XOR U3584 ( .A(n2736), .B(n2737), .Z(n2774) );
  XOR U3585 ( .A(n2775), .B(n2774), .Z(n2760) );
  XNOR U3586 ( .A(n2761), .B(n2760), .Z(n2762) );
  XOR U3587 ( .A(n2763), .B(n2762), .Z(n2779) );
  XNOR U3588 ( .A(n2778), .B(n2779), .Z(n2781) );
  NANDN U3589 ( .A(n2679), .B(n2678), .Z(n2683) );
  OR U3590 ( .A(n2681), .B(n2680), .Z(n2682) );
  AND U3591 ( .A(n2683), .B(n2682), .Z(n2769) );
  NANDN U3592 ( .A(n2685), .B(n2684), .Z(n2689) );
  NANDN U3593 ( .A(n2687), .B(n2686), .Z(n2688) );
  AND U3594 ( .A(n2689), .B(n2688), .Z(n2699) );
  XNOR U3595 ( .A(n2699), .B(n2698), .Z(n2701) );
  AND U3596 ( .A(x[11]), .B(y[56]), .Z(n2748) );
  AND U3597 ( .A(x[0]), .B(y[19]), .Z(n2746) );
  NAND U3598 ( .A(x[26]), .B(y[137]), .Z(n2745) );
  XNOR U3599 ( .A(n2746), .B(n2745), .Z(n2747) );
  XOR U3600 ( .A(n2748), .B(n2747), .Z(n2726) );
  AND U3601 ( .A(x[8]), .B(y[59]), .Z(n2721) );
  AND U3602 ( .A(x[10]), .B(y[57]), .Z(n2719) );
  NAND U3603 ( .A(x[27]), .B(y[136]), .Z(n2718) );
  XNOR U3604 ( .A(n2719), .B(n2718), .Z(n2720) );
  XOR U3605 ( .A(n2721), .B(n2720), .Z(n2724) );
  AND U3606 ( .A(x[9]), .B(y[58]), .Z(n2725) );
  XOR U3607 ( .A(n2724), .B(n2725), .Z(n2727) );
  XOR U3608 ( .A(n2726), .B(n2727), .Z(n2700) );
  XOR U3609 ( .A(n2701), .B(n2700), .Z(n2767) );
  NAND U3610 ( .A(n2693), .B(n2692), .Z(n2697) );
  NAND U3611 ( .A(n2695), .B(n2694), .Z(n2696) );
  AND U3612 ( .A(n2697), .B(n2696), .Z(n2766) );
  XNOR U3613 ( .A(n2767), .B(n2766), .Z(n2768) );
  XNOR U3614 ( .A(n2769), .B(n2768), .Z(n2780) );
  XOR U3615 ( .A(n2781), .B(n2780), .Z(o[19]) );
  NANDN U3616 ( .A(n2699), .B(n2698), .Z(n2703) );
  NAND U3617 ( .A(n2701), .B(n2700), .Z(n2702) );
  AND U3618 ( .A(n2703), .B(n2702), .Z(n2795) );
  AND U3619 ( .A(x[10]), .B(y[58]), .Z(n2928) );
  AND U3620 ( .A(y[60]), .B(x[8]), .Z(n2705) );
  NAND U3621 ( .A(y[57]), .B(x[11]), .Z(n2704) );
  XOR U3622 ( .A(n2705), .B(n2704), .Z(n2857) );
  XNOR U3623 ( .A(n2928), .B(n2857), .Z(n2860) );
  NAND U3624 ( .A(x[9]), .B(y[59]), .Z(n2861) );
  XNOR U3625 ( .A(n2860), .B(n2861), .Z(n2863) );
  AND U3626 ( .A(x[28]), .B(y[136]), .Z(n2817) );
  NAND U3627 ( .A(x[1]), .B(y[19]), .Z(n2818) );
  XNOR U3628 ( .A(n2817), .B(n2818), .Z(n2819) );
  NAND U3629 ( .A(x[0]), .B(y[20]), .Z(n2820) );
  XNOR U3630 ( .A(n2819), .B(n2820), .Z(n2862) );
  XOR U3631 ( .A(n2863), .B(n2862), .Z(n2875) );
  NANDN U3632 ( .A(n2707), .B(n2706), .Z(n2711) );
  OR U3633 ( .A(n2709), .B(n2708), .Z(n2710) );
  AND U3634 ( .A(n2711), .B(n2710), .Z(n2873) );
  AND U3635 ( .A(x[35]), .B(y[179]), .Z(n3070) );
  NANDN U3636 ( .A(n2712), .B(n3070), .Z(n2716) );
  NANDN U3637 ( .A(n2714), .B(n2713), .Z(n2715) );
  AND U3638 ( .A(n2716), .B(n2715), .Z(n2872) );
  XNOR U3639 ( .A(n2873), .B(n2872), .Z(n2874) );
  XNOR U3640 ( .A(n2875), .B(n2874), .Z(n2893) );
  NAND U3641 ( .A(x[4]), .B(y[16]), .Z(n2841) );
  NAND U3642 ( .A(x[26]), .B(y[138]), .Z(n2840) );
  NAND U3643 ( .A(x[16]), .B(y[100]), .Z(n2839) );
  XNOR U3644 ( .A(n2840), .B(n2839), .Z(n2842) );
  AND U3645 ( .A(y[178]), .B(x[34]), .Z(n2753) );
  AND U3646 ( .A(x[33]), .B(y[177]), .Z(n2717) );
  NAND U3647 ( .A(n2753), .B(n2717), .Z(n2837) );
  NAND U3648 ( .A(x[32]), .B(y[180]), .Z(n2998) );
  NAND U3649 ( .A(x[20]), .B(y[96]), .Z(n2935) );
  XNOR U3650 ( .A(n2998), .B(n2935), .Z(n2838) );
  XOR U3651 ( .A(n2837), .B(n2838), .Z(n2800) );
  XOR U3652 ( .A(n2801), .B(n2800), .Z(n2802) );
  NANDN U3653 ( .A(n2719), .B(n2718), .Z(n2723) );
  NANDN U3654 ( .A(n2721), .B(n2720), .Z(n2722) );
  NAND U3655 ( .A(n2723), .B(n2722), .Z(n2803) );
  XOR U3656 ( .A(n2802), .B(n2803), .Z(n2889) );
  XOR U3657 ( .A(n2889), .B(n2890), .Z(n2892) );
  XNOR U3658 ( .A(n2893), .B(n2892), .Z(n2794) );
  XNOR U3659 ( .A(n2795), .B(n2794), .Z(n2797) );
  NANDN U3660 ( .A(n2729), .B(n2728), .Z(n2733) );
  NANDN U3661 ( .A(n2731), .B(n2730), .Z(n2732) );
  NAND U3662 ( .A(n2733), .B(n2732), .Z(n2878) );
  NANDN U3663 ( .A(n2735), .B(n2734), .Z(n2739) );
  OR U3664 ( .A(n2737), .B(n2736), .Z(n2738) );
  NAND U3665 ( .A(n2739), .B(n2738), .Z(n2879) );
  XOR U3666 ( .A(n2878), .B(n2879), .Z(n2881) );
  AND U3667 ( .A(x[12]), .B(y[56]), .Z(n2823) );
  NAND U3668 ( .A(x[24]), .B(y[140]), .Z(n2824) );
  XNOR U3669 ( .A(n2823), .B(n2824), .Z(n2825) );
  NAND U3670 ( .A(x[25]), .B(y[139]), .Z(n2826) );
  XNOR U3671 ( .A(n2825), .B(n2826), .Z(n2866) );
  AND U3672 ( .A(y[98]), .B(x[18]), .Z(n2744) );
  NAND U3673 ( .A(y[97]), .B(x[19]), .Z(n2743) );
  XNOR U3674 ( .A(n2744), .B(n2743), .Z(n2813) );
  NAND U3675 ( .A(x[17]), .B(y[99]), .Z(n2814) );
  XOR U3676 ( .A(n2813), .B(n2814), .Z(n2867) );
  XNOR U3677 ( .A(n2866), .B(n2867), .Z(n2868) );
  NANDN U3678 ( .A(n2746), .B(n2745), .Z(n2750) );
  NANDN U3679 ( .A(n2748), .B(n2747), .Z(n2749) );
  NAND U3680 ( .A(n2750), .B(n2749), .Z(n2869) );
  XNOR U3681 ( .A(n2868), .B(n2869), .Z(n2883) );
  XOR U3682 ( .A(n2882), .B(n2883), .Z(n2886) );
  NAND U3683 ( .A(x[2]), .B(y[18]), .Z(n2852) );
  NAND U3684 ( .A(x[27]), .B(y[137]), .Z(n2851) );
  NAND U3685 ( .A(x[3]), .B(y[17]), .Z(n2850) );
  XNOR U3686 ( .A(n2851), .B(n2850), .Z(n2853) );
  AND U3687 ( .A(y[179]), .B(x[33]), .Z(n2752) );
  NAND U3688 ( .A(y[176]), .B(x[36]), .Z(n2751) );
  XNOR U3689 ( .A(n2752), .B(n2751), .Z(n2834) );
  AND U3690 ( .A(y[177]), .B(x[35]), .Z(n2940) );
  XOR U3691 ( .A(n2940), .B(n2753), .Z(n2833) );
  XOR U3692 ( .A(n2834), .B(n2833), .Z(n2806) );
  XOR U3693 ( .A(n2807), .B(n2806), .Z(n2808) );
  NANDN U3694 ( .A(n2755), .B(n2754), .Z(n2759) );
  OR U3695 ( .A(n2757), .B(n2756), .Z(n2758) );
  NAND U3696 ( .A(n2759), .B(n2758), .Z(n2809) );
  XNOR U3697 ( .A(n2808), .B(n2809), .Z(n2885) );
  XOR U3698 ( .A(n2886), .B(n2885), .Z(n2880) );
  XOR U3699 ( .A(n2881), .B(n2880), .Z(n2796) );
  XNOR U3700 ( .A(n2797), .B(n2796), .Z(n2787) );
  NANDN U3701 ( .A(n2761), .B(n2760), .Z(n2765) );
  NANDN U3702 ( .A(n2763), .B(n2762), .Z(n2764) );
  AND U3703 ( .A(n2765), .B(n2764), .Z(n2790) );
  NANDN U3704 ( .A(n2767), .B(n2766), .Z(n2771) );
  NAND U3705 ( .A(n2769), .B(n2768), .Z(n2770) );
  NAND U3706 ( .A(n2771), .B(n2770), .Z(n2788) );
  NAND U3707 ( .A(n2773), .B(n2772), .Z(n2777) );
  NAND U3708 ( .A(n2775), .B(n2774), .Z(n2776) );
  AND U3709 ( .A(n2777), .B(n2776), .Z(n2789) );
  XNOR U3710 ( .A(n2788), .B(n2789), .Z(n2791) );
  NANDN U3711 ( .A(n2779), .B(n2778), .Z(n2783) );
  NAND U3712 ( .A(n2781), .B(n2780), .Z(n2782) );
  NAND U3713 ( .A(n2783), .B(n2782), .Z(n2785) );
  XNOR U3714 ( .A(n2786), .B(n2785), .Z(n2784) );
  XNOR U3715 ( .A(n2787), .B(n2784), .Z(o[20]) );
  NAND U3716 ( .A(n2789), .B(n2788), .Z(n2793) );
  NANDN U3717 ( .A(n2791), .B(n2790), .Z(n2792) );
  AND U3718 ( .A(n2793), .B(n2792), .Z(n2896) );
  XNOR U3719 ( .A(n2897), .B(n2896), .Z(n2899) );
  NANDN U3720 ( .A(n2795), .B(n2794), .Z(n2799) );
  NAND U3721 ( .A(n2797), .B(n2796), .Z(n2798) );
  AND U3722 ( .A(n2799), .B(n2798), .Z(n2903) );
  NAND U3723 ( .A(n2801), .B(n2800), .Z(n2805) );
  NANDN U3724 ( .A(n2803), .B(n2802), .Z(n2804) );
  NAND U3725 ( .A(n2805), .B(n2804), .Z(n2952) );
  NAND U3726 ( .A(n2807), .B(n2806), .Z(n2811) );
  NANDN U3727 ( .A(n2809), .B(n2808), .Z(n2810) );
  NAND U3728 ( .A(n2811), .B(n2810), .Z(n2953) );
  XOR U3729 ( .A(n2952), .B(n2953), .Z(n2956) );
  AND U3730 ( .A(x[19]), .B(y[98]), .Z(n2937) );
  NAND U3731 ( .A(n2937), .B(n2812), .Z(n2816) );
  NANDN U3732 ( .A(n2814), .B(n2813), .Z(n2815) );
  NAND U3733 ( .A(n2816), .B(n2815), .Z(n2914) );
  NANDN U3734 ( .A(n2818), .B(n2817), .Z(n2822) );
  NANDN U3735 ( .A(n2820), .B(n2819), .Z(n2821) );
  NAND U3736 ( .A(n2822), .B(n2821), .Z(n2922) );
  AND U3737 ( .A(x[24]), .B(y[141]), .Z(n3245) );
  AND U3738 ( .A(x[13]), .B(y[56]), .Z(n2948) );
  AND U3739 ( .A(x[18]), .B(y[99]), .Z(n2947) );
  XOR U3740 ( .A(n2948), .B(n2947), .Z(n2949) );
  XOR U3741 ( .A(n3245), .B(n2949), .Z(n2921) );
  AND U3742 ( .A(x[4]), .B(y[17]), .Z(n3164) );
  AND U3743 ( .A(x[28]), .B(y[137]), .Z(n2943) );
  AND U3744 ( .A(x[5]), .B(y[16]), .Z(n2942) );
  XOR U3745 ( .A(n2943), .B(n2942), .Z(n2944) );
  XOR U3746 ( .A(n3164), .B(n2944), .Z(n2920) );
  XOR U3747 ( .A(n2921), .B(n2920), .Z(n2923) );
  XOR U3748 ( .A(n2922), .B(n2923), .Z(n2915) );
  XOR U3749 ( .A(n2914), .B(n2915), .Z(n2917) );
  NANDN U3750 ( .A(n2824), .B(n2823), .Z(n2828) );
  NANDN U3751 ( .A(n2826), .B(n2825), .Z(n2827) );
  NAND U3752 ( .A(n2828), .B(n2827), .Z(n3011) );
  AND U3753 ( .A(x[35]), .B(y[178]), .Z(n2847) );
  AND U3754 ( .A(n2847), .B(n2829), .Z(n3000) );
  AND U3755 ( .A(y[181]), .B(x[32]), .Z(n2831) );
  AND U3756 ( .A(y[180]), .B(x[33]), .Z(n2830) );
  XOR U3757 ( .A(n2831), .B(n2830), .Z(n2999) );
  XOR U3758 ( .A(n3000), .B(n2999), .Z(n3010) );
  AND U3759 ( .A(x[8]), .B(y[61]), .Z(n3018) );
  AND U3760 ( .A(x[1]), .B(y[20]), .Z(n3017) );
  XOR U3761 ( .A(n3018), .B(n3017), .Z(n3020) );
  AND U3762 ( .A(x[12]), .B(y[57]), .Z(n3019) );
  XOR U3763 ( .A(n3020), .B(n3019), .Z(n3009) );
  XOR U3764 ( .A(n3010), .B(n3009), .Z(n3012) );
  XOR U3765 ( .A(n3011), .B(n3012), .Z(n2916) );
  XOR U3766 ( .A(n2917), .B(n2916), .Z(n2955) );
  XOR U3767 ( .A(n2956), .B(n2955), .Z(n2908) );
  AND U3768 ( .A(x[36]), .B(y[179]), .Z(n3092) );
  NAND U3769 ( .A(n3092), .B(n2832), .Z(n2836) );
  NAND U3770 ( .A(n2834), .B(n2833), .Z(n2835) );
  NAND U3771 ( .A(n2836), .B(n2835), .Z(n2971) );
  XOR U3772 ( .A(n2971), .B(n2972), .Z(n2974) );
  NAND U3773 ( .A(n2840), .B(n2839), .Z(n2844) );
  NANDN U3774 ( .A(n2842), .B(n2841), .Z(n2843) );
  AND U3775 ( .A(n2844), .B(n2843), .Z(n2964) );
  AND U3776 ( .A(x[11]), .B(y[58]), .Z(n3150) );
  NAND U3777 ( .A(y[59]), .B(x[10]), .Z(n2845) );
  XNOR U3778 ( .A(n3150), .B(n2845), .Z(n2930) );
  AND U3779 ( .A(x[9]), .B(y[60]), .Z(n2929) );
  XOR U3780 ( .A(n2930), .B(n2929), .Z(n2962) );
  AND U3781 ( .A(x[34]), .B(y[179]), .Z(n2925) );
  AND U3782 ( .A(x[37]), .B(y[176]), .Z(n2924) );
  XOR U3783 ( .A(n2925), .B(n2924), .Z(n2927) );
  NAND U3784 ( .A(y[177]), .B(x[36]), .Z(n2846) );
  XNOR U3785 ( .A(n2847), .B(n2846), .Z(n2926) );
  XOR U3786 ( .A(n2927), .B(n2926), .Z(n2961) );
  XOR U3787 ( .A(n2962), .B(n2961), .Z(n2963) );
  XOR U3788 ( .A(n2964), .B(n2963), .Z(n2973) );
  XOR U3789 ( .A(n2974), .B(n2973), .Z(n2982) );
  AND U3790 ( .A(y[96]), .B(x[21]), .Z(n2849) );
  AND U3791 ( .A(y[97]), .B(x[20]), .Z(n2848) );
  XOR U3792 ( .A(n2849), .B(n2848), .Z(n2936) );
  XOR U3793 ( .A(n2937), .B(n2936), .Z(n3004) );
  AND U3794 ( .A(x[29]), .B(y[136]), .Z(n2932) );
  AND U3795 ( .A(x[3]), .B(y[18]), .Z(n2931) );
  XOR U3796 ( .A(n2932), .B(n2931), .Z(n2934) );
  AND U3797 ( .A(x[2]), .B(y[19]), .Z(n2933) );
  XOR U3798 ( .A(n2934), .B(n2933), .Z(n3003) );
  XOR U3799 ( .A(n3004), .B(n3003), .Z(n3006) );
  NAND U3800 ( .A(n2851), .B(n2850), .Z(n2855) );
  NANDN U3801 ( .A(n2853), .B(n2852), .Z(n2854) );
  AND U3802 ( .A(n2855), .B(n2854), .Z(n3005) );
  XOR U3803 ( .A(n3006), .B(n3005), .Z(n2980) );
  AND U3804 ( .A(x[11]), .B(y[60]), .Z(n3125) );
  NAND U3805 ( .A(n3125), .B(n2856), .Z(n2859) );
  NANDN U3806 ( .A(n2857), .B(n2928), .Z(n2858) );
  NAND U3807 ( .A(n2859), .B(n2858), .Z(n2967) );
  AND U3808 ( .A(x[17]), .B(y[100]), .Z(n3207) );
  AND U3809 ( .A(x[27]), .B(y[138]), .Z(n2985) );
  XOR U3810 ( .A(n3207), .B(n2985), .Z(n2987) );
  AND U3811 ( .A(x[16]), .B(y[101]), .Z(n2986) );
  XOR U3812 ( .A(n2987), .B(n2986), .Z(n2966) );
  AND U3813 ( .A(x[0]), .B(y[21]), .Z(n2991) );
  AND U3814 ( .A(x[25]), .B(y[140]), .Z(n2990) );
  XOR U3815 ( .A(n2991), .B(n2990), .Z(n2993) );
  AND U3816 ( .A(x[26]), .B(y[139]), .Z(n2992) );
  XOR U3817 ( .A(n2993), .B(n2992), .Z(n2965) );
  XNOR U3818 ( .A(n2966), .B(n2965), .Z(n2968) );
  XOR U3819 ( .A(n2967), .B(n2968), .Z(n2979) );
  XNOR U3820 ( .A(n2980), .B(n2979), .Z(n2981) );
  XOR U3821 ( .A(n2982), .B(n2981), .Z(n2907) );
  NANDN U3822 ( .A(n2861), .B(n2860), .Z(n2865) );
  NAND U3823 ( .A(n2863), .B(n2862), .Z(n2864) );
  NAND U3824 ( .A(n2865), .B(n2864), .Z(n2975) );
  NANDN U3825 ( .A(n2867), .B(n2866), .Z(n2871) );
  NANDN U3826 ( .A(n2869), .B(n2868), .Z(n2870) );
  NAND U3827 ( .A(n2871), .B(n2870), .Z(n2976) );
  XOR U3828 ( .A(n2975), .B(n2976), .Z(n2978) );
  NANDN U3829 ( .A(n2873), .B(n2872), .Z(n2877) );
  NANDN U3830 ( .A(n2875), .B(n2874), .Z(n2876) );
  AND U3831 ( .A(n2877), .B(n2876), .Z(n2977) );
  XOR U3832 ( .A(n2978), .B(n2977), .Z(n2906) );
  XNOR U3833 ( .A(n2907), .B(n2906), .Z(n2909) );
  XNOR U3834 ( .A(n2908), .B(n2909), .Z(n2902) );
  XNOR U3835 ( .A(n2903), .B(n2902), .Z(n2905) );
  IV U3836 ( .A(n2882), .Z(n2884) );
  NANDN U3837 ( .A(n2884), .B(n2883), .Z(n2888) );
  NAND U3838 ( .A(n2886), .B(n2885), .Z(n2887) );
  NAND U3839 ( .A(n2888), .B(n2887), .Z(n2910) );
  IV U3840 ( .A(n2889), .Z(n2891) );
  NANDN U3841 ( .A(n2891), .B(n2890), .Z(n2895) );
  NAND U3842 ( .A(n2893), .B(n2892), .Z(n2894) );
  AND U3843 ( .A(n2895), .B(n2894), .Z(n2911) );
  XOR U3844 ( .A(n2910), .B(n2911), .Z(n2913) );
  XOR U3845 ( .A(n2912), .B(n2913), .Z(n2904) );
  XOR U3846 ( .A(n2905), .B(n2904), .Z(n2898) );
  XOR U3847 ( .A(n2899), .B(n2898), .Z(o[21]) );
  NANDN U3848 ( .A(n2897), .B(n2896), .Z(n2901) );
  NAND U3849 ( .A(n2899), .B(n2898), .Z(n2900) );
  NAND U3850 ( .A(n2901), .B(n2900), .Z(n3318) );
  XOR U3851 ( .A(n3308), .B(n3307), .Z(n3306) );
  NAND U3852 ( .A(n2915), .B(n2914), .Z(n2919) );
  NAND U3853 ( .A(n2917), .B(n2916), .Z(n2918) );
  AND U3854 ( .A(n2919), .B(n2918), .Z(n3314) );
  AND U3855 ( .A(x[27]), .B(y[139]), .Z(n3198) );
  AND U3856 ( .A(x[19]), .B(y[99]), .Z(n3197) );
  XOR U3857 ( .A(n3198), .B(n3197), .Z(n3196) );
  AND U3858 ( .A(x[3]), .B(y[19]), .Z(n3195) );
  XOR U3859 ( .A(n3196), .B(n3195), .Z(n3273) );
  AND U3860 ( .A(x[26]), .B(y[140]), .Z(n3237) );
  AND U3861 ( .A(x[20]), .B(y[98]), .Z(n3236) );
  XOR U3862 ( .A(n3237), .B(n3236), .Z(n3235) );
  AND U3863 ( .A(x[2]), .B(y[20]), .Z(n3234) );
  XNOR U3864 ( .A(n3235), .B(n3234), .Z(n3272) );
  XNOR U3865 ( .A(n3270), .B(n3271), .Z(n3180) );
  XOR U3866 ( .A(n3177), .B(n3178), .Z(n3035) );
  XOR U3867 ( .A(n3034), .B(n3035), .Z(n3032) );
  AND U3868 ( .A(x[21]), .B(y[97]), .Z(n3145) );
  AND U3869 ( .A(y[17]), .B(x[5]), .Z(n2939) );
  NAND U3870 ( .A(y[18]), .B(x[4]), .Z(n2938) );
  XNOR U3871 ( .A(n2939), .B(n2938), .Z(n3162) );
  AND U3872 ( .A(x[30]), .B(y[136]), .Z(n3161) );
  XOR U3873 ( .A(n3162), .B(n3161), .Z(n3267) );
  AND U3874 ( .A(x[33]), .B(y[181]), .Z(n3156) );
  AND U3875 ( .A(x[36]), .B(y[178]), .Z(n2941) );
  AND U3876 ( .A(n2941), .B(n2940), .Z(n3158) );
  AND U3877 ( .A(x[34]), .B(y[180]), .Z(n3157) );
  XOR U3878 ( .A(n3158), .B(n3157), .Z(n3155) );
  XNOR U3879 ( .A(n3156), .B(n3155), .Z(n3266) );
  XOR U3880 ( .A(n3264), .B(n3265), .Z(n3057) );
  NAND U3881 ( .A(n2943), .B(n2942), .Z(n2946) );
  NAND U3882 ( .A(n3164), .B(n2944), .Z(n2945) );
  NAND U3883 ( .A(n2946), .B(n2945), .Z(n3060) );
  NAND U3884 ( .A(n2948), .B(n2947), .Z(n2951) );
  NAND U3885 ( .A(n3245), .B(n2949), .Z(n2950) );
  NAND U3886 ( .A(n2951), .B(n2950), .Z(n3059) );
  XNOR U3887 ( .A(n3060), .B(n3059), .Z(n3058) );
  XNOR U3888 ( .A(n3032), .B(n3033), .Z(n3031) );
  IV U3889 ( .A(n3031), .Z(n2960) );
  IV U3890 ( .A(n2952), .Z(n2954) );
  NANDN U3891 ( .A(n2954), .B(n2953), .Z(n2959) );
  IV U3892 ( .A(n2955), .Z(n2957) );
  NANDN U3893 ( .A(n2957), .B(n2956), .Z(n2958) );
  AND U3894 ( .A(n2959), .B(n2958), .Z(n3030) );
  XOR U3895 ( .A(n2960), .B(n3030), .Z(n3029) );
  NAND U3896 ( .A(n2966), .B(n2965), .Z(n2970) );
  NANDN U3897 ( .A(n2968), .B(n2967), .Z(n2969) );
  AND U3898 ( .A(n2970), .B(n2969), .Z(n3052) );
  XOR U3899 ( .A(n3052), .B(n3051), .Z(n3049) );
  XOR U3900 ( .A(n3050), .B(n3049), .Z(n3028) );
  XOR U3901 ( .A(n3029), .B(n3028), .Z(n3313) );
  XOR U3902 ( .A(n3314), .B(n3313), .Z(n3312) );
  NANDN U3903 ( .A(n2980), .B(n2979), .Z(n2984) );
  NANDN U3904 ( .A(n2982), .B(n2981), .Z(n2983) );
  NAND U3905 ( .A(n2984), .B(n2983), .Z(n3292) );
  AND U3906 ( .A(n3207), .B(n2985), .Z(n2989) );
  NAND U3907 ( .A(n2987), .B(n2986), .Z(n2988) );
  NANDN U3908 ( .A(n2989), .B(n2988), .Z(n3042) );
  NAND U3909 ( .A(n2991), .B(n2990), .Z(n2995) );
  NAND U3910 ( .A(n2993), .B(n2992), .Z(n2994) );
  AND U3911 ( .A(n2995), .B(n2994), .Z(n3183) );
  AND U3912 ( .A(x[1]), .B(y[21]), .Z(n3231) );
  AND U3913 ( .A(x[14]), .B(y[56]), .Z(n3230) );
  XOR U3914 ( .A(n3231), .B(n3230), .Z(n3229) );
  AND U3915 ( .A(x[8]), .B(y[62]), .Z(n3228) );
  XOR U3916 ( .A(n3229), .B(n3228), .Z(n3186) );
  AND U3917 ( .A(y[177]), .B(x[37]), .Z(n2997) );
  NAND U3918 ( .A(y[178]), .B(x[36]), .Z(n2996) );
  XNOR U3919 ( .A(n2997), .B(n2996), .Z(n3072) );
  AND U3920 ( .A(x[38]), .B(y[176]), .Z(n3071) );
  XOR U3921 ( .A(n3072), .B(n3071), .Z(n3069) );
  XNOR U3922 ( .A(n3070), .B(n3069), .Z(n3185) );
  XNOR U3923 ( .A(n3183), .B(n3184), .Z(n3046) );
  NANDN U3924 ( .A(n2998), .B(n3156), .Z(n3002) );
  NAND U3925 ( .A(n3000), .B(n2999), .Z(n3001) );
  NAND U3926 ( .A(n3002), .B(n3001), .Z(n3045) );
  XOR U3927 ( .A(n3042), .B(n3043), .Z(n3297) );
  NAND U3928 ( .A(n3004), .B(n3003), .Z(n3008) );
  NAND U3929 ( .A(n3006), .B(n3005), .Z(n3007) );
  AND U3930 ( .A(n3008), .B(n3007), .Z(n3299) );
  NAND U3931 ( .A(n3010), .B(n3009), .Z(n3014) );
  NAND U3932 ( .A(n3012), .B(n3011), .Z(n3013) );
  AND U3933 ( .A(n3014), .B(n3013), .Z(n3036) );
  AND U3934 ( .A(x[16]), .B(y[102]), .Z(n3192) );
  AND U3935 ( .A(x[6]), .B(y[16]), .Z(n3191) );
  XOR U3936 ( .A(n3192), .B(n3191), .Z(n3190) );
  AND U3937 ( .A(x[29]), .B(y[137]), .Z(n3189) );
  XOR U3938 ( .A(n3190), .B(n3189), .Z(n3066) );
  AND U3939 ( .A(x[13]), .B(y[57]), .Z(n3251) );
  AND U3940 ( .A(x[10]), .B(y[60]), .Z(n3250) );
  XOR U3941 ( .A(n3251), .B(n3250), .Z(n3249) );
  AND U3942 ( .A(x[9]), .B(y[61]), .Z(n3248) );
  XOR U3943 ( .A(n3249), .B(n3248), .Z(n3149) );
  AND U3944 ( .A(y[58]), .B(x[12]), .Z(n3016) );
  NAND U3945 ( .A(y[59]), .B(x[11]), .Z(n3015) );
  XNOR U3946 ( .A(n3016), .B(n3015), .Z(n3148) );
  XOR U3947 ( .A(n3149), .B(n3148), .Z(n3065) );
  XOR U3948 ( .A(n3066), .B(n3065), .Z(n3064) );
  AND U3949 ( .A(x[32]), .B(y[182]), .Z(n3144) );
  XOR U3950 ( .A(n3145), .B(n3144), .Z(n3143) );
  AND U3951 ( .A(x[22]), .B(y[96]), .Z(n3142) );
  XOR U3952 ( .A(n3143), .B(n3142), .Z(n3063) );
  XOR U3953 ( .A(n3064), .B(n3063), .Z(n3039) );
  NAND U3954 ( .A(n3018), .B(n3017), .Z(n3022) );
  NAND U3955 ( .A(n3020), .B(n3019), .Z(n3021) );
  AND U3956 ( .A(n3022), .B(n3021), .Z(n3137) );
  AND U3957 ( .A(y[100]), .B(x[18]), .Z(n3024) );
  NAND U3958 ( .A(y[101]), .B(x[17]), .Z(n3023) );
  XNOR U3959 ( .A(n3024), .B(n3023), .Z(n3206) );
  AND U3960 ( .A(x[28]), .B(y[138]), .Z(n3205) );
  XOR U3961 ( .A(n3206), .B(n3205), .Z(n3139) );
  AND U3962 ( .A(y[142]), .B(x[24]), .Z(n3026) );
  NAND U3963 ( .A(y[141]), .B(x[25]), .Z(n3025) );
  XNOR U3964 ( .A(n3026), .B(n3025), .Z(n3243) );
  AND U3965 ( .A(x[0]), .B(y[22]), .Z(n3242) );
  XNOR U3966 ( .A(n3243), .B(n3242), .Z(n3138) );
  XOR U3967 ( .A(n3137), .B(n3136), .Z(n3038) );
  XNOR U3968 ( .A(n3036), .B(n3037), .Z(n3298) );
  XOR U3969 ( .A(n3299), .B(n3298), .Z(n3296) );
  XOR U3970 ( .A(n3292), .B(n3293), .Z(n3291) );
  XNOR U3971 ( .A(n3290), .B(n3291), .Z(n3311) );
  XOR U3972 ( .A(n3312), .B(n3311), .Z(n3305) );
  XOR U3973 ( .A(n3306), .B(n3305), .Z(n3319) );
  XOR U3974 ( .A(n3317), .B(n3319), .Z(n3027) );
  XNOR U3975 ( .A(n3318), .B(n3027), .Z(o[22]) );
  NANDN U3976 ( .A(n3037), .B(n3036), .Z(n3041) );
  NANDN U3977 ( .A(n3039), .B(n3038), .Z(n3040) );
  AND U3978 ( .A(n3041), .B(n3040), .Z(n3289) );
  IV U3979 ( .A(n3042), .Z(n3044) );
  NANDN U3980 ( .A(n3044), .B(n3043), .Z(n3048) );
  NANDN U3981 ( .A(n3046), .B(n3045), .Z(n3047) );
  AND U3982 ( .A(n3048), .B(n3047), .Z(n3056) );
  NAND U3983 ( .A(n3050), .B(n3049), .Z(n3054) );
  NAND U3984 ( .A(n3052), .B(n3051), .Z(n3053) );
  NAND U3985 ( .A(n3054), .B(n3053), .Z(n3055) );
  XNOR U3986 ( .A(n3056), .B(n3055), .Z(n3287) );
  NANDN U3987 ( .A(n3058), .B(n3057), .Z(n3062) );
  NAND U3988 ( .A(n3060), .B(n3059), .Z(n3061) );
  AND U3989 ( .A(n3062), .B(n3061), .Z(n3285) );
  NAND U3990 ( .A(n3064), .B(n3063), .Z(n3068) );
  NAND U3991 ( .A(n3066), .B(n3065), .Z(n3067) );
  AND U3992 ( .A(n3068), .B(n3067), .Z(n3176) );
  NAND U3993 ( .A(n3070), .B(n3069), .Z(n3074) );
  NAND U3994 ( .A(n3072), .B(n3071), .Z(n3073) );
  AND U3995 ( .A(n3074), .B(n3073), .Z(n3135) );
  AND U3996 ( .A(y[177]), .B(x[38]), .Z(n3076) );
  NAND U3997 ( .A(y[19]), .B(x[4]), .Z(n3075) );
  XNOR U3998 ( .A(n3076), .B(n3075), .Z(n3080) );
  AND U3999 ( .A(y[176]), .B(x[39]), .Z(n3078) );
  NAND U4000 ( .A(y[103]), .B(x[16]), .Z(n3077) );
  XNOR U4001 ( .A(n3078), .B(n3077), .Z(n3079) );
  XOR U4002 ( .A(n3080), .B(n3079), .Z(n3088) );
  AND U4003 ( .A(y[138]), .B(x[29]), .Z(n3082) );
  NAND U4004 ( .A(y[98]), .B(x[21]), .Z(n3081) );
  XNOR U4005 ( .A(n3082), .B(n3081), .Z(n3086) );
  AND U4006 ( .A(y[180]), .B(x[35]), .Z(n3084) );
  NAND U4007 ( .A(y[181]), .B(x[34]), .Z(n3083) );
  XNOR U4008 ( .A(n3084), .B(n3083), .Z(n3085) );
  XNOR U4009 ( .A(n3086), .B(n3085), .Z(n3087) );
  XNOR U4010 ( .A(n3088), .B(n3087), .Z(n3133) );
  AND U4011 ( .A(y[140]), .B(x[27]), .Z(n3094) );
  AND U4012 ( .A(y[136]), .B(x[31]), .Z(n3090) );
  NAND U4013 ( .A(y[63]), .B(x[8]), .Z(n3089) );
  XNOR U4014 ( .A(n3090), .B(n3089), .Z(n3091) );
  XNOR U4015 ( .A(n3092), .B(n3091), .Z(n3093) );
  XNOR U4016 ( .A(n3094), .B(n3093), .Z(n3110) );
  AND U4017 ( .A(y[22]), .B(x[1]), .Z(n3096) );
  NAND U4018 ( .A(y[182]), .B(x[33]), .Z(n3095) );
  XNOR U4019 ( .A(n3096), .B(n3095), .Z(n3100) );
  AND U4020 ( .A(y[96]), .B(x[23]), .Z(n3098) );
  NAND U4021 ( .A(y[23]), .B(x[0]), .Z(n3097) );
  XNOR U4022 ( .A(n3098), .B(n3097), .Z(n3099) );
  XOR U4023 ( .A(n3100), .B(n3099), .Z(n3108) );
  AND U4024 ( .A(y[100]), .B(x[19]), .Z(n3102) );
  NAND U4025 ( .A(y[183]), .B(x[32]), .Z(n3101) );
  XNOR U4026 ( .A(n3102), .B(n3101), .Z(n3106) );
  AND U4027 ( .A(y[102]), .B(x[17]), .Z(n3104) );
  NAND U4028 ( .A(y[99]), .B(x[20]), .Z(n3103) );
  XNOR U4029 ( .A(n3104), .B(n3103), .Z(n3105) );
  XNOR U4030 ( .A(n3106), .B(n3105), .Z(n3107) );
  XNOR U4031 ( .A(n3108), .B(n3107), .Z(n3109) );
  XOR U4032 ( .A(n3110), .B(n3109), .Z(n3131) );
  AND U4033 ( .A(y[16]), .B(x[7]), .Z(n3112) );
  NAND U4034 ( .A(y[139]), .B(x[28]), .Z(n3111) );
  XNOR U4035 ( .A(n3112), .B(n3111), .Z(n3116) );
  AND U4036 ( .A(y[97]), .B(x[22]), .Z(n3114) );
  NAND U4037 ( .A(y[17]), .B(x[6]), .Z(n3113) );
  XNOR U4038 ( .A(n3114), .B(n3113), .Z(n3115) );
  XOR U4039 ( .A(n3116), .B(n3115), .Z(n3124) );
  AND U4040 ( .A(y[137]), .B(x[30]), .Z(n3118) );
  NAND U4041 ( .A(y[21]), .B(x[2]), .Z(n3117) );
  XNOR U4042 ( .A(n3118), .B(n3117), .Z(n3122) );
  AND U4043 ( .A(y[57]), .B(x[14]), .Z(n3120) );
  NAND U4044 ( .A(y[20]), .B(x[3]), .Z(n3119) );
  XNOR U4045 ( .A(n3120), .B(n3119), .Z(n3121) );
  XNOR U4046 ( .A(n3122), .B(n3121), .Z(n3123) );
  XNOR U4047 ( .A(n3124), .B(n3123), .Z(n3129) );
  AND U4048 ( .A(x[37]), .B(y[178]), .Z(n3220) );
  AND U4049 ( .A(x[25]), .B(y[142]), .Z(n3244) );
  XOR U4050 ( .A(n3220), .B(n3244), .Z(n3127) );
  AND U4051 ( .A(x[5]), .B(y[18]), .Z(n3163) );
  XNOR U4052 ( .A(n3163), .B(n3125), .Z(n3126) );
  XNOR U4053 ( .A(n3127), .B(n3126), .Z(n3128) );
  XNOR U4054 ( .A(n3129), .B(n3128), .Z(n3130) );
  XNOR U4055 ( .A(n3131), .B(n3130), .Z(n3132) );
  XNOR U4056 ( .A(n3133), .B(n3132), .Z(n3134) );
  XNOR U4057 ( .A(n3135), .B(n3134), .Z(n3174) );
  NAND U4058 ( .A(n3137), .B(n3136), .Z(n3141) );
  NANDN U4059 ( .A(n3139), .B(n3138), .Z(n3140) );
  AND U4060 ( .A(n3141), .B(n3140), .Z(n3172) );
  NAND U4061 ( .A(n3143), .B(n3142), .Z(n3147) );
  NAND U4062 ( .A(n3145), .B(n3144), .Z(n3146) );
  AND U4063 ( .A(n3147), .B(n3146), .Z(n3154) );
  NAND U4064 ( .A(n3149), .B(n3148), .Z(n3152) );
  AND U4065 ( .A(x[12]), .B(y[59]), .Z(n3222) );
  NAND U4066 ( .A(n3150), .B(n3222), .Z(n3151) );
  NAND U4067 ( .A(n3152), .B(n3151), .Z(n3153) );
  XNOR U4068 ( .A(n3154), .B(n3153), .Z(n3170) );
  NAND U4069 ( .A(n3156), .B(n3155), .Z(n3160) );
  NAND U4070 ( .A(n3158), .B(n3157), .Z(n3159) );
  AND U4071 ( .A(n3160), .B(n3159), .Z(n3168) );
  NAND U4072 ( .A(n3162), .B(n3161), .Z(n3166) );
  NAND U4073 ( .A(n3164), .B(n3163), .Z(n3165) );
  NAND U4074 ( .A(n3166), .B(n3165), .Z(n3167) );
  XNOR U4075 ( .A(n3168), .B(n3167), .Z(n3169) );
  XNOR U4076 ( .A(n3170), .B(n3169), .Z(n3171) );
  XNOR U4077 ( .A(n3172), .B(n3171), .Z(n3173) );
  XNOR U4078 ( .A(n3174), .B(n3173), .Z(n3175) );
  XNOR U4079 ( .A(n3176), .B(n3175), .Z(n3283) );
  NAND U4080 ( .A(n3178), .B(n3177), .Z(n3182) );
  NANDN U4081 ( .A(n3180), .B(n3179), .Z(n3181) );
  AND U4082 ( .A(n3182), .B(n3181), .Z(n3281) );
  NANDN U4083 ( .A(n3184), .B(n3183), .Z(n3188) );
  NANDN U4084 ( .A(n3186), .B(n3185), .Z(n3187) );
  AND U4085 ( .A(n3188), .B(n3187), .Z(n3263) );
  NAND U4086 ( .A(n3190), .B(n3189), .Z(n3194) );
  NAND U4087 ( .A(n3192), .B(n3191), .Z(n3193) );
  AND U4088 ( .A(n3194), .B(n3193), .Z(n3202) );
  NAND U4089 ( .A(n3196), .B(n3195), .Z(n3200) );
  NAND U4090 ( .A(n3198), .B(n3197), .Z(n3199) );
  NAND U4091 ( .A(n3200), .B(n3199), .Z(n3201) );
  XNOR U4092 ( .A(n3202), .B(n3201), .Z(n3261) );
  AND U4093 ( .A(y[56]), .B(x[15]), .Z(n3204) );
  NAND U4094 ( .A(y[141]), .B(x[26]), .Z(n3203) );
  XNOR U4095 ( .A(n3204), .B(n3203), .Z(n3227) );
  AND U4096 ( .A(x[18]), .B(y[101]), .Z(n3219) );
  NAND U4097 ( .A(n3206), .B(n3205), .Z(n3209) );
  NAND U4098 ( .A(n3207), .B(n3219), .Z(n3208) );
  AND U4099 ( .A(n3209), .B(n3208), .Z(n3217) );
  AND U4100 ( .A(y[58]), .B(x[13]), .Z(n3211) );
  NAND U4101 ( .A(y[61]), .B(x[10]), .Z(n3210) );
  XNOR U4102 ( .A(n3211), .B(n3210), .Z(n3215) );
  AND U4103 ( .A(y[143]), .B(x[24]), .Z(n3213) );
  NAND U4104 ( .A(y[62]), .B(x[9]), .Z(n3212) );
  XNOR U4105 ( .A(n3213), .B(n3212), .Z(n3214) );
  XNOR U4106 ( .A(n3215), .B(n3214), .Z(n3216) );
  XNOR U4107 ( .A(n3217), .B(n3216), .Z(n3218) );
  XOR U4108 ( .A(n3219), .B(n3218), .Z(n3225) );
  AND U4109 ( .A(x[36]), .B(y[177]), .Z(n3221) );
  AND U4110 ( .A(n3221), .B(n3220), .Z(n3223) );
  XNOR U4111 ( .A(n3223), .B(n3222), .Z(n3224) );
  XNOR U4112 ( .A(n3225), .B(n3224), .Z(n3226) );
  XOR U4113 ( .A(n3227), .B(n3226), .Z(n3259) );
  NAND U4114 ( .A(n3229), .B(n3228), .Z(n3233) );
  NAND U4115 ( .A(n3231), .B(n3230), .Z(n3232) );
  AND U4116 ( .A(n3233), .B(n3232), .Z(n3241) );
  NAND U4117 ( .A(n3235), .B(n3234), .Z(n3239) );
  NAND U4118 ( .A(n3237), .B(n3236), .Z(n3238) );
  NAND U4119 ( .A(n3239), .B(n3238), .Z(n3240) );
  XNOR U4120 ( .A(n3241), .B(n3240), .Z(n3257) );
  NAND U4121 ( .A(n3243), .B(n3242), .Z(n3247) );
  NAND U4122 ( .A(n3245), .B(n3244), .Z(n3246) );
  AND U4123 ( .A(n3247), .B(n3246), .Z(n3255) );
  NAND U4124 ( .A(n3249), .B(n3248), .Z(n3253) );
  NAND U4125 ( .A(n3251), .B(n3250), .Z(n3252) );
  NAND U4126 ( .A(n3253), .B(n3252), .Z(n3254) );
  XNOR U4127 ( .A(n3255), .B(n3254), .Z(n3256) );
  XNOR U4128 ( .A(n3257), .B(n3256), .Z(n3258) );
  XNOR U4129 ( .A(n3259), .B(n3258), .Z(n3260) );
  XNOR U4130 ( .A(n3261), .B(n3260), .Z(n3262) );
  XNOR U4131 ( .A(n3263), .B(n3262), .Z(n3279) );
  NANDN U4132 ( .A(n3265), .B(n3264), .Z(n3269) );
  NANDN U4133 ( .A(n3267), .B(n3266), .Z(n3268) );
  AND U4134 ( .A(n3269), .B(n3268), .Z(n3277) );
  NANDN U4135 ( .A(n3271), .B(n3270), .Z(n3275) );
  NANDN U4136 ( .A(n3273), .B(n3272), .Z(n3274) );
  NAND U4137 ( .A(n3275), .B(n3274), .Z(n3276) );
  XNOR U4138 ( .A(n3277), .B(n3276), .Z(n3278) );
  XNOR U4139 ( .A(n3279), .B(n3278), .Z(n3280) );
  XNOR U4140 ( .A(n3281), .B(n3280), .Z(n3282) );
  XNOR U4141 ( .A(n3283), .B(n3282), .Z(n3284) );
  XNOR U4142 ( .A(n3285), .B(n3284), .Z(n3286) );
  XNOR U4143 ( .A(n3287), .B(n3286), .Z(n3288) );
  NANDN U4144 ( .A(n3291), .B(n3290), .Z(n3295) );
  NANDN U4145 ( .A(n3293), .B(n3292), .Z(n3294) );
  AND U4146 ( .A(n3295), .B(n3294), .Z(n3303) );
  NANDN U4147 ( .A(n3297), .B(n3296), .Z(n3301) );
  NAND U4148 ( .A(n3299), .B(n3298), .Z(n3300) );
  NAND U4149 ( .A(n3301), .B(n3300), .Z(n3302) );
  XNOR U4150 ( .A(n3303), .B(n3302), .Z(n3304) );
  NAND U4151 ( .A(n3308), .B(n3307), .Z(n3309) );
  NAND U4152 ( .A(n3312), .B(n3311), .Z(n3316) );
  NAND U4153 ( .A(n3314), .B(n3313), .Z(n3315) );
  NAND U4154 ( .A(x[32]), .B(y[184]), .Z(n3458) );
  NAND U4155 ( .A(x[8]), .B(y[64]), .Z(n3322) );
  XOR U4156 ( .A(n3458), .B(n3322), .Z(n3323) );
  AND U4157 ( .A(x[0]), .B(y[24]), .Z(n3330) );
  AND U4158 ( .A(x[16]), .B(y[104]), .Z(n3327) );
  XOR U4159 ( .A(n3330), .B(n3327), .Z(n3326) );
  AND U4160 ( .A(x[24]), .B(y[144]), .Z(n3325) );
  XNOR U4161 ( .A(n3326), .B(n3325), .Z(n3324) );
  XNOR U4162 ( .A(n3323), .B(n3324), .Z(o[24]) );
  AND U4163 ( .A(y[24]), .B(x[1]), .Z(n3321) );
  NAND U4164 ( .A(y[25]), .B(x[0]), .Z(n3320) );
  XNOR U4165 ( .A(n3321), .B(n3320), .Z(n3332) );
  AND U4166 ( .A(x[9]), .B(y[64]), .Z(n3331) );
  XOR U4167 ( .A(n3332), .B(n3331), .Z(n3349) );
  AND U4168 ( .A(x[33]), .B(y[184]), .Z(n3561) );
  NAND U4169 ( .A(x[16]), .B(y[105]), .Z(n3335) );
  XNOR U4170 ( .A(n3561), .B(n3335), .Z(n3337) );
  AND U4171 ( .A(x[32]), .B(y[185]), .Z(n3360) );
  NAND U4172 ( .A(x[17]), .B(y[104]), .Z(n3359) );
  XNOR U4173 ( .A(n3360), .B(n3359), .Z(n3336) );
  XOR U4174 ( .A(n3337), .B(n3336), .Z(n3347) );
  AND U4175 ( .A(x[8]), .B(y[65]), .Z(n3584) );
  AND U4176 ( .A(x[24]), .B(y[145]), .Z(n3352) );
  XOR U4177 ( .A(n3584), .B(n3352), .Z(n3354) );
  AND U4178 ( .A(x[25]), .B(y[144]), .Z(n3353) );
  XNOR U4179 ( .A(n3354), .B(n3353), .Z(n3346) );
  XNOR U4180 ( .A(n3347), .B(n3346), .Z(n3348) );
  XNOR U4181 ( .A(n3349), .B(n3348), .Z(n3343) );
  NAND U4182 ( .A(n3326), .B(n3325), .Z(n3329) );
  AND U4183 ( .A(n3330), .B(n3327), .Z(n3328) );
  ANDN U4184 ( .B(n3329), .A(n3328), .Z(n3340) );
  XNOR U4185 ( .A(n3341), .B(n3340), .Z(n3342) );
  XNOR U4186 ( .A(n3343), .B(n3342), .Z(o[25]) );
  NAND U4187 ( .A(x[1]), .B(y[25]), .Z(n3382) );
  NANDN U4188 ( .A(n3382), .B(n3330), .Z(n3334) );
  NAND U4189 ( .A(n3332), .B(n3331), .Z(n3333) );
  AND U4190 ( .A(n3334), .B(n3333), .Z(n3402) );
  NANDN U4191 ( .A(n3335), .B(n3561), .Z(n3339) );
  NAND U4192 ( .A(n3337), .B(n3336), .Z(n3338) );
  AND U4193 ( .A(n3339), .B(n3338), .Z(n3401) );
  AND U4194 ( .A(x[24]), .B(y[146]), .Z(n3406) );
  NAND U4195 ( .A(x[0]), .B(y[26]), .Z(n3407) );
  XNOR U4196 ( .A(n3406), .B(n3407), .Z(n3408) );
  NAND U4197 ( .A(x[10]), .B(y[64]), .Z(n3409) );
  XNOR U4198 ( .A(n3408), .B(n3409), .Z(n3400) );
  XOR U4199 ( .A(n3401), .B(n3400), .Z(n3403) );
  XOR U4200 ( .A(n3402), .B(n3403), .Z(n3362) );
  NANDN U4201 ( .A(n3341), .B(n3340), .Z(n3345) );
  NAND U4202 ( .A(n3343), .B(n3342), .Z(n3344) );
  NAND U4203 ( .A(n3345), .B(n3344), .Z(n3361) );
  XNOR U4204 ( .A(n3362), .B(n3361), .Z(n3364) );
  NANDN U4205 ( .A(n3347), .B(n3346), .Z(n3351) );
  NANDN U4206 ( .A(n3349), .B(n3348), .Z(n3350) );
  AND U4207 ( .A(n3351), .B(n3350), .Z(n3370) );
  AND U4208 ( .A(x[2]), .B(y[24]), .Z(n3379) );
  NAND U4209 ( .A(x[16]), .B(y[106]), .Z(n3380) );
  XNOR U4210 ( .A(n3379), .B(n3380), .Z(n3381) );
  NAND U4211 ( .A(x[26]), .B(y[144]), .Z(n3415) );
  XNOR U4212 ( .A(n3414), .B(n3415), .Z(n3416) );
  AND U4213 ( .A(x[18]), .B(y[104]), .Z(n3498) );
  AND U4214 ( .A(x[32]), .B(y[186]), .Z(n3392) );
  XOR U4215 ( .A(n3498), .B(n3392), .Z(n3394) );
  NAND U4216 ( .A(x[17]), .B(y[105]), .Z(n3393) );
  XOR U4217 ( .A(n3394), .B(n3393), .Z(n3417) );
  XNOR U4218 ( .A(n3416), .B(n3417), .Z(n3367) );
  NAND U4219 ( .A(n3584), .B(n3352), .Z(n3356) );
  AND U4220 ( .A(n3354), .B(n3353), .Z(n3355) );
  ANDN U4221 ( .B(n3356), .A(n3355), .Z(n3376) );
  AND U4222 ( .A(y[184]), .B(x[34]), .Z(n3358) );
  NAND U4223 ( .A(y[185]), .B(x[33]), .Z(n3357) );
  XNOR U4224 ( .A(n3358), .B(n3357), .Z(n3413) );
  ANDN U4225 ( .B(n3360), .A(n3359), .Z(n3412) );
  XOR U4226 ( .A(n3413), .B(n3412), .Z(n3373) );
  AND U4227 ( .A(x[25]), .B(y[145]), .Z(n3385) );
  NAND U4228 ( .A(x[9]), .B(y[65]), .Z(n3386) );
  XNOR U4229 ( .A(n3385), .B(n3386), .Z(n3387) );
  NAND U4230 ( .A(x[8]), .B(y[66]), .Z(n3388) );
  XOR U4231 ( .A(n3387), .B(n3388), .Z(n3374) );
  XNOR U4232 ( .A(n3373), .B(n3374), .Z(n3375) );
  XOR U4233 ( .A(n3376), .B(n3375), .Z(n3368) );
  XNOR U4234 ( .A(n3367), .B(n3368), .Z(n3369) );
  XNOR U4235 ( .A(n3370), .B(n3369), .Z(n3363) );
  XNOR U4236 ( .A(n3364), .B(n3363), .Z(o[26]) );
  NANDN U4237 ( .A(n3362), .B(n3361), .Z(n3366) );
  NAND U4238 ( .A(n3364), .B(n3363), .Z(n3365) );
  AND U4239 ( .A(n3366), .B(n3365), .Z(n3420) );
  NANDN U4240 ( .A(n3368), .B(n3367), .Z(n3372) );
  NAND U4241 ( .A(n3370), .B(n3369), .Z(n3371) );
  AND U4242 ( .A(n3372), .B(n3371), .Z(n3429) );
  NANDN U4243 ( .A(n3374), .B(n3373), .Z(n3378) );
  NANDN U4244 ( .A(n3376), .B(n3375), .Z(n3377) );
  AND U4245 ( .A(n3378), .B(n3377), .Z(n3427) );
  NANDN U4246 ( .A(n3380), .B(n3379), .Z(n3384) );
  NANDN U4247 ( .A(n3382), .B(n3381), .Z(n3383) );
  AND U4248 ( .A(n3384), .B(n3383), .Z(n3439) );
  NANDN U4249 ( .A(n3386), .B(n3385), .Z(n3390) );
  NANDN U4250 ( .A(n3388), .B(n3387), .Z(n3389) );
  AND U4251 ( .A(n3390), .B(n3389), .Z(n3479) );
  AND U4252 ( .A(x[24]), .B(y[147]), .Z(n3493) );
  AND U4253 ( .A(x[16]), .B(y[107]), .Z(n3492) );
  NAND U4254 ( .A(x[3]), .B(y[24]), .Z(n3491) );
  XOR U4255 ( .A(n3492), .B(n3491), .Z(n3494) );
  XOR U4256 ( .A(n3493), .B(n3494), .Z(n3477) );
  AND U4257 ( .A(x[18]), .B(y[105]), .Z(n3529) );
  NAND U4258 ( .A(y[104]), .B(x[19]), .Z(n3391) );
  XNOR U4259 ( .A(n3529), .B(n3391), .Z(n3499) );
  NAND U4260 ( .A(x[17]), .B(y[106]), .Z(n3500) );
  XNOR U4261 ( .A(n3477), .B(n3476), .Z(n3478) );
  XNOR U4262 ( .A(n3479), .B(n3478), .Z(n3438) );
  XNOR U4263 ( .A(n3439), .B(n3438), .Z(n3440) );
  NAND U4264 ( .A(n3498), .B(n3392), .Z(n3396) );
  ANDN U4265 ( .B(n3394), .A(n3393), .Z(n3395) );
  ANDN U4266 ( .B(n3396), .A(n3395), .Z(n3485) );
  AND U4267 ( .A(x[1]), .B(y[26]), .Z(n3454) );
  AND U4268 ( .A(x[2]), .B(y[25]), .Z(n3453) );
  NAND U4269 ( .A(x[25]), .B(y[146]), .Z(n3452) );
  XOR U4270 ( .A(n3453), .B(n3452), .Z(n3455) );
  XOR U4271 ( .A(n3454), .B(n3455), .Z(n3483) );
  AND U4272 ( .A(y[187]), .B(x[32]), .Z(n3398) );
  NAND U4273 ( .A(y[184]), .B(x[35]), .Z(n3397) );
  XNOR U4274 ( .A(n3398), .B(n3397), .Z(n3459) );
  AND U4275 ( .A(y[185]), .B(x[34]), .Z(n3546) );
  NAND U4276 ( .A(y[186]), .B(x[33]), .Z(n3399) );
  XOR U4277 ( .A(n3546), .B(n3399), .Z(n3460) );
  XNOR U4278 ( .A(n3459), .B(n3460), .Z(n3482) );
  XNOR U4279 ( .A(n3483), .B(n3482), .Z(n3484) );
  XOR U4280 ( .A(n3485), .B(n3484), .Z(n3441) );
  XNOR U4281 ( .A(n3440), .B(n3441), .Z(n3426) );
  XNOR U4282 ( .A(n3427), .B(n3426), .Z(n3428) );
  XOR U4283 ( .A(n3429), .B(n3428), .Z(n3421) );
  XNOR U4284 ( .A(n3420), .B(n3421), .Z(n3423) );
  NANDN U4285 ( .A(n3401), .B(n3400), .Z(n3405) );
  OR U4286 ( .A(n3403), .B(n3402), .Z(n3404) );
  AND U4287 ( .A(n3405), .B(n3404), .Z(n3435) );
  NANDN U4288 ( .A(n3407), .B(n3406), .Z(n3411) );
  NANDN U4289 ( .A(n3409), .B(n3408), .Z(n3410) );
  AND U4290 ( .A(n3411), .B(n3410), .Z(n3445) );
  XNOR U4291 ( .A(n3445), .B(n3444), .Z(n3447) );
  AND U4292 ( .A(x[11]), .B(y[64]), .Z(n3507) );
  AND U4293 ( .A(x[0]), .B(y[27]), .Z(n3506) );
  NAND U4294 ( .A(x[26]), .B(y[145]), .Z(n3505) );
  XOR U4295 ( .A(n3506), .B(n3505), .Z(n3508) );
  XOR U4296 ( .A(n3507), .B(n3508), .Z(n3473) );
  AND U4297 ( .A(x[8]), .B(y[67]), .Z(n3466) );
  AND U4298 ( .A(x[10]), .B(y[65]), .Z(n3465) );
  NAND U4299 ( .A(x[27]), .B(y[144]), .Z(n3464) );
  XOR U4300 ( .A(n3465), .B(n3464), .Z(n3467) );
  XOR U4301 ( .A(n3466), .B(n3467), .Z(n3471) );
  AND U4302 ( .A(x[9]), .B(y[66]), .Z(n3470) );
  XOR U4303 ( .A(n3447), .B(n3446), .Z(n3433) );
  NANDN U4304 ( .A(n3415), .B(n3414), .Z(n3419) );
  NANDN U4305 ( .A(n3417), .B(n3416), .Z(n3418) );
  AND U4306 ( .A(n3419), .B(n3418), .Z(n3432) );
  XNOR U4307 ( .A(n3433), .B(n3432), .Z(n3434) );
  XNOR U4308 ( .A(n3435), .B(n3434), .Z(n3422) );
  XOR U4309 ( .A(n3423), .B(n3422), .Z(o[27]) );
  NANDN U4310 ( .A(n3421), .B(n3420), .Z(n3425) );
  NAND U4311 ( .A(n3423), .B(n3422), .Z(n3424) );
  AND U4312 ( .A(n3425), .B(n3424), .Z(n3517) );
  NANDN U4313 ( .A(n3427), .B(n3426), .Z(n3431) );
  NANDN U4314 ( .A(n3429), .B(n3428), .Z(n3430) );
  AND U4315 ( .A(n3431), .B(n3430), .Z(n3513) );
  NANDN U4316 ( .A(n3433), .B(n3432), .Z(n3437) );
  NAND U4317 ( .A(n3435), .B(n3434), .Z(n3436) );
  AND U4318 ( .A(n3437), .B(n3436), .Z(n3512) );
  NANDN U4319 ( .A(n3439), .B(n3438), .Z(n3443) );
  NANDN U4320 ( .A(n3441), .B(n3440), .Z(n3442) );
  AND U4321 ( .A(n3443), .B(n3442), .Z(n3511) );
  XOR U4322 ( .A(n3512), .B(n3511), .Z(n3514) );
  XOR U4323 ( .A(n3513), .B(n3514), .Z(n3518) );
  XNOR U4324 ( .A(n3517), .B(n3518), .Z(n3520) );
  NANDN U4325 ( .A(n3445), .B(n3444), .Z(n3449) );
  NAND U4326 ( .A(n3447), .B(n3446), .Z(n3448) );
  AND U4327 ( .A(n3449), .B(n3448), .Z(n3524) );
  AND U4328 ( .A(y[68]), .B(x[8]), .Z(n3451) );
  NAND U4329 ( .A(y[65]), .B(x[11]), .Z(n3450) );
  XNOR U4330 ( .A(n3451), .B(n3450), .Z(n3585) );
  NAND U4331 ( .A(x[10]), .B(y[66]), .Z(n3646) );
  NAND U4332 ( .A(x[9]), .B(y[67]), .Z(n3595) );
  AND U4333 ( .A(x[28]), .B(y[144]), .Z(n3534) );
  NAND U4334 ( .A(x[1]), .B(y[27]), .Z(n3535) );
  XNOR U4335 ( .A(n3534), .B(n3535), .Z(n3536) );
  NAND U4336 ( .A(x[0]), .B(y[28]), .Z(n3537) );
  XNOR U4337 ( .A(n3536), .B(n3537), .Z(n3596) );
  XOR U4338 ( .A(n3597), .B(n3596), .Z(n3591) );
  NANDN U4339 ( .A(n3453), .B(n3452), .Z(n3457) );
  OR U4340 ( .A(n3455), .B(n3454), .Z(n3456) );
  AND U4341 ( .A(n3457), .B(n3456), .Z(n3589) );
  AND U4342 ( .A(x[35]), .B(y[187]), .Z(n3800) );
  NANDN U4343 ( .A(n3458), .B(n3800), .Z(n3462) );
  NANDN U4344 ( .A(n3460), .B(n3459), .Z(n3461) );
  AND U4345 ( .A(n3462), .B(n3461), .Z(n3588) );
  XNOR U4346 ( .A(n3589), .B(n3588), .Z(n3590) );
  XNOR U4347 ( .A(n3591), .B(n3590), .Z(n3621) );
  NAND U4348 ( .A(x[4]), .B(y[24]), .Z(n3570) );
  NAND U4349 ( .A(x[26]), .B(y[146]), .Z(n3569) );
  NAND U4350 ( .A(x[16]), .B(y[108]), .Z(n3568) );
  XNOR U4351 ( .A(n3569), .B(n3568), .Z(n3571) );
  AND U4352 ( .A(y[186]), .B(x[34]), .Z(n3490) );
  AND U4353 ( .A(x[33]), .B(y[185]), .Z(n3463) );
  NAND U4354 ( .A(n3490), .B(n3463), .Z(n3566) );
  NAND U4355 ( .A(x[20]), .B(y[104]), .Z(n3667) );
  NAND U4356 ( .A(x[32]), .B(y[188]), .Z(n3729) );
  XNOR U4357 ( .A(n3667), .B(n3729), .Z(n3567) );
  XOR U4358 ( .A(n3566), .B(n3567), .Z(n3555) );
  XOR U4359 ( .A(n3556), .B(n3555), .Z(n3558) );
  NANDN U4360 ( .A(n3465), .B(n3464), .Z(n3469) );
  OR U4361 ( .A(n3467), .B(n3466), .Z(n3468) );
  AND U4362 ( .A(n3469), .B(n3468), .Z(n3557) );
  XOR U4363 ( .A(n3558), .B(n3557), .Z(n3619) );
  NANDN U4364 ( .A(n3471), .B(n3470), .Z(n3475) );
  NANDN U4365 ( .A(n3473), .B(n3472), .Z(n3474) );
  AND U4366 ( .A(n3475), .B(n3474), .Z(n3618) );
  XNOR U4367 ( .A(n3621), .B(n3620), .Z(n3523) );
  XNOR U4368 ( .A(n3524), .B(n3523), .Z(n3526) );
  NANDN U4369 ( .A(n3477), .B(n3476), .Z(n3481) );
  NANDN U4370 ( .A(n3479), .B(n3478), .Z(n3480) );
  AND U4371 ( .A(n3481), .B(n3480), .Z(n3607) );
  NANDN U4372 ( .A(n3483), .B(n3482), .Z(n3487) );
  NANDN U4373 ( .A(n3485), .B(n3484), .Z(n3486) );
  NAND U4374 ( .A(n3487), .B(n3486), .Z(n3606) );
  NAND U4375 ( .A(x[2]), .B(y[26]), .Z(n3580) );
  NAND U4376 ( .A(x[27]), .B(y[145]), .Z(n3579) );
  NAND U4377 ( .A(x[3]), .B(y[25]), .Z(n3578) );
  XNOR U4378 ( .A(n3579), .B(n3578), .Z(n3581) );
  AND U4379 ( .A(y[187]), .B(x[33]), .Z(n3489) );
  NAND U4380 ( .A(y[184]), .B(x[36]), .Z(n3488) );
  XNOR U4381 ( .A(n3489), .B(n3488), .Z(n3563) );
  AND U4382 ( .A(x[35]), .B(y[185]), .Z(n3674) );
  XOR U4383 ( .A(n3674), .B(n3490), .Z(n3562) );
  XOR U4384 ( .A(n3563), .B(n3562), .Z(n3549) );
  XOR U4385 ( .A(n3550), .B(n3549), .Z(n3551) );
  NANDN U4386 ( .A(n3492), .B(n3491), .Z(n3496) );
  OR U4387 ( .A(n3494), .B(n3493), .Z(n3495) );
  NAND U4388 ( .A(n3496), .B(n3495), .Z(n3552) );
  XNOR U4389 ( .A(n3551), .B(n3552), .Z(n3615) );
  AND U4390 ( .A(x[19]), .B(y[105]), .Z(n3497) );
  NAND U4391 ( .A(n3498), .B(n3497), .Z(n3502) );
  NANDN U4392 ( .A(n3500), .B(n3499), .Z(n3501) );
  AND U4393 ( .A(n3502), .B(n3501), .Z(n3613) );
  AND U4394 ( .A(x[12]), .B(y[64]), .Z(n3540) );
  NAND U4395 ( .A(x[24]), .B(y[148]), .Z(n3541) );
  XNOR U4396 ( .A(n3540), .B(n3541), .Z(n3542) );
  NAND U4397 ( .A(x[25]), .B(y[147]), .Z(n3543) );
  XNOR U4398 ( .A(n3542), .B(n3543), .Z(n3600) );
  AND U4399 ( .A(y[106]), .B(x[18]), .Z(n3504) );
  NAND U4400 ( .A(y[105]), .B(x[19]), .Z(n3503) );
  XNOR U4401 ( .A(n3504), .B(n3503), .Z(n3530) );
  NAND U4402 ( .A(x[17]), .B(y[107]), .Z(n3531) );
  XOR U4403 ( .A(n3530), .B(n3531), .Z(n3601) );
  XNOR U4404 ( .A(n3600), .B(n3601), .Z(n3602) );
  NANDN U4405 ( .A(n3506), .B(n3505), .Z(n3510) );
  OR U4406 ( .A(n3508), .B(n3507), .Z(n3509) );
  NAND U4407 ( .A(n3510), .B(n3509), .Z(n3603) );
  XNOR U4408 ( .A(n3602), .B(n3603), .Z(n3612) );
  XOR U4409 ( .A(n3615), .B(n3614), .Z(n3608) );
  XOR U4410 ( .A(n3609), .B(n3608), .Z(n3525) );
  XNOR U4411 ( .A(n3526), .B(n3525), .Z(n3519) );
  XNOR U4412 ( .A(n3520), .B(n3519), .Z(o[28]) );
  NANDN U4413 ( .A(n3512), .B(n3511), .Z(n3516) );
  NANDN U4414 ( .A(n3514), .B(n3513), .Z(n3515) );
  AND U4415 ( .A(n3516), .B(n3515), .Z(n3765) );
  NANDN U4416 ( .A(n3518), .B(n3517), .Z(n3522) );
  NAND U4417 ( .A(n3520), .B(n3519), .Z(n3521) );
  NAND U4418 ( .A(n3522), .B(n3521), .Z(n3766) );
  XNOR U4419 ( .A(n3765), .B(n3766), .Z(n3768) );
  NANDN U4420 ( .A(n3524), .B(n3523), .Z(n3528) );
  NAND U4421 ( .A(n3526), .B(n3525), .Z(n3527) );
  AND U4422 ( .A(n3528), .B(n3527), .Z(n3625) );
  AND U4423 ( .A(x[19]), .B(y[106]), .Z(n3668) );
  NAND U4424 ( .A(n3529), .B(n3668), .Z(n3533) );
  NANDN U4425 ( .A(n3531), .B(n3530), .Z(n3532) );
  AND U4426 ( .A(n3533), .B(n3532), .Z(n3629) );
  NANDN U4427 ( .A(n3535), .B(n3534), .Z(n3539) );
  NANDN U4428 ( .A(n3537), .B(n3536), .Z(n3538) );
  NAND U4429 ( .A(n3539), .B(n3538), .Z(n3653) );
  AND U4430 ( .A(x[24]), .B(y[149]), .Z(n3975) );
  AND U4431 ( .A(x[13]), .B(y[64]), .Z(n3658) );
  AND U4432 ( .A(x[18]), .B(y[107]), .Z(n3657) );
  XOR U4433 ( .A(n3658), .B(n3657), .Z(n3659) );
  XOR U4434 ( .A(n3975), .B(n3659), .Z(n3652) );
  AND U4435 ( .A(x[28]), .B(y[145]), .Z(n3663) );
  AND U4436 ( .A(x[5]), .B(y[24]), .Z(n3662) );
  XOR U4437 ( .A(n3663), .B(n3662), .Z(n3664) );
  AND U4438 ( .A(x[4]), .B(y[25]), .Z(n3995) );
  XOR U4439 ( .A(n3664), .B(n3995), .Z(n3651) );
  XOR U4440 ( .A(n3652), .B(n3651), .Z(n3654) );
  XOR U4441 ( .A(n3653), .B(n3654), .Z(n3628) );
  NANDN U4442 ( .A(n3541), .B(n3540), .Z(n3545) );
  NANDN U4443 ( .A(n3543), .B(n3542), .Z(n3544) );
  NAND U4444 ( .A(n3545), .B(n3544), .Z(n3707) );
  AND U4445 ( .A(y[186]), .B(x[35]), .Z(n3575) );
  AND U4446 ( .A(n3575), .B(n3546), .Z(n3731) );
  AND U4447 ( .A(y[189]), .B(x[32]), .Z(n3548) );
  AND U4448 ( .A(y[188]), .B(x[33]), .Z(n3547) );
  XOR U4449 ( .A(n3548), .B(n3547), .Z(n3730) );
  XOR U4450 ( .A(n3731), .B(n3730), .Z(n3706) );
  AND U4451 ( .A(x[8]), .B(y[69]), .Z(n3714) );
  AND U4452 ( .A(x[1]), .B(y[28]), .Z(n3713) );
  XOR U4453 ( .A(n3714), .B(n3713), .Z(n3716) );
  AND U4454 ( .A(x[12]), .B(y[65]), .Z(n3715) );
  XOR U4455 ( .A(n3716), .B(n3715), .Z(n3705) );
  XOR U4456 ( .A(n3706), .B(n3705), .Z(n3708) );
  XOR U4457 ( .A(n3707), .B(n3708), .Z(n3630) );
  XOR U4458 ( .A(n3631), .B(n3630), .Z(n3678) );
  NAND U4459 ( .A(n3550), .B(n3549), .Z(n3554) );
  NANDN U4460 ( .A(n3552), .B(n3551), .Z(n3553) );
  AND U4461 ( .A(n3554), .B(n3553), .Z(n3675) );
  NAND U4462 ( .A(n3556), .B(n3555), .Z(n3560) );
  NAND U4463 ( .A(n3558), .B(n3557), .Z(n3559) );
  NAND U4464 ( .A(n3560), .B(n3559), .Z(n3676) );
  AND U4465 ( .A(x[36]), .B(y[187]), .Z(n3866) );
  NAND U4466 ( .A(n3866), .B(n3561), .Z(n3565) );
  NAND U4467 ( .A(n3563), .B(n3562), .Z(n3564) );
  AND U4468 ( .A(n3565), .B(n3564), .Z(n3688) );
  NAND U4469 ( .A(n3569), .B(n3568), .Z(n3573) );
  NANDN U4470 ( .A(n3571), .B(n3570), .Z(n3572) );
  AND U4471 ( .A(n3573), .B(n3572), .Z(n3696) );
  AND U4472 ( .A(x[9]), .B(y[68]), .Z(n3647) );
  AND U4473 ( .A(x[11]), .B(y[66]), .Z(n3796) );
  NAND U4474 ( .A(y[67]), .B(x[10]), .Z(n3574) );
  XOR U4475 ( .A(n3796), .B(n3574), .Z(n3648) );
  NAND U4476 ( .A(x[36]), .B(y[185]), .Z(n3821) );
  XNOR U4477 ( .A(n3575), .B(n3821), .Z(n3637) );
  AND U4478 ( .A(x[37]), .B(y[184]), .Z(n3634) );
  NAND U4479 ( .A(x[34]), .B(y[187]), .Z(n3635) );
  XOR U4480 ( .A(n3637), .B(n3636), .Z(n3693) );
  XOR U4481 ( .A(n3694), .B(n3693), .Z(n3695) );
  XOR U4482 ( .A(n3696), .B(n3695), .Z(n3689) );
  XOR U4483 ( .A(n3690), .B(n3689), .Z(n3750) );
  AND U4484 ( .A(y[104]), .B(x[21]), .Z(n3577) );
  NAND U4485 ( .A(y[105]), .B(x[20]), .Z(n3576) );
  XOR U4486 ( .A(n3577), .B(n3576), .Z(n3669) );
  AND U4487 ( .A(x[29]), .B(y[144]), .Z(n3640) );
  NAND U4488 ( .A(x[3]), .B(y[26]), .Z(n3641) );
  NAND U4489 ( .A(x[2]), .B(y[27]), .Z(n3643) );
  XOR U4490 ( .A(n3724), .B(n3723), .Z(n3726) );
  NAND U4491 ( .A(n3579), .B(n3578), .Z(n3583) );
  NANDN U4492 ( .A(n3581), .B(n3580), .Z(n3582) );
  AND U4493 ( .A(n3583), .B(n3582), .Z(n3725) );
  XOR U4494 ( .A(n3726), .B(n3725), .Z(n3748) );
  AND U4495 ( .A(x[11]), .B(y[68]), .Z(n3869) );
  NAND U4496 ( .A(n3869), .B(n3584), .Z(n3587) );
  NANDN U4497 ( .A(n3646), .B(n3585), .Z(n3586) );
  AND U4498 ( .A(n3587), .B(n3586), .Z(n3684) );
  AND U4499 ( .A(x[27]), .B(y[146]), .Z(n3742) );
  AND U4500 ( .A(x[17]), .B(y[108]), .Z(n3927) );
  XOR U4501 ( .A(n3742), .B(n3927), .Z(n3744) );
  AND U4502 ( .A(x[16]), .B(y[109]), .Z(n3743) );
  XOR U4503 ( .A(n3744), .B(n3743), .Z(n3682) );
  AND U4504 ( .A(x[0]), .B(y[29]), .Z(n3735) );
  AND U4505 ( .A(x[25]), .B(y[148]), .Z(n3734) );
  XOR U4506 ( .A(n3735), .B(n3734), .Z(n3737) );
  AND U4507 ( .A(x[26]), .B(y[147]), .Z(n3736) );
  XOR U4508 ( .A(n3737), .B(n3736), .Z(n3681) );
  XOR U4509 ( .A(n3682), .B(n3681), .Z(n3683) );
  XOR U4510 ( .A(n3684), .B(n3683), .Z(n3747) );
  NANDN U4511 ( .A(n3589), .B(n3588), .Z(n3593) );
  NANDN U4512 ( .A(n3591), .B(n3590), .Z(n3592) );
  AND U4513 ( .A(n3593), .B(n3592), .Z(n3702) );
  NANDN U4514 ( .A(n3595), .B(n3594), .Z(n3599) );
  NAND U4515 ( .A(n3597), .B(n3596), .Z(n3598) );
  AND U4516 ( .A(n3599), .B(n3598), .Z(n3700) );
  NANDN U4517 ( .A(n3601), .B(n3600), .Z(n3605) );
  NANDN U4518 ( .A(n3603), .B(n3602), .Z(n3604) );
  NAND U4519 ( .A(n3605), .B(n3604), .Z(n3699) );
  XOR U4520 ( .A(n3702), .B(n3701), .Z(n3760) );
  XOR U4521 ( .A(n3759), .B(n3760), .Z(n3762) );
  XOR U4522 ( .A(n3761), .B(n3762), .Z(n3624) );
  XNOR U4523 ( .A(n3625), .B(n3624), .Z(n3627) );
  NANDN U4524 ( .A(n3607), .B(n3606), .Z(n3611) );
  NAND U4525 ( .A(n3609), .B(n3608), .Z(n3610) );
  AND U4526 ( .A(n3611), .B(n3610), .Z(n3756) );
  NANDN U4527 ( .A(n3613), .B(n3612), .Z(n3617) );
  NAND U4528 ( .A(n3615), .B(n3614), .Z(n3616) );
  AND U4529 ( .A(n3617), .B(n3616), .Z(n3754) );
  NANDN U4530 ( .A(n3619), .B(n3618), .Z(n3623) );
  NAND U4531 ( .A(n3621), .B(n3620), .Z(n3622) );
  AND U4532 ( .A(n3623), .B(n3622), .Z(n3753) );
  XOR U4533 ( .A(n3627), .B(n3626), .Z(n3767) );
  XOR U4534 ( .A(n3768), .B(n3767), .Z(o[29]) );
  NANDN U4535 ( .A(n3629), .B(n3628), .Z(n3633) );
  NAND U4536 ( .A(n3631), .B(n3630), .Z(n3632) );
  AND U4537 ( .A(n3633), .B(n3632), .Z(n4045) );
  NANDN U4538 ( .A(n3635), .B(n3634), .Z(n3639) );
  NAND U4539 ( .A(n3637), .B(n3636), .Z(n3638) );
  NAND U4540 ( .A(n3639), .B(n3638), .Z(n3906) );
  NANDN U4541 ( .A(n3641), .B(n3640), .Z(n3645) );
  NANDN U4542 ( .A(n3643), .B(n3642), .Z(n3644) );
  NAND U4543 ( .A(n3645), .B(n3644), .Z(n3909) );
  AND U4544 ( .A(y[67]), .B(x[11]), .Z(n3711) );
  NANDN U4545 ( .A(n3646), .B(n3711), .Z(n3650) );
  NANDN U4546 ( .A(n3648), .B(n3647), .Z(n3649) );
  AND U4547 ( .A(n3650), .B(n3649), .Z(n3791) );
  AND U4548 ( .A(x[27]), .B(y[147]), .Z(n3933) );
  AND U4549 ( .A(x[19]), .B(y[107]), .Z(n3932) );
  XOR U4550 ( .A(n3933), .B(n3932), .Z(n3931) );
  AND U4551 ( .A(x[3]), .B(y[27]), .Z(n3930) );
  XOR U4552 ( .A(n3931), .B(n3930), .Z(n3793) );
  AND U4553 ( .A(x[26]), .B(y[148]), .Z(n3816) );
  AND U4554 ( .A(x[20]), .B(y[106]), .Z(n3815) );
  XOR U4555 ( .A(n3816), .B(n3815), .Z(n3814) );
  AND U4556 ( .A(x[2]), .B(y[28]), .Z(n3813) );
  XNOR U4557 ( .A(n3814), .B(n3813), .Z(n3792) );
  XNOR U4558 ( .A(n3791), .B(n3790), .Z(n3908) );
  XOR U4559 ( .A(n3909), .B(n3908), .Z(n3907) );
  XOR U4560 ( .A(n3906), .B(n3907), .Z(n4013) );
  NAND U4561 ( .A(n3652), .B(n3651), .Z(n3656) );
  NAND U4562 ( .A(n3654), .B(n3653), .Z(n3655) );
  NAND U4563 ( .A(n3656), .B(n3655), .Z(n4012) );
  XOR U4564 ( .A(n4013), .B(n4012), .Z(n4011) );
  NAND U4565 ( .A(n3658), .B(n3657), .Z(n3661) );
  NAND U4566 ( .A(n3975), .B(n3659), .Z(n3660) );
  NAND U4567 ( .A(n3661), .B(n3660), .Z(n3915) );
  NAND U4568 ( .A(n3663), .B(n3662), .Z(n3666) );
  NAND U4569 ( .A(n3664), .B(n3995), .Z(n3665) );
  NAND U4570 ( .A(n3666), .B(n3665), .Z(n3914) );
  XOR U4571 ( .A(n3915), .B(n3914), .Z(n3913) );
  AND U4572 ( .A(x[21]), .B(y[105]), .Z(n3941) );
  NANDN U4573 ( .A(n3667), .B(n3941), .Z(n3671) );
  NANDN U4574 ( .A(n3669), .B(n3668), .Z(n3670) );
  AND U4575 ( .A(n3671), .B(n3670), .Z(n3784) );
  AND U4576 ( .A(y[25]), .B(x[5]), .Z(n3673) );
  NAND U4577 ( .A(y[26]), .B(x[4]), .Z(n3672) );
  XNOR U4578 ( .A(n3673), .B(n3672), .Z(n3993) );
  AND U4579 ( .A(x[30]), .B(y[144]), .Z(n3992) );
  XOR U4580 ( .A(n3993), .B(n3992), .Z(n3786) );
  AND U4581 ( .A(x[33]), .B(y[189]), .Z(n3808) );
  AND U4582 ( .A(x[36]), .B(y[186]), .Z(n3741) );
  AND U4583 ( .A(n3674), .B(n3741), .Z(n3806) );
  AND U4584 ( .A(x[34]), .B(y[188]), .Z(n3805) );
  XOR U4585 ( .A(n3806), .B(n3805), .Z(n3807) );
  XNOR U4586 ( .A(n3808), .B(n3807), .Z(n3785) );
  XNOR U4587 ( .A(n3784), .B(n3783), .Z(n3912) );
  XOR U4588 ( .A(n3913), .B(n3912), .Z(n4010) );
  XOR U4589 ( .A(n4011), .B(n4010), .Z(n3780) );
  NANDN U4590 ( .A(n3676), .B(n3675), .Z(n3680) );
  NANDN U4591 ( .A(n3678), .B(n3677), .Z(n3679) );
  NAND U4592 ( .A(n3680), .B(n3679), .Z(n3779) );
  NAND U4593 ( .A(n3682), .B(n3681), .Z(n3686) );
  NANDN U4594 ( .A(n3684), .B(n3683), .Z(n3685) );
  AND U4595 ( .A(n3686), .B(n3685), .Z(n4007) );
  NANDN U4596 ( .A(n3688), .B(n3687), .Z(n3692) );
  NAND U4597 ( .A(n3690), .B(n3689), .Z(n3691) );
  AND U4598 ( .A(n3692), .B(n3691), .Z(n4006) );
  XOR U4599 ( .A(n4007), .B(n4006), .Z(n4005) );
  NAND U4600 ( .A(n3694), .B(n3693), .Z(n3698) );
  NAND U4601 ( .A(n3696), .B(n3695), .Z(n3697) );
  AND U4602 ( .A(n3698), .B(n3697), .Z(n4004) );
  XOR U4603 ( .A(n4005), .B(n4004), .Z(n3777) );
  XOR U4604 ( .A(n3778), .B(n3777), .Z(n4044) );
  XOR U4605 ( .A(n4045), .B(n4044), .Z(n4047) );
  NANDN U4606 ( .A(n3700), .B(n3699), .Z(n3704) );
  NAND U4607 ( .A(n3702), .B(n3701), .Z(n3703) );
  AND U4608 ( .A(n3704), .B(n3703), .Z(n4027) );
  NAND U4609 ( .A(n3706), .B(n3705), .Z(n3710) );
  NAND U4610 ( .A(n3708), .B(n3707), .Z(n3709) );
  AND U4611 ( .A(n3710), .B(n3709), .Z(n3900) );
  AND U4612 ( .A(x[32]), .B(y[190]), .Z(n3940) );
  XOR U4613 ( .A(n3941), .B(n3940), .Z(n3939) );
  AND U4614 ( .A(x[22]), .B(y[104]), .Z(n3938) );
  XOR U4615 ( .A(n3939), .B(n3938), .Z(n3789) );
  AND U4616 ( .A(x[16]), .B(y[110]), .Z(n3947) );
  AND U4617 ( .A(x[6]), .B(y[24]), .Z(n3946) );
  XOR U4618 ( .A(n3947), .B(n3946), .Z(n3945) );
  AND U4619 ( .A(x[29]), .B(y[145]), .Z(n3944) );
  XNOR U4620 ( .A(n3945), .B(n3944), .Z(n3788) );
  AND U4621 ( .A(x[13]), .B(y[65]), .Z(n3981) );
  AND U4622 ( .A(x[10]), .B(y[68]), .Z(n3980) );
  XOR U4623 ( .A(n3981), .B(n3980), .Z(n3979) );
  AND U4624 ( .A(x[9]), .B(y[69]), .Z(n3978) );
  XOR U4625 ( .A(n3979), .B(n3978), .Z(n3795) );
  AND U4626 ( .A(y[66]), .B(x[12]), .Z(n3712) );
  XOR U4627 ( .A(n3712), .B(n3711), .Z(n3794) );
  XOR U4628 ( .A(n3795), .B(n3794), .Z(n3787) );
  NAND U4629 ( .A(n3714), .B(n3713), .Z(n3718) );
  NAND U4630 ( .A(n3716), .B(n3715), .Z(n3717) );
  AND U4631 ( .A(n3718), .B(n3717), .Z(n3919) );
  AND U4632 ( .A(x[28]), .B(y[146]), .Z(n3925) );
  AND U4633 ( .A(x[18]), .B(y[108]), .Z(n3720) );
  AND U4634 ( .A(y[109]), .B(x[17]), .Z(n3719) );
  XOR U4635 ( .A(n3720), .B(n3719), .Z(n3924) );
  XOR U4636 ( .A(n3925), .B(n3924), .Z(n3921) );
  AND U4637 ( .A(x[0]), .B(y[30]), .Z(n3973) );
  AND U4638 ( .A(y[150]), .B(x[24]), .Z(n3722) );
  NAND U4639 ( .A(y[149]), .B(x[25]), .Z(n3721) );
  XNOR U4640 ( .A(n3722), .B(n3721), .Z(n3972) );
  XNOR U4641 ( .A(n3973), .B(n3972), .Z(n3920) );
  XOR U4642 ( .A(n3919), .B(n3918), .Z(n3902) );
  XNOR U4643 ( .A(n3900), .B(n3901), .Z(n4034) );
  NAND U4644 ( .A(n3724), .B(n3723), .Z(n3728) );
  NAND U4645 ( .A(n3726), .B(n3725), .Z(n3727) );
  NAND U4646 ( .A(n3728), .B(n3727), .Z(n4032) );
  NANDN U4647 ( .A(n3729), .B(n3808), .Z(n3733) );
  NAND U4648 ( .A(n3731), .B(n3730), .Z(n3732) );
  NAND U4649 ( .A(n3733), .B(n3732), .Z(n3959) );
  NAND U4650 ( .A(n3735), .B(n3734), .Z(n3739) );
  NAND U4651 ( .A(n3737), .B(n3736), .Z(n3738) );
  AND U4652 ( .A(n3739), .B(n3738), .Z(n3963) );
  AND U4653 ( .A(x[1]), .B(y[29]), .Z(n3989) );
  AND U4654 ( .A(x[14]), .B(y[64]), .Z(n3988) );
  XOR U4655 ( .A(n3989), .B(n3988), .Z(n3987) );
  AND U4656 ( .A(x[8]), .B(y[70]), .Z(n3986) );
  XOR U4657 ( .A(n3987), .B(n3986), .Z(n3965) );
  NAND U4658 ( .A(y[185]), .B(x[37]), .Z(n3740) );
  XNOR U4659 ( .A(n3741), .B(n3740), .Z(n3802) );
  AND U4660 ( .A(x[38]), .B(y[184]), .Z(n3801) );
  XOR U4661 ( .A(n3802), .B(n3801), .Z(n3799) );
  XNOR U4662 ( .A(n3800), .B(n3799), .Z(n3964) );
  XNOR U4663 ( .A(n3963), .B(n3962), .Z(n3958) );
  XOR U4664 ( .A(n3959), .B(n3958), .Z(n3957) );
  NAND U4665 ( .A(n3742), .B(n3927), .Z(n3746) );
  NAND U4666 ( .A(n3744), .B(n3743), .Z(n3745) );
  NAND U4667 ( .A(n3746), .B(n3745), .Z(n3956) );
  XOR U4668 ( .A(n3957), .B(n3956), .Z(n4033) );
  XOR U4669 ( .A(n4032), .B(n4033), .Z(n4035) );
  NANDN U4670 ( .A(n3748), .B(n3747), .Z(n3752) );
  NANDN U4671 ( .A(n3750), .B(n3749), .Z(n3751) );
  NAND U4672 ( .A(n3752), .B(n3751), .Z(n4029) );
  XOR U4673 ( .A(n4027), .B(n4026), .Z(n4046) );
  XOR U4674 ( .A(n4047), .B(n4046), .Z(n4053) );
  NANDN U4675 ( .A(n3754), .B(n3753), .Z(n3758) );
  NANDN U4676 ( .A(n3756), .B(n3755), .Z(n3757) );
  NAND U4677 ( .A(n3758), .B(n3757), .Z(n4051) );
  NAND U4678 ( .A(n3760), .B(n3759), .Z(n3764) );
  NAND U4679 ( .A(n3762), .B(n3761), .Z(n3763) );
  NAND U4680 ( .A(n3764), .B(n3763), .Z(n4050) );
  XOR U4681 ( .A(n4051), .B(n4050), .Z(n4052) );
  NANDN U4682 ( .A(n3766), .B(n3765), .Z(n3770) );
  NAND U4683 ( .A(n3768), .B(n3767), .Z(n3769) );
  NAND U4684 ( .A(n3770), .B(n3769), .Z(n3771) );
  XOR U4685 ( .A(n3772), .B(n3771), .Z(o[30]) );
  NAND U4686 ( .A(n3772), .B(n3771), .Z(n3776) );
  NANDN U4687 ( .A(n3774), .B(n3773), .Z(n3775) );
  AND U4688 ( .A(n3776), .B(n3775), .Z(n4043) );
  NAND U4689 ( .A(n3778), .B(n3777), .Z(n3782) );
  NANDN U4690 ( .A(n3780), .B(n3779), .Z(n3781) );
  AND U4691 ( .A(n3782), .B(n3781), .Z(n4025) );
  NAND U4692 ( .A(n3795), .B(n3794), .Z(n3798) );
  AND U4693 ( .A(x[12]), .B(y[67]), .Z(n3865) );
  NAND U4694 ( .A(n3796), .B(n3865), .Z(n3797) );
  NAND U4695 ( .A(n3800), .B(n3799), .Z(n3804) );
  AND U4696 ( .A(n3802), .B(n3801), .Z(n3803) );
  ANDN U4697 ( .B(n3804), .A(n3803), .Z(n3812) );
  AND U4698 ( .A(n3806), .B(n3805), .Z(n3810) );
  AND U4699 ( .A(n3808), .B(n3807), .Z(n3809) );
  OR U4700 ( .A(n3810), .B(n3809), .Z(n3811) );
  XNOR U4701 ( .A(n3812), .B(n3811), .Z(n3899) );
  NAND U4702 ( .A(n3814), .B(n3813), .Z(n3818) );
  NAND U4703 ( .A(n3816), .B(n3815), .Z(n3817) );
  AND U4704 ( .A(n3818), .B(n3817), .Z(n3897) );
  AND U4705 ( .A(y[188]), .B(x[35]), .Z(n3820) );
  NAND U4706 ( .A(y[189]), .B(x[34]), .Z(n3819) );
  XNOR U4707 ( .A(n3820), .B(n3819), .Z(n3826) );
  AND U4708 ( .A(y[186]), .B(n3821), .Z(n3822) );
  AND U4709 ( .A(n3822), .B(x[37]), .Z(n3824) );
  NAND U4710 ( .A(y[27]), .B(x[4]), .Z(n3823) );
  XNOR U4711 ( .A(n3824), .B(n3823), .Z(n3825) );
  XOR U4712 ( .A(n3826), .B(n3825), .Z(n3834) );
  AND U4713 ( .A(y[105]), .B(x[22]), .Z(n3828) );
  NAND U4714 ( .A(y[25]), .B(x[6]), .Z(n3827) );
  XNOR U4715 ( .A(n3828), .B(n3827), .Z(n3832) );
  AND U4716 ( .A(y[24]), .B(x[7]), .Z(n3830) );
  NAND U4717 ( .A(y[147]), .B(x[28]), .Z(n3829) );
  XNOR U4718 ( .A(n3830), .B(n3829), .Z(n3831) );
  XNOR U4719 ( .A(n3832), .B(n3831), .Z(n3833) );
  XNOR U4720 ( .A(n3834), .B(n3833), .Z(n3895) );
  AND U4721 ( .A(y[104]), .B(x[23]), .Z(n3836) );
  NAND U4722 ( .A(y[191]), .B(x[32]), .Z(n3835) );
  XNOR U4723 ( .A(n3836), .B(n3835), .Z(n3840) );
  AND U4724 ( .A(y[31]), .B(x[0]), .Z(n3838) );
  NAND U4725 ( .A(y[190]), .B(x[33]), .Z(n3837) );
  XNOR U4726 ( .A(n3838), .B(n3837), .Z(n3839) );
  XOR U4727 ( .A(n3840), .B(n3839), .Z(n3848) );
  AND U4728 ( .A(y[30]), .B(x[1]), .Z(n3842) );
  NAND U4729 ( .A(y[106]), .B(x[21]), .Z(n3841) );
  XNOR U4730 ( .A(n3842), .B(n3841), .Z(n3846) );
  AND U4731 ( .A(y[146]), .B(x[29]), .Z(n3844) );
  NAND U4732 ( .A(y[111]), .B(x[16]), .Z(n3843) );
  XNOR U4733 ( .A(n3844), .B(n3843), .Z(n3845) );
  XNOR U4734 ( .A(n3846), .B(n3845), .Z(n3847) );
  XNOR U4735 ( .A(n3848), .B(n3847), .Z(n3864) );
  AND U4736 ( .A(y[184]), .B(x[39]), .Z(n3850) );
  NAND U4737 ( .A(y[148]), .B(x[27]), .Z(n3849) );
  XNOR U4738 ( .A(n3850), .B(n3849), .Z(n3854) );
  AND U4739 ( .A(y[110]), .B(x[17]), .Z(n3852) );
  NAND U4740 ( .A(y[108]), .B(x[19]), .Z(n3851) );
  XNOR U4741 ( .A(n3852), .B(n3851), .Z(n3853) );
  XOR U4742 ( .A(n3854), .B(n3853), .Z(n3862) );
  AND U4743 ( .A(y[144]), .B(x[31]), .Z(n3856) );
  NAND U4744 ( .A(y[107]), .B(x[20]), .Z(n3855) );
  XNOR U4745 ( .A(n3856), .B(n3855), .Z(n3860) );
  AND U4746 ( .A(y[71]), .B(x[8]), .Z(n3858) );
  NAND U4747 ( .A(y[29]), .B(x[2]), .Z(n3857) );
  XNOR U4748 ( .A(n3858), .B(n3857), .Z(n3859) );
  XNOR U4749 ( .A(n3860), .B(n3859), .Z(n3861) );
  XNOR U4750 ( .A(n3862), .B(n3861), .Z(n3863) );
  XOR U4751 ( .A(n3864), .B(n3863), .Z(n3893) );
  AND U4752 ( .A(x[18]), .B(y[109]), .Z(n3926) );
  AND U4753 ( .A(x[25]), .B(y[150]), .Z(n3974) );
  XOR U4754 ( .A(n3926), .B(n3974), .Z(n3868) );
  XNOR U4755 ( .A(n3866), .B(n3865), .Z(n3867) );
  XNOR U4756 ( .A(n3868), .B(n3867), .Z(n3891) );
  AND U4757 ( .A(y[70]), .B(x[9]), .Z(n3889) );
  AND U4758 ( .A(y[151]), .B(x[24]), .Z(n3871) );
  AND U4759 ( .A(x[5]), .B(y[26]), .Z(n3994) );
  XNOR U4760 ( .A(n3994), .B(n3869), .Z(n3870) );
  XNOR U4761 ( .A(n3871), .B(n3870), .Z(n3887) );
  AND U4762 ( .A(y[185]), .B(x[38]), .Z(n3873) );
  NAND U4763 ( .A(y[145]), .B(x[30]), .Z(n3872) );
  XNOR U4764 ( .A(n3873), .B(n3872), .Z(n3877) );
  AND U4765 ( .A(y[65]), .B(x[14]), .Z(n3875) );
  NAND U4766 ( .A(y[28]), .B(x[3]), .Z(n3874) );
  XNOR U4767 ( .A(n3875), .B(n3874), .Z(n3876) );
  XOR U4768 ( .A(n3877), .B(n3876), .Z(n3885) );
  AND U4769 ( .A(y[64]), .B(x[15]), .Z(n3879) );
  NAND U4770 ( .A(y[149]), .B(x[26]), .Z(n3878) );
  XNOR U4771 ( .A(n3879), .B(n3878), .Z(n3883) );
  AND U4772 ( .A(y[66]), .B(x[13]), .Z(n3881) );
  NAND U4773 ( .A(y[69]), .B(x[10]), .Z(n3880) );
  XNOR U4774 ( .A(n3881), .B(n3880), .Z(n3882) );
  XNOR U4775 ( .A(n3883), .B(n3882), .Z(n3884) );
  XNOR U4776 ( .A(n3885), .B(n3884), .Z(n3886) );
  XNOR U4777 ( .A(n3887), .B(n3886), .Z(n3888) );
  XNOR U4778 ( .A(n3889), .B(n3888), .Z(n3890) );
  XNOR U4779 ( .A(n3891), .B(n3890), .Z(n3892) );
  XNOR U4780 ( .A(n3893), .B(n3892), .Z(n3894) );
  XNOR U4781 ( .A(n3895), .B(n3894), .Z(n3896) );
  XNOR U4782 ( .A(n3897), .B(n3896), .Z(n3898) );
  NANDN U4783 ( .A(n3901), .B(n3900), .Z(n3905) );
  NANDN U4784 ( .A(n3903), .B(n3902), .Z(n3904) );
  NAND U4785 ( .A(n3907), .B(n3906), .Z(n3911) );
  NAND U4786 ( .A(n3909), .B(n3908), .Z(n3910) );
  NAND U4787 ( .A(n3913), .B(n3912), .Z(n3917) );
  NAND U4788 ( .A(n3915), .B(n3914), .Z(n3916) );
  AND U4789 ( .A(n3917), .B(n3916), .Z(n4021) );
  NAND U4790 ( .A(n3919), .B(n3918), .Z(n3923) );
  NANDN U4791 ( .A(n3921), .B(n3920), .Z(n3922) );
  AND U4792 ( .A(n3923), .B(n3922), .Z(n3955) );
  NAND U4793 ( .A(n3925), .B(n3924), .Z(n3929) );
  NAND U4794 ( .A(n3927), .B(n3926), .Z(n3928) );
  AND U4795 ( .A(n3929), .B(n3928), .Z(n3937) );
  NAND U4796 ( .A(n3931), .B(n3930), .Z(n3935) );
  NAND U4797 ( .A(n3933), .B(n3932), .Z(n3934) );
  NAND U4798 ( .A(n3935), .B(n3934), .Z(n3936) );
  XNOR U4799 ( .A(n3937), .B(n3936), .Z(n3953) );
  NAND U4800 ( .A(n3939), .B(n3938), .Z(n3943) );
  NAND U4801 ( .A(n3941), .B(n3940), .Z(n3942) );
  AND U4802 ( .A(n3943), .B(n3942), .Z(n3951) );
  NAND U4803 ( .A(n3945), .B(n3944), .Z(n3949) );
  NAND U4804 ( .A(n3947), .B(n3946), .Z(n3948) );
  NAND U4805 ( .A(n3949), .B(n3948), .Z(n3950) );
  XNOR U4806 ( .A(n3951), .B(n3950), .Z(n3952) );
  XNOR U4807 ( .A(n3953), .B(n3952), .Z(n3954) );
  XNOR U4808 ( .A(n3955), .B(n3954), .Z(n3971) );
  NAND U4809 ( .A(n3957), .B(n3956), .Z(n3961) );
  NAND U4810 ( .A(n3959), .B(n3958), .Z(n3960) );
  AND U4811 ( .A(n3961), .B(n3960), .Z(n3969) );
  NAND U4812 ( .A(n3963), .B(n3962), .Z(n3967) );
  NANDN U4813 ( .A(n3965), .B(n3964), .Z(n3966) );
  NAND U4814 ( .A(n3967), .B(n3966), .Z(n3968) );
  XNOR U4815 ( .A(n3969), .B(n3968), .Z(n3970) );
  XOR U4816 ( .A(n3971), .B(n3970), .Z(n4003) );
  NAND U4817 ( .A(n3973), .B(n3972), .Z(n3977) );
  NAND U4818 ( .A(n3975), .B(n3974), .Z(n3976) );
  AND U4819 ( .A(n3977), .B(n3976), .Z(n3985) );
  NAND U4820 ( .A(n3979), .B(n3978), .Z(n3983) );
  NAND U4821 ( .A(n3981), .B(n3980), .Z(n3982) );
  NAND U4822 ( .A(n3983), .B(n3982), .Z(n3984) );
  XNOR U4823 ( .A(n3985), .B(n3984), .Z(n4001) );
  NAND U4824 ( .A(n3987), .B(n3986), .Z(n3991) );
  NAND U4825 ( .A(n3989), .B(n3988), .Z(n3990) );
  AND U4826 ( .A(n3991), .B(n3990), .Z(n3999) );
  NAND U4827 ( .A(n3993), .B(n3992), .Z(n3997) );
  NAND U4828 ( .A(n3995), .B(n3994), .Z(n3996) );
  NAND U4829 ( .A(n3997), .B(n3996), .Z(n3998) );
  XNOR U4830 ( .A(n3999), .B(n3998), .Z(n4000) );
  XNOR U4831 ( .A(n4001), .B(n4000), .Z(n4002) );
  XNOR U4832 ( .A(n4003), .B(n4002), .Z(n4019) );
  NAND U4833 ( .A(n4005), .B(n4004), .Z(n4009) );
  NAND U4834 ( .A(n4007), .B(n4006), .Z(n4008) );
  AND U4835 ( .A(n4009), .B(n4008), .Z(n4017) );
  NAND U4836 ( .A(n4011), .B(n4010), .Z(n4015) );
  NAND U4837 ( .A(n4013), .B(n4012), .Z(n4014) );
  NAND U4838 ( .A(n4015), .B(n4014), .Z(n4016) );
  XNOR U4839 ( .A(n4017), .B(n4016), .Z(n4018) );
  XNOR U4840 ( .A(n4019), .B(n4018), .Z(n4020) );
  XNOR U4841 ( .A(n4021), .B(n4020), .Z(n4022) );
  XNOR U4842 ( .A(n4023), .B(n4022), .Z(n4024) );
  XNOR U4843 ( .A(n4025), .B(n4024), .Z(n4041) );
  NAND U4844 ( .A(n4027), .B(n4026), .Z(n4031) );
  ANDN U4845 ( .B(n4029), .A(n4028), .Z(n4030) );
  ANDN U4846 ( .B(n4031), .A(n4030), .Z(n4039) );
  AND U4847 ( .A(n4033), .B(n4032), .Z(n4037) );
  ANDN U4848 ( .B(n4035), .A(n4034), .Z(n4036) );
  OR U4849 ( .A(n4037), .B(n4036), .Z(n4038) );
  XNOR U4850 ( .A(n4039), .B(n4038), .Z(n4040) );
  XNOR U4851 ( .A(n4041), .B(n4040), .Z(n4042) );
  XNOR U4852 ( .A(n4043), .B(n4042), .Z(n4059) );
  AND U4853 ( .A(n4045), .B(n4044), .Z(n4049) );
  AND U4854 ( .A(n4047), .B(n4046), .Z(n4048) );
  NOR U4855 ( .A(n4049), .B(n4048), .Z(n4057) );
  NAND U4856 ( .A(n4051), .B(n4050), .Z(n4055) );
  NANDN U4857 ( .A(n4053), .B(n4052), .Z(n4054) );
  AND U4858 ( .A(n4055), .B(n4054), .Z(n4056) );
  XNOR U4859 ( .A(n4057), .B(n4056), .Z(n4058) );
  XNOR U4860 ( .A(n4059), .B(n4058), .Z(o[31]) );
  NAND U4861 ( .A(x[32]), .B(y[192]), .Z(n4194) );
  NAND U4862 ( .A(x[8]), .B(y[72]), .Z(n4062) );
  XOR U4863 ( .A(n4194), .B(n4062), .Z(n4063) );
  AND U4864 ( .A(x[0]), .B(y[32]), .Z(n4070) );
  AND U4865 ( .A(x[16]), .B(y[112]), .Z(n4067) );
  XOR U4866 ( .A(n4070), .B(n4067), .Z(n4066) );
  AND U4867 ( .A(x[24]), .B(y[152]), .Z(n4065) );
  XNOR U4868 ( .A(n4066), .B(n4065), .Z(n4064) );
  XNOR U4869 ( .A(n4063), .B(n4064), .Z(o[32]) );
  AND U4870 ( .A(y[32]), .B(x[1]), .Z(n4061) );
  NAND U4871 ( .A(y[33]), .B(x[0]), .Z(n4060) );
  XNOR U4872 ( .A(n4061), .B(n4060), .Z(n4071) );
  NAND U4873 ( .A(x[9]), .B(y[72]), .Z(n4072) );
  XOR U4874 ( .A(n4071), .B(n4072), .Z(n4088) );
  AND U4875 ( .A(x[33]), .B(y[192]), .Z(n4285) );
  NAND U4876 ( .A(x[16]), .B(y[113]), .Z(n4075) );
  XNOR U4877 ( .A(n4285), .B(n4075), .Z(n4076) );
  AND U4878 ( .A(x[32]), .B(y[193]), .Z(n4100) );
  NAND U4879 ( .A(x[17]), .B(y[112]), .Z(n4099) );
  XOR U4880 ( .A(n4100), .B(n4099), .Z(n4077) );
  XOR U4881 ( .A(n4076), .B(n4077), .Z(n4087) );
  AND U4882 ( .A(x[8]), .B(y[73]), .Z(n4309) );
  AND U4883 ( .A(x[24]), .B(y[153]), .Z(n4092) );
  XOR U4884 ( .A(n4309), .B(n4092), .Z(n4094) );
  AND U4885 ( .A(x[25]), .B(y[152]), .Z(n4093) );
  XNOR U4886 ( .A(n4094), .B(n4093), .Z(n4086) );
  XOR U4887 ( .A(n4087), .B(n4086), .Z(n4089) );
  XOR U4888 ( .A(n4088), .B(n4089), .Z(n4083) );
  NAND U4889 ( .A(n4066), .B(n4065), .Z(n4069) );
  AND U4890 ( .A(n4070), .B(n4067), .Z(n4068) );
  ANDN U4891 ( .B(n4069), .A(n4068), .Z(n4080) );
  XNOR U4892 ( .A(n4081), .B(n4080), .Z(n4082) );
  XNOR U4893 ( .A(n4083), .B(n4082), .Z(o[33]) );
  AND U4894 ( .A(x[1]), .B(y[33]), .Z(n4122) );
  NAND U4895 ( .A(n4122), .B(n4070), .Z(n4074) );
  NANDN U4896 ( .A(n4072), .B(n4071), .Z(n4073) );
  NAND U4897 ( .A(n4074), .B(n4073), .Z(n4142) );
  NANDN U4898 ( .A(n4075), .B(n4285), .Z(n4079) );
  NANDN U4899 ( .A(n4077), .B(n4076), .Z(n4078) );
  NAND U4900 ( .A(n4079), .B(n4078), .Z(n4140) );
  AND U4901 ( .A(x[24]), .B(y[154]), .Z(n4146) );
  NAND U4902 ( .A(x[0]), .B(y[34]), .Z(n4147) );
  XNOR U4903 ( .A(n4146), .B(n4147), .Z(n4149) );
  AND U4904 ( .A(x[10]), .B(y[72]), .Z(n4148) );
  XOR U4905 ( .A(n4149), .B(n4148), .Z(n4141) );
  XOR U4906 ( .A(n4140), .B(n4141), .Z(n4143) );
  XNOR U4907 ( .A(n4142), .B(n4143), .Z(n4102) );
  NANDN U4908 ( .A(n4081), .B(n4080), .Z(n4085) );
  NAND U4909 ( .A(n4083), .B(n4082), .Z(n4084) );
  NAND U4910 ( .A(n4085), .B(n4084), .Z(n4101) );
  XOR U4911 ( .A(n4102), .B(n4101), .Z(n4104) );
  NAND U4912 ( .A(n4087), .B(n4086), .Z(n4091) );
  NAND U4913 ( .A(n4089), .B(n4088), .Z(n4090) );
  AND U4914 ( .A(n4091), .B(n4090), .Z(n4110) );
  AND U4915 ( .A(x[2]), .B(y[32]), .Z(n4120) );
  AND U4916 ( .A(x[16]), .B(y[114]), .Z(n4119) );
  XOR U4917 ( .A(n4120), .B(n4119), .Z(n4121) );
  XOR U4918 ( .A(n4122), .B(n4121), .Z(n4155) );
  AND U4919 ( .A(x[26]), .B(y[152]), .Z(n4154) );
  XOR U4920 ( .A(n4155), .B(n4154), .Z(n4157) );
  AND U4921 ( .A(x[18]), .B(y[112]), .Z(n4223) );
  AND U4922 ( .A(x[32]), .B(y[194]), .Z(n4132) );
  XOR U4923 ( .A(n4223), .B(n4132), .Z(n4134) );
  AND U4924 ( .A(x[17]), .B(y[113]), .Z(n4133) );
  XOR U4925 ( .A(n4134), .B(n4133), .Z(n4156) );
  XOR U4926 ( .A(n4157), .B(n4156), .Z(n4107) );
  AND U4927 ( .A(n4309), .B(n4092), .Z(n4096) );
  NAND U4928 ( .A(n4094), .B(n4093), .Z(n4095) );
  NANDN U4929 ( .A(n4096), .B(n4095), .Z(n4115) );
  AND U4930 ( .A(y[192]), .B(x[34]), .Z(n4098) );
  NAND U4931 ( .A(y[193]), .B(x[33]), .Z(n4097) );
  XNOR U4932 ( .A(n4098), .B(n4097), .Z(n4153) );
  ANDN U4933 ( .B(n4100), .A(n4099), .Z(n4152) );
  XOR U4934 ( .A(n4153), .B(n4152), .Z(n4114) );
  AND U4935 ( .A(x[25]), .B(y[153]), .Z(n4125) );
  NAND U4936 ( .A(x[9]), .B(y[73]), .Z(n4126) );
  XNOR U4937 ( .A(n4125), .B(n4126), .Z(n4127) );
  NAND U4938 ( .A(x[8]), .B(y[74]), .Z(n4128) );
  XNOR U4939 ( .A(n4127), .B(n4128), .Z(n4113) );
  XOR U4940 ( .A(n4114), .B(n4113), .Z(n4116) );
  XOR U4941 ( .A(n4115), .B(n4116), .Z(n4108) );
  XOR U4942 ( .A(n4107), .B(n4108), .Z(n4109) );
  XNOR U4943 ( .A(n4110), .B(n4109), .Z(n4103) );
  XNOR U4944 ( .A(n4104), .B(n4103), .Z(o[34]) );
  NAND U4945 ( .A(n4102), .B(n4101), .Z(n4106) );
  NAND U4946 ( .A(n4104), .B(n4103), .Z(n4105) );
  AND U4947 ( .A(n4106), .B(n4105), .Z(n4161) );
  NAND U4948 ( .A(n4108), .B(n4107), .Z(n4112) );
  NAND U4949 ( .A(n4110), .B(n4109), .Z(n4111) );
  NAND U4950 ( .A(n4112), .B(n4111), .Z(n4166) );
  NAND U4951 ( .A(n4114), .B(n4113), .Z(n4118) );
  NAND U4952 ( .A(n4116), .B(n4115), .Z(n4117) );
  NAND U4953 ( .A(n4118), .B(n4117), .Z(n4164) );
  NAND U4954 ( .A(n4120), .B(n4119), .Z(n4124) );
  NAND U4955 ( .A(n4122), .B(n4121), .Z(n4123) );
  NAND U4956 ( .A(n4124), .B(n4123), .Z(n4176) );
  NANDN U4957 ( .A(n4126), .B(n4125), .Z(n4130) );
  NANDN U4958 ( .A(n4128), .B(n4127), .Z(n4129) );
  AND U4959 ( .A(n4130), .B(n4129), .Z(n4213) );
  AND U4960 ( .A(x[24]), .B(y[155]), .Z(n4239) );
  AND U4961 ( .A(x[16]), .B(y[115]), .Z(n4238) );
  NAND U4962 ( .A(x[3]), .B(y[32]), .Z(n4237) );
  XOR U4963 ( .A(n4238), .B(n4237), .Z(n4240) );
  XOR U4964 ( .A(n4239), .B(n4240), .Z(n4211) );
  AND U4965 ( .A(y[113]), .B(x[18]), .Z(n4269) );
  NAND U4966 ( .A(y[112]), .B(x[19]), .Z(n4131) );
  XNOR U4967 ( .A(n4269), .B(n4131), .Z(n4224) );
  NAND U4968 ( .A(x[17]), .B(y[114]), .Z(n4225) );
  XNOR U4969 ( .A(n4211), .B(n4210), .Z(n4212) );
  XNOR U4970 ( .A(n4213), .B(n4212), .Z(n4177) );
  XOR U4971 ( .A(n4176), .B(n4177), .Z(n4179) );
  NAND U4972 ( .A(n4223), .B(n4132), .Z(n4136) );
  AND U4973 ( .A(n4134), .B(n4133), .Z(n4135) );
  ANDN U4974 ( .B(n4136), .A(n4135), .Z(n4218) );
  AND U4975 ( .A(x[1]), .B(y[34]), .Z(n4190) );
  AND U4976 ( .A(x[2]), .B(y[33]), .Z(n4189) );
  NAND U4977 ( .A(x[25]), .B(y[154]), .Z(n4188) );
  XOR U4978 ( .A(n4189), .B(n4188), .Z(n4191) );
  XOR U4979 ( .A(n4190), .B(n4191), .Z(n4217) );
  AND U4980 ( .A(y[195]), .B(x[32]), .Z(n4138) );
  NAND U4981 ( .A(y[192]), .B(x[35]), .Z(n4137) );
  XNOR U4982 ( .A(n4138), .B(n4137), .Z(n4195) );
  AND U4983 ( .A(y[193]), .B(x[34]), .Z(n4282) );
  NAND U4984 ( .A(y[194]), .B(x[33]), .Z(n4139) );
  XOR U4985 ( .A(n4282), .B(n4139), .Z(n4196) );
  XNOR U4986 ( .A(n4195), .B(n4196), .Z(n4216) );
  XOR U4987 ( .A(n4217), .B(n4216), .Z(n4219) );
  XOR U4988 ( .A(n4218), .B(n4219), .Z(n4178) );
  XOR U4989 ( .A(n4179), .B(n4178), .Z(n4165) );
  XOR U4990 ( .A(n4164), .B(n4165), .Z(n4167) );
  XOR U4991 ( .A(n4166), .B(n4167), .Z(n4160) );
  XOR U4992 ( .A(n4161), .B(n4160), .Z(n4163) );
  NAND U4993 ( .A(n4141), .B(n4140), .Z(n4145) );
  NAND U4994 ( .A(n4143), .B(n4142), .Z(n4144) );
  AND U4995 ( .A(n4145), .B(n4144), .Z(n4173) );
  NANDN U4996 ( .A(n4147), .B(n4146), .Z(n4151) );
  NAND U4997 ( .A(n4149), .B(n4148), .Z(n4150) );
  AND U4998 ( .A(n4151), .B(n4150), .Z(n4183) );
  XNOR U4999 ( .A(n4183), .B(n4182), .Z(n4185) );
  NAND U5000 ( .A(x[11]), .B(y[72]), .Z(n4232) );
  NAND U5001 ( .A(x[0]), .B(y[35]), .Z(n4230) );
  NAND U5002 ( .A(x[26]), .B(y[153]), .Z(n4231) );
  XNOR U5003 ( .A(n4230), .B(n4231), .Z(n4233) );
  XOR U5004 ( .A(n4232), .B(n4233), .Z(n4206) );
  NAND U5005 ( .A(x[8]), .B(y[75]), .Z(n4202) );
  NAND U5006 ( .A(x[10]), .B(y[73]), .Z(n4200) );
  NAND U5007 ( .A(x[27]), .B(y[152]), .Z(n4201) );
  XNOR U5008 ( .A(n4200), .B(n4201), .Z(n4203) );
  XOR U5009 ( .A(n4202), .B(n4203), .Z(n4204) );
  AND U5010 ( .A(x[9]), .B(y[74]), .Z(n4205) );
  XOR U5011 ( .A(n4204), .B(n4205), .Z(n4207) );
  XOR U5012 ( .A(n4206), .B(n4207), .Z(n4184) );
  XNOR U5013 ( .A(n4185), .B(n4184), .Z(n4171) );
  NAND U5014 ( .A(n4155), .B(n4154), .Z(n4159) );
  NAND U5015 ( .A(n4157), .B(n4156), .Z(n4158) );
  AND U5016 ( .A(n4159), .B(n4158), .Z(n4170) );
  XOR U5017 ( .A(n4171), .B(n4170), .Z(n4172) );
  XNOR U5018 ( .A(n4173), .B(n4172), .Z(n4162) );
  XOR U5019 ( .A(n4163), .B(n4162), .Z(o[35]) );
  NAND U5020 ( .A(n4165), .B(n4164), .Z(n4169) );
  NAND U5021 ( .A(n4167), .B(n4166), .Z(n4168) );
  AND U5022 ( .A(n4169), .B(n4168), .Z(n4249) );
  NAND U5023 ( .A(n4171), .B(n4170), .Z(n4175) );
  NAND U5024 ( .A(n4173), .B(n4172), .Z(n4174) );
  NAND U5025 ( .A(n4175), .B(n4174), .Z(n4247) );
  NAND U5026 ( .A(n4177), .B(n4176), .Z(n4181) );
  NAND U5027 ( .A(n4179), .B(n4178), .Z(n4180) );
  AND U5028 ( .A(n4181), .B(n4180), .Z(n4248) );
  XOR U5029 ( .A(n4247), .B(n4248), .Z(n4250) );
  XOR U5030 ( .A(n4249), .B(n4250), .Z(n4243) );
  XOR U5031 ( .A(n4244), .B(n4243), .Z(n4246) );
  AND U5032 ( .A(x[10]), .B(y[74]), .Z(n4376) );
  AND U5033 ( .A(y[76]), .B(x[8]), .Z(n4187) );
  AND U5034 ( .A(y[73]), .B(x[11]), .Z(n4186) );
  XOR U5035 ( .A(n4187), .B(n4186), .Z(n4310) );
  XOR U5036 ( .A(n4376), .B(n4310), .Z(n4316) );
  AND U5037 ( .A(x[9]), .B(y[75]), .Z(n4315) );
  XOR U5038 ( .A(n4316), .B(n4315), .Z(n4318) );
  AND U5039 ( .A(x[28]), .B(y[152]), .Z(n4275) );
  AND U5040 ( .A(x[1]), .B(y[35]), .Z(n4274) );
  XOR U5041 ( .A(n4275), .B(n4274), .Z(n4277) );
  AND U5042 ( .A(x[0]), .B(y[36]), .Z(n4276) );
  XOR U5043 ( .A(n4277), .B(n4276), .Z(n4317) );
  XOR U5044 ( .A(n4318), .B(n4317), .Z(n4314) );
  NANDN U5045 ( .A(n4189), .B(n4188), .Z(n4193) );
  OR U5046 ( .A(n4191), .B(n4190), .Z(n4192) );
  NAND U5047 ( .A(n4193), .B(n4192), .Z(n4311) );
  AND U5048 ( .A(x[35]), .B(y[195]), .Z(n4593) );
  NANDN U5049 ( .A(n4194), .B(n4593), .Z(n4198) );
  NANDN U5050 ( .A(n4196), .B(n4195), .Z(n4197) );
  AND U5051 ( .A(n4198), .B(n4197), .Z(n4312) );
  XOR U5052 ( .A(n4311), .B(n4312), .Z(n4313) );
  XNOR U5053 ( .A(n4314), .B(n4313), .Z(n4338) );
  AND U5054 ( .A(x[4]), .B(y[32]), .Z(n4295) );
  AND U5055 ( .A(x[26]), .B(y[154]), .Z(n4293) );
  NAND U5056 ( .A(x[16]), .B(y[116]), .Z(n4292) );
  XNOR U5057 ( .A(n4293), .B(n4292), .Z(n4294) );
  XNOR U5058 ( .A(n4295), .B(n4294), .Z(n4260) );
  AND U5059 ( .A(y[194]), .B(x[34]), .Z(n4236) );
  AND U5060 ( .A(x[33]), .B(y[193]), .Z(n4199) );
  NAND U5061 ( .A(n4236), .B(n4199), .Z(n4290) );
  NAND U5062 ( .A(x[32]), .B(y[196]), .Z(n4445) );
  NAND U5063 ( .A(x[20]), .B(y[112]), .Z(n4397) );
  XNOR U5064 ( .A(n4445), .B(n4397), .Z(n4291) );
  XOR U5065 ( .A(n4290), .B(n4291), .Z(n4259) );
  XNOR U5066 ( .A(n4260), .B(n4259), .Z(n4262) );
  XOR U5067 ( .A(n4262), .B(n4261), .Z(n4336) );
  NAND U5068 ( .A(n4205), .B(n4204), .Z(n4209) );
  NAND U5069 ( .A(n4207), .B(n4206), .Z(n4208) );
  AND U5070 ( .A(n4209), .B(n4208), .Z(n4335) );
  XNOR U5071 ( .A(n4338), .B(n4337), .Z(n4253) );
  XNOR U5072 ( .A(n4254), .B(n4253), .Z(n4256) );
  NANDN U5073 ( .A(n4211), .B(n4210), .Z(n4215) );
  NANDN U5074 ( .A(n4213), .B(n4212), .Z(n4214) );
  AND U5075 ( .A(n4215), .B(n4214), .Z(n4324) );
  NANDN U5076 ( .A(n4217), .B(n4216), .Z(n4221) );
  OR U5077 ( .A(n4219), .B(n4218), .Z(n4220) );
  NAND U5078 ( .A(n4221), .B(n4220), .Z(n4323) );
  AND U5079 ( .A(x[19]), .B(y[113]), .Z(n4222) );
  NAND U5080 ( .A(n4223), .B(n4222), .Z(n4227) );
  NANDN U5081 ( .A(n4225), .B(n4224), .Z(n4226) );
  AND U5082 ( .A(n4227), .B(n4226), .Z(n4330) );
  AND U5083 ( .A(x[12]), .B(y[72]), .Z(n4279) );
  AND U5084 ( .A(x[24]), .B(y[156]), .Z(n4278) );
  XOR U5085 ( .A(n4279), .B(n4278), .Z(n4281) );
  AND U5086 ( .A(x[25]), .B(y[155]), .Z(n4280) );
  XOR U5087 ( .A(n4281), .B(n4280), .Z(n4320) );
  AND U5088 ( .A(y[114]), .B(x[18]), .Z(n4229) );
  NAND U5089 ( .A(y[113]), .B(x[19]), .Z(n4228) );
  XNOR U5090 ( .A(n4229), .B(n4228), .Z(n4271) );
  AND U5091 ( .A(x[17]), .B(y[115]), .Z(n4270) );
  XOR U5092 ( .A(n4271), .B(n4270), .Z(n4319) );
  XOR U5093 ( .A(n4320), .B(n4319), .Z(n4322) );
  XOR U5094 ( .A(n4322), .B(n4321), .Z(n4329) );
  NAND U5095 ( .A(x[2]), .B(y[34]), .Z(n4305) );
  NAND U5096 ( .A(x[27]), .B(y[153]), .Z(n4304) );
  NAND U5097 ( .A(x[3]), .B(y[33]), .Z(n4303) );
  XOR U5098 ( .A(n4304), .B(n4303), .Z(n4306) );
  XOR U5099 ( .A(n4305), .B(n4306), .Z(n4266) );
  AND U5100 ( .A(y[195]), .B(x[33]), .Z(n4235) );
  NAND U5101 ( .A(y[192]), .B(x[36]), .Z(n4234) );
  XNOR U5102 ( .A(n4235), .B(n4234), .Z(n4286) );
  AND U5103 ( .A(x[35]), .B(y[193]), .Z(n4403) );
  XNOR U5104 ( .A(n4403), .B(n4236), .Z(n4287) );
  XNOR U5105 ( .A(n4286), .B(n4287), .Z(n4265) );
  XNOR U5106 ( .A(n4266), .B(n4265), .Z(n4268) );
  NANDN U5107 ( .A(n4238), .B(n4237), .Z(n4242) );
  OR U5108 ( .A(n4240), .B(n4239), .Z(n4241) );
  AND U5109 ( .A(n4242), .B(n4241), .Z(n4267) );
  XOR U5110 ( .A(n4268), .B(n4267), .Z(n4331) );
  XOR U5111 ( .A(n4332), .B(n4331), .Z(n4325) );
  XOR U5112 ( .A(n4326), .B(n4325), .Z(n4255) );
  XNOR U5113 ( .A(n4256), .B(n4255), .Z(n4245) );
  XNOR U5114 ( .A(n4246), .B(n4245), .Z(o[36]) );
  NAND U5115 ( .A(n4248), .B(n4247), .Z(n4252) );
  NAND U5116 ( .A(n4250), .B(n4249), .Z(n4251) );
  NAND U5117 ( .A(n4252), .B(n4251), .Z(n4476) );
  XNOR U5118 ( .A(n4475), .B(n4476), .Z(n4478) );
  NANDN U5119 ( .A(n4254), .B(n4253), .Z(n4258) );
  NAND U5120 ( .A(n4256), .B(n4255), .Z(n4257) );
  AND U5121 ( .A(n4258), .B(n4257), .Z(n4342) );
  NANDN U5122 ( .A(n4260), .B(n4259), .Z(n4264) );
  NAND U5123 ( .A(n4262), .B(n4261), .Z(n4263) );
  NAND U5124 ( .A(n4264), .B(n4263), .Z(n4345) );
  XOR U5125 ( .A(n4345), .B(n4346), .Z(n4349) );
  AND U5126 ( .A(x[19]), .B(y[114]), .Z(n4399) );
  NAND U5127 ( .A(n4269), .B(n4399), .Z(n4273) );
  NAND U5128 ( .A(n4271), .B(n4270), .Z(n4272) );
  NAND U5129 ( .A(n4273), .B(n4272), .Z(n4405) );
  AND U5130 ( .A(x[13]), .B(y[72]), .Z(n4388) );
  AND U5131 ( .A(x[18]), .B(y[115]), .Z(n4387) );
  XOR U5132 ( .A(n4388), .B(n4387), .Z(n4389) );
  AND U5133 ( .A(x[24]), .B(y[157]), .Z(n4643) );
  XOR U5134 ( .A(n4389), .B(n4643), .Z(n4381) );
  AND U5135 ( .A(x[28]), .B(y[153]), .Z(n4393) );
  AND U5136 ( .A(x[5]), .B(y[32]), .Z(n4392) );
  XOR U5137 ( .A(n4393), .B(n4392), .Z(n4394) );
  AND U5138 ( .A(x[4]), .B(y[33]), .Z(n4703) );
  XNOR U5139 ( .A(n4394), .B(n4703), .Z(n4382) );
  XNOR U5140 ( .A(n4381), .B(n4382), .Z(n4383) );
  XNOR U5141 ( .A(n4384), .B(n4383), .Z(n4406) );
  XOR U5142 ( .A(n4405), .B(n4406), .Z(n4408) );
  AND U5143 ( .A(y[194]), .B(x[35]), .Z(n4300) );
  AND U5144 ( .A(n4282), .B(n4300), .Z(n4447) );
  AND U5145 ( .A(y[197]), .B(x[32]), .Z(n4284) );
  AND U5146 ( .A(y[196]), .B(x[33]), .Z(n4283) );
  XOR U5147 ( .A(n4284), .B(n4283), .Z(n4446) );
  XOR U5148 ( .A(n4447), .B(n4446), .Z(n4440) );
  AND U5149 ( .A(x[12]), .B(y[73]), .Z(n4432) );
  AND U5150 ( .A(x[8]), .B(y[77]), .Z(n4430) );
  AND U5151 ( .A(x[1]), .B(y[36]), .Z(n4429) );
  XOR U5152 ( .A(n4430), .B(n4429), .Z(n4431) );
  XOR U5153 ( .A(n4432), .B(n4431), .Z(n4439) );
  XOR U5154 ( .A(n4440), .B(n4439), .Z(n4442) );
  XOR U5155 ( .A(n4441), .B(n4442), .Z(n4407) );
  XOR U5156 ( .A(n4408), .B(n4407), .Z(n4348) );
  XOR U5157 ( .A(n4349), .B(n4348), .Z(n4472) );
  AND U5158 ( .A(x[36]), .B(y[195]), .Z(n4675) );
  NAND U5159 ( .A(n4675), .B(n4285), .Z(n4289) );
  NANDN U5160 ( .A(n4287), .B(n4286), .Z(n4288) );
  NAND U5161 ( .A(n4289), .B(n4288), .Z(n4361) );
  XOR U5162 ( .A(n4361), .B(n4362), .Z(n4364) );
  NANDN U5163 ( .A(n4293), .B(n4292), .Z(n4297) );
  NANDN U5164 ( .A(n4295), .B(n4294), .Z(n4296) );
  AND U5165 ( .A(n4297), .B(n4296), .Z(n4356) );
  AND U5166 ( .A(x[11]), .B(y[74]), .Z(n4523) );
  NAND U5167 ( .A(y[75]), .B(x[10]), .Z(n4298) );
  XNOR U5168 ( .A(n4523), .B(n4298), .Z(n4378) );
  AND U5169 ( .A(x[9]), .B(y[76]), .Z(n4377) );
  XOR U5170 ( .A(n4378), .B(n4377), .Z(n4354) );
  AND U5171 ( .A(x[34]), .B(y[195]), .Z(n4366) );
  AND U5172 ( .A(x[37]), .B(y[192]), .Z(n4365) );
  XOR U5173 ( .A(n4366), .B(n4365), .Z(n4368) );
  NAND U5174 ( .A(y[193]), .B(x[36]), .Z(n4299) );
  XNOR U5175 ( .A(n4300), .B(n4299), .Z(n4367) );
  XOR U5176 ( .A(n4368), .B(n4367), .Z(n4353) );
  XOR U5177 ( .A(n4354), .B(n4353), .Z(n4355) );
  XOR U5178 ( .A(n4356), .B(n4355), .Z(n4363) );
  XOR U5179 ( .A(n4364), .B(n4363), .Z(n4418) );
  AND U5180 ( .A(x[21]), .B(y[112]), .Z(n4302) );
  AND U5181 ( .A(y[113]), .B(x[20]), .Z(n4301) );
  XOR U5182 ( .A(n4302), .B(n4301), .Z(n4398) );
  XOR U5183 ( .A(n4399), .B(n4398), .Z(n4422) );
  AND U5184 ( .A(x[29]), .B(y[152]), .Z(n4372) );
  AND U5185 ( .A(x[3]), .B(y[34]), .Z(n4371) );
  XOR U5186 ( .A(n4372), .B(n4371), .Z(n4374) );
  AND U5187 ( .A(x[2]), .B(y[35]), .Z(n4373) );
  XOR U5188 ( .A(n4374), .B(n4373), .Z(n4421) );
  XOR U5189 ( .A(n4422), .B(n4421), .Z(n4424) );
  NAND U5190 ( .A(n4304), .B(n4303), .Z(n4308) );
  NAND U5191 ( .A(n4306), .B(n4305), .Z(n4307) );
  AND U5192 ( .A(n4308), .B(n4307), .Z(n4423) );
  XOR U5193 ( .A(n4424), .B(n4423), .Z(n4416) );
  AND U5194 ( .A(x[11]), .B(y[76]), .Z(n4674) );
  AND U5195 ( .A(x[27]), .B(y[154]), .Z(n4458) );
  AND U5196 ( .A(x[17]), .B(y[116]), .Z(n4689) );
  XOR U5197 ( .A(n4458), .B(n4689), .Z(n4460) );
  AND U5198 ( .A(x[16]), .B(y[117]), .Z(n4459) );
  XOR U5199 ( .A(n4460), .B(n4459), .Z(n4358) );
  AND U5200 ( .A(x[0]), .B(y[37]), .Z(n4451) );
  AND U5201 ( .A(x[25]), .B(y[156]), .Z(n4450) );
  XOR U5202 ( .A(n4451), .B(n4450), .Z(n4453) );
  AND U5203 ( .A(x[26]), .B(y[155]), .Z(n4452) );
  XOR U5204 ( .A(n4453), .B(n4452), .Z(n4357) );
  XOR U5205 ( .A(n4358), .B(n4357), .Z(n4360) );
  XOR U5206 ( .A(n4359), .B(n4360), .Z(n4415) );
  XOR U5207 ( .A(n4416), .B(n4415), .Z(n4417) );
  XOR U5208 ( .A(n4418), .B(n4417), .Z(n4469) );
  XNOR U5209 ( .A(n4411), .B(n4412), .Z(n4414) );
  XNOR U5210 ( .A(n4413), .B(n4414), .Z(n4470) );
  XOR U5211 ( .A(n4469), .B(n4470), .Z(n4471) );
  XOR U5212 ( .A(n4472), .B(n4471), .Z(n4341) );
  XNOR U5213 ( .A(n4342), .B(n4341), .Z(n4344) );
  NANDN U5214 ( .A(n4324), .B(n4323), .Z(n4328) );
  NAND U5215 ( .A(n4326), .B(n4325), .Z(n4327) );
  AND U5216 ( .A(n4328), .B(n4327), .Z(n4466) );
  NANDN U5217 ( .A(n4330), .B(n4329), .Z(n4334) );
  NAND U5218 ( .A(n4332), .B(n4331), .Z(n4333) );
  AND U5219 ( .A(n4334), .B(n4333), .Z(n4464) );
  NANDN U5220 ( .A(n4336), .B(n4335), .Z(n4340) );
  NAND U5221 ( .A(n4338), .B(n4337), .Z(n4339) );
  AND U5222 ( .A(n4340), .B(n4339), .Z(n4463) );
  XOR U5223 ( .A(n4344), .B(n4343), .Z(n4477) );
  XOR U5224 ( .A(n4478), .B(n4477), .Z(o[37]) );
  IV U5225 ( .A(n4345), .Z(n4347) );
  NANDN U5226 ( .A(n4347), .B(n4346), .Z(n4352) );
  IV U5227 ( .A(n4348), .Z(n4350) );
  NANDN U5228 ( .A(n4350), .B(n4349), .Z(n4351) );
  NAND U5229 ( .A(n4352), .B(n4351), .Z(n4481) );
  XOR U5230 ( .A(n4488), .B(n4487), .Z(n4485) );
  XOR U5231 ( .A(n4486), .B(n4485), .Z(n4484) );
  IV U5232 ( .A(n4484), .Z(n4404) );
  NAND U5233 ( .A(n4366), .B(n4365), .Z(n4370) );
  NAND U5234 ( .A(n4368), .B(n4367), .Z(n4369) );
  NAND U5235 ( .A(n4370), .B(n4369), .Z(n4628) );
  AND U5236 ( .A(x[11]), .B(y[75]), .Z(n4375) );
  NAND U5237 ( .A(n4376), .B(n4375), .Z(n4380) );
  NAND U5238 ( .A(n4378), .B(n4377), .Z(n4379) );
  AND U5239 ( .A(n4380), .B(n4379), .Z(n4723) );
  AND U5240 ( .A(x[27]), .B(y[155]), .Z(n4615) );
  AND U5241 ( .A(x[19]), .B(y[115]), .Z(n4614) );
  XOR U5242 ( .A(n4615), .B(n4614), .Z(n4613) );
  AND U5243 ( .A(x[3]), .B(y[35]), .Z(n4612) );
  XOR U5244 ( .A(n4613), .B(n4612), .Z(n4725) );
  AND U5245 ( .A(x[26]), .B(y[156]), .Z(n4649) );
  AND U5246 ( .A(x[20]), .B(y[114]), .Z(n4648) );
  XOR U5247 ( .A(n4649), .B(n4648), .Z(n4647) );
  AND U5248 ( .A(x[2]), .B(y[36]), .Z(n4646) );
  XNOR U5249 ( .A(n4647), .B(n4646), .Z(n4724) );
  XNOR U5250 ( .A(n4723), .B(n4722), .Z(n4630) );
  XOR U5251 ( .A(n4631), .B(n4630), .Z(n4629) );
  XOR U5252 ( .A(n4628), .B(n4629), .Z(n4492) );
  NANDN U5253 ( .A(n4382), .B(n4381), .Z(n4386) );
  NANDN U5254 ( .A(n4384), .B(n4383), .Z(n4385) );
  NAND U5255 ( .A(n4386), .B(n4385), .Z(n4491) );
  XOR U5256 ( .A(n4492), .B(n4491), .Z(n4490) );
  NAND U5257 ( .A(n4388), .B(n4387), .Z(n4391) );
  NAND U5258 ( .A(n4389), .B(n4643), .Z(n4390) );
  NAND U5259 ( .A(n4391), .B(n4390), .Z(n4512) );
  NAND U5260 ( .A(n4393), .B(n4392), .Z(n4396) );
  NAND U5261 ( .A(n4394), .B(n4703), .Z(n4395) );
  NAND U5262 ( .A(n4396), .B(n4395), .Z(n4511) );
  XOR U5263 ( .A(n4512), .B(n4511), .Z(n4510) );
  AND U5264 ( .A(x[21]), .B(y[113]), .Z(n4661) );
  AND U5265 ( .A(y[33]), .B(x[5]), .Z(n4401) );
  NAND U5266 ( .A(y[34]), .B(x[4]), .Z(n4400) );
  XNOR U5267 ( .A(n4401), .B(n4400), .Z(n4701) );
  AND U5268 ( .A(x[30]), .B(y[152]), .Z(n4700) );
  XOR U5269 ( .A(n4701), .B(n4700), .Z(n4637) );
  AND U5270 ( .A(x[33]), .B(y[197]), .Z(n4601) );
  AND U5271 ( .A(x[36]), .B(y[194]), .Z(n4402) );
  AND U5272 ( .A(n4403), .B(n4402), .Z(n4599) );
  AND U5273 ( .A(x[34]), .B(y[196]), .Z(n4598) );
  XOR U5274 ( .A(n4599), .B(n4598), .Z(n4600) );
  XNOR U5275 ( .A(n4601), .B(n4600), .Z(n4636) );
  XNOR U5276 ( .A(n4635), .B(n4634), .Z(n4509) );
  XOR U5277 ( .A(n4510), .B(n4509), .Z(n4489) );
  XOR U5278 ( .A(n4490), .B(n4489), .Z(n4483) );
  XOR U5279 ( .A(n4404), .B(n4483), .Z(n4482) );
  XOR U5280 ( .A(n4481), .B(n4482), .Z(n4765) );
  NAND U5281 ( .A(n4406), .B(n4405), .Z(n4410) );
  NAND U5282 ( .A(n4408), .B(n4407), .Z(n4409) );
  AND U5283 ( .A(n4410), .B(n4409), .Z(n4764) );
  OR U5284 ( .A(n4416), .B(n4415), .Z(n4420) );
  NANDN U5285 ( .A(n4418), .B(n4417), .Z(n4419) );
  NAND U5286 ( .A(n4420), .B(n4419), .Z(n4744) );
  NAND U5287 ( .A(n4422), .B(n4421), .Z(n4426) );
  NAND U5288 ( .A(n4424), .B(n4423), .Z(n4425) );
  AND U5289 ( .A(n4426), .B(n4425), .Z(n4749) );
  AND U5290 ( .A(x[16]), .B(y[118]), .Z(n4609) );
  AND U5291 ( .A(x[6]), .B(y[32]), .Z(n4608) );
  XOR U5292 ( .A(n4609), .B(n4608), .Z(n4607) );
  AND U5293 ( .A(x[29]), .B(y[153]), .Z(n4606) );
  XOR U5294 ( .A(n4607), .B(n4606), .Z(n4719) );
  AND U5295 ( .A(x[13]), .B(y[73]), .Z(n4697) );
  AND U5296 ( .A(x[10]), .B(y[76]), .Z(n4696) );
  XOR U5297 ( .A(n4697), .B(n4696), .Z(n4695) );
  AND U5298 ( .A(x[9]), .B(y[77]), .Z(n4694) );
  XOR U5299 ( .A(n4695), .B(n4694), .Z(n4522) );
  AND U5300 ( .A(y[74]), .B(x[12]), .Z(n4428) );
  NAND U5301 ( .A(y[75]), .B(x[11]), .Z(n4427) );
  XNOR U5302 ( .A(n4428), .B(n4427), .Z(n4521) );
  XOR U5303 ( .A(n4522), .B(n4521), .Z(n4718) );
  XOR U5304 ( .A(n4719), .B(n4718), .Z(n4717) );
  AND U5305 ( .A(x[32]), .B(y[198]), .Z(n4660) );
  XOR U5306 ( .A(n4661), .B(n4660), .Z(n4659) );
  AND U5307 ( .A(x[22]), .B(y[112]), .Z(n4658) );
  XOR U5308 ( .A(n4659), .B(n4658), .Z(n4716) );
  XOR U5309 ( .A(n4717), .B(n4716), .Z(n4501) );
  NAND U5310 ( .A(n4430), .B(n4429), .Z(n4434) );
  NAND U5311 ( .A(n4432), .B(n4431), .Z(n4433) );
  AND U5312 ( .A(n4434), .B(n4433), .Z(n4586) );
  AND U5313 ( .A(x[28]), .B(y[154]), .Z(n4687) );
  AND U5314 ( .A(x[18]), .B(y[116]), .Z(n4436) );
  AND U5315 ( .A(y[117]), .B(x[17]), .Z(n4435) );
  XOR U5316 ( .A(n4436), .B(n4435), .Z(n4686) );
  XOR U5317 ( .A(n4687), .B(n4686), .Z(n4589) );
  AND U5318 ( .A(x[0]), .B(y[38]), .Z(n4641) );
  AND U5319 ( .A(y[158]), .B(x[24]), .Z(n4438) );
  AND U5320 ( .A(y[157]), .B(x[25]), .Z(n4437) );
  XOR U5321 ( .A(n4438), .B(n4437), .Z(n4640) );
  XNOR U5322 ( .A(n4641), .B(n4640), .Z(n4588) );
  XNOR U5323 ( .A(n4586), .B(n4587), .Z(n4502) );
  XNOR U5324 ( .A(n4501), .B(n4502), .Z(n4504) );
  NAND U5325 ( .A(n4440), .B(n4439), .Z(n4444) );
  NAND U5326 ( .A(n4442), .B(n4441), .Z(n4443) );
  AND U5327 ( .A(n4444), .B(n4443), .Z(n4503) );
  XOR U5328 ( .A(n4504), .B(n4503), .Z(n4748) );
  XOR U5329 ( .A(n4749), .B(n4748), .Z(n4751) );
  NANDN U5330 ( .A(n4445), .B(n4601), .Z(n4449) );
  NAND U5331 ( .A(n4447), .B(n4446), .Z(n4448) );
  NAND U5332 ( .A(n4449), .B(n4448), .Z(n4498) );
  NAND U5333 ( .A(n4451), .B(n4450), .Z(n4455) );
  NAND U5334 ( .A(n4453), .B(n4452), .Z(n4454) );
  AND U5335 ( .A(n4455), .B(n4454), .Z(n4516) );
  AND U5336 ( .A(x[1]), .B(y[37]), .Z(n4683) );
  AND U5337 ( .A(x[14]), .B(y[72]), .Z(n4682) );
  XOR U5338 ( .A(n4683), .B(n4682), .Z(n4681) );
  AND U5339 ( .A(x[8]), .B(y[78]), .Z(n4680) );
  XOR U5340 ( .A(n4681), .B(n4680), .Z(n4518) );
  AND U5341 ( .A(y[193]), .B(x[37]), .Z(n4457) );
  NAND U5342 ( .A(y[194]), .B(x[36]), .Z(n4456) );
  XNOR U5343 ( .A(n4457), .B(n4456), .Z(n4595) );
  AND U5344 ( .A(x[38]), .B(y[192]), .Z(n4594) );
  XOR U5345 ( .A(n4595), .B(n4594), .Z(n4592) );
  XNOR U5346 ( .A(n4593), .B(n4592), .Z(n4517) );
  XNOR U5347 ( .A(n4516), .B(n4515), .Z(n4497) );
  XOR U5348 ( .A(n4498), .B(n4497), .Z(n4496) );
  NAND U5349 ( .A(n4458), .B(n4689), .Z(n4462) );
  NAND U5350 ( .A(n4460), .B(n4459), .Z(n4461) );
  NAND U5351 ( .A(n4462), .B(n4461), .Z(n4495) );
  XNOR U5352 ( .A(n4496), .B(n4495), .Z(n4750) );
  XOR U5353 ( .A(n4751), .B(n4750), .Z(n4745) );
  XNOR U5354 ( .A(n4744), .B(n4745), .Z(n4743) );
  XNOR U5355 ( .A(n4742), .B(n4743), .Z(n4762) );
  XOR U5356 ( .A(n4763), .B(n4762), .Z(n4769) );
  NANDN U5357 ( .A(n4464), .B(n4463), .Z(n4468) );
  NANDN U5358 ( .A(n4466), .B(n4465), .Z(n4467) );
  AND U5359 ( .A(n4468), .B(n4467), .Z(n4771) );
  NAND U5360 ( .A(n4470), .B(n4469), .Z(n4474) );
  NAND U5361 ( .A(n4472), .B(n4471), .Z(n4473) );
  NAND U5362 ( .A(n4474), .B(n4473), .Z(n4770) );
  NANDN U5363 ( .A(n4476), .B(n4475), .Z(n4480) );
  NAND U5364 ( .A(n4478), .B(n4477), .Z(n4479) );
  NAND U5365 ( .A(n4480), .B(n4479), .Z(n4756) );
  XOR U5366 ( .A(n4757), .B(n4756), .Z(o[38]) );
  NAND U5367 ( .A(n4490), .B(n4489), .Z(n4494) );
  NAND U5368 ( .A(n4492), .B(n4491), .Z(n4493) );
  AND U5369 ( .A(n4494), .B(n4493), .Z(n4741) );
  NAND U5370 ( .A(n4496), .B(n4495), .Z(n4500) );
  AND U5371 ( .A(n4498), .B(n4497), .Z(n4499) );
  ANDN U5372 ( .B(n4500), .A(n4499), .Z(n4508) );
  ANDN U5373 ( .B(n4502), .A(n4501), .Z(n4506) );
  AND U5374 ( .A(n4504), .B(n4503), .Z(n4505) );
  OR U5375 ( .A(n4506), .B(n4505), .Z(n4507) );
  XNOR U5376 ( .A(n4508), .B(n4507), .Z(n4739) );
  NAND U5377 ( .A(n4510), .B(n4509), .Z(n4514) );
  NAND U5378 ( .A(n4512), .B(n4511), .Z(n4513) );
  AND U5379 ( .A(n4514), .B(n4513), .Z(n4737) );
  NAND U5380 ( .A(n4516), .B(n4515), .Z(n4520) );
  NANDN U5381 ( .A(n4518), .B(n4517), .Z(n4519) );
  AND U5382 ( .A(n4520), .B(n4519), .Z(n4627) );
  NAND U5383 ( .A(n4522), .B(n4521), .Z(n4525) );
  AND U5384 ( .A(x[12]), .B(y[75]), .Z(n4575) );
  NAND U5385 ( .A(n4523), .B(n4575), .Z(n4524) );
  AND U5386 ( .A(n4525), .B(n4524), .Z(n4585) );
  AND U5387 ( .A(y[116]), .B(x[19]), .Z(n4527) );
  NAND U5388 ( .A(y[115]), .B(x[20]), .Z(n4526) );
  XNOR U5389 ( .A(n4527), .B(n4526), .Z(n4531) );
  AND U5390 ( .A(y[36]), .B(x[3]), .Z(n4529) );
  NAND U5391 ( .A(y[119]), .B(x[16]), .Z(n4528) );
  XNOR U5392 ( .A(n4529), .B(n4528), .Z(n4530) );
  XOR U5393 ( .A(n4531), .B(n4530), .Z(n4539) );
  AND U5394 ( .A(y[112]), .B(x[23]), .Z(n4533) );
  NAND U5395 ( .A(y[38]), .B(x[1]), .Z(n4532) );
  XNOR U5396 ( .A(n4533), .B(n4532), .Z(n4537) );
  AND U5397 ( .A(y[154]), .B(x[29]), .Z(n4535) );
  NAND U5398 ( .A(y[114]), .B(x[21]), .Z(n4534) );
  XNOR U5399 ( .A(n4535), .B(n4534), .Z(n4536) );
  XNOR U5400 ( .A(n4537), .B(n4536), .Z(n4538) );
  XNOR U5401 ( .A(n4539), .B(n4538), .Z(n4583) );
  AND U5402 ( .A(y[157]), .B(x[26]), .Z(n4544) );
  AND U5403 ( .A(x[37]), .B(y[194]), .Z(n4656) );
  AND U5404 ( .A(y[159]), .B(x[24]), .Z(n4541) );
  NAND U5405 ( .A(y[78]), .B(x[9]), .Z(n4540) );
  XNOR U5406 ( .A(n4541), .B(n4540), .Z(n4542) );
  XNOR U5407 ( .A(n4656), .B(n4542), .Z(n4543) );
  XNOR U5408 ( .A(n4544), .B(n4543), .Z(n4560) );
  AND U5409 ( .A(y[199]), .B(x[32]), .Z(n4546) );
  NAND U5410 ( .A(y[198]), .B(x[33]), .Z(n4545) );
  XNOR U5411 ( .A(n4546), .B(n4545), .Z(n4550) );
  AND U5412 ( .A(y[73]), .B(x[14]), .Z(n4548) );
  NAND U5413 ( .A(y[39]), .B(x[0]), .Z(n4547) );
  XNOR U5414 ( .A(n4548), .B(n4547), .Z(n4549) );
  XOR U5415 ( .A(n4550), .B(n4549), .Z(n4558) );
  AND U5416 ( .A(y[118]), .B(x[17]), .Z(n4552) );
  NAND U5417 ( .A(y[77]), .B(x[10]), .Z(n4551) );
  XNOR U5418 ( .A(n4552), .B(n4551), .Z(n4556) );
  AND U5419 ( .A(y[72]), .B(x[15]), .Z(n4554) );
  NAND U5420 ( .A(y[74]), .B(x[13]), .Z(n4553) );
  XNOR U5421 ( .A(n4554), .B(n4553), .Z(n4555) );
  XNOR U5422 ( .A(n4556), .B(n4555), .Z(n4557) );
  XNOR U5423 ( .A(n4558), .B(n4557), .Z(n4559) );
  XOR U5424 ( .A(n4560), .B(n4559), .Z(n4581) );
  AND U5425 ( .A(y[35]), .B(x[4]), .Z(n4562) );
  NAND U5426 ( .A(y[197]), .B(x[34]), .Z(n4561) );
  XNOR U5427 ( .A(n4562), .B(n4561), .Z(n4566) );
  AND U5428 ( .A(y[192]), .B(x[39]), .Z(n4564) );
  NAND U5429 ( .A(y[196]), .B(x[35]), .Z(n4563) );
  XNOR U5430 ( .A(n4564), .B(n4563), .Z(n4565) );
  XOR U5431 ( .A(n4566), .B(n4565), .Z(n4574) );
  AND U5432 ( .A(y[32]), .B(x[7]), .Z(n4568) );
  NAND U5433 ( .A(y[155]), .B(x[28]), .Z(n4567) );
  XNOR U5434 ( .A(n4568), .B(n4567), .Z(n4572) );
  AND U5435 ( .A(y[113]), .B(x[22]), .Z(n4570) );
  NAND U5436 ( .A(y[33]), .B(x[6]), .Z(n4569) );
  XNOR U5437 ( .A(n4570), .B(n4569), .Z(n4571) );
  XNOR U5438 ( .A(n4572), .B(n4571), .Z(n4573) );
  XNOR U5439 ( .A(n4574), .B(n4573), .Z(n4579) );
  AND U5440 ( .A(x[18]), .B(y[117]), .Z(n4688) );
  AND U5441 ( .A(x[25]), .B(y[158]), .Z(n4642) );
  XOR U5442 ( .A(n4688), .B(n4642), .Z(n4577) );
  AND U5443 ( .A(x[5]), .B(y[34]), .Z(n4702) );
  XNOR U5444 ( .A(n4702), .B(n4575), .Z(n4576) );
  XNOR U5445 ( .A(n4577), .B(n4576), .Z(n4578) );
  XNOR U5446 ( .A(n4579), .B(n4578), .Z(n4580) );
  XNOR U5447 ( .A(n4581), .B(n4580), .Z(n4582) );
  XNOR U5448 ( .A(n4583), .B(n4582), .Z(n4584) );
  XNOR U5449 ( .A(n4585), .B(n4584), .Z(n4625) );
  NANDN U5450 ( .A(n4587), .B(n4586), .Z(n4591) );
  NANDN U5451 ( .A(n4589), .B(n4588), .Z(n4590) );
  AND U5452 ( .A(n4591), .B(n4590), .Z(n4623) );
  NAND U5453 ( .A(n4593), .B(n4592), .Z(n4597) );
  AND U5454 ( .A(n4595), .B(n4594), .Z(n4596) );
  ANDN U5455 ( .B(n4597), .A(n4596), .Z(n4605) );
  AND U5456 ( .A(n4599), .B(n4598), .Z(n4603) );
  AND U5457 ( .A(n4601), .B(n4600), .Z(n4602) );
  OR U5458 ( .A(n4603), .B(n4602), .Z(n4604) );
  XNOR U5459 ( .A(n4605), .B(n4604), .Z(n4621) );
  NAND U5460 ( .A(n4607), .B(n4606), .Z(n4611) );
  NAND U5461 ( .A(n4609), .B(n4608), .Z(n4610) );
  AND U5462 ( .A(n4611), .B(n4610), .Z(n4619) );
  NAND U5463 ( .A(n4613), .B(n4612), .Z(n4617) );
  NAND U5464 ( .A(n4615), .B(n4614), .Z(n4616) );
  NAND U5465 ( .A(n4617), .B(n4616), .Z(n4618) );
  XNOR U5466 ( .A(n4619), .B(n4618), .Z(n4620) );
  XNOR U5467 ( .A(n4621), .B(n4620), .Z(n4622) );
  XNOR U5468 ( .A(n4623), .B(n4622), .Z(n4624) );
  XNOR U5469 ( .A(n4625), .B(n4624), .Z(n4626) );
  XNOR U5470 ( .A(n4627), .B(n4626), .Z(n4735) );
  NAND U5471 ( .A(n4629), .B(n4628), .Z(n4633) );
  NAND U5472 ( .A(n4631), .B(n4630), .Z(n4632) );
  AND U5473 ( .A(n4633), .B(n4632), .Z(n4733) );
  NAND U5474 ( .A(n4635), .B(n4634), .Z(n4639) );
  NANDN U5475 ( .A(n4637), .B(n4636), .Z(n4638) );
  AND U5476 ( .A(n4639), .B(n4638), .Z(n4715) );
  NAND U5477 ( .A(n4641), .B(n4640), .Z(n4645) );
  NAND U5478 ( .A(n4643), .B(n4642), .Z(n4644) );
  AND U5479 ( .A(n4645), .B(n4644), .Z(n4653) );
  NAND U5480 ( .A(n4647), .B(n4646), .Z(n4651) );
  NAND U5481 ( .A(n4649), .B(n4648), .Z(n4650) );
  NAND U5482 ( .A(n4651), .B(n4650), .Z(n4652) );
  XNOR U5483 ( .A(n4653), .B(n4652), .Z(n4713) );
  AND U5484 ( .A(y[153]), .B(x[30]), .Z(n4655) );
  NAND U5485 ( .A(y[156]), .B(x[27]), .Z(n4654) );
  XNOR U5486 ( .A(n4655), .B(n4654), .Z(n4679) );
  AND U5487 ( .A(x[36]), .B(y[193]), .Z(n4657) );
  AND U5488 ( .A(n4657), .B(n4656), .Z(n4673) );
  NAND U5489 ( .A(n4659), .B(n4658), .Z(n4663) );
  NAND U5490 ( .A(n4661), .B(n4660), .Z(n4662) );
  AND U5491 ( .A(n4663), .B(n4662), .Z(n4671) );
  AND U5492 ( .A(y[152]), .B(x[31]), .Z(n4665) );
  NAND U5493 ( .A(y[37]), .B(x[2]), .Z(n4664) );
  XNOR U5494 ( .A(n4665), .B(n4664), .Z(n4669) );
  AND U5495 ( .A(y[193]), .B(x[38]), .Z(n4667) );
  NAND U5496 ( .A(y[79]), .B(x[8]), .Z(n4666) );
  XNOR U5497 ( .A(n4667), .B(n4666), .Z(n4668) );
  XNOR U5498 ( .A(n4669), .B(n4668), .Z(n4670) );
  XNOR U5499 ( .A(n4671), .B(n4670), .Z(n4672) );
  XOR U5500 ( .A(n4673), .B(n4672), .Z(n4677) );
  XNOR U5501 ( .A(n4675), .B(n4674), .Z(n4676) );
  XNOR U5502 ( .A(n4677), .B(n4676), .Z(n4678) );
  XOR U5503 ( .A(n4679), .B(n4678), .Z(n4711) );
  NAND U5504 ( .A(n4681), .B(n4680), .Z(n4685) );
  NAND U5505 ( .A(n4683), .B(n4682), .Z(n4684) );
  AND U5506 ( .A(n4685), .B(n4684), .Z(n4693) );
  NAND U5507 ( .A(n4687), .B(n4686), .Z(n4691) );
  NAND U5508 ( .A(n4689), .B(n4688), .Z(n4690) );
  NAND U5509 ( .A(n4691), .B(n4690), .Z(n4692) );
  XNOR U5510 ( .A(n4693), .B(n4692), .Z(n4709) );
  NAND U5511 ( .A(n4695), .B(n4694), .Z(n4699) );
  NAND U5512 ( .A(n4697), .B(n4696), .Z(n4698) );
  AND U5513 ( .A(n4699), .B(n4698), .Z(n4707) );
  NAND U5514 ( .A(n4701), .B(n4700), .Z(n4705) );
  NAND U5515 ( .A(n4703), .B(n4702), .Z(n4704) );
  NAND U5516 ( .A(n4705), .B(n4704), .Z(n4706) );
  XNOR U5517 ( .A(n4707), .B(n4706), .Z(n4708) );
  XNOR U5518 ( .A(n4709), .B(n4708), .Z(n4710) );
  XNOR U5519 ( .A(n4711), .B(n4710), .Z(n4712) );
  XNOR U5520 ( .A(n4713), .B(n4712), .Z(n4714) );
  XNOR U5521 ( .A(n4715), .B(n4714), .Z(n4731) );
  NAND U5522 ( .A(n4717), .B(n4716), .Z(n4721) );
  NAND U5523 ( .A(n4719), .B(n4718), .Z(n4720) );
  AND U5524 ( .A(n4721), .B(n4720), .Z(n4729) );
  NAND U5525 ( .A(n4723), .B(n4722), .Z(n4727) );
  NANDN U5526 ( .A(n4725), .B(n4724), .Z(n4726) );
  NAND U5527 ( .A(n4727), .B(n4726), .Z(n4728) );
  XNOR U5528 ( .A(n4729), .B(n4728), .Z(n4730) );
  XNOR U5529 ( .A(n4731), .B(n4730), .Z(n4732) );
  XNOR U5530 ( .A(n4733), .B(n4732), .Z(n4734) );
  XNOR U5531 ( .A(n4735), .B(n4734), .Z(n4736) );
  XNOR U5532 ( .A(n4737), .B(n4736), .Z(n4738) );
  XNOR U5533 ( .A(n4739), .B(n4738), .Z(n4740) );
  NANDN U5534 ( .A(n4743), .B(n4742), .Z(n4747) );
  AND U5535 ( .A(n4745), .B(n4744), .Z(n4746) );
  ANDN U5536 ( .B(n4747), .A(n4746), .Z(n4755) );
  AND U5537 ( .A(n4749), .B(n4748), .Z(n4753) );
  AND U5538 ( .A(n4751), .B(n4750), .Z(n4752) );
  OR U5539 ( .A(n4753), .B(n4752), .Z(n4754) );
  NAND U5540 ( .A(n4757), .B(n4756), .Z(n4761) );
  NANDN U5541 ( .A(n4759), .B(n4758), .Z(n4760) );
  NAND U5542 ( .A(n4763), .B(n4762), .Z(n4767) );
  NANDN U5543 ( .A(n4765), .B(n4764), .Z(n4766) );
  NAND U5544 ( .A(y[160]), .B(x[72]), .Z(n4906) );
  NAND U5545 ( .A(y[40]), .B(x[48]), .Z(n4774) );
  XOR U5546 ( .A(n4906), .B(n4774), .Z(n4775) );
  AND U5547 ( .A(y[0]), .B(x[40]), .Z(n4782) );
  AND U5548 ( .A(y[80]), .B(x[56]), .Z(n4779) );
  XOR U5549 ( .A(n4782), .B(n4779), .Z(n4778) );
  AND U5550 ( .A(y[120]), .B(x[64]), .Z(n4777) );
  XNOR U5551 ( .A(n4778), .B(n4777), .Z(n4776) );
  XNOR U5552 ( .A(n4775), .B(n4776), .Z(o[40]) );
  AND U5553 ( .A(x[40]), .B(y[1]), .Z(n4773) );
  NAND U5554 ( .A(x[41]), .B(y[0]), .Z(n4772) );
  XNOR U5555 ( .A(n4773), .B(n4772), .Z(n4783) );
  NAND U5556 ( .A(y[40]), .B(x[49]), .Z(n4784) );
  XOR U5557 ( .A(n4783), .B(n4784), .Z(n4800) );
  AND U5558 ( .A(y[160]), .B(x[73]), .Z(n5005) );
  NAND U5559 ( .A(y[81]), .B(x[56]), .Z(n4787) );
  XNOR U5560 ( .A(n5005), .B(n4787), .Z(n4788) );
  AND U5561 ( .A(y[161]), .B(x[72]), .Z(n4811) );
  NAND U5562 ( .A(y[80]), .B(x[57]), .Z(n4810) );
  XOR U5563 ( .A(n4811), .B(n4810), .Z(n4789) );
  XOR U5564 ( .A(n4788), .B(n4789), .Z(n4799) );
  AND U5565 ( .A(y[41]), .B(x[48]), .Z(n5030) );
  AND U5566 ( .A(y[121]), .B(x[64]), .Z(n4804) );
  XOR U5567 ( .A(n5030), .B(n4804), .Z(n4806) );
  AND U5568 ( .A(y[120]), .B(x[65]), .Z(n4805) );
  XNOR U5569 ( .A(n4806), .B(n4805), .Z(n4798) );
  XOR U5570 ( .A(n4799), .B(n4798), .Z(n4801) );
  XOR U5571 ( .A(n4800), .B(n4801), .Z(n4795) );
  NAND U5572 ( .A(n4778), .B(n4777), .Z(n4781) );
  AND U5573 ( .A(n4782), .B(n4779), .Z(n4780) );
  ANDN U5574 ( .B(n4781), .A(n4780), .Z(n4792) );
  XNOR U5575 ( .A(n4793), .B(n4792), .Z(n4794) );
  XNOR U5576 ( .A(n4795), .B(n4794), .Z(o[41]) );
  AND U5577 ( .A(y[1]), .B(x[41]), .Z(n4833) );
  NAND U5578 ( .A(n4833), .B(n4782), .Z(n4786) );
  NANDN U5579 ( .A(n4784), .B(n4783), .Z(n4785) );
  NAND U5580 ( .A(n4786), .B(n4785), .Z(n4854) );
  NANDN U5581 ( .A(n4787), .B(n5005), .Z(n4791) );
  NANDN U5582 ( .A(n4789), .B(n4788), .Z(n4790) );
  NAND U5583 ( .A(n4791), .B(n4790), .Z(n4852) );
  AND U5584 ( .A(y[122]), .B(x[64]), .Z(n4858) );
  NAND U5585 ( .A(y[2]), .B(x[40]), .Z(n4859) );
  XNOR U5586 ( .A(n4858), .B(n4859), .Z(n4861) );
  AND U5587 ( .A(y[40]), .B(x[50]), .Z(n4860) );
  XOR U5588 ( .A(n4861), .B(n4860), .Z(n4853) );
  XOR U5589 ( .A(n4852), .B(n4853), .Z(n4855) );
  XNOR U5590 ( .A(n4854), .B(n4855), .Z(n4813) );
  NANDN U5591 ( .A(n4793), .B(n4792), .Z(n4797) );
  NAND U5592 ( .A(n4795), .B(n4794), .Z(n4796) );
  NAND U5593 ( .A(n4797), .B(n4796), .Z(n4812) );
  XOR U5594 ( .A(n4813), .B(n4812), .Z(n4815) );
  NAND U5595 ( .A(n4799), .B(n4798), .Z(n4803) );
  NAND U5596 ( .A(n4801), .B(n4800), .Z(n4802) );
  AND U5597 ( .A(n4803), .B(n4802), .Z(n4821) );
  AND U5598 ( .A(y[0]), .B(x[42]), .Z(n4831) );
  AND U5599 ( .A(y[82]), .B(x[56]), .Z(n4830) );
  XOR U5600 ( .A(n4831), .B(n4830), .Z(n4832) );
  XOR U5601 ( .A(n4833), .B(n4832), .Z(n4867) );
  AND U5602 ( .A(y[120]), .B(x[66]), .Z(n4866) );
  XOR U5603 ( .A(n4867), .B(n4866), .Z(n4869) );
  AND U5604 ( .A(y[80]), .B(x[58]), .Z(n4936) );
  AND U5605 ( .A(y[162]), .B(x[72]), .Z(n4843) );
  XOR U5606 ( .A(n4936), .B(n4843), .Z(n4845) );
  AND U5607 ( .A(y[81]), .B(x[57]), .Z(n4844) );
  XOR U5608 ( .A(n4845), .B(n4844), .Z(n4868) );
  XOR U5609 ( .A(n4869), .B(n4868), .Z(n4818) );
  AND U5610 ( .A(n5030), .B(n4804), .Z(n4808) );
  NAND U5611 ( .A(n4806), .B(n4805), .Z(n4807) );
  NANDN U5612 ( .A(n4808), .B(n4807), .Z(n4826) );
  AND U5613 ( .A(x[73]), .B(y[161]), .Z(n4911) );
  NAND U5614 ( .A(x[74]), .B(y[160]), .Z(n4809) );
  XNOR U5615 ( .A(n4911), .B(n4809), .Z(n4865) );
  ANDN U5616 ( .B(n4811), .A(n4810), .Z(n4864) );
  XOR U5617 ( .A(n4865), .B(n4864), .Z(n4825) );
  AND U5618 ( .A(y[121]), .B(x[65]), .Z(n4836) );
  NAND U5619 ( .A(y[41]), .B(x[49]), .Z(n4837) );
  XNOR U5620 ( .A(n4836), .B(n4837), .Z(n4838) );
  NAND U5621 ( .A(y[42]), .B(x[48]), .Z(n4839) );
  XNOR U5622 ( .A(n4838), .B(n4839), .Z(n4824) );
  XOR U5623 ( .A(n4825), .B(n4824), .Z(n4827) );
  XOR U5624 ( .A(n4826), .B(n4827), .Z(n4819) );
  XOR U5625 ( .A(n4818), .B(n4819), .Z(n4820) );
  XNOR U5626 ( .A(n4821), .B(n4820), .Z(n4814) );
  XNOR U5627 ( .A(n4815), .B(n4814), .Z(o[42]) );
  NAND U5628 ( .A(n4813), .B(n4812), .Z(n4817) );
  NAND U5629 ( .A(n4815), .B(n4814), .Z(n4816) );
  AND U5630 ( .A(n4817), .B(n4816), .Z(n4873) );
  NAND U5631 ( .A(n4819), .B(n4818), .Z(n4823) );
  NAND U5632 ( .A(n4821), .B(n4820), .Z(n4822) );
  NAND U5633 ( .A(n4823), .B(n4822), .Z(n4878) );
  NAND U5634 ( .A(n4825), .B(n4824), .Z(n4829) );
  NAND U5635 ( .A(n4827), .B(n4826), .Z(n4828) );
  NAND U5636 ( .A(n4829), .B(n4828), .Z(n4876) );
  NAND U5637 ( .A(n4831), .B(n4830), .Z(n4835) );
  NAND U5638 ( .A(n4833), .B(n4832), .Z(n4834) );
  NAND U5639 ( .A(n4835), .B(n4834), .Z(n4888) );
  NANDN U5640 ( .A(n4837), .B(n4836), .Z(n4841) );
  NANDN U5641 ( .A(n4839), .B(n4838), .Z(n4840) );
  AND U5642 ( .A(n4841), .B(n4840), .Z(n4927) );
  AND U5643 ( .A(y[123]), .B(x[64]), .Z(n4952) );
  AND U5644 ( .A(y[83]), .B(x[56]), .Z(n4951) );
  NAND U5645 ( .A(y[0]), .B(x[43]), .Z(n4950) );
  XOR U5646 ( .A(n4951), .B(n4950), .Z(n4953) );
  XOR U5647 ( .A(n4952), .B(n4953), .Z(n4925) );
  AND U5648 ( .A(x[58]), .B(y[81]), .Z(n4985) );
  NAND U5649 ( .A(x[59]), .B(y[80]), .Z(n4842) );
  XNOR U5650 ( .A(n4985), .B(n4842), .Z(n4938) );
  NAND U5651 ( .A(y[82]), .B(x[57]), .Z(n4939) );
  XNOR U5652 ( .A(n4925), .B(n4924), .Z(n4926) );
  XNOR U5653 ( .A(n4927), .B(n4926), .Z(n4889) );
  XOR U5654 ( .A(n4888), .B(n4889), .Z(n4891) );
  NAND U5655 ( .A(n4936), .B(n4843), .Z(n4847) );
  AND U5656 ( .A(n4845), .B(n4844), .Z(n4846) );
  ANDN U5657 ( .B(n4847), .A(n4846), .Z(n4932) );
  AND U5658 ( .A(y[2]), .B(x[41]), .Z(n4902) );
  AND U5659 ( .A(y[1]), .B(x[42]), .Z(n4901) );
  NAND U5660 ( .A(y[122]), .B(x[65]), .Z(n4900) );
  XOR U5661 ( .A(n4901), .B(n4900), .Z(n4903) );
  XOR U5662 ( .A(n4902), .B(n4903), .Z(n4931) );
  AND U5663 ( .A(x[75]), .B(y[160]), .Z(n4849) );
  NAND U5664 ( .A(x[72]), .B(y[163]), .Z(n4848) );
  XNOR U5665 ( .A(n4849), .B(n4848), .Z(n4907) );
  AND U5666 ( .A(x[73]), .B(y[162]), .Z(n4851) );
  NAND U5667 ( .A(x[74]), .B(y[161]), .Z(n4850) );
  XOR U5668 ( .A(n4851), .B(n4850), .Z(n4908) );
  XNOR U5669 ( .A(n4907), .B(n4908), .Z(n4930) );
  XOR U5670 ( .A(n4931), .B(n4930), .Z(n4933) );
  XOR U5671 ( .A(n4932), .B(n4933), .Z(n4890) );
  XOR U5672 ( .A(n4891), .B(n4890), .Z(n4877) );
  XOR U5673 ( .A(n4876), .B(n4877), .Z(n4879) );
  XOR U5674 ( .A(n4878), .B(n4879), .Z(n4872) );
  XOR U5675 ( .A(n4873), .B(n4872), .Z(n4875) );
  NAND U5676 ( .A(n4853), .B(n4852), .Z(n4857) );
  NAND U5677 ( .A(n4855), .B(n4854), .Z(n4856) );
  AND U5678 ( .A(n4857), .B(n4856), .Z(n4885) );
  NANDN U5679 ( .A(n4859), .B(n4858), .Z(n4863) );
  NAND U5680 ( .A(n4861), .B(n4860), .Z(n4862) );
  AND U5681 ( .A(n4863), .B(n4862), .Z(n4895) );
  AND U5682 ( .A(y[161]), .B(x[74]), .Z(n5002) );
  XNOR U5683 ( .A(n4895), .B(n4894), .Z(n4897) );
  AND U5684 ( .A(y[40]), .B(x[51]), .Z(n4946) );
  AND U5685 ( .A(y[3]), .B(x[40]), .Z(n4945) );
  NAND U5686 ( .A(y[121]), .B(x[66]), .Z(n4944) );
  XOR U5687 ( .A(n4945), .B(n4944), .Z(n4947) );
  XOR U5688 ( .A(n4946), .B(n4947), .Z(n4921) );
  AND U5689 ( .A(y[43]), .B(x[48]), .Z(n4914) );
  AND U5690 ( .A(y[41]), .B(x[50]), .Z(n4913) );
  NAND U5691 ( .A(y[120]), .B(x[67]), .Z(n4912) );
  XOR U5692 ( .A(n4913), .B(n4912), .Z(n4915) );
  XOR U5693 ( .A(n4914), .B(n4915), .Z(n4919) );
  AND U5694 ( .A(y[42]), .B(x[49]), .Z(n4918) );
  XNOR U5695 ( .A(n4897), .B(n4896), .Z(n4883) );
  NAND U5696 ( .A(n4867), .B(n4866), .Z(n4871) );
  NAND U5697 ( .A(n4869), .B(n4868), .Z(n4870) );
  AND U5698 ( .A(n4871), .B(n4870), .Z(n4882) );
  XOR U5699 ( .A(n4883), .B(n4882), .Z(n4884) );
  XNOR U5700 ( .A(n4885), .B(n4884), .Z(n4874) );
  XOR U5701 ( .A(n4875), .B(n4874), .Z(o[43]) );
  NAND U5702 ( .A(n4877), .B(n4876), .Z(n4881) );
  NAND U5703 ( .A(n4879), .B(n4878), .Z(n4880) );
  AND U5704 ( .A(n4881), .B(n4880), .Z(n4965) );
  NAND U5705 ( .A(n4883), .B(n4882), .Z(n4887) );
  NAND U5706 ( .A(n4885), .B(n4884), .Z(n4886) );
  NAND U5707 ( .A(n4887), .B(n4886), .Z(n4963) );
  NAND U5708 ( .A(n4889), .B(n4888), .Z(n4893) );
  NAND U5709 ( .A(n4891), .B(n4890), .Z(n4892) );
  AND U5710 ( .A(n4893), .B(n4892), .Z(n4964) );
  XOR U5711 ( .A(n4963), .B(n4964), .Z(n4966) );
  XOR U5712 ( .A(n4965), .B(n4966), .Z(n4959) );
  XOR U5713 ( .A(n4960), .B(n4959), .Z(n4962) );
  AND U5714 ( .A(y[42]), .B(x[50]), .Z(n5098) );
  AND U5715 ( .A(x[51]), .B(y[41]), .Z(n4899) );
  NAND U5716 ( .A(x[48]), .B(y[44]), .Z(n4898) );
  XOR U5717 ( .A(n4899), .B(n4898), .Z(n5031) );
  XNOR U5718 ( .A(n5098), .B(n5031), .Z(n5040) );
  NAND U5719 ( .A(y[43]), .B(x[49]), .Z(n5041) );
  XNOR U5720 ( .A(n5040), .B(n5041), .Z(n5043) );
  AND U5721 ( .A(y[120]), .B(x[68]), .Z(n4990) );
  NAND U5722 ( .A(y[3]), .B(x[41]), .Z(n4991) );
  XNOR U5723 ( .A(n4990), .B(n4991), .Z(n4992) );
  NAND U5724 ( .A(y[4]), .B(x[40]), .Z(n4993) );
  XNOR U5725 ( .A(n4992), .B(n4993), .Z(n5042) );
  XOR U5726 ( .A(n5043), .B(n5042), .Z(n5037) );
  NANDN U5727 ( .A(n4901), .B(n4900), .Z(n4905) );
  OR U5728 ( .A(n4903), .B(n4902), .Z(n4904) );
  AND U5729 ( .A(n4905), .B(n4904), .Z(n5035) );
  AND U5730 ( .A(y[163]), .B(x[75]), .Z(n5319) );
  NANDN U5731 ( .A(n4906), .B(n5319), .Z(n4910) );
  NANDN U5732 ( .A(n4908), .B(n4907), .Z(n4909) );
  AND U5733 ( .A(n4910), .B(n4909), .Z(n5034) );
  XNOR U5734 ( .A(n5035), .B(n5034), .Z(n5036) );
  XNOR U5735 ( .A(n5037), .B(n5036), .Z(n5067) );
  NAND U5736 ( .A(y[0]), .B(x[44]), .Z(n5014) );
  NAND U5737 ( .A(y[122]), .B(x[66]), .Z(n5013) );
  NAND U5738 ( .A(y[84]), .B(x[56]), .Z(n5012) );
  XOR U5739 ( .A(n5013), .B(n5012), .Z(n5015) );
  XNOR U5740 ( .A(n5014), .B(n5015), .Z(n4976) );
  AND U5741 ( .A(y[162]), .B(x[74]), .Z(n4958) );
  NAND U5742 ( .A(n4911), .B(n4958), .Z(n5010) );
  NAND U5743 ( .A(y[164]), .B(x[72]), .Z(n5171) );
  NAND U5744 ( .A(y[80]), .B(x[60]), .Z(n5113) );
  XNOR U5745 ( .A(n5171), .B(n5113), .Z(n5011) );
  XOR U5746 ( .A(n5010), .B(n5011), .Z(n4975) );
  XOR U5747 ( .A(n4976), .B(n4975), .Z(n4978) );
  NANDN U5748 ( .A(n4913), .B(n4912), .Z(n4917) );
  OR U5749 ( .A(n4915), .B(n4914), .Z(n4916) );
  AND U5750 ( .A(n4917), .B(n4916), .Z(n4977) );
  XOR U5751 ( .A(n4978), .B(n4977), .Z(n5065) );
  NANDN U5752 ( .A(n4919), .B(n4918), .Z(n4923) );
  NANDN U5753 ( .A(n4921), .B(n4920), .Z(n4922) );
  AND U5754 ( .A(n4923), .B(n4922), .Z(n5064) );
  XNOR U5755 ( .A(n5067), .B(n5066), .Z(n4969) );
  XNOR U5756 ( .A(n4970), .B(n4969), .Z(n4972) );
  NANDN U5757 ( .A(n4925), .B(n4924), .Z(n4929) );
  NANDN U5758 ( .A(n4927), .B(n4926), .Z(n4928) );
  AND U5759 ( .A(n4929), .B(n4928), .Z(n5053) );
  NANDN U5760 ( .A(n4931), .B(n4930), .Z(n4935) );
  OR U5761 ( .A(n4933), .B(n4932), .Z(n4934) );
  NAND U5762 ( .A(n4935), .B(n4934), .Z(n5052) );
  AND U5763 ( .A(y[81]), .B(x[59]), .Z(n4937) );
  NAND U5764 ( .A(n4937), .B(n4936), .Z(n4941) );
  NANDN U5765 ( .A(n4939), .B(n4938), .Z(n4940) );
  AND U5766 ( .A(n4941), .B(n4940), .Z(n5059) );
  AND U5767 ( .A(y[40]), .B(x[52]), .Z(n4996) );
  NAND U5768 ( .A(y[124]), .B(x[64]), .Z(n4997) );
  XNOR U5769 ( .A(n4996), .B(n4997), .Z(n4998) );
  NAND U5770 ( .A(y[123]), .B(x[65]), .Z(n4999) );
  XNOR U5771 ( .A(n4998), .B(n4999), .Z(n5046) );
  AND U5772 ( .A(x[58]), .B(y[82]), .Z(n4943) );
  NAND U5773 ( .A(x[59]), .B(y[81]), .Z(n4942) );
  XNOR U5774 ( .A(n4943), .B(n4942), .Z(n4986) );
  NAND U5775 ( .A(y[83]), .B(x[57]), .Z(n4987) );
  XOR U5776 ( .A(n4986), .B(n4987), .Z(n5047) );
  XNOR U5777 ( .A(n5046), .B(n5047), .Z(n5048) );
  NANDN U5778 ( .A(n4945), .B(n4944), .Z(n4949) );
  OR U5779 ( .A(n4947), .B(n4946), .Z(n4948) );
  NAND U5780 ( .A(n4949), .B(n4948), .Z(n5049) );
  XNOR U5781 ( .A(n5048), .B(n5049), .Z(n5058) );
  NAND U5782 ( .A(y[2]), .B(x[42]), .Z(n5026) );
  NAND U5783 ( .A(y[121]), .B(x[67]), .Z(n5025) );
  NAND U5784 ( .A(y[1]), .B(x[43]), .Z(n5024) );
  XNOR U5785 ( .A(n5025), .B(n5024), .Z(n5027) );
  NANDN U5786 ( .A(n4951), .B(n4950), .Z(n4955) );
  OR U5787 ( .A(n4953), .B(n4952), .Z(n4954) );
  AND U5788 ( .A(n4955), .B(n4954), .Z(n4981) );
  XOR U5789 ( .A(n4982), .B(n4981), .Z(n4984) );
  AND U5790 ( .A(x[76]), .B(y[160]), .Z(n4957) );
  NAND U5791 ( .A(x[73]), .B(y[163]), .Z(n4956) );
  XNOR U5792 ( .A(n4957), .B(n4956), .Z(n5007) );
  AND U5793 ( .A(y[161]), .B(x[75]), .Z(n5120) );
  XOR U5794 ( .A(n4958), .B(n5120), .Z(n5006) );
  XOR U5795 ( .A(n5007), .B(n5006), .Z(n4983) );
  XOR U5796 ( .A(n4984), .B(n4983), .Z(n5060) );
  XOR U5797 ( .A(n5061), .B(n5060), .Z(n5054) );
  XOR U5798 ( .A(n5055), .B(n5054), .Z(n4971) );
  XNOR U5799 ( .A(n4972), .B(n4971), .Z(n4961) );
  XNOR U5800 ( .A(n4962), .B(n4961), .Z(o[44]) );
  NAND U5801 ( .A(n4964), .B(n4963), .Z(n4968) );
  NAND U5802 ( .A(n4966), .B(n4965), .Z(n4967) );
  NAND U5803 ( .A(n4968), .B(n4967), .Z(n5209) );
  XNOR U5804 ( .A(n5208), .B(n5209), .Z(n5211) );
  NANDN U5805 ( .A(n4970), .B(n4969), .Z(n4974) );
  NAND U5806 ( .A(n4972), .B(n4971), .Z(n4973) );
  AND U5807 ( .A(n4974), .B(n4973), .Z(n5071) );
  NAND U5808 ( .A(n4976), .B(n4975), .Z(n4980) );
  NAND U5809 ( .A(n4978), .B(n4977), .Z(n4979) );
  AND U5810 ( .A(n4980), .B(n4979), .Z(n5132) );
  XNOR U5811 ( .A(n5132), .B(n5131), .Z(n5134) );
  AND U5812 ( .A(y[82]), .B(x[59]), .Z(n5114) );
  NAND U5813 ( .A(n5114), .B(n4985), .Z(n4989) );
  NANDN U5814 ( .A(n4987), .B(n4986), .Z(n4988) );
  AND U5815 ( .A(n4989), .B(n4988), .Z(n5087) );
  NANDN U5816 ( .A(n4991), .B(n4990), .Z(n4995) );
  NANDN U5817 ( .A(n4993), .B(n4992), .Z(n4994) );
  NAND U5818 ( .A(n4995), .B(n4994), .Z(n5111) );
  AND U5819 ( .A(y[125]), .B(x[64]), .Z(n5420) );
  AND U5820 ( .A(y[83]), .B(x[58]), .Z(n5127) );
  AND U5821 ( .A(y[40]), .B(x[53]), .Z(n5126) );
  XOR U5822 ( .A(n5127), .B(n5126), .Z(n5128) );
  XOR U5823 ( .A(n5420), .B(n5128), .Z(n5110) );
  AND U5824 ( .A(y[121]), .B(x[68]), .Z(n5122) );
  AND U5825 ( .A(y[0]), .B(x[45]), .Z(n5121) );
  XOR U5826 ( .A(n5122), .B(n5121), .Z(n5123) );
  AND U5827 ( .A(y[1]), .B(x[44]), .Z(n5426) );
  XOR U5828 ( .A(n5123), .B(n5426), .Z(n5109) );
  XOR U5829 ( .A(n5110), .B(n5109), .Z(n5112) );
  XOR U5830 ( .A(n5111), .B(n5112), .Z(n5086) );
  NANDN U5831 ( .A(n4997), .B(n4996), .Z(n5001) );
  NANDN U5832 ( .A(n4999), .B(n4998), .Z(n5000) );
  NAND U5833 ( .A(n5001), .B(n5000), .Z(n5204) );
  AND U5834 ( .A(y[162]), .B(x[75]), .Z(n5021) );
  AND U5835 ( .A(n5021), .B(n5002), .Z(n5173) );
  AND U5836 ( .A(x[72]), .B(y[165]), .Z(n5004) );
  AND U5837 ( .A(x[73]), .B(y[164]), .Z(n5003) );
  XOR U5838 ( .A(n5004), .B(n5003), .Z(n5172) );
  XOR U5839 ( .A(n5173), .B(n5172), .Z(n5203) );
  AND U5840 ( .A(y[41]), .B(x[52]), .Z(n5195) );
  AND U5841 ( .A(y[45]), .B(x[48]), .Z(n5193) );
  AND U5842 ( .A(y[4]), .B(x[41]), .Z(n5192) );
  XOR U5843 ( .A(n5193), .B(n5192), .Z(n5194) );
  XOR U5844 ( .A(n5195), .B(n5194), .Z(n5202) );
  XOR U5845 ( .A(n5203), .B(n5202), .Z(n5205) );
  XOR U5846 ( .A(n5204), .B(n5205), .Z(n5088) );
  XOR U5847 ( .A(n5089), .B(n5088), .Z(n5133) );
  XOR U5848 ( .A(n5134), .B(n5133), .Z(n5077) );
  AND U5849 ( .A(y[163]), .B(x[76]), .Z(n5412) );
  NAND U5850 ( .A(n5412), .B(n5005), .Z(n5009) );
  NAND U5851 ( .A(n5007), .B(n5006), .Z(n5008) );
  AND U5852 ( .A(n5009), .B(n5008), .Z(n5143) );
  XNOR U5853 ( .A(n5143), .B(n5142), .Z(n5145) );
  NAND U5854 ( .A(n5013), .B(n5012), .Z(n5017) );
  NAND U5855 ( .A(n5015), .B(n5014), .Z(n5016) );
  AND U5856 ( .A(n5017), .B(n5016), .Z(n5151) );
  AND U5857 ( .A(x[50]), .B(y[43]), .Z(n5019) );
  NAND U5858 ( .A(x[51]), .B(y[42]), .Z(n5018) );
  XNOR U5859 ( .A(n5019), .B(n5018), .Z(n5099) );
  NAND U5860 ( .A(y[44]), .B(x[49]), .Z(n5100) );
  XNOR U5861 ( .A(n5099), .B(n5100), .Z(n5149) );
  AND U5862 ( .A(y[163]), .B(x[74]), .Z(n5092) );
  NAND U5863 ( .A(y[160]), .B(x[77]), .Z(n5093) );
  XNOR U5864 ( .A(n5092), .B(n5093), .Z(n5094) );
  NAND U5865 ( .A(x[76]), .B(y[161]), .Z(n5020) );
  XOR U5866 ( .A(n5021), .B(n5020), .Z(n5095) );
  XNOR U5867 ( .A(n5094), .B(n5095), .Z(n5148) );
  XOR U5868 ( .A(n5149), .B(n5148), .Z(n5150) );
  XOR U5869 ( .A(n5151), .B(n5150), .Z(n5144) );
  XOR U5870 ( .A(n5145), .B(n5144), .Z(n5162) );
  AND U5871 ( .A(x[60]), .B(y[81]), .Z(n5023) );
  NAND U5872 ( .A(x[61]), .B(y[80]), .Z(n5022) );
  XOR U5873 ( .A(n5023), .B(n5022), .Z(n5115) );
  XNOR U5874 ( .A(n5114), .B(n5115), .Z(n5185) );
  AND U5875 ( .A(y[120]), .B(x[69]), .Z(n5103) );
  NAND U5876 ( .A(y[2]), .B(x[43]), .Z(n5104) );
  XNOR U5877 ( .A(n5103), .B(n5104), .Z(n5106) );
  AND U5878 ( .A(y[3]), .B(x[42]), .Z(n5105) );
  XOR U5879 ( .A(n5106), .B(n5105), .Z(n5184) );
  XOR U5880 ( .A(n5185), .B(n5184), .Z(n5187) );
  NAND U5881 ( .A(n5025), .B(n5024), .Z(n5029) );
  NANDN U5882 ( .A(n5027), .B(n5026), .Z(n5028) );
  AND U5883 ( .A(n5029), .B(n5028), .Z(n5186) );
  XOR U5884 ( .A(n5187), .B(n5186), .Z(n5161) );
  AND U5885 ( .A(y[44]), .B(x[51]), .Z(n5301) );
  NAND U5886 ( .A(n5301), .B(n5030), .Z(n5033) );
  NANDN U5887 ( .A(n5031), .B(n5098), .Z(n5032) );
  AND U5888 ( .A(n5033), .B(n5032), .Z(n5141) );
  AND U5889 ( .A(y[122]), .B(x[67]), .Z(n5166) );
  AND U5890 ( .A(y[84]), .B(x[57]), .Z(n5335) );
  XOR U5891 ( .A(n5166), .B(n5335), .Z(n5168) );
  AND U5892 ( .A(y[85]), .B(x[56]), .Z(n5167) );
  XOR U5893 ( .A(n5168), .B(n5167), .Z(n5139) );
  AND U5894 ( .A(y[5]), .B(x[40]), .Z(n5177) );
  AND U5895 ( .A(y[124]), .B(x[65]), .Z(n5176) );
  XOR U5896 ( .A(n5177), .B(n5176), .Z(n5179) );
  AND U5897 ( .A(y[123]), .B(x[66]), .Z(n5178) );
  XOR U5898 ( .A(n5179), .B(n5178), .Z(n5138) );
  XOR U5899 ( .A(n5139), .B(n5138), .Z(n5140) );
  XOR U5900 ( .A(n5141), .B(n5140), .Z(n5160) );
  XOR U5901 ( .A(n5161), .B(n5160), .Z(n5163) );
  XOR U5902 ( .A(n5162), .B(n5163), .Z(n5075) );
  NANDN U5903 ( .A(n5035), .B(n5034), .Z(n5039) );
  NANDN U5904 ( .A(n5037), .B(n5036), .Z(n5038) );
  AND U5905 ( .A(n5039), .B(n5038), .Z(n5156) );
  NANDN U5906 ( .A(n5041), .B(n5040), .Z(n5045) );
  NAND U5907 ( .A(n5043), .B(n5042), .Z(n5044) );
  AND U5908 ( .A(n5045), .B(n5044), .Z(n5155) );
  NANDN U5909 ( .A(n5047), .B(n5046), .Z(n5051) );
  NANDN U5910 ( .A(n5049), .B(n5048), .Z(n5050) );
  NAND U5911 ( .A(n5051), .B(n5050), .Z(n5154) );
  XOR U5912 ( .A(n5155), .B(n5154), .Z(n5157) );
  XNOR U5913 ( .A(n5156), .B(n5157), .Z(n5074) );
  XOR U5914 ( .A(n5077), .B(n5076), .Z(n5070) );
  XNOR U5915 ( .A(n5071), .B(n5070), .Z(n5073) );
  NANDN U5916 ( .A(n5053), .B(n5052), .Z(n5057) );
  NAND U5917 ( .A(n5055), .B(n5054), .Z(n5056) );
  AND U5918 ( .A(n5057), .B(n5056), .Z(n5083) );
  NANDN U5919 ( .A(n5059), .B(n5058), .Z(n5063) );
  NAND U5920 ( .A(n5061), .B(n5060), .Z(n5062) );
  AND U5921 ( .A(n5063), .B(n5062), .Z(n5081) );
  NANDN U5922 ( .A(n5065), .B(n5064), .Z(n5069) );
  NAND U5923 ( .A(n5067), .B(n5066), .Z(n5068) );
  AND U5924 ( .A(n5069), .B(n5068), .Z(n5080) );
  XOR U5925 ( .A(n5073), .B(n5072), .Z(n5210) );
  XOR U5926 ( .A(n5211), .B(n5210), .Z(o[45]) );
  NANDN U5927 ( .A(n5075), .B(n5074), .Z(n5079) );
  NAND U5928 ( .A(n5077), .B(n5076), .Z(n5078) );
  AND U5929 ( .A(n5079), .B(n5078), .Z(n5480) );
  NANDN U5930 ( .A(n5081), .B(n5080), .Z(n5085) );
  NANDN U5931 ( .A(n5083), .B(n5082), .Z(n5084) );
  NAND U5932 ( .A(n5085), .B(n5084), .Z(n5481) );
  NANDN U5933 ( .A(n5087), .B(n5086), .Z(n5091) );
  NAND U5934 ( .A(n5089), .B(n5088), .Z(n5090) );
  AND U5935 ( .A(n5091), .B(n5090), .Z(n5487) );
  NANDN U5936 ( .A(n5093), .B(n5092), .Z(n5097) );
  NANDN U5937 ( .A(n5095), .B(n5094), .Z(n5096) );
  NAND U5938 ( .A(n5097), .B(n5096), .Z(n5236) );
  AND U5939 ( .A(x[51]), .B(y[43]), .Z(n5191) );
  NAND U5940 ( .A(n5098), .B(n5191), .Z(n5102) );
  NANDN U5941 ( .A(n5100), .B(n5099), .Z(n5101) );
  AND U5942 ( .A(n5102), .B(n5101), .Z(n5372) );
  AND U5943 ( .A(y[123]), .B(x[67]), .Z(n5399) );
  AND U5944 ( .A(y[83]), .B(x[59]), .Z(n5398) );
  XOR U5945 ( .A(n5399), .B(n5398), .Z(n5397) );
  AND U5946 ( .A(y[3]), .B(x[43]), .Z(n5396) );
  XOR U5947 ( .A(n5397), .B(n5396), .Z(n5375) );
  AND U5948 ( .A(y[124]), .B(x[66]), .Z(n5341) );
  AND U5949 ( .A(y[82]), .B(x[60]), .Z(n5340) );
  XOR U5950 ( .A(n5341), .B(n5340), .Z(n5339) );
  AND U5951 ( .A(y[4]), .B(x[42]), .Z(n5338) );
  XNOR U5952 ( .A(n5339), .B(n5338), .Z(n5374) );
  XNOR U5953 ( .A(n5372), .B(n5373), .Z(n5239) );
  NANDN U5954 ( .A(n5104), .B(n5103), .Z(n5108) );
  NAND U5955 ( .A(n5106), .B(n5105), .Z(n5107) );
  NAND U5956 ( .A(n5108), .B(n5107), .Z(n5238) );
  XOR U5957 ( .A(n5236), .B(n5237), .Z(n5221) );
  XOR U5958 ( .A(n5221), .B(n5220), .Z(n5218) );
  AND U5959 ( .A(y[81]), .B(x[61]), .Z(n5381) );
  NANDN U5960 ( .A(n5113), .B(n5381), .Z(n5117) );
  NANDN U5961 ( .A(n5115), .B(n5114), .Z(n5116) );
  AND U5962 ( .A(n5117), .B(n5116), .Z(n5367) );
  AND U5963 ( .A(x[45]), .B(y[1]), .Z(n5119) );
  NAND U5964 ( .A(x[44]), .B(y[2]), .Z(n5118) );
  XNOR U5965 ( .A(n5119), .B(n5118), .Z(n5424) );
  AND U5966 ( .A(y[120]), .B(x[70]), .Z(n5423) );
  XNOR U5967 ( .A(n5424), .B(n5423), .Z(n5365) );
  AND U5968 ( .A(y[165]), .B(x[73]), .Z(n5327) );
  AND U5969 ( .A(x[76]), .B(y[162]), .Z(n5183) );
  AND U5970 ( .A(n5183), .B(n5120), .Z(n5325) );
  AND U5971 ( .A(y[164]), .B(x[74]), .Z(n5324) );
  XOR U5972 ( .A(n5325), .B(n5324), .Z(n5326) );
  XOR U5973 ( .A(n5327), .B(n5326), .Z(n5364) );
  XOR U5974 ( .A(n5367), .B(n5366), .Z(n5352) );
  NAND U5975 ( .A(n5122), .B(n5121), .Z(n5125) );
  NAND U5976 ( .A(n5123), .B(n5426), .Z(n5124) );
  NAND U5977 ( .A(n5125), .B(n5124), .Z(n5355) );
  NAND U5978 ( .A(n5127), .B(n5126), .Z(n5130) );
  NAND U5979 ( .A(n5420), .B(n5128), .Z(n5129) );
  NAND U5980 ( .A(n5130), .B(n5129), .Z(n5354) );
  XNOR U5981 ( .A(n5355), .B(n5354), .Z(n5353) );
  XNOR U5982 ( .A(n5218), .B(n5219), .Z(n5217) );
  NANDN U5983 ( .A(n5132), .B(n5131), .Z(n5137) );
  IV U5984 ( .A(n5133), .Z(n5135) );
  NANDN U5985 ( .A(n5135), .B(n5134), .Z(n5136) );
  AND U5986 ( .A(n5137), .B(n5136), .Z(n5216) );
  NANDN U5987 ( .A(n5143), .B(n5142), .Z(n5147) );
  NAND U5988 ( .A(n5145), .B(n5144), .Z(n5146) );
  AND U5989 ( .A(n5147), .B(n5146), .Z(n5224) );
  XOR U5990 ( .A(n5225), .B(n5224), .Z(n5223) );
  NAND U5991 ( .A(n5149), .B(n5148), .Z(n5153) );
  NAND U5992 ( .A(n5151), .B(n5150), .Z(n5152) );
  AND U5993 ( .A(n5153), .B(n5152), .Z(n5222) );
  XOR U5994 ( .A(n5223), .B(n5222), .Z(n5214) );
  XOR U5995 ( .A(n5215), .B(n5214), .Z(n5486) );
  XOR U5996 ( .A(n5487), .B(n5486), .Z(n5484) );
  NANDN U5997 ( .A(n5155), .B(n5154), .Z(n5159) );
  NANDN U5998 ( .A(n5157), .B(n5156), .Z(n5158) );
  AND U5999 ( .A(n5159), .B(n5158), .Z(n5458) );
  NANDN U6000 ( .A(n5161), .B(n5160), .Z(n5165) );
  OR U6001 ( .A(n5163), .B(n5162), .Z(n5164) );
  NAND U6002 ( .A(n5165), .B(n5164), .Z(n5461) );
  NAND U6003 ( .A(n5166), .B(n5335), .Z(n5170) );
  NAND U6004 ( .A(n5168), .B(n5167), .Z(n5169) );
  NAND U6005 ( .A(n5170), .B(n5169), .Z(n5232) );
  NANDN U6006 ( .A(n5171), .B(n5327), .Z(n5175) );
  NAND U6007 ( .A(n5173), .B(n5172), .Z(n5174) );
  NAND U6008 ( .A(n5175), .B(n5174), .Z(n5235) );
  NAND U6009 ( .A(n5177), .B(n5176), .Z(n5181) );
  NAND U6010 ( .A(n5179), .B(n5178), .Z(n5180) );
  AND U6011 ( .A(n5181), .B(n5180), .Z(n5359) );
  AND U6012 ( .A(y[5]), .B(x[41]), .Z(n5440) );
  AND U6013 ( .A(y[40]), .B(x[54]), .Z(n5439) );
  XOR U6014 ( .A(n5440), .B(n5439), .Z(n5438) );
  AND U6015 ( .A(y[46]), .B(x[48]), .Z(n5437) );
  XOR U6016 ( .A(n5438), .B(n5437), .Z(n5360) );
  NAND U6017 ( .A(x[77]), .B(y[161]), .Z(n5182) );
  XNOR U6018 ( .A(n5183), .B(n5182), .Z(n5321) );
  AND U6019 ( .A(y[160]), .B(x[78]), .Z(n5320) );
  XOR U6020 ( .A(n5321), .B(n5320), .Z(n5318) );
  XNOR U6021 ( .A(n5319), .B(n5318), .Z(n5361) );
  XNOR U6022 ( .A(n5359), .B(n5358), .Z(n5234) );
  XOR U6023 ( .A(n5235), .B(n5234), .Z(n5233) );
  XOR U6024 ( .A(n5232), .B(n5233), .Z(n5466) );
  NAND U6025 ( .A(n5185), .B(n5184), .Z(n5189) );
  NAND U6026 ( .A(n5187), .B(n5186), .Z(n5188) );
  AND U6027 ( .A(n5189), .B(n5188), .Z(n5465) );
  AND U6028 ( .A(y[86]), .B(x[56]), .Z(n5434) );
  AND U6029 ( .A(y[0]), .B(x[46]), .Z(n5433) );
  XOR U6030 ( .A(n5434), .B(n5433), .Z(n5432) );
  AND U6031 ( .A(y[121]), .B(x[69]), .Z(n5431) );
  XOR U6032 ( .A(n5432), .B(n5431), .Z(n5315) );
  AND U6033 ( .A(y[41]), .B(x[53]), .Z(n5387) );
  AND U6034 ( .A(y[44]), .B(x[50]), .Z(n5386) );
  XOR U6035 ( .A(n5387), .B(n5386), .Z(n5385) );
  AND U6036 ( .A(y[45]), .B(x[49]), .Z(n5384) );
  XOR U6037 ( .A(n5385), .B(n5384), .Z(n5247) );
  NAND U6038 ( .A(x[52]), .B(y[42]), .Z(n5190) );
  XNOR U6039 ( .A(n5191), .B(n5190), .Z(n5246) );
  XOR U6040 ( .A(n5247), .B(n5246), .Z(n5314) );
  XOR U6041 ( .A(n5315), .B(n5314), .Z(n5313) );
  AND U6042 ( .A(y[166]), .B(x[72]), .Z(n5380) );
  XOR U6043 ( .A(n5381), .B(n5380), .Z(n5379) );
  AND U6044 ( .A(y[80]), .B(x[62]), .Z(n5378) );
  XOR U6045 ( .A(n5379), .B(n5378), .Z(n5312) );
  XOR U6046 ( .A(n5313), .B(n5312), .Z(n5231) );
  NAND U6047 ( .A(n5193), .B(n5192), .Z(n5197) );
  NAND U6048 ( .A(n5195), .B(n5194), .Z(n5196) );
  AND U6049 ( .A(n5197), .B(n5196), .Z(n5240) );
  AND U6050 ( .A(x[57]), .B(y[85]), .Z(n5199) );
  NAND U6051 ( .A(x[58]), .B(y[84]), .Z(n5198) );
  XNOR U6052 ( .A(n5199), .B(n5198), .Z(n5333) );
  AND U6053 ( .A(y[122]), .B(x[68]), .Z(n5332) );
  XOR U6054 ( .A(n5333), .B(n5332), .Z(n5243) );
  AND U6055 ( .A(x[64]), .B(y[126]), .Z(n5201) );
  NAND U6056 ( .A(x[65]), .B(y[125]), .Z(n5200) );
  XNOR U6057 ( .A(n5201), .B(n5200), .Z(n5418) );
  AND U6058 ( .A(y[6]), .B(x[40]), .Z(n5417) );
  XNOR U6059 ( .A(n5418), .B(n5417), .Z(n5242) );
  XNOR U6060 ( .A(n5240), .B(n5241), .Z(n5230) );
  NAND U6061 ( .A(n5203), .B(n5202), .Z(n5207) );
  NAND U6062 ( .A(n5205), .B(n5204), .Z(n5206) );
  AND U6063 ( .A(n5207), .B(n5206), .Z(n5228) );
  XOR U6064 ( .A(n5229), .B(n5228), .Z(n5464) );
  XOR U6065 ( .A(n5465), .B(n5464), .Z(n5467) );
  XOR U6066 ( .A(n5461), .B(n5460), .Z(n5459) );
  XOR U6067 ( .A(n5458), .B(n5459), .Z(n5485) );
  XNOR U6068 ( .A(n5479), .B(n5478), .Z(n5474) );
  NANDN U6069 ( .A(n5209), .B(n5208), .Z(n5213) );
  NAND U6070 ( .A(n5211), .B(n5210), .Z(n5212) );
  NAND U6071 ( .A(n5213), .B(n5212), .Z(n5472) );
  XOR U6072 ( .A(n5473), .B(n5472), .Z(o[46]) );
  NAND U6073 ( .A(n5223), .B(n5222), .Z(n5227) );
  NAND U6074 ( .A(n5225), .B(n5224), .Z(n5226) );
  AND U6075 ( .A(n5227), .B(n5226), .Z(n5457) );
  NANDN U6076 ( .A(n5241), .B(n5240), .Z(n5245) );
  NANDN U6077 ( .A(n5243), .B(n5242), .Z(n5244) );
  NAND U6078 ( .A(n5247), .B(n5246), .Z(n5250) );
  AND U6079 ( .A(y[42]), .B(x[51]), .Z(n5248) );
  AND U6080 ( .A(y[43]), .B(x[52]), .Z(n5300) );
  NAND U6081 ( .A(n5248), .B(n5300), .Z(n5249) );
  AND U6082 ( .A(n5250), .B(n5249), .Z(n5311) );
  AND U6083 ( .A(x[68]), .B(y[123]), .Z(n5252) );
  NAND U6084 ( .A(x[46]), .B(y[1]), .Z(n5251) );
  XNOR U6085 ( .A(n5252), .B(n5251), .Z(n5256) );
  AND U6086 ( .A(x[47]), .B(y[0]), .Z(n5254) );
  NAND U6087 ( .A(x[59]), .B(y[84]), .Z(n5253) );
  XNOR U6088 ( .A(n5254), .B(n5253), .Z(n5255) );
  XOR U6089 ( .A(n5256), .B(n5255), .Z(n5264) );
  AND U6090 ( .A(x[42]), .B(y[5]), .Z(n5258) );
  NAND U6091 ( .A(x[79]), .B(y[160]), .Z(n5257) );
  XNOR U6092 ( .A(n5258), .B(n5257), .Z(n5262) );
  AND U6093 ( .A(x[70]), .B(y[121]), .Z(n5260) );
  NAND U6094 ( .A(x[62]), .B(y[81]), .Z(n5259) );
  XNOR U6095 ( .A(n5260), .B(n5259), .Z(n5261) );
  XNOR U6096 ( .A(n5262), .B(n5261), .Z(n5263) );
  XNOR U6097 ( .A(n5264), .B(n5263), .Z(n5309) );
  AND U6098 ( .A(x[71]), .B(y[120]), .Z(n5269) );
  AND U6099 ( .A(y[162]), .B(x[77]), .Z(n5394) );
  AND U6100 ( .A(x[48]), .B(y[47]), .Z(n5266) );
  NAND U6101 ( .A(x[56]), .B(y[87]), .Z(n5265) );
  XNOR U6102 ( .A(n5266), .B(n5265), .Z(n5267) );
  XNOR U6103 ( .A(n5394), .B(n5267), .Z(n5268) );
  XNOR U6104 ( .A(n5269), .B(n5268), .Z(n5285) );
  AND U6105 ( .A(x[64]), .B(y[127]), .Z(n5271) );
  NAND U6106 ( .A(x[49]), .B(y[46]), .Z(n5270) );
  XNOR U6107 ( .A(n5271), .B(n5270), .Z(n5275) );
  AND U6108 ( .A(x[66]), .B(y[125]), .Z(n5273) );
  NAND U6109 ( .A(x[55]), .B(y[40]), .Z(n5272) );
  XNOR U6110 ( .A(n5273), .B(n5272), .Z(n5274) );
  XOR U6111 ( .A(n5275), .B(n5274), .Z(n5283) );
  AND U6112 ( .A(x[50]), .B(y[45]), .Z(n5277) );
  NAND U6113 ( .A(x[53]), .B(y[42]), .Z(n5276) );
  XNOR U6114 ( .A(n5277), .B(n5276), .Z(n5281) );
  AND U6115 ( .A(x[67]), .B(y[124]), .Z(n5279) );
  NAND U6116 ( .A(x[78]), .B(y[161]), .Z(n5278) );
  XNOR U6117 ( .A(n5279), .B(n5278), .Z(n5280) );
  XNOR U6118 ( .A(n5281), .B(n5280), .Z(n5282) );
  XNOR U6119 ( .A(n5283), .B(n5282), .Z(n5284) );
  XOR U6120 ( .A(n5285), .B(n5284), .Z(n5307) );
  AND U6121 ( .A(x[40]), .B(y[7]), .Z(n5287) );
  NAND U6122 ( .A(x[75]), .B(y[164]), .Z(n5286) );
  XNOR U6123 ( .A(n5287), .B(n5286), .Z(n5291) );
  AND U6124 ( .A(x[41]), .B(y[6]), .Z(n5289) );
  NAND U6125 ( .A(x[73]), .B(y[166]), .Z(n5288) );
  XNOR U6126 ( .A(n5289), .B(n5288), .Z(n5290) );
  XOR U6127 ( .A(n5291), .B(n5290), .Z(n5299) );
  AND U6128 ( .A(x[57]), .B(y[86]), .Z(n5293) );
  NAND U6129 ( .A(x[60]), .B(y[83]), .Z(n5292) );
  XNOR U6130 ( .A(n5293), .B(n5292), .Z(n5297) );
  AND U6131 ( .A(x[74]), .B(y[165]), .Z(n5295) );
  NAND U6132 ( .A(x[44]), .B(y[3]), .Z(n5294) );
  XNOR U6133 ( .A(n5295), .B(n5294), .Z(n5296) );
  XNOR U6134 ( .A(n5297), .B(n5296), .Z(n5298) );
  XNOR U6135 ( .A(n5299), .B(n5298), .Z(n5305) );
  AND U6136 ( .A(y[85]), .B(x[58]), .Z(n5334) );
  AND U6137 ( .A(y[126]), .B(x[65]), .Z(n5419) );
  XOR U6138 ( .A(n5334), .B(n5419), .Z(n5303) );
  XNOR U6139 ( .A(n5301), .B(n5300), .Z(n5302) );
  XNOR U6140 ( .A(n5303), .B(n5302), .Z(n5304) );
  XNOR U6141 ( .A(n5305), .B(n5304), .Z(n5306) );
  XNOR U6142 ( .A(n5307), .B(n5306), .Z(n5308) );
  XNOR U6143 ( .A(n5309), .B(n5308), .Z(n5310) );
  XNOR U6144 ( .A(n5311), .B(n5310), .Z(n5351) );
  NAND U6145 ( .A(n5313), .B(n5312), .Z(n5317) );
  NAND U6146 ( .A(n5315), .B(n5314), .Z(n5316) );
  AND U6147 ( .A(n5317), .B(n5316), .Z(n5349) );
  NAND U6148 ( .A(n5319), .B(n5318), .Z(n5323) );
  AND U6149 ( .A(n5321), .B(n5320), .Z(n5322) );
  ANDN U6150 ( .B(n5323), .A(n5322), .Z(n5331) );
  AND U6151 ( .A(n5325), .B(n5324), .Z(n5329) );
  AND U6152 ( .A(n5327), .B(n5326), .Z(n5328) );
  OR U6153 ( .A(n5329), .B(n5328), .Z(n5330) );
  XNOR U6154 ( .A(n5331), .B(n5330), .Z(n5347) );
  NAND U6155 ( .A(n5333), .B(n5332), .Z(n5337) );
  NAND U6156 ( .A(n5335), .B(n5334), .Z(n5336) );
  AND U6157 ( .A(n5337), .B(n5336), .Z(n5345) );
  NAND U6158 ( .A(n5339), .B(n5338), .Z(n5343) );
  NAND U6159 ( .A(n5341), .B(n5340), .Z(n5342) );
  NAND U6160 ( .A(n5343), .B(n5342), .Z(n5344) );
  XNOR U6161 ( .A(n5345), .B(n5344), .Z(n5346) );
  XNOR U6162 ( .A(n5347), .B(n5346), .Z(n5348) );
  XNOR U6163 ( .A(n5349), .B(n5348), .Z(n5350) );
  NANDN U6164 ( .A(n5353), .B(n5352), .Z(n5357) );
  NAND U6165 ( .A(n5355), .B(n5354), .Z(n5356) );
  NAND U6166 ( .A(n5359), .B(n5358), .Z(n5363) );
  ANDN U6167 ( .B(n5361), .A(n5360), .Z(n5362) );
  ANDN U6168 ( .B(n5363), .A(n5362), .Z(n5371) );
  ANDN U6169 ( .B(n5365), .A(n5364), .Z(n5369) );
  ANDN U6170 ( .B(n5367), .A(n5366), .Z(n5368) );
  OR U6171 ( .A(n5369), .B(n5368), .Z(n5370) );
  XNOR U6172 ( .A(n5371), .B(n5370), .Z(n5454) );
  NANDN U6173 ( .A(n5373), .B(n5372), .Z(n5377) );
  NANDN U6174 ( .A(n5375), .B(n5374), .Z(n5376) );
  AND U6175 ( .A(n5377), .B(n5376), .Z(n5452) );
  NAND U6176 ( .A(n5379), .B(n5378), .Z(n5383) );
  NAND U6177 ( .A(n5381), .B(n5380), .Z(n5382) );
  AND U6178 ( .A(n5383), .B(n5382), .Z(n5391) );
  NAND U6179 ( .A(n5385), .B(n5384), .Z(n5389) );
  NAND U6180 ( .A(n5387), .B(n5386), .Z(n5388) );
  NAND U6181 ( .A(n5389), .B(n5388), .Z(n5390) );
  XNOR U6182 ( .A(n5391), .B(n5390), .Z(n5450) );
  AND U6183 ( .A(x[43]), .B(y[4]), .Z(n5393) );
  NAND U6184 ( .A(x[54]), .B(y[41]), .Z(n5392) );
  XNOR U6185 ( .A(n5393), .B(n5392), .Z(n5416) );
  AND U6186 ( .A(y[161]), .B(x[76]), .Z(n5395) );
  AND U6187 ( .A(n5395), .B(n5394), .Z(n5411) );
  NAND U6188 ( .A(n5397), .B(n5396), .Z(n5401) );
  NAND U6189 ( .A(n5399), .B(n5398), .Z(n5400) );
  AND U6190 ( .A(n5401), .B(n5400), .Z(n5409) );
  AND U6191 ( .A(x[72]), .B(y[167]), .Z(n5403) );
  NAND U6192 ( .A(x[63]), .B(y[80]), .Z(n5402) );
  XNOR U6193 ( .A(n5403), .B(n5402), .Z(n5407) );
  AND U6194 ( .A(x[61]), .B(y[82]), .Z(n5405) );
  NAND U6195 ( .A(x[69]), .B(y[122]), .Z(n5404) );
  XNOR U6196 ( .A(n5405), .B(n5404), .Z(n5406) );
  XNOR U6197 ( .A(n5407), .B(n5406), .Z(n5408) );
  XNOR U6198 ( .A(n5409), .B(n5408), .Z(n5410) );
  XOR U6199 ( .A(n5411), .B(n5410), .Z(n5414) );
  AND U6200 ( .A(y[2]), .B(x[45]), .Z(n5425) );
  XNOR U6201 ( .A(n5425), .B(n5412), .Z(n5413) );
  XNOR U6202 ( .A(n5414), .B(n5413), .Z(n5415) );
  XOR U6203 ( .A(n5416), .B(n5415), .Z(n5448) );
  NAND U6204 ( .A(n5418), .B(n5417), .Z(n5422) );
  NAND U6205 ( .A(n5420), .B(n5419), .Z(n5421) );
  AND U6206 ( .A(n5422), .B(n5421), .Z(n5430) );
  NAND U6207 ( .A(n5424), .B(n5423), .Z(n5428) );
  NAND U6208 ( .A(n5426), .B(n5425), .Z(n5427) );
  NAND U6209 ( .A(n5428), .B(n5427), .Z(n5429) );
  XNOR U6210 ( .A(n5430), .B(n5429), .Z(n5446) );
  NAND U6211 ( .A(n5432), .B(n5431), .Z(n5436) );
  NAND U6212 ( .A(n5434), .B(n5433), .Z(n5435) );
  AND U6213 ( .A(n5436), .B(n5435), .Z(n5444) );
  NAND U6214 ( .A(n5438), .B(n5437), .Z(n5442) );
  NAND U6215 ( .A(n5440), .B(n5439), .Z(n5441) );
  NAND U6216 ( .A(n5442), .B(n5441), .Z(n5443) );
  XNOR U6217 ( .A(n5444), .B(n5443), .Z(n5445) );
  XNOR U6218 ( .A(n5446), .B(n5445), .Z(n5447) );
  XNOR U6219 ( .A(n5448), .B(n5447), .Z(n5449) );
  XNOR U6220 ( .A(n5450), .B(n5449), .Z(n5451) );
  XNOR U6221 ( .A(n5452), .B(n5451), .Z(n5453) );
  XNOR U6222 ( .A(n5454), .B(n5453), .Z(n5455) );
  NANDN U6223 ( .A(n5459), .B(n5458), .Z(n5463) );
  ANDN U6224 ( .B(n5461), .A(n5460), .Z(n5462) );
  ANDN U6225 ( .B(n5463), .A(n5462), .Z(n5471) );
  AND U6226 ( .A(n5465), .B(n5464), .Z(n5469) );
  ANDN U6227 ( .B(n5467), .A(n5466), .Z(n5468) );
  OR U6228 ( .A(n5469), .B(n5468), .Z(n5470) );
  NAND U6229 ( .A(n5473), .B(n5472), .Z(n5477) );
  NANDN U6230 ( .A(n5475), .B(n5474), .Z(n5476) );
  NAND U6231 ( .A(n5479), .B(n5478), .Z(n5483) );
  NANDN U6232 ( .A(n5481), .B(n5480), .Z(n5482) );
  NAND U6233 ( .A(y[168]), .B(x[72]), .Z(n5626) );
  NAND U6234 ( .A(y[48]), .B(x[48]), .Z(n5490) );
  XOR U6235 ( .A(n5626), .B(n5490), .Z(n5491) );
  AND U6236 ( .A(y[8]), .B(x[40]), .Z(n5498) );
  AND U6237 ( .A(y[88]), .B(x[56]), .Z(n5495) );
  XOR U6238 ( .A(n5498), .B(n5495), .Z(n5494) );
  AND U6239 ( .A(y[128]), .B(x[64]), .Z(n5493) );
  XNOR U6240 ( .A(n5494), .B(n5493), .Z(n5492) );
  XNOR U6241 ( .A(n5491), .B(n5492), .Z(o[48]) );
  AND U6242 ( .A(x[40]), .B(y[9]), .Z(n5489) );
  NAND U6243 ( .A(x[41]), .B(y[8]), .Z(n5488) );
  XNOR U6244 ( .A(n5489), .B(n5488), .Z(n5500) );
  AND U6245 ( .A(y[48]), .B(x[49]), .Z(n5499) );
  XOR U6246 ( .A(n5500), .B(n5499), .Z(n5517) );
  AND U6247 ( .A(y[168]), .B(x[73]), .Z(n5729) );
  AND U6248 ( .A(y[89]), .B(x[56]), .Z(n5503) );
  XOR U6249 ( .A(n5729), .B(n5503), .Z(n5505) );
  AND U6250 ( .A(y[169]), .B(x[72]), .Z(n5527) );
  NAND U6251 ( .A(y[88]), .B(x[57]), .Z(n5526) );
  XNOR U6252 ( .A(n5527), .B(n5526), .Z(n5504) );
  XOR U6253 ( .A(n5505), .B(n5504), .Z(n5515) );
  AND U6254 ( .A(y[49]), .B(x[48]), .Z(n5753) );
  AND U6255 ( .A(y[129]), .B(x[64]), .Z(n5520) );
  XOR U6256 ( .A(n5753), .B(n5520), .Z(n5522) );
  AND U6257 ( .A(y[128]), .B(x[65]), .Z(n5521) );
  XNOR U6258 ( .A(n5522), .B(n5521), .Z(n5514) );
  XNOR U6259 ( .A(n5515), .B(n5514), .Z(n5516) );
  XNOR U6260 ( .A(n5517), .B(n5516), .Z(n5511) );
  NAND U6261 ( .A(n5494), .B(n5493), .Z(n5497) );
  AND U6262 ( .A(n5498), .B(n5495), .Z(n5496) );
  ANDN U6263 ( .B(n5497), .A(n5496), .Z(n5508) );
  XNOR U6264 ( .A(n5509), .B(n5508), .Z(n5510) );
  XNOR U6265 ( .A(n5511), .B(n5510), .Z(o[49]) );
  NAND U6266 ( .A(y[9]), .B(x[41]), .Z(n5549) );
  NANDN U6267 ( .A(n5549), .B(n5498), .Z(n5502) );
  NAND U6268 ( .A(n5500), .B(n5499), .Z(n5501) );
  AND U6269 ( .A(n5502), .B(n5501), .Z(n5583) );
  NAND U6270 ( .A(n5729), .B(n5503), .Z(n5507) );
  NAND U6271 ( .A(n5505), .B(n5504), .Z(n5506) );
  AND U6272 ( .A(n5507), .B(n5506), .Z(n5582) );
  AND U6273 ( .A(y[130]), .B(x[64]), .Z(n5567) );
  NAND U6274 ( .A(y[10]), .B(x[40]), .Z(n5568) );
  XNOR U6275 ( .A(n5567), .B(n5568), .Z(n5569) );
  NAND U6276 ( .A(y[48]), .B(x[50]), .Z(n5570) );
  XNOR U6277 ( .A(n5569), .B(n5570), .Z(n5581) );
  XOR U6278 ( .A(n5582), .B(n5581), .Z(n5584) );
  XOR U6279 ( .A(n5583), .B(n5584), .Z(n5529) );
  NANDN U6280 ( .A(n5509), .B(n5508), .Z(n5513) );
  NAND U6281 ( .A(n5511), .B(n5510), .Z(n5512) );
  NAND U6282 ( .A(n5513), .B(n5512), .Z(n5528) );
  XNOR U6283 ( .A(n5529), .B(n5528), .Z(n5531) );
  NANDN U6284 ( .A(n5515), .B(n5514), .Z(n5519) );
  NANDN U6285 ( .A(n5517), .B(n5516), .Z(n5518) );
  AND U6286 ( .A(n5519), .B(n5518), .Z(n5537) );
  AND U6287 ( .A(y[8]), .B(x[42]), .Z(n5546) );
  NAND U6288 ( .A(y[90]), .B(x[56]), .Z(n5547) );
  XNOR U6289 ( .A(n5546), .B(n5547), .Z(n5548) );
  AND U6290 ( .A(y[128]), .B(x[66]), .Z(n5575) );
  XOR U6291 ( .A(n5576), .B(n5575), .Z(n5578) );
  AND U6292 ( .A(y[88]), .B(x[58]), .Z(n5656) );
  AND U6293 ( .A(y[170]), .B(x[72]), .Z(n5559) );
  XOR U6294 ( .A(n5656), .B(n5559), .Z(n5561) );
  AND U6295 ( .A(y[89]), .B(x[57]), .Z(n5560) );
  XOR U6296 ( .A(n5561), .B(n5560), .Z(n5577) );
  XOR U6297 ( .A(n5578), .B(n5577), .Z(n5534) );
  NAND U6298 ( .A(n5753), .B(n5520), .Z(n5524) );
  AND U6299 ( .A(n5522), .B(n5521), .Z(n5523) );
  ANDN U6300 ( .B(n5524), .A(n5523), .Z(n5543) );
  AND U6301 ( .A(x[73]), .B(y[169]), .Z(n5631) );
  NAND U6302 ( .A(x[74]), .B(y[168]), .Z(n5525) );
  XNOR U6303 ( .A(n5631), .B(n5525), .Z(n5574) );
  ANDN U6304 ( .B(n5527), .A(n5526), .Z(n5573) );
  XOR U6305 ( .A(n5574), .B(n5573), .Z(n5540) );
  AND U6306 ( .A(y[129]), .B(x[65]), .Z(n5552) );
  NAND U6307 ( .A(y[49]), .B(x[49]), .Z(n5553) );
  XNOR U6308 ( .A(n5552), .B(n5553), .Z(n5554) );
  NAND U6309 ( .A(y[50]), .B(x[48]), .Z(n5555) );
  XOR U6310 ( .A(n5554), .B(n5555), .Z(n5541) );
  XNOR U6311 ( .A(n5540), .B(n5541), .Z(n5542) );
  XOR U6312 ( .A(n5543), .B(n5542), .Z(n5535) );
  XNOR U6313 ( .A(n5534), .B(n5535), .Z(n5536) );
  XNOR U6314 ( .A(n5537), .B(n5536), .Z(n5530) );
  XNOR U6315 ( .A(n5531), .B(n5530), .Z(o[50]) );
  NANDN U6316 ( .A(n5529), .B(n5528), .Z(n5533) );
  NAND U6317 ( .A(n5531), .B(n5530), .Z(n5532) );
  AND U6318 ( .A(n5533), .B(n5532), .Z(n5605) );
  NANDN U6319 ( .A(n5535), .B(n5534), .Z(n5539) );
  NAND U6320 ( .A(n5537), .B(n5536), .Z(n5538) );
  AND U6321 ( .A(n5539), .B(n5538), .Z(n5590) );
  NANDN U6322 ( .A(n5541), .B(n5540), .Z(n5545) );
  NANDN U6323 ( .A(n5543), .B(n5542), .Z(n5544) );
  AND U6324 ( .A(n5545), .B(n5544), .Z(n5588) );
  NANDN U6325 ( .A(n5547), .B(n5546), .Z(n5551) );
  NANDN U6326 ( .A(n5549), .B(n5548), .Z(n5550) );
  NAND U6327 ( .A(n5551), .B(n5550), .Z(n5599) );
  NANDN U6328 ( .A(n5553), .B(n5552), .Z(n5557) );
  NANDN U6329 ( .A(n5555), .B(n5554), .Z(n5556) );
  AND U6330 ( .A(n5557), .B(n5556), .Z(n5647) );
  AND U6331 ( .A(y[131]), .B(x[64]), .Z(n5674) );
  AND U6332 ( .A(y[91]), .B(x[56]), .Z(n5673) );
  NAND U6333 ( .A(y[8]), .B(x[43]), .Z(n5672) );
  XOR U6334 ( .A(n5673), .B(n5672), .Z(n5675) );
  XOR U6335 ( .A(n5674), .B(n5675), .Z(n5645) );
  AND U6336 ( .A(y[89]), .B(x[58]), .Z(n5696) );
  NAND U6337 ( .A(x[59]), .B(y[88]), .Z(n5558) );
  XNOR U6338 ( .A(n5696), .B(n5558), .Z(n5657) );
  NAND U6339 ( .A(y[90]), .B(x[57]), .Z(n5658) );
  XNOR U6340 ( .A(n5657), .B(n5658), .Z(n5644) );
  XNOR U6341 ( .A(n5645), .B(n5644), .Z(n5646) );
  XNOR U6342 ( .A(n5647), .B(n5646), .Z(n5600) );
  XOR U6343 ( .A(n5599), .B(n5600), .Z(n5602) );
  NAND U6344 ( .A(n5656), .B(n5559), .Z(n5563) );
  AND U6345 ( .A(n5561), .B(n5560), .Z(n5562) );
  ANDN U6346 ( .B(n5563), .A(n5562), .Z(n5652) );
  AND U6347 ( .A(y[10]), .B(x[41]), .Z(n5622) );
  AND U6348 ( .A(y[9]), .B(x[42]), .Z(n5621) );
  NAND U6349 ( .A(y[130]), .B(x[65]), .Z(n5620) );
  XOR U6350 ( .A(n5621), .B(n5620), .Z(n5623) );
  XOR U6351 ( .A(n5622), .B(n5623), .Z(n5651) );
  AND U6352 ( .A(x[75]), .B(y[168]), .Z(n5565) );
  NAND U6353 ( .A(x[72]), .B(y[171]), .Z(n5564) );
  XNOR U6354 ( .A(n5565), .B(n5564), .Z(n5627) );
  AND U6355 ( .A(y[169]), .B(x[74]), .Z(n5713) );
  NAND U6356 ( .A(x[73]), .B(y[170]), .Z(n5566) );
  XOR U6357 ( .A(n5713), .B(n5566), .Z(n5628) );
  XNOR U6358 ( .A(n5627), .B(n5628), .Z(n5650) );
  XOR U6359 ( .A(n5651), .B(n5650), .Z(n5653) );
  XOR U6360 ( .A(n5652), .B(n5653), .Z(n5601) );
  XOR U6361 ( .A(n5602), .B(n5601), .Z(n5587) );
  XNOR U6362 ( .A(n5588), .B(n5587), .Z(n5589) );
  XOR U6363 ( .A(n5590), .B(n5589), .Z(n5606) );
  XNOR U6364 ( .A(n5605), .B(n5606), .Z(n5608) );
  NANDN U6365 ( .A(n5568), .B(n5567), .Z(n5572) );
  NANDN U6366 ( .A(n5570), .B(n5569), .Z(n5571) );
  AND U6367 ( .A(n5572), .B(n5571), .Z(n5612) );
  XNOR U6368 ( .A(n5612), .B(n5611), .Z(n5614) );
  NAND U6369 ( .A(y[48]), .B(x[51]), .Z(n5666) );
  NAND U6370 ( .A(y[11]), .B(x[40]), .Z(n5664) );
  NAND U6371 ( .A(y[129]), .B(x[66]), .Z(n5663) );
  XOR U6372 ( .A(n5664), .B(n5663), .Z(n5665) );
  XNOR U6373 ( .A(n5666), .B(n5665), .Z(n5641) );
  NAND U6374 ( .A(y[51]), .B(x[48]), .Z(n5635) );
  NAND U6375 ( .A(y[49]), .B(x[50]), .Z(n5633) );
  NAND U6376 ( .A(y[128]), .B(x[67]), .Z(n5632) );
  XOR U6377 ( .A(n5633), .B(n5632), .Z(n5634) );
  XNOR U6378 ( .A(n5635), .B(n5634), .Z(n5639) );
  AND U6379 ( .A(y[50]), .B(x[49]), .Z(n5638) );
  XOR U6380 ( .A(n5639), .B(n5638), .Z(n5640) );
  XOR U6381 ( .A(n5641), .B(n5640), .Z(n5613) );
  XOR U6382 ( .A(n5614), .B(n5613), .Z(n5594) );
  NAND U6383 ( .A(n5576), .B(n5575), .Z(n5580) );
  NAND U6384 ( .A(n5578), .B(n5577), .Z(n5579) );
  AND U6385 ( .A(n5580), .B(n5579), .Z(n5593) );
  XNOR U6386 ( .A(n5594), .B(n5593), .Z(n5596) );
  NANDN U6387 ( .A(n5582), .B(n5581), .Z(n5586) );
  OR U6388 ( .A(n5584), .B(n5583), .Z(n5585) );
  AND U6389 ( .A(n5586), .B(n5585), .Z(n5595) );
  XNOR U6390 ( .A(n5596), .B(n5595), .Z(n5607) );
  XOR U6391 ( .A(n5608), .B(n5607), .Z(o[51]) );
  NANDN U6392 ( .A(n5588), .B(n5587), .Z(n5592) );
  NANDN U6393 ( .A(n5590), .B(n5589), .Z(n5591) );
  AND U6394 ( .A(n5592), .B(n5591), .Z(n5686) );
  NANDN U6395 ( .A(n5594), .B(n5593), .Z(n5598) );
  NAND U6396 ( .A(n5596), .B(n5595), .Z(n5597) );
  NAND U6397 ( .A(n5598), .B(n5597), .Z(n5684) );
  NAND U6398 ( .A(n5600), .B(n5599), .Z(n5604) );
  NAND U6399 ( .A(n5602), .B(n5601), .Z(n5603) );
  AND U6400 ( .A(n5604), .B(n5603), .Z(n5685) );
  XOR U6401 ( .A(n5684), .B(n5685), .Z(n5687) );
  XOR U6402 ( .A(n5686), .B(n5687), .Z(n5678) );
  NANDN U6403 ( .A(n5606), .B(n5605), .Z(n5610) );
  NAND U6404 ( .A(n5608), .B(n5607), .Z(n5609) );
  NAND U6405 ( .A(n5610), .B(n5609), .Z(n5679) );
  XNOR U6406 ( .A(n5678), .B(n5679), .Z(n5681) );
  NANDN U6407 ( .A(n5612), .B(n5611), .Z(n5616) );
  NAND U6408 ( .A(n5614), .B(n5613), .Z(n5615) );
  AND U6409 ( .A(n5616), .B(n5615), .Z(n5691) );
  AND U6410 ( .A(x[51]), .B(y[49]), .Z(n5618) );
  NAND U6411 ( .A(x[48]), .B(y[52]), .Z(n5617) );
  XNOR U6412 ( .A(n5618), .B(n5617), .Z(n5754) );
  NAND U6413 ( .A(y[50]), .B(x[50]), .Z(n5813) );
  IV U6414 ( .A(n5813), .Z(n5619) );
  XOR U6415 ( .A(n5754), .B(n5619), .Z(n5757) );
  NAND U6416 ( .A(y[51]), .B(x[49]), .Z(n5758) );
  AND U6417 ( .A(y[128]), .B(x[68]), .Z(n5701) );
  NAND U6418 ( .A(y[11]), .B(x[41]), .Z(n5702) );
  NAND U6419 ( .A(y[12]), .B(x[40]), .Z(n5704) );
  XOR U6420 ( .A(n5760), .B(n5759), .Z(n5772) );
  NANDN U6421 ( .A(n5621), .B(n5620), .Z(n5625) );
  OR U6422 ( .A(n5623), .B(n5622), .Z(n5624) );
  AND U6423 ( .A(n5625), .B(n5624), .Z(n5770) );
  AND U6424 ( .A(y[171]), .B(x[75]), .Z(n6053) );
  NANDN U6425 ( .A(n5626), .B(n6053), .Z(n5630) );
  NANDN U6426 ( .A(n5628), .B(n5627), .Z(n5629) );
  AND U6427 ( .A(n5630), .B(n5629), .Z(n5769) );
  NAND U6428 ( .A(y[8]), .B(x[44]), .Z(n5738) );
  NAND U6429 ( .A(y[130]), .B(x[66]), .Z(n5737) );
  NAND U6430 ( .A(y[92]), .B(x[56]), .Z(n5736) );
  XNOR U6431 ( .A(n5737), .B(n5736), .Z(n5739) );
  AND U6432 ( .A(y[170]), .B(x[74]), .Z(n5671) );
  NAND U6433 ( .A(n5671), .B(n5631), .Z(n5734) );
  NAND U6434 ( .A(y[172]), .B(x[72]), .Z(n5908) );
  NAND U6435 ( .A(y[88]), .B(x[60]), .Z(n5834) );
  XNOR U6436 ( .A(n5908), .B(n5834), .Z(n5735) );
  XOR U6437 ( .A(n5734), .B(n5735), .Z(n5717) );
  XOR U6438 ( .A(n5718), .B(n5717), .Z(n5720) );
  NAND U6439 ( .A(n5633), .B(n5632), .Z(n5637) );
  NAND U6440 ( .A(n5635), .B(n5634), .Z(n5636) );
  AND U6441 ( .A(n5637), .B(n5636), .Z(n5719) );
  XOR U6442 ( .A(n5720), .B(n5719), .Z(n5784) );
  NAND U6443 ( .A(n5639), .B(n5638), .Z(n5643) );
  NAND U6444 ( .A(n5641), .B(n5640), .Z(n5642) );
  AND U6445 ( .A(n5643), .B(n5642), .Z(n5783) );
  XNOR U6446 ( .A(n5784), .B(n5783), .Z(n5785) );
  XNOR U6447 ( .A(n5786), .B(n5785), .Z(n5690) );
  XNOR U6448 ( .A(n5691), .B(n5690), .Z(n5693) );
  NANDN U6449 ( .A(n5645), .B(n5644), .Z(n5649) );
  NANDN U6450 ( .A(n5647), .B(n5646), .Z(n5648) );
  AND U6451 ( .A(n5649), .B(n5648), .Z(n5776) );
  NANDN U6452 ( .A(n5651), .B(n5650), .Z(n5655) );
  OR U6453 ( .A(n5653), .B(n5652), .Z(n5654) );
  NAND U6454 ( .A(n5655), .B(n5654), .Z(n5775) );
  XNOR U6455 ( .A(n5776), .B(n5775), .Z(n5778) );
  AND U6456 ( .A(x[59]), .B(y[89]), .Z(n5662) );
  NAND U6457 ( .A(n5656), .B(n5662), .Z(n5660) );
  NANDN U6458 ( .A(n5658), .B(n5657), .Z(n5659) );
  AND U6459 ( .A(n5660), .B(n5659), .Z(n5780) );
  AND U6460 ( .A(y[48]), .B(x[52]), .Z(n5707) );
  NAND U6461 ( .A(y[132]), .B(x[64]), .Z(n5708) );
  NAND U6462 ( .A(y[131]), .B(x[65]), .Z(n5710) );
  NAND U6463 ( .A(x[58]), .B(y[90]), .Z(n5661) );
  XNOR U6464 ( .A(n5662), .B(n5661), .Z(n5697) );
  NAND U6465 ( .A(y[91]), .B(x[57]), .Z(n5698) );
  XOR U6466 ( .A(n5764), .B(n5763), .Z(n5765) );
  NAND U6467 ( .A(n5664), .B(n5663), .Z(n5668) );
  NAND U6468 ( .A(n5666), .B(n5665), .Z(n5667) );
  NAND U6469 ( .A(n5668), .B(n5667), .Z(n5766) );
  XNOR U6470 ( .A(n5780), .B(n5779), .Z(n5782) );
  NAND U6471 ( .A(y[10]), .B(x[42]), .Z(n5749) );
  NAND U6472 ( .A(y[129]), .B(x[67]), .Z(n5748) );
  NAND U6473 ( .A(y[9]), .B(x[43]), .Z(n5747) );
  XNOR U6474 ( .A(n5748), .B(n5747), .Z(n5750) );
  AND U6475 ( .A(x[76]), .B(y[168]), .Z(n5670) );
  NAND U6476 ( .A(x[73]), .B(y[171]), .Z(n5669) );
  XNOR U6477 ( .A(n5670), .B(n5669), .Z(n5731) );
  AND U6478 ( .A(y[169]), .B(x[75]), .Z(n5842) );
  XOR U6479 ( .A(n5842), .B(n5671), .Z(n5730) );
  XOR U6480 ( .A(n5731), .B(n5730), .Z(n5724) );
  XOR U6481 ( .A(n5723), .B(n5724), .Z(n5725) );
  NANDN U6482 ( .A(n5673), .B(n5672), .Z(n5677) );
  OR U6483 ( .A(n5675), .B(n5674), .Z(n5676) );
  NAND U6484 ( .A(n5677), .B(n5676), .Z(n5726) );
  XOR U6485 ( .A(n5782), .B(n5781), .Z(n5777) );
  XOR U6486 ( .A(n5778), .B(n5777), .Z(n5692) );
  XNOR U6487 ( .A(n5693), .B(n5692), .Z(n5680) );
  XNOR U6488 ( .A(n5681), .B(n5680), .Z(o[52]) );
  NANDN U6489 ( .A(n5679), .B(n5678), .Z(n5683) );
  NAND U6490 ( .A(n5681), .B(n5680), .Z(n5682) );
  AND U6491 ( .A(n5683), .B(n5682), .Z(n5932) );
  NAND U6492 ( .A(n5685), .B(n5684), .Z(n5689) );
  NAND U6493 ( .A(n5687), .B(n5686), .Z(n5688) );
  NAND U6494 ( .A(n5689), .B(n5688), .Z(n5933) );
  XNOR U6495 ( .A(n5932), .B(n5933), .Z(n5935) );
  NANDN U6496 ( .A(n5691), .B(n5690), .Z(n5695) );
  NAND U6497 ( .A(n5693), .B(n5692), .Z(n5694) );
  AND U6498 ( .A(n5695), .B(n5694), .Z(n5790) );
  AND U6499 ( .A(y[90]), .B(x[59]), .Z(n5835) );
  NAND U6500 ( .A(n5696), .B(n5835), .Z(n5700) );
  NANDN U6501 ( .A(n5698), .B(n5697), .Z(n5699) );
  AND U6502 ( .A(n5700), .B(n5699), .Z(n5796) );
  AND U6503 ( .A(y[133]), .B(x[64]), .Z(n6143) );
  AND U6504 ( .A(y[48]), .B(x[53]), .Z(n5825) );
  AND U6505 ( .A(y[91]), .B(x[58]), .Z(n5824) );
  XOR U6506 ( .A(n5825), .B(n5824), .Z(n5826) );
  XOR U6507 ( .A(n6143), .B(n5826), .Z(n5819) );
  AND U6508 ( .A(y[9]), .B(x[44]), .Z(n6121) );
  AND U6509 ( .A(y[129]), .B(x[68]), .Z(n5830) );
  AND U6510 ( .A(y[8]), .B(x[45]), .Z(n5829) );
  XOR U6511 ( .A(n5830), .B(n5829), .Z(n5831) );
  XOR U6512 ( .A(n6121), .B(n5831), .Z(n5818) );
  XOR U6513 ( .A(n5819), .B(n5818), .Z(n5821) );
  NANDN U6514 ( .A(n5702), .B(n5701), .Z(n5706) );
  NANDN U6515 ( .A(n5704), .B(n5703), .Z(n5705) );
  NAND U6516 ( .A(n5706), .B(n5705), .Z(n5820) );
  XOR U6517 ( .A(n5821), .B(n5820), .Z(n5795) );
  NANDN U6518 ( .A(n5708), .B(n5707), .Z(n5712) );
  NANDN U6519 ( .A(n5710), .B(n5709), .Z(n5711) );
  NAND U6520 ( .A(n5712), .B(n5711), .Z(n5899) );
  AND U6521 ( .A(y[170]), .B(x[75]), .Z(n5714) );
  AND U6522 ( .A(n5714), .B(n5713), .Z(n5910) );
  AND U6523 ( .A(x[72]), .B(y[173]), .Z(n5716) );
  AND U6524 ( .A(x[73]), .B(y[172]), .Z(n5715) );
  XOR U6525 ( .A(n5716), .B(n5715), .Z(n5909) );
  XOR U6526 ( .A(n5910), .B(n5909), .Z(n5898) );
  AND U6527 ( .A(y[49]), .B(x[52]), .Z(n5890) );
  AND U6528 ( .A(y[53]), .B(x[48]), .Z(n5888) );
  AND U6529 ( .A(y[12]), .B(x[41]), .Z(n5887) );
  XOR U6530 ( .A(n5888), .B(n5887), .Z(n5889) );
  XOR U6531 ( .A(n5890), .B(n5889), .Z(n5897) );
  XOR U6532 ( .A(n5898), .B(n5897), .Z(n5900) );
  XOR U6533 ( .A(n5899), .B(n5900), .Z(n5797) );
  XOR U6534 ( .A(n5798), .B(n5797), .Z(n5846) );
  NAND U6535 ( .A(n5718), .B(n5717), .Z(n5722) );
  NAND U6536 ( .A(n5720), .B(n5719), .Z(n5721) );
  AND U6537 ( .A(n5722), .B(n5721), .Z(n5844) );
  NAND U6538 ( .A(n5724), .B(n5723), .Z(n5728) );
  NANDN U6539 ( .A(n5726), .B(n5725), .Z(n5727) );
  NAND U6540 ( .A(n5728), .B(n5727), .Z(n5843) );
  XOR U6541 ( .A(n5846), .B(n5845), .Z(n5930) );
  AND U6542 ( .A(y[171]), .B(x[76]), .Z(n6135) );
  NAND U6543 ( .A(n6135), .B(n5729), .Z(n5733) );
  NAND U6544 ( .A(n5731), .B(n5730), .Z(n5732) );
  AND U6545 ( .A(n5733), .B(n5732), .Z(n5856) );
  NAND U6546 ( .A(n5737), .B(n5736), .Z(n5741) );
  NANDN U6547 ( .A(n5739), .B(n5738), .Z(n5740) );
  AND U6548 ( .A(n5741), .B(n5740), .Z(n5864) );
  AND U6549 ( .A(y[52]), .B(x[49]), .Z(n5814) );
  AND U6550 ( .A(x[50]), .B(y[51]), .Z(n5743) );
  NAND U6551 ( .A(x[51]), .B(y[50]), .Z(n5742) );
  XOR U6552 ( .A(n5743), .B(n5742), .Z(n5815) );
  AND U6553 ( .A(y[169]), .B(x[76]), .Z(n6117) );
  NAND U6554 ( .A(x[75]), .B(y[170]), .Z(n5744) );
  XNOR U6555 ( .A(n6117), .B(n5744), .Z(n5804) );
  AND U6556 ( .A(y[168]), .B(x[77]), .Z(n5801) );
  NAND U6557 ( .A(y[171]), .B(x[74]), .Z(n5802) );
  XOR U6558 ( .A(n5804), .B(n5803), .Z(n5861) );
  XOR U6559 ( .A(n5862), .B(n5861), .Z(n5863) );
  XOR U6560 ( .A(n5864), .B(n5863), .Z(n5857) );
  XOR U6561 ( .A(n5858), .B(n5857), .Z(n5876) );
  AND U6562 ( .A(x[60]), .B(y[89]), .Z(n5746) );
  NAND U6563 ( .A(x[61]), .B(y[88]), .Z(n5745) );
  XOR U6564 ( .A(n5746), .B(n5745), .Z(n5836) );
  AND U6565 ( .A(y[128]), .B(x[69]), .Z(n5807) );
  NAND U6566 ( .A(y[10]), .B(x[43]), .Z(n5808) );
  AND U6567 ( .A(y[11]), .B(x[42]), .Z(n5809) );
  XOR U6568 ( .A(n5810), .B(n5809), .Z(n5879) );
  XOR U6569 ( .A(n5880), .B(n5879), .Z(n5882) );
  NAND U6570 ( .A(n5748), .B(n5747), .Z(n5752) );
  NANDN U6571 ( .A(n5750), .B(n5749), .Z(n5751) );
  AND U6572 ( .A(n5752), .B(n5751), .Z(n5881) );
  XOR U6573 ( .A(n5882), .B(n5881), .Z(n5874) );
  AND U6574 ( .A(y[13]), .B(x[40]), .Z(n5914) );
  AND U6575 ( .A(y[132]), .B(x[65]), .Z(n5913) );
  XOR U6576 ( .A(n5914), .B(n5913), .Z(n5916) );
  AND U6577 ( .A(y[131]), .B(x[66]), .Z(n5915) );
  XOR U6578 ( .A(n5916), .B(n5915), .Z(n5850) );
  AND U6579 ( .A(y[130]), .B(x[67]), .Z(n5903) );
  AND U6580 ( .A(y[92]), .B(x[57]), .Z(n6069) );
  XOR U6581 ( .A(n5903), .B(n6069), .Z(n5905) );
  AND U6582 ( .A(y[93]), .B(x[56]), .Z(n5904) );
  XOR U6583 ( .A(n5905), .B(n5904), .Z(n5849) );
  XOR U6584 ( .A(n5850), .B(n5849), .Z(n5852) );
  AND U6585 ( .A(y[52]), .B(x[51]), .Z(n6134) );
  NAND U6586 ( .A(n6134), .B(n5753), .Z(n5756) );
  NANDN U6587 ( .A(n5813), .B(n5754), .Z(n5755) );
  NAND U6588 ( .A(n5756), .B(n5755), .Z(n5851) );
  XNOR U6589 ( .A(n5852), .B(n5851), .Z(n5873) );
  NANDN U6590 ( .A(n5758), .B(n5757), .Z(n5762) );
  NAND U6591 ( .A(n5760), .B(n5759), .Z(n5761) );
  AND U6592 ( .A(n5762), .B(n5761), .Z(n5868) );
  NAND U6593 ( .A(n5764), .B(n5763), .Z(n5768) );
  NANDN U6594 ( .A(n5766), .B(n5765), .Z(n5767) );
  NAND U6595 ( .A(n5768), .B(n5767), .Z(n5867) );
  NANDN U6596 ( .A(n5770), .B(n5769), .Z(n5774) );
  NANDN U6597 ( .A(n5772), .B(n5771), .Z(n5773) );
  NAND U6598 ( .A(n5774), .B(n5773), .Z(n5870) );
  XOR U6599 ( .A(n5928), .B(n5927), .Z(n5929) );
  XOR U6600 ( .A(n5930), .B(n5929), .Z(n5789) );
  XNOR U6601 ( .A(n5790), .B(n5789), .Z(n5791) );
  NANDN U6602 ( .A(n5784), .B(n5783), .Z(n5788) );
  NAND U6603 ( .A(n5786), .B(n5785), .Z(n5787) );
  AND U6604 ( .A(n5788), .B(n5787), .Z(n5921) );
  XNOR U6605 ( .A(n5922), .B(n5921), .Z(n5923) );
  XOR U6606 ( .A(n5924), .B(n5923), .Z(n5792) );
  XNOR U6607 ( .A(n5791), .B(n5792), .Z(n5934) );
  XOR U6608 ( .A(n5935), .B(n5934), .Z(o[53]) );
  NANDN U6609 ( .A(n5790), .B(n5789), .Z(n5794) );
  NANDN U6610 ( .A(n5792), .B(n5791), .Z(n5793) );
  AND U6611 ( .A(n5794), .B(n5793), .Z(n6219) );
  NANDN U6612 ( .A(n5796), .B(n5795), .Z(n5800) );
  NAND U6613 ( .A(n5798), .B(n5797), .Z(n5799) );
  AND U6614 ( .A(n5800), .B(n5799), .Z(n6224) );
  NANDN U6615 ( .A(n5802), .B(n5801), .Z(n5806) );
  NAND U6616 ( .A(n5804), .B(n5803), .Z(n5805) );
  NAND U6617 ( .A(n5806), .B(n5805), .Z(n6088) );
  NANDN U6618 ( .A(n5808), .B(n5807), .Z(n5812) );
  NAND U6619 ( .A(n5810), .B(n5809), .Z(n5811) );
  NAND U6620 ( .A(n5812), .B(n5811), .Z(n6091) );
  AND U6621 ( .A(x[51]), .B(y[51]), .Z(n5886) );
  NANDN U6622 ( .A(n5813), .B(n5886), .Z(n5817) );
  NANDN U6623 ( .A(n5815), .B(n5814), .Z(n5816) );
  AND U6624 ( .A(n5817), .B(n5816), .Z(n6047) );
  AND U6625 ( .A(y[131]), .B(x[67]), .Z(n6109) );
  AND U6626 ( .A(y[91]), .B(x[59]), .Z(n6108) );
  XOR U6627 ( .A(n6109), .B(n6108), .Z(n6107) );
  AND U6628 ( .A(y[11]), .B(x[43]), .Z(n6106) );
  XOR U6629 ( .A(n6107), .B(n6106), .Z(n6049) );
  AND U6630 ( .A(y[132]), .B(x[66]), .Z(n6149) );
  AND U6631 ( .A(y[90]), .B(x[60]), .Z(n6148) );
  XOR U6632 ( .A(n6149), .B(n6148), .Z(n6147) );
  AND U6633 ( .A(y[12]), .B(x[42]), .Z(n6146) );
  XNOR U6634 ( .A(n6147), .B(n6146), .Z(n6048) );
  XNOR U6635 ( .A(n6047), .B(n6046), .Z(n6090) );
  XOR U6636 ( .A(n6091), .B(n6090), .Z(n6089) );
  XOR U6637 ( .A(n6088), .B(n6089), .Z(n5948) );
  NAND U6638 ( .A(n5819), .B(n5818), .Z(n5823) );
  NAND U6639 ( .A(n5821), .B(n5820), .Z(n5822) );
  NAND U6640 ( .A(n5823), .B(n5822), .Z(n5947) );
  XOR U6641 ( .A(n5948), .B(n5947), .Z(n5946) );
  NAND U6642 ( .A(n5825), .B(n5824), .Z(n5828) );
  NAND U6643 ( .A(n6143), .B(n5826), .Z(n5827) );
  NAND U6644 ( .A(n5828), .B(n5827), .Z(n5972) );
  NAND U6645 ( .A(n5830), .B(n5829), .Z(n5833) );
  NAND U6646 ( .A(n6121), .B(n5831), .Z(n5832) );
  NAND U6647 ( .A(n5833), .B(n5832), .Z(n5971) );
  XOR U6648 ( .A(n5972), .B(n5971), .Z(n5970) );
  AND U6649 ( .A(y[89]), .B(x[61]), .Z(n6075) );
  NANDN U6650 ( .A(n5834), .B(n6075), .Z(n5838) );
  NANDN U6651 ( .A(n5836), .B(n5835), .Z(n5837) );
  AND U6652 ( .A(n5838), .B(n5837), .Z(n6095) );
  AND U6653 ( .A(x[45]), .B(y[9]), .Z(n5840) );
  NAND U6654 ( .A(x[44]), .B(y[10]), .Z(n5839) );
  XNOR U6655 ( .A(n5840), .B(n5839), .Z(n6119) );
  AND U6656 ( .A(y[128]), .B(x[70]), .Z(n6118) );
  XOR U6657 ( .A(n6119), .B(n6118), .Z(n6097) );
  AND U6658 ( .A(y[173]), .B(x[73]), .Z(n6061) );
  AND U6659 ( .A(y[170]), .B(x[76]), .Z(n5841) );
  AND U6660 ( .A(n5842), .B(n5841), .Z(n6059) );
  AND U6661 ( .A(y[172]), .B(x[74]), .Z(n6058) );
  XOR U6662 ( .A(n6059), .B(n6058), .Z(n6060) );
  XNOR U6663 ( .A(n6061), .B(n6060), .Z(n6096) );
  XNOR U6664 ( .A(n6095), .B(n6094), .Z(n5969) );
  XOR U6665 ( .A(n5970), .B(n5969), .Z(n5945) );
  XOR U6666 ( .A(n5946), .B(n5945), .Z(n5944) );
  NANDN U6667 ( .A(n5844), .B(n5843), .Z(n5848) );
  NAND U6668 ( .A(n5846), .B(n5845), .Z(n5847) );
  AND U6669 ( .A(n5848), .B(n5847), .Z(n5943) );
  NAND U6670 ( .A(n5850), .B(n5849), .Z(n5854) );
  NAND U6671 ( .A(n5852), .B(n5851), .Z(n5853) );
  AND U6672 ( .A(n5854), .B(n5853), .Z(n5952) );
  NANDN U6673 ( .A(n5856), .B(n5855), .Z(n5860) );
  NAND U6674 ( .A(n5858), .B(n5857), .Z(n5859) );
  AND U6675 ( .A(n5860), .B(n5859), .Z(n5951) );
  XOR U6676 ( .A(n5952), .B(n5951), .Z(n5950) );
  NAND U6677 ( .A(n5862), .B(n5861), .Z(n5866) );
  NAND U6678 ( .A(n5864), .B(n5863), .Z(n5865) );
  AND U6679 ( .A(n5866), .B(n5865), .Z(n5949) );
  XOR U6680 ( .A(n5950), .B(n5949), .Z(n5941) );
  XOR U6681 ( .A(n5942), .B(n5941), .Z(n6223) );
  XOR U6682 ( .A(n6224), .B(n6223), .Z(n6226) );
  NANDN U6683 ( .A(n5868), .B(n5867), .Z(n5872) );
  NANDN U6684 ( .A(n5870), .B(n5869), .Z(n5871) );
  AND U6685 ( .A(n5872), .B(n5871), .Z(n6203) );
  NANDN U6686 ( .A(n5874), .B(n5873), .Z(n5878) );
  NANDN U6687 ( .A(n5876), .B(n5875), .Z(n5877) );
  NAND U6688 ( .A(n5878), .B(n5877), .Z(n6204) );
  NAND U6689 ( .A(n5880), .B(n5879), .Z(n5884) );
  NAND U6690 ( .A(n5882), .B(n5881), .Z(n5883) );
  AND U6691 ( .A(n5884), .B(n5883), .Z(n6209) );
  AND U6692 ( .A(y[94]), .B(x[56]), .Z(n6103) );
  AND U6693 ( .A(y[8]), .B(x[46]), .Z(n6102) );
  XOR U6694 ( .A(n6103), .B(n6102), .Z(n6101) );
  AND U6695 ( .A(y[129]), .B(x[69]), .Z(n6100) );
  XOR U6696 ( .A(n6101), .B(n6100), .Z(n5978) );
  AND U6697 ( .A(y[49]), .B(x[53]), .Z(n6163) );
  AND U6698 ( .A(y[52]), .B(x[50]), .Z(n6162) );
  XOR U6699 ( .A(n6163), .B(n6162), .Z(n6161) );
  AND U6700 ( .A(y[53]), .B(x[49]), .Z(n6160) );
  XOR U6701 ( .A(n6161), .B(n6160), .Z(n5982) );
  NAND U6702 ( .A(x[52]), .B(y[50]), .Z(n5885) );
  XNOR U6703 ( .A(n5886), .B(n5885), .Z(n5981) );
  XOR U6704 ( .A(n5982), .B(n5981), .Z(n5977) );
  XOR U6705 ( .A(n5978), .B(n5977), .Z(n5976) );
  AND U6706 ( .A(y[174]), .B(x[72]), .Z(n6074) );
  XOR U6707 ( .A(n6075), .B(n6074), .Z(n6073) );
  AND U6708 ( .A(y[88]), .B(x[62]), .Z(n6072) );
  XOR U6709 ( .A(n6073), .B(n6072), .Z(n5975) );
  XOR U6710 ( .A(n5976), .B(n5975), .Z(n5961) );
  NAND U6711 ( .A(n5888), .B(n5887), .Z(n5892) );
  NAND U6712 ( .A(n5890), .B(n5889), .Z(n5891) );
  AND U6713 ( .A(n5892), .B(n5891), .Z(n6185) );
  AND U6714 ( .A(y[130]), .B(x[68]), .Z(n6067) );
  AND U6715 ( .A(x[57]), .B(y[93]), .Z(n5894) );
  AND U6716 ( .A(x[58]), .B(y[92]), .Z(n5893) );
  XOR U6717 ( .A(n5894), .B(n5893), .Z(n6066) );
  XNOR U6718 ( .A(n6067), .B(n6066), .Z(n6183) );
  AND U6719 ( .A(y[14]), .B(x[40]), .Z(n6141) );
  AND U6720 ( .A(y[134]), .B(x[64]), .Z(n5896) );
  AND U6721 ( .A(x[65]), .B(y[133]), .Z(n5895) );
  XOR U6722 ( .A(n5896), .B(n5895), .Z(n6140) );
  XOR U6723 ( .A(n6141), .B(n6140), .Z(n6182) );
  XNOR U6724 ( .A(n6185), .B(n6184), .Z(n5962) );
  NAND U6725 ( .A(n5898), .B(n5897), .Z(n5902) );
  NAND U6726 ( .A(n5900), .B(n5899), .Z(n5901) );
  AND U6727 ( .A(n5902), .B(n5901), .Z(n5963) );
  XOR U6728 ( .A(n5964), .B(n5963), .Z(n6208) );
  XOR U6729 ( .A(n6209), .B(n6208), .Z(n6211) );
  NAND U6730 ( .A(n5903), .B(n6069), .Z(n5907) );
  NAND U6731 ( .A(n5905), .B(n5904), .Z(n5906) );
  NAND U6732 ( .A(n5907), .B(n5906), .Z(n5955) );
  NANDN U6733 ( .A(n5908), .B(n6061), .Z(n5912) );
  NAND U6734 ( .A(n5910), .B(n5909), .Z(n5911) );
  NAND U6735 ( .A(n5912), .B(n5911), .Z(n5958) );
  NAND U6736 ( .A(n5914), .B(n5913), .Z(n5918) );
  NAND U6737 ( .A(n5916), .B(n5915), .Z(n5917) );
  AND U6738 ( .A(n5918), .B(n5917), .Z(n6177) );
  AND U6739 ( .A(y[13]), .B(x[41]), .Z(n6157) );
  AND U6740 ( .A(y[48]), .B(x[54]), .Z(n6156) );
  XOR U6741 ( .A(n6157), .B(n6156), .Z(n6155) );
  AND U6742 ( .A(y[54]), .B(x[48]), .Z(n6154) );
  XOR U6743 ( .A(n6155), .B(n6154), .Z(n6178) );
  AND U6744 ( .A(x[77]), .B(y[169]), .Z(n5920) );
  NAND U6745 ( .A(x[76]), .B(y[170]), .Z(n5919) );
  XNOR U6746 ( .A(n5920), .B(n5919), .Z(n6055) );
  AND U6747 ( .A(y[168]), .B(x[78]), .Z(n6054) );
  XOR U6748 ( .A(n6055), .B(n6054), .Z(n6052) );
  XNOR U6749 ( .A(n6053), .B(n6052), .Z(n6179) );
  XNOR U6750 ( .A(n6177), .B(n6176), .Z(n5957) );
  XOR U6751 ( .A(n5958), .B(n5957), .Z(n5956) );
  XOR U6752 ( .A(n5955), .B(n5956), .Z(n6210) );
  XOR U6753 ( .A(n6204), .B(n6205), .Z(n6202) );
  XOR U6754 ( .A(n6203), .B(n6202), .Z(n6225) );
  XOR U6755 ( .A(n6226), .B(n6225), .Z(n5940) );
  NANDN U6756 ( .A(n5922), .B(n5921), .Z(n5926) );
  NANDN U6757 ( .A(n5924), .B(n5923), .Z(n5925) );
  AND U6758 ( .A(n5926), .B(n5925), .Z(n5939) );
  XOR U6759 ( .A(n5939), .B(n5938), .Z(n5931) );
  XOR U6760 ( .A(n5940), .B(n5931), .Z(n6220) );
  NANDN U6761 ( .A(n5933), .B(n5932), .Z(n5937) );
  NAND U6762 ( .A(n5935), .B(n5934), .Z(n5936) );
  NAND U6763 ( .A(n5937), .B(n5936), .Z(n6217) );
  XOR U6764 ( .A(n6218), .B(n6217), .Z(o[54]) );
  NAND U6765 ( .A(n5950), .B(n5949), .Z(n5954) );
  NAND U6766 ( .A(n5952), .B(n5951), .Z(n5953) );
  AND U6767 ( .A(n5954), .B(n5953), .Z(n6201) );
  NAND U6768 ( .A(n5956), .B(n5955), .Z(n5960) );
  AND U6769 ( .A(n5958), .B(n5957), .Z(n5959) );
  ANDN U6770 ( .B(n5960), .A(n5959), .Z(n5968) );
  ANDN U6771 ( .B(n5962), .A(n5961), .Z(n5966) );
  AND U6772 ( .A(n5964), .B(n5963), .Z(n5965) );
  OR U6773 ( .A(n5966), .B(n5965), .Z(n5967) );
  XNOR U6774 ( .A(n5968), .B(n5967), .Z(n6199) );
  NAND U6775 ( .A(n5970), .B(n5969), .Z(n5974) );
  NAND U6776 ( .A(n5972), .B(n5971), .Z(n5973) );
  AND U6777 ( .A(n5974), .B(n5973), .Z(n6197) );
  NAND U6778 ( .A(n5976), .B(n5975), .Z(n5980) );
  NAND U6779 ( .A(n5978), .B(n5977), .Z(n5979) );
  AND U6780 ( .A(n5980), .B(n5979), .Z(n6087) );
  NAND U6781 ( .A(n5982), .B(n5981), .Z(n5985) );
  AND U6782 ( .A(y[50]), .B(x[51]), .Z(n5983) );
  AND U6783 ( .A(y[51]), .B(x[52]), .Z(n6035) );
  NAND U6784 ( .A(n5983), .B(n6035), .Z(n5984) );
  AND U6785 ( .A(n5985), .B(n5984), .Z(n6045) );
  AND U6786 ( .A(x[40]), .B(y[15]), .Z(n5987) );
  NAND U6787 ( .A(x[73]), .B(y[174]), .Z(n5986) );
  XNOR U6788 ( .A(n5987), .B(n5986), .Z(n5991) );
  AND U6789 ( .A(x[41]), .B(y[14]), .Z(n5989) );
  NAND U6790 ( .A(x[69]), .B(y[130]), .Z(n5988) );
  XNOR U6791 ( .A(n5989), .B(n5988), .Z(n5990) );
  XOR U6792 ( .A(n5991), .B(n5990), .Z(n5999) );
  AND U6793 ( .A(x[68]), .B(y[131]), .Z(n5993) );
  NAND U6794 ( .A(x[47]), .B(y[8]), .Z(n5992) );
  XNOR U6795 ( .A(n5993), .B(n5992), .Z(n5997) );
  AND U6796 ( .A(x[46]), .B(y[9]), .Z(n5995) );
  NAND U6797 ( .A(x[62]), .B(y[89]), .Z(n5994) );
  XNOR U6798 ( .A(n5995), .B(n5994), .Z(n5996) );
  XNOR U6799 ( .A(n5997), .B(n5996), .Z(n5998) );
  XNOR U6800 ( .A(n5999), .B(n5998), .Z(n6043) );
  AND U6801 ( .A(x[79]), .B(y[168]), .Z(n6004) );
  AND U6802 ( .A(y[170]), .B(x[77]), .Z(n6116) );
  AND U6803 ( .A(x[57]), .B(y[94]), .Z(n6001) );
  NAND U6804 ( .A(x[78]), .B(y[169]), .Z(n6000) );
  XNOR U6805 ( .A(n6001), .B(n6000), .Z(n6002) );
  XNOR U6806 ( .A(n6116), .B(n6002), .Z(n6003) );
  XNOR U6807 ( .A(n6004), .B(n6003), .Z(n6020) );
  AND U6808 ( .A(x[72]), .B(y[175]), .Z(n6006) );
  NAND U6809 ( .A(x[63]), .B(y[88]), .Z(n6005) );
  XNOR U6810 ( .A(n6006), .B(n6005), .Z(n6010) );
  AND U6811 ( .A(x[60]), .B(y[91]), .Z(n6008) );
  NAND U6812 ( .A(x[59]), .B(y[92]), .Z(n6007) );
  XNOR U6813 ( .A(n6008), .B(n6007), .Z(n6009) );
  XOR U6814 ( .A(n6010), .B(n6009), .Z(n6018) );
  AND U6815 ( .A(x[43]), .B(y[12]), .Z(n6012) );
  NAND U6816 ( .A(x[54]), .B(y[49]), .Z(n6011) );
  XNOR U6817 ( .A(n6012), .B(n6011), .Z(n6016) );
  AND U6818 ( .A(x[42]), .B(y[13]), .Z(n6014) );
  NAND U6819 ( .A(x[70]), .B(y[129]), .Z(n6013) );
  XNOR U6820 ( .A(n6014), .B(n6013), .Z(n6015) );
  XNOR U6821 ( .A(n6016), .B(n6015), .Z(n6017) );
  XNOR U6822 ( .A(n6018), .B(n6017), .Z(n6019) );
  XOR U6823 ( .A(n6020), .B(n6019), .Z(n6041) );
  AND U6824 ( .A(x[64]), .B(y[135]), .Z(n6022) );
  NAND U6825 ( .A(x[49]), .B(y[54]), .Z(n6021) );
  XNOR U6826 ( .A(n6022), .B(n6021), .Z(n6026) );
  AND U6827 ( .A(x[66]), .B(y[133]), .Z(n6024) );
  NAND U6828 ( .A(x[55]), .B(y[48]), .Z(n6023) );
  XNOR U6829 ( .A(n6024), .B(n6023), .Z(n6025) );
  XOR U6830 ( .A(n6026), .B(n6025), .Z(n6034) );
  AND U6831 ( .A(x[74]), .B(y[173]), .Z(n6028) );
  NAND U6832 ( .A(x[61]), .B(y[90]), .Z(n6027) );
  XNOR U6833 ( .A(n6028), .B(n6027), .Z(n6032) );
  AND U6834 ( .A(x[44]), .B(y[11]), .Z(n6030) );
  NAND U6835 ( .A(x[75]), .B(y[172]), .Z(n6029) );
  XNOR U6836 ( .A(n6030), .B(n6029), .Z(n6031) );
  XNOR U6837 ( .A(n6032), .B(n6031), .Z(n6033) );
  XNOR U6838 ( .A(n6034), .B(n6033), .Z(n6039) );
  AND U6839 ( .A(y[93]), .B(x[58]), .Z(n6068) );
  AND U6840 ( .A(y[134]), .B(x[65]), .Z(n6142) );
  XOR U6841 ( .A(n6068), .B(n6142), .Z(n6037) );
  AND U6842 ( .A(y[10]), .B(x[45]), .Z(n6120) );
  XNOR U6843 ( .A(n6120), .B(n6035), .Z(n6036) );
  XNOR U6844 ( .A(n6037), .B(n6036), .Z(n6038) );
  XNOR U6845 ( .A(n6039), .B(n6038), .Z(n6040) );
  XNOR U6846 ( .A(n6041), .B(n6040), .Z(n6042) );
  XNOR U6847 ( .A(n6043), .B(n6042), .Z(n6044) );
  XNOR U6848 ( .A(n6045), .B(n6044), .Z(n6085) );
  NAND U6849 ( .A(n6047), .B(n6046), .Z(n6051) );
  NANDN U6850 ( .A(n6049), .B(n6048), .Z(n6050) );
  AND U6851 ( .A(n6051), .B(n6050), .Z(n6083) );
  NAND U6852 ( .A(n6053), .B(n6052), .Z(n6057) );
  AND U6853 ( .A(n6055), .B(n6054), .Z(n6056) );
  ANDN U6854 ( .B(n6057), .A(n6056), .Z(n6065) );
  AND U6855 ( .A(n6059), .B(n6058), .Z(n6063) );
  AND U6856 ( .A(n6061), .B(n6060), .Z(n6062) );
  OR U6857 ( .A(n6063), .B(n6062), .Z(n6064) );
  XNOR U6858 ( .A(n6065), .B(n6064), .Z(n6081) );
  NAND U6859 ( .A(n6067), .B(n6066), .Z(n6071) );
  NAND U6860 ( .A(n6069), .B(n6068), .Z(n6070) );
  AND U6861 ( .A(n6071), .B(n6070), .Z(n6079) );
  NAND U6862 ( .A(n6073), .B(n6072), .Z(n6077) );
  NAND U6863 ( .A(n6075), .B(n6074), .Z(n6076) );
  NAND U6864 ( .A(n6077), .B(n6076), .Z(n6078) );
  XNOR U6865 ( .A(n6079), .B(n6078), .Z(n6080) );
  XNOR U6866 ( .A(n6081), .B(n6080), .Z(n6082) );
  XNOR U6867 ( .A(n6083), .B(n6082), .Z(n6084) );
  XNOR U6868 ( .A(n6085), .B(n6084), .Z(n6086) );
  XNOR U6869 ( .A(n6087), .B(n6086), .Z(n6195) );
  NAND U6870 ( .A(n6089), .B(n6088), .Z(n6093) );
  NAND U6871 ( .A(n6091), .B(n6090), .Z(n6092) );
  AND U6872 ( .A(n6093), .B(n6092), .Z(n6193) );
  NAND U6873 ( .A(n6095), .B(n6094), .Z(n6099) );
  NANDN U6874 ( .A(n6097), .B(n6096), .Z(n6098) );
  AND U6875 ( .A(n6099), .B(n6098), .Z(n6175) );
  NAND U6876 ( .A(n6101), .B(n6100), .Z(n6105) );
  NAND U6877 ( .A(n6103), .B(n6102), .Z(n6104) );
  AND U6878 ( .A(n6105), .B(n6104), .Z(n6113) );
  NAND U6879 ( .A(n6107), .B(n6106), .Z(n6111) );
  NAND U6880 ( .A(n6109), .B(n6108), .Z(n6110) );
  NAND U6881 ( .A(n6111), .B(n6110), .Z(n6112) );
  XNOR U6882 ( .A(n6113), .B(n6112), .Z(n6173) );
  AND U6883 ( .A(x[56]), .B(y[95]), .Z(n6115) );
  NAND U6884 ( .A(x[67]), .B(y[132]), .Z(n6114) );
  XNOR U6885 ( .A(n6115), .B(n6114), .Z(n6139) );
  AND U6886 ( .A(n6117), .B(n6116), .Z(n6133) );
  NAND U6887 ( .A(n6119), .B(n6118), .Z(n6123) );
  NAND U6888 ( .A(n6121), .B(n6120), .Z(n6122) );
  AND U6889 ( .A(n6123), .B(n6122), .Z(n6131) );
  AND U6890 ( .A(x[48]), .B(y[55]), .Z(n6125) );
  NAND U6891 ( .A(x[71]), .B(y[128]), .Z(n6124) );
  XNOR U6892 ( .A(n6125), .B(n6124), .Z(n6129) );
  AND U6893 ( .A(x[50]), .B(y[53]), .Z(n6127) );
  NAND U6894 ( .A(x[53]), .B(y[50]), .Z(n6126) );
  XNOR U6895 ( .A(n6127), .B(n6126), .Z(n6128) );
  XNOR U6896 ( .A(n6129), .B(n6128), .Z(n6130) );
  XNOR U6897 ( .A(n6131), .B(n6130), .Z(n6132) );
  XOR U6898 ( .A(n6133), .B(n6132), .Z(n6137) );
  XNOR U6899 ( .A(n6135), .B(n6134), .Z(n6136) );
  XNOR U6900 ( .A(n6137), .B(n6136), .Z(n6138) );
  XOR U6901 ( .A(n6139), .B(n6138), .Z(n6171) );
  NAND U6902 ( .A(n6141), .B(n6140), .Z(n6145) );
  NAND U6903 ( .A(n6143), .B(n6142), .Z(n6144) );
  AND U6904 ( .A(n6145), .B(n6144), .Z(n6153) );
  NAND U6905 ( .A(n6147), .B(n6146), .Z(n6151) );
  NAND U6906 ( .A(n6149), .B(n6148), .Z(n6150) );
  NAND U6907 ( .A(n6151), .B(n6150), .Z(n6152) );
  XNOR U6908 ( .A(n6153), .B(n6152), .Z(n6169) );
  NAND U6909 ( .A(n6155), .B(n6154), .Z(n6159) );
  NAND U6910 ( .A(n6157), .B(n6156), .Z(n6158) );
  AND U6911 ( .A(n6159), .B(n6158), .Z(n6167) );
  NAND U6912 ( .A(n6161), .B(n6160), .Z(n6165) );
  NAND U6913 ( .A(n6163), .B(n6162), .Z(n6164) );
  NAND U6914 ( .A(n6165), .B(n6164), .Z(n6166) );
  XNOR U6915 ( .A(n6167), .B(n6166), .Z(n6168) );
  XNOR U6916 ( .A(n6169), .B(n6168), .Z(n6170) );
  XNOR U6917 ( .A(n6171), .B(n6170), .Z(n6172) );
  XNOR U6918 ( .A(n6173), .B(n6172), .Z(n6174) );
  XNOR U6919 ( .A(n6175), .B(n6174), .Z(n6191) );
  NAND U6920 ( .A(n6177), .B(n6176), .Z(n6181) );
  ANDN U6921 ( .B(n6179), .A(n6178), .Z(n6180) );
  ANDN U6922 ( .B(n6181), .A(n6180), .Z(n6189) );
  ANDN U6923 ( .B(n6183), .A(n6182), .Z(n6187) );
  ANDN U6924 ( .B(n6185), .A(n6184), .Z(n6186) );
  OR U6925 ( .A(n6187), .B(n6186), .Z(n6188) );
  XNOR U6926 ( .A(n6189), .B(n6188), .Z(n6190) );
  XNOR U6927 ( .A(n6191), .B(n6190), .Z(n6192) );
  XNOR U6928 ( .A(n6193), .B(n6192), .Z(n6194) );
  XNOR U6929 ( .A(n6195), .B(n6194), .Z(n6196) );
  XNOR U6930 ( .A(n6197), .B(n6196), .Z(n6198) );
  XNOR U6931 ( .A(n6199), .B(n6198), .Z(n6200) );
  NAND U6932 ( .A(n6203), .B(n6202), .Z(n6207) );
  AND U6933 ( .A(n6205), .B(n6204), .Z(n6206) );
  ANDN U6934 ( .B(n6207), .A(n6206), .Z(n6215) );
  AND U6935 ( .A(n6209), .B(n6208), .Z(n6213) );
  ANDN U6936 ( .B(n6211), .A(n6210), .Z(n6212) );
  OR U6937 ( .A(n6213), .B(n6212), .Z(n6214) );
  XNOR U6938 ( .A(n6215), .B(n6214), .Z(n6216) );
  NAND U6939 ( .A(n6218), .B(n6217), .Z(n6222) );
  ANDN U6940 ( .B(n6220), .A(n6219), .Z(n6221) );
  AND U6941 ( .A(n6224), .B(n6223), .Z(n6228) );
  AND U6942 ( .A(n6226), .B(n6225), .Z(n6227) );
  NAND U6943 ( .A(y[176]), .B(x[72]), .Z(n6364) );
  NAND U6944 ( .A(y[56]), .B(x[48]), .Z(n6231) );
  XOR U6945 ( .A(n6364), .B(n6231), .Z(n6232) );
  AND U6946 ( .A(y[16]), .B(x[40]), .Z(n6239) );
  AND U6947 ( .A(y[96]), .B(x[56]), .Z(n6236) );
  XOR U6948 ( .A(n6239), .B(n6236), .Z(n6235) );
  AND U6949 ( .A(y[136]), .B(x[64]), .Z(n6234) );
  XNOR U6950 ( .A(n6235), .B(n6234), .Z(n6233) );
  XNOR U6951 ( .A(n6232), .B(n6233), .Z(o[56]) );
  AND U6952 ( .A(x[41]), .B(y[16]), .Z(n6230) );
  NAND U6953 ( .A(x[40]), .B(y[17]), .Z(n6229) );
  XNOR U6954 ( .A(n6230), .B(n6229), .Z(n6240) );
  NAND U6955 ( .A(y[56]), .B(x[49]), .Z(n6241) );
  XOR U6956 ( .A(n6240), .B(n6241), .Z(n6257) );
  AND U6957 ( .A(y[176]), .B(x[73]), .Z(n6465) );
  NAND U6958 ( .A(y[97]), .B(x[56]), .Z(n6244) );
  XNOR U6959 ( .A(n6465), .B(n6244), .Z(n6245) );
  AND U6960 ( .A(y[177]), .B(x[72]), .Z(n6269) );
  NAND U6961 ( .A(y[96]), .B(x[57]), .Z(n6268) );
  XOR U6962 ( .A(n6269), .B(n6268), .Z(n6246) );
  XOR U6963 ( .A(n6245), .B(n6246), .Z(n6256) );
  AND U6964 ( .A(y[57]), .B(x[48]), .Z(n6488) );
  AND U6965 ( .A(y[137]), .B(x[64]), .Z(n6261) );
  XOR U6966 ( .A(n6488), .B(n6261), .Z(n6263) );
  AND U6967 ( .A(y[136]), .B(x[65]), .Z(n6262) );
  XNOR U6968 ( .A(n6263), .B(n6262), .Z(n6255) );
  XOR U6969 ( .A(n6256), .B(n6255), .Z(n6258) );
  XOR U6970 ( .A(n6257), .B(n6258), .Z(n6252) );
  NAND U6971 ( .A(n6235), .B(n6234), .Z(n6238) );
  AND U6972 ( .A(n6239), .B(n6236), .Z(n6237) );
  ANDN U6973 ( .B(n6238), .A(n6237), .Z(n6249) );
  XNOR U6974 ( .A(n6250), .B(n6249), .Z(n6251) );
  XNOR U6975 ( .A(n6252), .B(n6251), .Z(o[57]) );
  AND U6976 ( .A(y[17]), .B(x[41]), .Z(n6299) );
  NAND U6977 ( .A(n6299), .B(n6239), .Z(n6243) );
  NANDN U6978 ( .A(n6241), .B(n6240), .Z(n6242) );
  NAND U6979 ( .A(n6243), .B(n6242), .Z(n6312) );
  NANDN U6980 ( .A(n6244), .B(n6465), .Z(n6248) );
  NANDN U6981 ( .A(n6246), .B(n6245), .Z(n6247) );
  NAND U6982 ( .A(n6248), .B(n6247), .Z(n6310) );
  AND U6983 ( .A(y[138]), .B(x[64]), .Z(n6316) );
  NAND U6984 ( .A(y[18]), .B(x[40]), .Z(n6317) );
  XNOR U6985 ( .A(n6316), .B(n6317), .Z(n6319) );
  AND U6986 ( .A(y[56]), .B(x[50]), .Z(n6318) );
  XOR U6987 ( .A(n6319), .B(n6318), .Z(n6311) );
  XOR U6988 ( .A(n6310), .B(n6311), .Z(n6313) );
  XNOR U6989 ( .A(n6312), .B(n6313), .Z(n6271) );
  NANDN U6990 ( .A(n6250), .B(n6249), .Z(n6254) );
  NAND U6991 ( .A(n6252), .B(n6251), .Z(n6253) );
  NAND U6992 ( .A(n6254), .B(n6253), .Z(n6270) );
  XOR U6993 ( .A(n6271), .B(n6270), .Z(n6273) );
  NAND U6994 ( .A(n6256), .B(n6255), .Z(n6260) );
  NAND U6995 ( .A(n6258), .B(n6257), .Z(n6259) );
  AND U6996 ( .A(n6260), .B(n6259), .Z(n6279) );
  AND U6997 ( .A(y[16]), .B(x[42]), .Z(n6297) );
  AND U6998 ( .A(y[98]), .B(x[56]), .Z(n6296) );
  XOR U6999 ( .A(n6297), .B(n6296), .Z(n6298) );
  XOR U7000 ( .A(n6299), .B(n6298), .Z(n6325) );
  AND U7001 ( .A(y[136]), .B(x[66]), .Z(n6324) );
  XOR U7002 ( .A(n6325), .B(n6324), .Z(n6327) );
  AND U7003 ( .A(y[96]), .B(x[58]), .Z(n6394) );
  AND U7004 ( .A(y[178]), .B(x[72]), .Z(n6288) );
  XOR U7005 ( .A(n6394), .B(n6288), .Z(n6290) );
  AND U7006 ( .A(y[97]), .B(x[57]), .Z(n6289) );
  XOR U7007 ( .A(n6290), .B(n6289), .Z(n6326) );
  XOR U7008 ( .A(n6327), .B(n6326), .Z(n6276) );
  AND U7009 ( .A(n6488), .B(n6261), .Z(n6265) );
  NAND U7010 ( .A(n6263), .B(n6262), .Z(n6264) );
  NANDN U7011 ( .A(n6265), .B(n6264), .Z(n6284) );
  AND U7012 ( .A(x[74]), .B(y[176]), .Z(n6267) );
  NAND U7013 ( .A(x[73]), .B(y[177]), .Z(n6266) );
  XNOR U7014 ( .A(n6267), .B(n6266), .Z(n6323) );
  ANDN U7015 ( .B(n6269), .A(n6268), .Z(n6322) );
  XOR U7016 ( .A(n6323), .B(n6322), .Z(n6283) );
  AND U7017 ( .A(y[137]), .B(x[65]), .Z(n6302) );
  NAND U7018 ( .A(y[57]), .B(x[49]), .Z(n6303) );
  XNOR U7019 ( .A(n6302), .B(n6303), .Z(n6304) );
  NAND U7020 ( .A(y[58]), .B(x[48]), .Z(n6305) );
  XNOR U7021 ( .A(n6304), .B(n6305), .Z(n6282) );
  XOR U7022 ( .A(n6283), .B(n6282), .Z(n6285) );
  XOR U7023 ( .A(n6284), .B(n6285), .Z(n6277) );
  XOR U7024 ( .A(n6276), .B(n6277), .Z(n6278) );
  XNOR U7025 ( .A(n6279), .B(n6278), .Z(n6272) );
  XNOR U7026 ( .A(n6273), .B(n6272), .Z(o[58]) );
  NAND U7027 ( .A(n6271), .B(n6270), .Z(n6275) );
  NAND U7028 ( .A(n6273), .B(n6272), .Z(n6274) );
  AND U7029 ( .A(n6275), .B(n6274), .Z(n6331) );
  NAND U7030 ( .A(n6277), .B(n6276), .Z(n6281) );
  NAND U7031 ( .A(n6279), .B(n6278), .Z(n6280) );
  NAND U7032 ( .A(n6281), .B(n6280), .Z(n6336) );
  NAND U7033 ( .A(n6283), .B(n6282), .Z(n6287) );
  NAND U7034 ( .A(n6285), .B(n6284), .Z(n6286) );
  NAND U7035 ( .A(n6287), .B(n6286), .Z(n6334) );
  AND U7036 ( .A(y[18]), .B(x[41]), .Z(n6360) );
  AND U7037 ( .A(y[17]), .B(x[42]), .Z(n6359) );
  NAND U7038 ( .A(y[138]), .B(x[65]), .Z(n6358) );
  XOR U7039 ( .A(n6359), .B(n6358), .Z(n6361) );
  XOR U7040 ( .A(n6360), .B(n6361), .Z(n6391) );
  NAND U7041 ( .A(n6394), .B(n6288), .Z(n6292) );
  AND U7042 ( .A(n6290), .B(n6289), .Z(n6291) );
  ANDN U7043 ( .B(n6292), .A(n6291), .Z(n6389) );
  AND U7044 ( .A(x[75]), .B(y[176]), .Z(n6294) );
  NAND U7045 ( .A(x[72]), .B(y[179]), .Z(n6293) );
  XNOR U7046 ( .A(n6294), .B(n6293), .Z(n6365) );
  AND U7047 ( .A(x[74]), .B(y[177]), .Z(n6461) );
  NAND U7048 ( .A(x[73]), .B(y[178]), .Z(n6295) );
  XOR U7049 ( .A(n6461), .B(n6295), .Z(n6366) );
  XNOR U7050 ( .A(n6365), .B(n6366), .Z(n6388) );
  XNOR U7051 ( .A(n6389), .B(n6388), .Z(n6390) );
  XNOR U7052 ( .A(n6391), .B(n6390), .Z(n6348) );
  NAND U7053 ( .A(n6297), .B(n6296), .Z(n6301) );
  NAND U7054 ( .A(n6299), .B(n6298), .Z(n6300) );
  NAND U7055 ( .A(n6301), .B(n6300), .Z(n6346) );
  NANDN U7056 ( .A(n6303), .B(n6302), .Z(n6307) );
  NANDN U7057 ( .A(n6305), .B(n6304), .Z(n6306) );
  AND U7058 ( .A(n6307), .B(n6306), .Z(n6384) );
  AND U7059 ( .A(y[139]), .B(x[64]), .Z(n6412) );
  AND U7060 ( .A(y[99]), .B(x[56]), .Z(n6411) );
  NAND U7061 ( .A(y[16]), .B(x[43]), .Z(n6410) );
  XOR U7062 ( .A(n6411), .B(n6410), .Z(n6413) );
  XOR U7063 ( .A(n6412), .B(n6413), .Z(n6383) );
  AND U7064 ( .A(x[59]), .B(y[96]), .Z(n6309) );
  NAND U7065 ( .A(x[58]), .B(y[97]), .Z(n6308) );
  XNOR U7066 ( .A(n6309), .B(n6308), .Z(n6395) );
  NAND U7067 ( .A(y[98]), .B(x[57]), .Z(n6396) );
  XOR U7068 ( .A(n6383), .B(n6382), .Z(n6385) );
  XOR U7069 ( .A(n6384), .B(n6385), .Z(n6347) );
  XOR U7070 ( .A(n6346), .B(n6347), .Z(n6349) );
  XOR U7071 ( .A(n6348), .B(n6349), .Z(n6335) );
  XOR U7072 ( .A(n6334), .B(n6335), .Z(n6337) );
  XOR U7073 ( .A(n6336), .B(n6337), .Z(n6330) );
  XOR U7074 ( .A(n6331), .B(n6330), .Z(n6333) );
  NAND U7075 ( .A(n6311), .B(n6310), .Z(n6315) );
  NAND U7076 ( .A(n6313), .B(n6312), .Z(n6314) );
  AND U7077 ( .A(n6315), .B(n6314), .Z(n6343) );
  NANDN U7078 ( .A(n6317), .B(n6316), .Z(n6321) );
  NAND U7079 ( .A(n6319), .B(n6318), .Z(n6320) );
  AND U7080 ( .A(n6321), .B(n6320), .Z(n6353) );
  XNOR U7081 ( .A(n6353), .B(n6352), .Z(n6355) );
  AND U7082 ( .A(y[56]), .B(x[51]), .Z(n6403) );
  AND U7083 ( .A(y[19]), .B(x[40]), .Z(n6402) );
  NAND U7084 ( .A(y[137]), .B(x[66]), .Z(n6401) );
  XOR U7085 ( .A(n6402), .B(n6401), .Z(n6404) );
  XOR U7086 ( .A(n6403), .B(n6404), .Z(n6379) );
  AND U7087 ( .A(y[59]), .B(x[48]), .Z(n6372) );
  AND U7088 ( .A(y[57]), .B(x[50]), .Z(n6371) );
  NAND U7089 ( .A(y[136]), .B(x[67]), .Z(n6370) );
  XOR U7090 ( .A(n6371), .B(n6370), .Z(n6373) );
  XOR U7091 ( .A(n6372), .B(n6373), .Z(n6377) );
  AND U7092 ( .A(y[58]), .B(x[49]), .Z(n6376) );
  XNOR U7093 ( .A(n6355), .B(n6354), .Z(n6341) );
  NAND U7094 ( .A(n6325), .B(n6324), .Z(n6329) );
  NAND U7095 ( .A(n6327), .B(n6326), .Z(n6328) );
  AND U7096 ( .A(n6329), .B(n6328), .Z(n6340) );
  XOR U7097 ( .A(n6341), .B(n6340), .Z(n6342) );
  XNOR U7098 ( .A(n6343), .B(n6342), .Z(n6332) );
  XOR U7099 ( .A(n6333), .B(n6332), .Z(o[59]) );
  NAND U7100 ( .A(n6335), .B(n6334), .Z(n6339) );
  NAND U7101 ( .A(n6337), .B(n6336), .Z(n6338) );
  AND U7102 ( .A(n6339), .B(n6338), .Z(n6422) );
  NAND U7103 ( .A(n6341), .B(n6340), .Z(n6345) );
  NAND U7104 ( .A(n6343), .B(n6342), .Z(n6344) );
  NAND U7105 ( .A(n6345), .B(n6344), .Z(n6420) );
  NAND U7106 ( .A(n6347), .B(n6346), .Z(n6351) );
  NAND U7107 ( .A(n6349), .B(n6348), .Z(n6350) );
  AND U7108 ( .A(n6351), .B(n6350), .Z(n6421) );
  XOR U7109 ( .A(n6420), .B(n6421), .Z(n6423) );
  XOR U7110 ( .A(n6422), .B(n6423), .Z(n6416) );
  XOR U7111 ( .A(n6417), .B(n6416), .Z(n6419) );
  AND U7112 ( .A(y[58]), .B(x[50]), .Z(n6563) );
  AND U7113 ( .A(x[48]), .B(y[60]), .Z(n6357) );
  NAND U7114 ( .A(x[51]), .B(y[57]), .Z(n6356) );
  XOR U7115 ( .A(n6357), .B(n6356), .Z(n6489) );
  XNOR U7116 ( .A(n6563), .B(n6489), .Z(n6498) );
  NAND U7117 ( .A(y[59]), .B(x[49]), .Z(n6499) );
  XNOR U7118 ( .A(n6498), .B(n6499), .Z(n6501) );
  AND U7119 ( .A(y[136]), .B(x[68]), .Z(n6449) );
  NAND U7120 ( .A(y[19]), .B(x[41]), .Z(n6450) );
  XNOR U7121 ( .A(n6449), .B(n6450), .Z(n6451) );
  NAND U7122 ( .A(y[20]), .B(x[40]), .Z(n6452) );
  XNOR U7123 ( .A(n6451), .B(n6452), .Z(n6500) );
  XOR U7124 ( .A(n6501), .B(n6500), .Z(n6495) );
  NANDN U7125 ( .A(n6359), .B(n6358), .Z(n6363) );
  OR U7126 ( .A(n6361), .B(n6360), .Z(n6362) );
  AND U7127 ( .A(n6363), .B(n6362), .Z(n6493) );
  AND U7128 ( .A(y[179]), .B(x[75]), .Z(n6788) );
  NANDN U7129 ( .A(n6364), .B(n6788), .Z(n6368) );
  NANDN U7130 ( .A(n6366), .B(n6365), .Z(n6367) );
  AND U7131 ( .A(n6368), .B(n6367), .Z(n6492) );
  XNOR U7132 ( .A(n6493), .B(n6492), .Z(n6494) );
  XNOR U7133 ( .A(n6495), .B(n6494), .Z(n6525) );
  NAND U7134 ( .A(y[16]), .B(x[44]), .Z(n6474) );
  NAND U7135 ( .A(y[138]), .B(x[66]), .Z(n6473) );
  NAND U7136 ( .A(y[100]), .B(x[56]), .Z(n6472) );
  XNOR U7137 ( .A(n6473), .B(n6472), .Z(n6475) );
  AND U7138 ( .A(y[177]), .B(x[73]), .Z(n6369) );
  AND U7139 ( .A(x[74]), .B(y[178]), .Z(n6409) );
  NAND U7140 ( .A(n6369), .B(n6409), .Z(n6470) );
  NAND U7141 ( .A(y[180]), .B(x[72]), .Z(n6623) );
  NAND U7142 ( .A(y[96]), .B(x[60]), .Z(n6582) );
  XNOR U7143 ( .A(n6623), .B(n6582), .Z(n6471) );
  XOR U7144 ( .A(n6470), .B(n6471), .Z(n6432) );
  XOR U7145 ( .A(n6433), .B(n6432), .Z(n6435) );
  NANDN U7146 ( .A(n6371), .B(n6370), .Z(n6375) );
  OR U7147 ( .A(n6373), .B(n6372), .Z(n6374) );
  AND U7148 ( .A(n6375), .B(n6374), .Z(n6434) );
  XOR U7149 ( .A(n6435), .B(n6434), .Z(n6523) );
  NANDN U7150 ( .A(n6377), .B(n6376), .Z(n6381) );
  NANDN U7151 ( .A(n6379), .B(n6378), .Z(n6380) );
  AND U7152 ( .A(n6381), .B(n6380), .Z(n6522) );
  XNOR U7153 ( .A(n6525), .B(n6524), .Z(n6426) );
  XNOR U7154 ( .A(n6427), .B(n6426), .Z(n6429) );
  NANDN U7155 ( .A(n6383), .B(n6382), .Z(n6387) );
  OR U7156 ( .A(n6385), .B(n6384), .Z(n6386) );
  AND U7157 ( .A(n6387), .B(n6386), .Z(n6511) );
  NANDN U7158 ( .A(n6389), .B(n6388), .Z(n6393) );
  NANDN U7159 ( .A(n6391), .B(n6390), .Z(n6392) );
  NAND U7160 ( .A(n6393), .B(n6392), .Z(n6510) );
  AND U7161 ( .A(y[97]), .B(x[59]), .Z(n6400) );
  NAND U7162 ( .A(n6400), .B(n6394), .Z(n6398) );
  NANDN U7163 ( .A(n6396), .B(n6395), .Z(n6397) );
  AND U7164 ( .A(n6398), .B(n6397), .Z(n6517) );
  AND U7165 ( .A(y[56]), .B(x[52]), .Z(n6455) );
  NAND U7166 ( .A(y[140]), .B(x[64]), .Z(n6456) );
  XNOR U7167 ( .A(n6455), .B(n6456), .Z(n6457) );
  NAND U7168 ( .A(y[139]), .B(x[65]), .Z(n6458) );
  XNOR U7169 ( .A(n6457), .B(n6458), .Z(n6504) );
  NAND U7170 ( .A(x[58]), .B(y[98]), .Z(n6399) );
  XNOR U7171 ( .A(n6400), .B(n6399), .Z(n6445) );
  NAND U7172 ( .A(y[99]), .B(x[57]), .Z(n6446) );
  XOR U7173 ( .A(n6445), .B(n6446), .Z(n6505) );
  XNOR U7174 ( .A(n6504), .B(n6505), .Z(n6506) );
  NANDN U7175 ( .A(n6402), .B(n6401), .Z(n6406) );
  OR U7176 ( .A(n6404), .B(n6403), .Z(n6405) );
  NAND U7177 ( .A(n6406), .B(n6405), .Z(n6507) );
  XNOR U7178 ( .A(n6506), .B(n6507), .Z(n6516) );
  NAND U7179 ( .A(y[18]), .B(x[42]), .Z(n6484) );
  NAND U7180 ( .A(y[137]), .B(x[67]), .Z(n6483) );
  NAND U7181 ( .A(y[17]), .B(x[43]), .Z(n6482) );
  XNOR U7182 ( .A(n6483), .B(n6482), .Z(n6485) );
  AND U7183 ( .A(x[76]), .B(y[176]), .Z(n6408) );
  NAND U7184 ( .A(x[73]), .B(y[179]), .Z(n6407) );
  XNOR U7185 ( .A(n6408), .B(n6407), .Z(n6467) );
  AND U7186 ( .A(y[177]), .B(x[75]), .Z(n6589) );
  XOR U7187 ( .A(n6589), .B(n6409), .Z(n6466) );
  XOR U7188 ( .A(n6467), .B(n6466), .Z(n6438) );
  XOR U7189 ( .A(n6439), .B(n6438), .Z(n6440) );
  NANDN U7190 ( .A(n6411), .B(n6410), .Z(n6415) );
  OR U7191 ( .A(n6413), .B(n6412), .Z(n6414) );
  NAND U7192 ( .A(n6415), .B(n6414), .Z(n6441) );
  XOR U7193 ( .A(n6440), .B(n6441), .Z(n6519) );
  XOR U7194 ( .A(n6513), .B(n6512), .Z(n6428) );
  XNOR U7195 ( .A(n6429), .B(n6428), .Z(n6418) );
  XNOR U7196 ( .A(n6419), .B(n6418), .Z(o[60]) );
  NAND U7197 ( .A(n6421), .B(n6420), .Z(n6425) );
  NAND U7198 ( .A(n6423), .B(n6422), .Z(n6424) );
  NAND U7199 ( .A(n6425), .B(n6424), .Z(n6666) );
  XNOR U7200 ( .A(n6665), .B(n6666), .Z(n6668) );
  NANDN U7201 ( .A(n6427), .B(n6426), .Z(n6431) );
  NAND U7202 ( .A(n6429), .B(n6428), .Z(n6430) );
  AND U7203 ( .A(n6431), .B(n6430), .Z(n6529) );
  NAND U7204 ( .A(n6433), .B(n6432), .Z(n6437) );
  NAND U7205 ( .A(n6435), .B(n6434), .Z(n6436) );
  AND U7206 ( .A(n6437), .B(n6436), .Z(n6592) );
  NAND U7207 ( .A(n6439), .B(n6438), .Z(n6443) );
  NANDN U7208 ( .A(n6441), .B(n6440), .Z(n6442) );
  NAND U7209 ( .A(n6443), .B(n6442), .Z(n6591) );
  XNOR U7210 ( .A(n6592), .B(n6591), .Z(n6594) );
  AND U7211 ( .A(y[97]), .B(x[58]), .Z(n6444) );
  AND U7212 ( .A(y[98]), .B(x[59]), .Z(n6583) );
  NAND U7213 ( .A(n6444), .B(n6583), .Z(n6448) );
  NANDN U7214 ( .A(n6446), .B(n6445), .Z(n6447) );
  NAND U7215 ( .A(n6448), .B(n6447), .Z(n6544) );
  NANDN U7216 ( .A(n6450), .B(n6449), .Z(n6454) );
  NANDN U7217 ( .A(n6452), .B(n6451), .Z(n6453) );
  NAND U7218 ( .A(n6454), .B(n6453), .Z(n6570) );
  AND U7219 ( .A(y[56]), .B(x[53]), .Z(n6573) );
  AND U7220 ( .A(y[99]), .B(x[58]), .Z(n6572) );
  XOR U7221 ( .A(n6573), .B(n6572), .Z(n6574) );
  AND U7222 ( .A(y[141]), .B(x[64]), .Z(n6852) );
  XOR U7223 ( .A(n6574), .B(n6852), .Z(n6569) );
  AND U7224 ( .A(y[137]), .B(x[68]), .Z(n6578) );
  AND U7225 ( .A(y[16]), .B(x[45]), .Z(n6577) );
  XOR U7226 ( .A(n6578), .B(n6577), .Z(n6579) );
  AND U7227 ( .A(y[17]), .B(x[44]), .Z(n6869) );
  XOR U7228 ( .A(n6579), .B(n6869), .Z(n6568) );
  XOR U7229 ( .A(n6569), .B(n6568), .Z(n6571) );
  XOR U7230 ( .A(n6570), .B(n6571), .Z(n6545) );
  XOR U7231 ( .A(n6544), .B(n6545), .Z(n6546) );
  NANDN U7232 ( .A(n6456), .B(n6455), .Z(n6460) );
  NANDN U7233 ( .A(n6458), .B(n6457), .Z(n6459) );
  NAND U7234 ( .A(n6460), .B(n6459), .Z(n6643) );
  AND U7235 ( .A(y[178]), .B(x[75]), .Z(n6462) );
  AND U7236 ( .A(n6462), .B(n6461), .Z(n6625) );
  AND U7237 ( .A(x[72]), .B(y[181]), .Z(n6464) );
  AND U7238 ( .A(x[73]), .B(y[180]), .Z(n6463) );
  XOR U7239 ( .A(n6464), .B(n6463), .Z(n6624) );
  XOR U7240 ( .A(n6625), .B(n6624), .Z(n6642) );
  AND U7241 ( .A(y[61]), .B(x[48]), .Z(n6650) );
  AND U7242 ( .A(y[20]), .B(x[41]), .Z(n6649) );
  XOR U7243 ( .A(n6650), .B(n6649), .Z(n6652) );
  AND U7244 ( .A(y[57]), .B(x[52]), .Z(n6651) );
  XOR U7245 ( .A(n6652), .B(n6651), .Z(n6641) );
  XOR U7246 ( .A(n6642), .B(n6641), .Z(n6644) );
  XNOR U7247 ( .A(n6643), .B(n6644), .Z(n6547) );
  XOR U7248 ( .A(n6594), .B(n6593), .Z(n6535) );
  AND U7249 ( .A(y[179]), .B(x[76]), .Z(n6882) );
  NAND U7250 ( .A(n6882), .B(n6465), .Z(n6469) );
  NAND U7251 ( .A(n6467), .B(n6466), .Z(n6468) );
  AND U7252 ( .A(n6469), .B(n6468), .Z(n6600) );
  XNOR U7253 ( .A(n6600), .B(n6599), .Z(n6602) );
  NAND U7254 ( .A(n6473), .B(n6472), .Z(n6477) );
  NANDN U7255 ( .A(n6475), .B(n6474), .Z(n6476) );
  AND U7256 ( .A(n6477), .B(n6476), .Z(n6608) );
  AND U7257 ( .A(y[58]), .B(x[51]), .Z(n6717) );
  NAND U7258 ( .A(x[50]), .B(y[59]), .Z(n6478) );
  XNOR U7259 ( .A(n6717), .B(n6478), .Z(n6564) );
  NAND U7260 ( .A(y[60]), .B(x[49]), .Z(n6565) );
  XNOR U7261 ( .A(n6564), .B(n6565), .Z(n6606) );
  AND U7262 ( .A(y[179]), .B(x[74]), .Z(n6550) );
  NAND U7263 ( .A(y[176]), .B(x[77]), .Z(n6551) );
  XNOR U7264 ( .A(n6550), .B(n6551), .Z(n6552) );
  AND U7265 ( .A(y[177]), .B(x[76]), .Z(n6866) );
  NAND U7266 ( .A(x[75]), .B(y[178]), .Z(n6479) );
  XOR U7267 ( .A(n6866), .B(n6479), .Z(n6553) );
  XNOR U7268 ( .A(n6552), .B(n6553), .Z(n6605) );
  XOR U7269 ( .A(n6606), .B(n6605), .Z(n6607) );
  XOR U7270 ( .A(n6608), .B(n6607), .Z(n6601) );
  XOR U7271 ( .A(n6602), .B(n6601), .Z(n6619) );
  AND U7272 ( .A(x[61]), .B(y[96]), .Z(n6481) );
  NAND U7273 ( .A(x[60]), .B(y[97]), .Z(n6480) );
  XOR U7274 ( .A(n6481), .B(n6480), .Z(n6584) );
  XNOR U7275 ( .A(n6583), .B(n6584), .Z(n6660) );
  AND U7276 ( .A(y[136]), .B(x[69]), .Z(n6556) );
  NAND U7277 ( .A(y[18]), .B(x[43]), .Z(n6557) );
  XNOR U7278 ( .A(n6556), .B(n6557), .Z(n6559) );
  AND U7279 ( .A(y[19]), .B(x[42]), .Z(n6558) );
  XOR U7280 ( .A(n6559), .B(n6558), .Z(n6659) );
  XOR U7281 ( .A(n6660), .B(n6659), .Z(n6662) );
  NAND U7282 ( .A(n6483), .B(n6482), .Z(n6487) );
  NANDN U7283 ( .A(n6485), .B(n6484), .Z(n6486) );
  AND U7284 ( .A(n6487), .B(n6486), .Z(n6661) );
  XOR U7285 ( .A(n6662), .B(n6661), .Z(n6618) );
  AND U7286 ( .A(y[60]), .B(x[51]), .Z(n6770) );
  NAND U7287 ( .A(n6770), .B(n6488), .Z(n6491) );
  NANDN U7288 ( .A(n6489), .B(n6563), .Z(n6490) );
  AND U7289 ( .A(n6491), .B(n6490), .Z(n6598) );
  AND U7290 ( .A(y[138]), .B(x[67]), .Z(n6636) );
  AND U7291 ( .A(y[100]), .B(x[57]), .Z(n6804) );
  XOR U7292 ( .A(n6636), .B(n6804), .Z(n6638) );
  AND U7293 ( .A(y[101]), .B(x[56]), .Z(n6637) );
  XOR U7294 ( .A(n6638), .B(n6637), .Z(n6596) );
  AND U7295 ( .A(y[21]), .B(x[40]), .Z(n6629) );
  AND U7296 ( .A(y[140]), .B(x[65]), .Z(n6628) );
  XOR U7297 ( .A(n6629), .B(n6628), .Z(n6631) );
  AND U7298 ( .A(y[139]), .B(x[66]), .Z(n6630) );
  XOR U7299 ( .A(n6631), .B(n6630), .Z(n6595) );
  XOR U7300 ( .A(n6596), .B(n6595), .Z(n6597) );
  XOR U7301 ( .A(n6598), .B(n6597), .Z(n6617) );
  XOR U7302 ( .A(n6618), .B(n6617), .Z(n6620) );
  XOR U7303 ( .A(n6619), .B(n6620), .Z(n6533) );
  NANDN U7304 ( .A(n6493), .B(n6492), .Z(n6497) );
  NANDN U7305 ( .A(n6495), .B(n6494), .Z(n6496) );
  AND U7306 ( .A(n6497), .B(n6496), .Z(n6613) );
  NANDN U7307 ( .A(n6499), .B(n6498), .Z(n6503) );
  NAND U7308 ( .A(n6501), .B(n6500), .Z(n6502) );
  AND U7309 ( .A(n6503), .B(n6502), .Z(n6612) );
  NANDN U7310 ( .A(n6505), .B(n6504), .Z(n6509) );
  NANDN U7311 ( .A(n6507), .B(n6506), .Z(n6508) );
  NAND U7312 ( .A(n6509), .B(n6508), .Z(n6611) );
  XOR U7313 ( .A(n6612), .B(n6611), .Z(n6614) );
  XNOR U7314 ( .A(n6613), .B(n6614), .Z(n6532) );
  XOR U7315 ( .A(n6535), .B(n6534), .Z(n6528) );
  XNOR U7316 ( .A(n6529), .B(n6528), .Z(n6531) );
  NANDN U7317 ( .A(n6511), .B(n6510), .Z(n6515) );
  NAND U7318 ( .A(n6513), .B(n6512), .Z(n6514) );
  AND U7319 ( .A(n6515), .B(n6514), .Z(n6541) );
  NANDN U7320 ( .A(n6517), .B(n6516), .Z(n6521) );
  NANDN U7321 ( .A(n6519), .B(n6518), .Z(n6520) );
  AND U7322 ( .A(n6521), .B(n6520), .Z(n6539) );
  NANDN U7323 ( .A(n6523), .B(n6522), .Z(n6527) );
  NAND U7324 ( .A(n6525), .B(n6524), .Z(n6526) );
  AND U7325 ( .A(n6527), .B(n6526), .Z(n6538) );
  XOR U7326 ( .A(n6531), .B(n6530), .Z(n6667) );
  XOR U7327 ( .A(n6668), .B(n6667), .Z(o[61]) );
  NANDN U7328 ( .A(n6533), .B(n6532), .Z(n6537) );
  NAND U7329 ( .A(n6535), .B(n6534), .Z(n6536) );
  AND U7330 ( .A(n6537), .B(n6536), .Z(n6962) );
  NANDN U7331 ( .A(n6539), .B(n6538), .Z(n6543) );
  NANDN U7332 ( .A(n6541), .B(n6540), .Z(n6542) );
  NAND U7333 ( .A(n6543), .B(n6542), .Z(n6963) );
  NAND U7334 ( .A(n6545), .B(n6544), .Z(n6549) );
  NANDN U7335 ( .A(n6547), .B(n6546), .Z(n6548) );
  AND U7336 ( .A(n6549), .B(n6548), .Z(n6973) );
  NANDN U7337 ( .A(n6551), .B(n6550), .Z(n6555) );
  NANDN U7338 ( .A(n6553), .B(n6552), .Z(n6554) );
  NAND U7339 ( .A(n6555), .B(n6554), .Z(n6703) );
  NANDN U7340 ( .A(n6557), .B(n6556), .Z(n6561) );
  NAND U7341 ( .A(n6559), .B(n6558), .Z(n6560) );
  NAND U7342 ( .A(n6561), .B(n6560), .Z(n6706) );
  AND U7343 ( .A(y[59]), .B(x[51]), .Z(n6562) );
  NAND U7344 ( .A(n6563), .B(n6562), .Z(n6567) );
  NANDN U7345 ( .A(n6565), .B(n6564), .Z(n6566) );
  AND U7346 ( .A(n6567), .B(n6566), .Z(n6782) );
  AND U7347 ( .A(y[139]), .B(x[67]), .Z(n6911) );
  AND U7348 ( .A(y[99]), .B(x[59]), .Z(n6910) );
  XOR U7349 ( .A(n6911), .B(n6910), .Z(n6909) );
  AND U7350 ( .A(y[19]), .B(x[43]), .Z(n6908) );
  XOR U7351 ( .A(n6909), .B(n6908), .Z(n6784) );
  AND U7352 ( .A(y[140]), .B(x[66]), .Z(n6897) );
  AND U7353 ( .A(y[98]), .B(x[60]), .Z(n6896) );
  XOR U7354 ( .A(n6897), .B(n6896), .Z(n6895) );
  AND U7355 ( .A(y[20]), .B(x[42]), .Z(n6894) );
  XNOR U7356 ( .A(n6895), .B(n6894), .Z(n6783) );
  XNOR U7357 ( .A(n6782), .B(n6781), .Z(n6705) );
  XOR U7358 ( .A(n6706), .B(n6705), .Z(n6704) );
  XOR U7359 ( .A(n6703), .B(n6704), .Z(n6680) );
  XOR U7360 ( .A(n6680), .B(n6679), .Z(n6678) );
  NAND U7361 ( .A(n6573), .B(n6572), .Z(n6576) );
  NAND U7362 ( .A(n6574), .B(n6852), .Z(n6575) );
  NAND U7363 ( .A(n6576), .B(n6575), .Z(n6826) );
  NAND U7364 ( .A(n6578), .B(n6577), .Z(n6581) );
  NAND U7365 ( .A(n6579), .B(n6869), .Z(n6580) );
  NAND U7366 ( .A(n6581), .B(n6580), .Z(n6825) );
  XOR U7367 ( .A(n6826), .B(n6825), .Z(n6823) );
  AND U7368 ( .A(y[97]), .B(x[61]), .Z(n6810) );
  NANDN U7369 ( .A(n6582), .B(n6810), .Z(n6586) );
  NANDN U7370 ( .A(n6584), .B(n6583), .Z(n6585) );
  AND U7371 ( .A(n6586), .B(n6585), .Z(n6838) );
  AND U7372 ( .A(x[44]), .B(y[18]), .Z(n6588) );
  NAND U7373 ( .A(x[45]), .B(y[17]), .Z(n6587) );
  XNOR U7374 ( .A(n6588), .B(n6587), .Z(n6868) );
  AND U7375 ( .A(y[136]), .B(x[70]), .Z(n6867) );
  XNOR U7376 ( .A(n6868), .B(n6867), .Z(n6836) );
  AND U7377 ( .A(y[181]), .B(x[73]), .Z(n6796) );
  AND U7378 ( .A(y[178]), .B(x[76]), .Z(n6590) );
  AND U7379 ( .A(n6590), .B(n6589), .Z(n6794) );
  AND U7380 ( .A(y[180]), .B(x[74]), .Z(n6793) );
  XOR U7381 ( .A(n6794), .B(n6793), .Z(n6795) );
  XOR U7382 ( .A(n6796), .B(n6795), .Z(n6835) );
  XNOR U7383 ( .A(n6838), .B(n6837), .Z(n6824) );
  XOR U7384 ( .A(n6678), .B(n6677), .Z(n6674) );
  NANDN U7385 ( .A(n6600), .B(n6599), .Z(n6604) );
  NAND U7386 ( .A(n6602), .B(n6601), .Z(n6603) );
  AND U7387 ( .A(n6604), .B(n6603), .Z(n6697) );
  XOR U7388 ( .A(n6698), .B(n6697), .Z(n6696) );
  NAND U7389 ( .A(n6606), .B(n6605), .Z(n6610) );
  NAND U7390 ( .A(n6608), .B(n6607), .Z(n6609) );
  AND U7391 ( .A(n6610), .B(n6609), .Z(n6695) );
  XOR U7392 ( .A(n6696), .B(n6695), .Z(n6671) );
  XOR U7393 ( .A(n6672), .B(n6671), .Z(n6972) );
  XOR U7394 ( .A(n6973), .B(n6972), .Z(n6975) );
  NANDN U7395 ( .A(n6612), .B(n6611), .Z(n6616) );
  NANDN U7396 ( .A(n6614), .B(n6613), .Z(n6615) );
  AND U7397 ( .A(n6616), .B(n6615), .Z(n6937) );
  NANDN U7398 ( .A(n6618), .B(n6617), .Z(n6622) );
  OR U7399 ( .A(n6620), .B(n6619), .Z(n6621) );
  AND U7400 ( .A(n6622), .B(n6621), .Z(n6939) );
  NANDN U7401 ( .A(n6623), .B(n6796), .Z(n6627) );
  NAND U7402 ( .A(n6625), .B(n6624), .Z(n6626) );
  AND U7403 ( .A(n6627), .B(n6626), .Z(n6692) );
  NAND U7404 ( .A(n6629), .B(n6628), .Z(n6633) );
  NAND U7405 ( .A(n6631), .B(n6630), .Z(n6632) );
  AND U7406 ( .A(n6633), .B(n6632), .Z(n6830) );
  AND U7407 ( .A(y[21]), .B(x[41]), .Z(n6891) );
  AND U7408 ( .A(y[56]), .B(x[54]), .Z(n6890) );
  XOR U7409 ( .A(n6891), .B(n6890), .Z(n6889) );
  AND U7410 ( .A(y[62]), .B(x[48]), .Z(n6888) );
  XOR U7411 ( .A(n6889), .B(n6888), .Z(n6831) );
  AND U7412 ( .A(x[77]), .B(y[177]), .Z(n6635) );
  NAND U7413 ( .A(x[76]), .B(y[178]), .Z(n6634) );
  XNOR U7414 ( .A(n6635), .B(n6634), .Z(n6790) );
  AND U7415 ( .A(y[176]), .B(x[78]), .Z(n6789) );
  XOR U7416 ( .A(n6790), .B(n6789), .Z(n6787) );
  XNOR U7417 ( .A(n6788), .B(n6787), .Z(n6832) );
  XNOR U7418 ( .A(n6830), .B(n6829), .Z(n6691) );
  NAND U7419 ( .A(n6636), .B(n6804), .Z(n6640) );
  NAND U7420 ( .A(n6638), .B(n6637), .Z(n6639) );
  AND U7421 ( .A(n6640), .B(n6639), .Z(n6690) );
  XNOR U7422 ( .A(n6689), .B(n6690), .Z(n6944) );
  NAND U7423 ( .A(n6642), .B(n6641), .Z(n6646) );
  NAND U7424 ( .A(n6644), .B(n6643), .Z(n6645) );
  AND U7425 ( .A(n6646), .B(n6645), .Z(n6684) );
  AND U7426 ( .A(y[102]), .B(x[56]), .Z(n6905) );
  AND U7427 ( .A(y[16]), .B(x[46]), .Z(n6904) );
  XOR U7428 ( .A(n6905), .B(n6904), .Z(n6903) );
  AND U7429 ( .A(y[137]), .B(x[69]), .Z(n6902) );
  XOR U7430 ( .A(n6903), .B(n6902), .Z(n6712) );
  AND U7431 ( .A(y[57]), .B(x[53]), .Z(n6858) );
  AND U7432 ( .A(y[60]), .B(x[50]), .Z(n6857) );
  XOR U7433 ( .A(n6858), .B(n6857), .Z(n6856) );
  AND U7434 ( .A(y[61]), .B(x[49]), .Z(n6855) );
  XOR U7435 ( .A(n6856), .B(n6855), .Z(n6716) );
  AND U7436 ( .A(x[52]), .B(y[58]), .Z(n6648) );
  NAND U7437 ( .A(x[51]), .B(y[59]), .Z(n6647) );
  XNOR U7438 ( .A(n6648), .B(n6647), .Z(n6715) );
  XOR U7439 ( .A(n6716), .B(n6715), .Z(n6711) );
  XOR U7440 ( .A(n6712), .B(n6711), .Z(n6710) );
  AND U7441 ( .A(y[182]), .B(x[72]), .Z(n6809) );
  XOR U7442 ( .A(n6810), .B(n6809), .Z(n6808) );
  AND U7443 ( .A(y[96]), .B(x[62]), .Z(n6807) );
  XOR U7444 ( .A(n6808), .B(n6807), .Z(n6709) );
  XOR U7445 ( .A(n6710), .B(n6709), .Z(n6686) );
  NAND U7446 ( .A(n6650), .B(n6649), .Z(n6654) );
  NAND U7447 ( .A(n6652), .B(n6651), .Z(n6653) );
  AND U7448 ( .A(n6654), .B(n6653), .Z(n6843) );
  AND U7449 ( .A(y[138]), .B(x[68]), .Z(n6802) );
  AND U7450 ( .A(x[57]), .B(y[101]), .Z(n6656) );
  AND U7451 ( .A(x[58]), .B(y[100]), .Z(n6655) );
  XOR U7452 ( .A(n6656), .B(n6655), .Z(n6801) );
  XOR U7453 ( .A(n6802), .B(n6801), .Z(n6846) );
  AND U7454 ( .A(y[22]), .B(x[40]), .Z(n6850) );
  AND U7455 ( .A(y[142]), .B(x[64]), .Z(n6658) );
  AND U7456 ( .A(x[65]), .B(y[141]), .Z(n6657) );
  XOR U7457 ( .A(n6658), .B(n6657), .Z(n6849) );
  XNOR U7458 ( .A(n6850), .B(n6849), .Z(n6845) );
  XNOR U7459 ( .A(n6843), .B(n6844), .Z(n6685) );
  XOR U7460 ( .A(n6684), .B(n6683), .Z(n6945) );
  NAND U7461 ( .A(n6660), .B(n6659), .Z(n6664) );
  NAND U7462 ( .A(n6662), .B(n6661), .Z(n6663) );
  NAND U7463 ( .A(n6664), .B(n6663), .Z(n6942) );
  XNOR U7464 ( .A(n6943), .B(n6942), .Z(n6938) );
  XOR U7465 ( .A(n6937), .B(n6936), .Z(n6974) );
  XOR U7466 ( .A(n6975), .B(n6974), .Z(n6960) );
  XNOR U7467 ( .A(n6961), .B(n6960), .Z(n6956) );
  NANDN U7468 ( .A(n6666), .B(n6665), .Z(n6670) );
  NAND U7469 ( .A(n6668), .B(n6667), .Z(n6669) );
  NAND U7470 ( .A(n6670), .B(n6669), .Z(n6954) );
  XOR U7471 ( .A(n6955), .B(n6954), .Z(o[62]) );
  NAND U7472 ( .A(n6672), .B(n6671), .Z(n6676) );
  NANDN U7473 ( .A(n6674), .B(n6673), .Z(n6675) );
  AND U7474 ( .A(n6676), .B(n6675), .Z(n6971) );
  NAND U7475 ( .A(n6678), .B(n6677), .Z(n6682) );
  NAND U7476 ( .A(n6680), .B(n6679), .Z(n6681) );
  AND U7477 ( .A(n6682), .B(n6681), .Z(n6953) );
  NAND U7478 ( .A(n6684), .B(n6683), .Z(n6688) );
  NANDN U7479 ( .A(n6686), .B(n6685), .Z(n6687) );
  AND U7480 ( .A(n6688), .B(n6687), .Z(n6935) );
  NANDN U7481 ( .A(n6690), .B(n6689), .Z(n6694) );
  NANDN U7482 ( .A(n6692), .B(n6691), .Z(n6693) );
  AND U7483 ( .A(n6694), .B(n6693), .Z(n6702) );
  NAND U7484 ( .A(n6696), .B(n6695), .Z(n6700) );
  NAND U7485 ( .A(n6698), .B(n6697), .Z(n6699) );
  NAND U7486 ( .A(n6700), .B(n6699), .Z(n6701) );
  XNOR U7487 ( .A(n6702), .B(n6701), .Z(n6933) );
  NAND U7488 ( .A(n6704), .B(n6703), .Z(n6708) );
  NAND U7489 ( .A(n6706), .B(n6705), .Z(n6707) );
  AND U7490 ( .A(n6708), .B(n6707), .Z(n6931) );
  NAND U7491 ( .A(n6710), .B(n6709), .Z(n6714) );
  NAND U7492 ( .A(n6712), .B(n6711), .Z(n6713) );
  AND U7493 ( .A(n6714), .B(n6713), .Z(n6822) );
  NAND U7494 ( .A(n6716), .B(n6715), .Z(n6719) );
  AND U7495 ( .A(y[59]), .B(x[52]), .Z(n6769) );
  NAND U7496 ( .A(n6717), .B(n6769), .Z(n6718) );
  AND U7497 ( .A(n6719), .B(n6718), .Z(n6780) );
  AND U7498 ( .A(x[72]), .B(y[183]), .Z(n6721) );
  NAND U7499 ( .A(x[42]), .B(y[21]), .Z(n6720) );
  XNOR U7500 ( .A(n6721), .B(n6720), .Z(n6725) );
  AND U7501 ( .A(x[73]), .B(y[182]), .Z(n6723) );
  NAND U7502 ( .A(x[70]), .B(y[137]), .Z(n6722) );
  XNOR U7503 ( .A(n6723), .B(n6722), .Z(n6724) );
  XOR U7504 ( .A(n6725), .B(n6724), .Z(n6733) );
  AND U7505 ( .A(x[68]), .B(y[139]), .Z(n6727) );
  NAND U7506 ( .A(x[47]), .B(y[16]), .Z(n6726) );
  XNOR U7507 ( .A(n6727), .B(n6726), .Z(n6731) );
  AND U7508 ( .A(x[63]), .B(y[96]), .Z(n6729) );
  NAND U7509 ( .A(x[54]), .B(y[57]), .Z(n6728) );
  XNOR U7510 ( .A(n6729), .B(n6728), .Z(n6730) );
  XNOR U7511 ( .A(n6731), .B(n6730), .Z(n6732) );
  XNOR U7512 ( .A(n6733), .B(n6732), .Z(n6778) );
  AND U7513 ( .A(x[53]), .B(y[58]), .Z(n6738) );
  AND U7514 ( .A(y[142]), .B(x[65]), .Z(n6851) );
  AND U7515 ( .A(x[64]), .B(y[143]), .Z(n6735) );
  NAND U7516 ( .A(x[49]), .B(y[62]), .Z(n6734) );
  XNOR U7517 ( .A(n6735), .B(n6734), .Z(n6736) );
  XNOR U7518 ( .A(n6851), .B(n6736), .Z(n6737) );
  XNOR U7519 ( .A(n6738), .B(n6737), .Z(n6754) );
  AND U7520 ( .A(x[46]), .B(y[17]), .Z(n6740) );
  NAND U7521 ( .A(x[62]), .B(y[97]), .Z(n6739) );
  XNOR U7522 ( .A(n6740), .B(n6739), .Z(n6744) );
  AND U7523 ( .A(x[79]), .B(y[176]), .Z(n6742) );
  NAND U7524 ( .A(x[78]), .B(y[177]), .Z(n6741) );
  XNOR U7525 ( .A(n6742), .B(n6741), .Z(n6743) );
  XOR U7526 ( .A(n6744), .B(n6743), .Z(n6752) );
  AND U7527 ( .A(x[40]), .B(y[23]), .Z(n6746) );
  NAND U7528 ( .A(x[55]), .B(y[56]), .Z(n6745) );
  XNOR U7529 ( .A(n6746), .B(n6745), .Z(n6750) );
  AND U7530 ( .A(x[50]), .B(y[61]), .Z(n6748) );
  NAND U7531 ( .A(x[66]), .B(y[141]), .Z(n6747) );
  XNOR U7532 ( .A(n6748), .B(n6747), .Z(n6749) );
  XNOR U7533 ( .A(n6750), .B(n6749), .Z(n6751) );
  XNOR U7534 ( .A(n6752), .B(n6751), .Z(n6753) );
  XOR U7535 ( .A(n6754), .B(n6753), .Z(n6776) );
  AND U7536 ( .A(x[48]), .B(y[63]), .Z(n6756) );
  NAND U7537 ( .A(x[41]), .B(y[22]), .Z(n6755) );
  XNOR U7538 ( .A(n6756), .B(n6755), .Z(n6760) );
  AND U7539 ( .A(x[59]), .B(y[100]), .Z(n6758) );
  NAND U7540 ( .A(x[60]), .B(y[99]), .Z(n6757) );
  XNOR U7541 ( .A(n6758), .B(n6757), .Z(n6759) );
  XOR U7542 ( .A(n6760), .B(n6759), .Z(n6768) );
  AND U7543 ( .A(x[67]), .B(y[140]), .Z(n6762) );
  NAND U7544 ( .A(x[43]), .B(y[20]), .Z(n6761) );
  XNOR U7545 ( .A(n6762), .B(n6761), .Z(n6766) );
  AND U7546 ( .A(x[56]), .B(y[103]), .Z(n6764) );
  NAND U7547 ( .A(x[71]), .B(y[136]), .Z(n6763) );
  XNOR U7548 ( .A(n6764), .B(n6763), .Z(n6765) );
  XNOR U7549 ( .A(n6766), .B(n6765), .Z(n6767) );
  XNOR U7550 ( .A(n6768), .B(n6767), .Z(n6774) );
  AND U7551 ( .A(y[101]), .B(x[58]), .Z(n6803) );
  XOR U7552 ( .A(n6769), .B(n6803), .Z(n6772) );
  AND U7553 ( .A(y[178]), .B(x[77]), .Z(n6865) );
  XNOR U7554 ( .A(n6770), .B(n6865), .Z(n6771) );
  XNOR U7555 ( .A(n6772), .B(n6771), .Z(n6773) );
  XNOR U7556 ( .A(n6774), .B(n6773), .Z(n6775) );
  XNOR U7557 ( .A(n6776), .B(n6775), .Z(n6777) );
  XNOR U7558 ( .A(n6778), .B(n6777), .Z(n6779) );
  XNOR U7559 ( .A(n6780), .B(n6779), .Z(n6820) );
  NAND U7560 ( .A(n6782), .B(n6781), .Z(n6786) );
  NANDN U7561 ( .A(n6784), .B(n6783), .Z(n6785) );
  AND U7562 ( .A(n6786), .B(n6785), .Z(n6818) );
  NAND U7563 ( .A(n6788), .B(n6787), .Z(n6792) );
  AND U7564 ( .A(n6790), .B(n6789), .Z(n6791) );
  ANDN U7565 ( .B(n6792), .A(n6791), .Z(n6800) );
  AND U7566 ( .A(n6794), .B(n6793), .Z(n6798) );
  AND U7567 ( .A(n6796), .B(n6795), .Z(n6797) );
  OR U7568 ( .A(n6798), .B(n6797), .Z(n6799) );
  XNOR U7569 ( .A(n6800), .B(n6799), .Z(n6816) );
  NAND U7570 ( .A(n6802), .B(n6801), .Z(n6806) );
  NAND U7571 ( .A(n6804), .B(n6803), .Z(n6805) );
  AND U7572 ( .A(n6806), .B(n6805), .Z(n6814) );
  NAND U7573 ( .A(n6808), .B(n6807), .Z(n6812) );
  NAND U7574 ( .A(n6810), .B(n6809), .Z(n6811) );
  NAND U7575 ( .A(n6812), .B(n6811), .Z(n6813) );
  XNOR U7576 ( .A(n6814), .B(n6813), .Z(n6815) );
  XNOR U7577 ( .A(n6816), .B(n6815), .Z(n6817) );
  XNOR U7578 ( .A(n6818), .B(n6817), .Z(n6819) );
  XNOR U7579 ( .A(n6820), .B(n6819), .Z(n6821) );
  XNOR U7580 ( .A(n6822), .B(n6821), .Z(n6929) );
  NANDN U7581 ( .A(n6824), .B(n6823), .Z(n6828) );
  NAND U7582 ( .A(n6826), .B(n6825), .Z(n6827) );
  AND U7583 ( .A(n6828), .B(n6827), .Z(n6927) );
  NAND U7584 ( .A(n6830), .B(n6829), .Z(n6834) );
  ANDN U7585 ( .B(n6832), .A(n6831), .Z(n6833) );
  ANDN U7586 ( .B(n6834), .A(n6833), .Z(n6842) );
  ANDN U7587 ( .B(n6836), .A(n6835), .Z(n6840) );
  ANDN U7588 ( .B(n6838), .A(n6837), .Z(n6839) );
  OR U7589 ( .A(n6840), .B(n6839), .Z(n6841) );
  XNOR U7590 ( .A(n6842), .B(n6841), .Z(n6925) );
  NANDN U7591 ( .A(n6844), .B(n6843), .Z(n6848) );
  NANDN U7592 ( .A(n6846), .B(n6845), .Z(n6847) );
  AND U7593 ( .A(n6848), .B(n6847), .Z(n6923) );
  NAND U7594 ( .A(n6850), .B(n6849), .Z(n6854) );
  NAND U7595 ( .A(n6852), .B(n6851), .Z(n6853) );
  AND U7596 ( .A(n6854), .B(n6853), .Z(n6862) );
  NAND U7597 ( .A(n6856), .B(n6855), .Z(n6860) );
  NAND U7598 ( .A(n6858), .B(n6857), .Z(n6859) );
  NAND U7599 ( .A(n6860), .B(n6859), .Z(n6861) );
  XNOR U7600 ( .A(n6862), .B(n6861), .Z(n6921) );
  AND U7601 ( .A(x[69]), .B(y[138]), .Z(n6864) );
  NAND U7602 ( .A(x[61]), .B(y[98]), .Z(n6863) );
  XNOR U7603 ( .A(n6864), .B(n6863), .Z(n6887) );
  AND U7604 ( .A(n6866), .B(n6865), .Z(n6881) );
  NAND U7605 ( .A(n6868), .B(n6867), .Z(n6871) );
  AND U7606 ( .A(y[18]), .B(x[45]), .Z(n6883) );
  NAND U7607 ( .A(n6869), .B(n6883), .Z(n6870) );
  AND U7608 ( .A(n6871), .B(n6870), .Z(n6879) );
  AND U7609 ( .A(x[57]), .B(y[102]), .Z(n6873) );
  NAND U7610 ( .A(x[74]), .B(y[181]), .Z(n6872) );
  XNOR U7611 ( .A(n6873), .B(n6872), .Z(n6877) );
  AND U7612 ( .A(x[75]), .B(y[180]), .Z(n6875) );
  NAND U7613 ( .A(x[44]), .B(y[19]), .Z(n6874) );
  XNOR U7614 ( .A(n6875), .B(n6874), .Z(n6876) );
  XNOR U7615 ( .A(n6877), .B(n6876), .Z(n6878) );
  XNOR U7616 ( .A(n6879), .B(n6878), .Z(n6880) );
  XOR U7617 ( .A(n6881), .B(n6880), .Z(n6885) );
  XNOR U7618 ( .A(n6883), .B(n6882), .Z(n6884) );
  XNOR U7619 ( .A(n6885), .B(n6884), .Z(n6886) );
  XOR U7620 ( .A(n6887), .B(n6886), .Z(n6919) );
  NAND U7621 ( .A(n6889), .B(n6888), .Z(n6893) );
  NAND U7622 ( .A(n6891), .B(n6890), .Z(n6892) );
  AND U7623 ( .A(n6893), .B(n6892), .Z(n6901) );
  NAND U7624 ( .A(n6895), .B(n6894), .Z(n6899) );
  NAND U7625 ( .A(n6897), .B(n6896), .Z(n6898) );
  NAND U7626 ( .A(n6899), .B(n6898), .Z(n6900) );
  XNOR U7627 ( .A(n6901), .B(n6900), .Z(n6917) );
  NAND U7628 ( .A(n6903), .B(n6902), .Z(n6907) );
  NAND U7629 ( .A(n6905), .B(n6904), .Z(n6906) );
  AND U7630 ( .A(n6907), .B(n6906), .Z(n6915) );
  NAND U7631 ( .A(n6909), .B(n6908), .Z(n6913) );
  NAND U7632 ( .A(n6911), .B(n6910), .Z(n6912) );
  NAND U7633 ( .A(n6913), .B(n6912), .Z(n6914) );
  XNOR U7634 ( .A(n6915), .B(n6914), .Z(n6916) );
  XNOR U7635 ( .A(n6917), .B(n6916), .Z(n6918) );
  XNOR U7636 ( .A(n6919), .B(n6918), .Z(n6920) );
  XNOR U7637 ( .A(n6921), .B(n6920), .Z(n6922) );
  XNOR U7638 ( .A(n6923), .B(n6922), .Z(n6924) );
  XNOR U7639 ( .A(n6925), .B(n6924), .Z(n6926) );
  XNOR U7640 ( .A(n6927), .B(n6926), .Z(n6928) );
  XNOR U7641 ( .A(n6929), .B(n6928), .Z(n6930) );
  XNOR U7642 ( .A(n6931), .B(n6930), .Z(n6932) );
  XNOR U7643 ( .A(n6933), .B(n6932), .Z(n6934) );
  XNOR U7644 ( .A(n6935), .B(n6934), .Z(n6951) );
  NAND U7645 ( .A(n6937), .B(n6936), .Z(n6941) );
  NANDN U7646 ( .A(n6939), .B(n6938), .Z(n6940) );
  AND U7647 ( .A(n6941), .B(n6940), .Z(n6949) );
  NAND U7648 ( .A(n6943), .B(n6942), .Z(n6947) );
  NANDN U7649 ( .A(n6945), .B(n6944), .Z(n6946) );
  NAND U7650 ( .A(n6947), .B(n6946), .Z(n6948) );
  XNOR U7651 ( .A(n6949), .B(n6948), .Z(n6950) );
  XNOR U7652 ( .A(n6951), .B(n6950), .Z(n6952) );
  XNOR U7653 ( .A(n6953), .B(n6952), .Z(n6969) );
  NAND U7654 ( .A(n6955), .B(n6954), .Z(n6959) );
  NANDN U7655 ( .A(n6957), .B(n6956), .Z(n6958) );
  AND U7656 ( .A(n6959), .B(n6958), .Z(n6967) );
  NAND U7657 ( .A(n6961), .B(n6960), .Z(n6965) );
  NANDN U7658 ( .A(n6963), .B(n6962), .Z(n6964) );
  NAND U7659 ( .A(n6965), .B(n6964), .Z(n6966) );
  XNOR U7660 ( .A(n6967), .B(n6966), .Z(n6968) );
  XNOR U7661 ( .A(n6969), .B(n6968), .Z(n6970) );
  XNOR U7662 ( .A(n6971), .B(n6970), .Z(n6979) );
  AND U7663 ( .A(n6973), .B(n6972), .Z(n6977) );
  AND U7664 ( .A(n6975), .B(n6974), .Z(n6976) );
  NOR U7665 ( .A(n6977), .B(n6976), .Z(n6978) );
  XNOR U7666 ( .A(n6979), .B(n6978), .Z(o[63]) );
  NAND U7667 ( .A(y[184]), .B(x[72]), .Z(n7093) );
  NAND U7668 ( .A(y[64]), .B(x[48]), .Z(n6982) );
  XOR U7669 ( .A(n7093), .B(n6982), .Z(n6983) );
  AND U7670 ( .A(y[24]), .B(x[40]), .Z(n6990) );
  AND U7671 ( .A(y[104]), .B(x[56]), .Z(n6987) );
  XOR U7672 ( .A(n6990), .B(n6987), .Z(n6986) );
  AND U7673 ( .A(y[144]), .B(x[64]), .Z(n6985) );
  XNOR U7674 ( .A(n6986), .B(n6985), .Z(n6984) );
  XNOR U7675 ( .A(n6983), .B(n6984), .Z(o[64]) );
  AND U7676 ( .A(x[41]), .B(y[24]), .Z(n6981) );
  NAND U7677 ( .A(x[40]), .B(y[25]), .Z(n6980) );
  XNOR U7678 ( .A(n6981), .B(n6980), .Z(n6992) );
  AND U7679 ( .A(y[64]), .B(x[49]), .Z(n6991) );
  XOR U7680 ( .A(n6992), .B(n6991), .Z(n7009) );
  AND U7681 ( .A(y[184]), .B(x[73]), .Z(n7211) );
  AND U7682 ( .A(y[105]), .B(x[56]), .Z(n6995) );
  XOR U7683 ( .A(n7211), .B(n6995), .Z(n6997) );
  AND U7684 ( .A(y[185]), .B(x[72]), .Z(n7019) );
  NAND U7685 ( .A(y[104]), .B(x[57]), .Z(n7018) );
  XNOR U7686 ( .A(n7019), .B(n7018), .Z(n6996) );
  XOR U7687 ( .A(n6997), .B(n6996), .Z(n7007) );
  AND U7688 ( .A(y[65]), .B(x[48]), .Z(n7230) );
  AND U7689 ( .A(y[145]), .B(x[64]), .Z(n7012) );
  XOR U7690 ( .A(n7230), .B(n7012), .Z(n7014) );
  AND U7691 ( .A(y[144]), .B(x[65]), .Z(n7013) );
  XNOR U7692 ( .A(n7014), .B(n7013), .Z(n7006) );
  XNOR U7693 ( .A(n7007), .B(n7006), .Z(n7008) );
  XNOR U7694 ( .A(n7009), .B(n7008), .Z(n7003) );
  NAND U7695 ( .A(n6986), .B(n6985), .Z(n6989) );
  AND U7696 ( .A(n6990), .B(n6987), .Z(n6988) );
  ANDN U7697 ( .B(n6989), .A(n6988), .Z(n7000) );
  XNOR U7698 ( .A(n7001), .B(n7000), .Z(n7002) );
  XNOR U7699 ( .A(n7003), .B(n7002), .Z(o[65]) );
  NAND U7700 ( .A(y[25]), .B(x[41]), .Z(n7041) );
  NANDN U7701 ( .A(n7041), .B(n6990), .Z(n6994) );
  NAND U7702 ( .A(n6992), .B(n6991), .Z(n6993) );
  AND U7703 ( .A(n6994), .B(n6993), .Z(n7061) );
  NAND U7704 ( .A(n7211), .B(n6995), .Z(n6999) );
  NAND U7705 ( .A(n6997), .B(n6996), .Z(n6998) );
  AND U7706 ( .A(n6999), .B(n6998), .Z(n7060) );
  AND U7707 ( .A(y[146]), .B(x[64]), .Z(n7065) );
  NAND U7708 ( .A(y[26]), .B(x[40]), .Z(n7066) );
  XNOR U7709 ( .A(n7065), .B(n7066), .Z(n7067) );
  NAND U7710 ( .A(y[64]), .B(x[50]), .Z(n7068) );
  XNOR U7711 ( .A(n7067), .B(n7068), .Z(n7059) );
  XOR U7712 ( .A(n7060), .B(n7059), .Z(n7062) );
  XOR U7713 ( .A(n7061), .B(n7062), .Z(n7021) );
  NANDN U7714 ( .A(n7001), .B(n7000), .Z(n7005) );
  NAND U7715 ( .A(n7003), .B(n7002), .Z(n7004) );
  NAND U7716 ( .A(n7005), .B(n7004), .Z(n7020) );
  XNOR U7717 ( .A(n7021), .B(n7020), .Z(n7023) );
  NANDN U7718 ( .A(n7007), .B(n7006), .Z(n7011) );
  NANDN U7719 ( .A(n7009), .B(n7008), .Z(n7010) );
  AND U7720 ( .A(n7011), .B(n7010), .Z(n7029) );
  AND U7721 ( .A(y[24]), .B(x[42]), .Z(n7038) );
  NAND U7722 ( .A(y[106]), .B(x[56]), .Z(n7039) );
  XNOR U7723 ( .A(n7038), .B(n7039), .Z(n7040) );
  AND U7724 ( .A(y[144]), .B(x[66]), .Z(n7073) );
  XOR U7725 ( .A(n7074), .B(n7073), .Z(n7076) );
  AND U7726 ( .A(y[104]), .B(x[58]), .Z(n7121) );
  AND U7727 ( .A(y[186]), .B(x[72]), .Z(n7051) );
  XOR U7728 ( .A(n7121), .B(n7051), .Z(n7053) );
  AND U7729 ( .A(y[105]), .B(x[57]), .Z(n7052) );
  XOR U7730 ( .A(n7053), .B(n7052), .Z(n7075) );
  XOR U7731 ( .A(n7076), .B(n7075), .Z(n7026) );
  NAND U7732 ( .A(n7230), .B(n7012), .Z(n7016) );
  AND U7733 ( .A(n7014), .B(n7013), .Z(n7015) );
  ANDN U7734 ( .B(n7016), .A(n7015), .Z(n7035) );
  AND U7735 ( .A(x[73]), .B(y[185]), .Z(n7098) );
  NAND U7736 ( .A(x[74]), .B(y[184]), .Z(n7017) );
  XNOR U7737 ( .A(n7098), .B(n7017), .Z(n7072) );
  ANDN U7738 ( .B(n7019), .A(n7018), .Z(n7071) );
  XOR U7739 ( .A(n7072), .B(n7071), .Z(n7032) );
  AND U7740 ( .A(y[145]), .B(x[65]), .Z(n7044) );
  NAND U7741 ( .A(y[65]), .B(x[49]), .Z(n7045) );
  XNOR U7742 ( .A(n7044), .B(n7045), .Z(n7046) );
  NAND U7743 ( .A(y[66]), .B(x[48]), .Z(n7047) );
  XOR U7744 ( .A(n7046), .B(n7047), .Z(n7033) );
  XNOR U7745 ( .A(n7032), .B(n7033), .Z(n7034) );
  XOR U7746 ( .A(n7035), .B(n7034), .Z(n7027) );
  XNOR U7747 ( .A(n7026), .B(n7027), .Z(n7028) );
  XNOR U7748 ( .A(n7029), .B(n7028), .Z(n7022) );
  XNOR U7749 ( .A(n7023), .B(n7022), .Z(o[66]) );
  NANDN U7750 ( .A(n7021), .B(n7020), .Z(n7025) );
  NAND U7751 ( .A(n7023), .B(n7022), .Z(n7024) );
  AND U7752 ( .A(n7025), .B(n7024), .Z(n7159) );
  NANDN U7753 ( .A(n7027), .B(n7026), .Z(n7031) );
  NAND U7754 ( .A(n7029), .B(n7028), .Z(n7030) );
  AND U7755 ( .A(n7031), .B(n7030), .Z(n7144) );
  NANDN U7756 ( .A(n7033), .B(n7032), .Z(n7037) );
  NANDN U7757 ( .A(n7035), .B(n7034), .Z(n7036) );
  AND U7758 ( .A(n7037), .B(n7036), .Z(n7142) );
  NANDN U7759 ( .A(n7039), .B(n7038), .Z(n7043) );
  NANDN U7760 ( .A(n7041), .B(n7040), .Z(n7042) );
  NAND U7761 ( .A(n7043), .B(n7042), .Z(n7153) );
  NANDN U7762 ( .A(n7045), .B(n7044), .Z(n7049) );
  NANDN U7763 ( .A(n7047), .B(n7046), .Z(n7048) );
  AND U7764 ( .A(n7049), .B(n7048), .Z(n7112) );
  AND U7765 ( .A(y[147]), .B(x[64]), .Z(n7137) );
  AND U7766 ( .A(y[107]), .B(x[56]), .Z(n7136) );
  NAND U7767 ( .A(y[24]), .B(x[43]), .Z(n7135) );
  XOR U7768 ( .A(n7136), .B(n7135), .Z(n7138) );
  XOR U7769 ( .A(n7137), .B(n7138), .Z(n7110) );
  AND U7770 ( .A(x[58]), .B(y[105]), .Z(n7191) );
  NAND U7771 ( .A(x[59]), .B(y[104]), .Z(n7050) );
  XNOR U7772 ( .A(n7191), .B(n7050), .Z(n7123) );
  AND U7773 ( .A(y[106]), .B(x[57]), .Z(n7122) );
  XOR U7774 ( .A(n7123), .B(n7122), .Z(n7109) );
  XNOR U7775 ( .A(n7110), .B(n7109), .Z(n7111) );
  XNOR U7776 ( .A(n7112), .B(n7111), .Z(n7154) );
  XOR U7777 ( .A(n7153), .B(n7154), .Z(n7156) );
  NAND U7778 ( .A(n7121), .B(n7051), .Z(n7055) );
  AND U7779 ( .A(n7053), .B(n7052), .Z(n7054) );
  ANDN U7780 ( .B(n7055), .A(n7054), .Z(n7117) );
  AND U7781 ( .A(y[26]), .B(x[41]), .Z(n7089) );
  AND U7782 ( .A(y[25]), .B(x[42]), .Z(n7088) );
  NAND U7783 ( .A(y[146]), .B(x[65]), .Z(n7087) );
  XOR U7784 ( .A(n7088), .B(n7087), .Z(n7090) );
  XOR U7785 ( .A(n7089), .B(n7090), .Z(n7116) );
  AND U7786 ( .A(x[75]), .B(y[184]), .Z(n7057) );
  NAND U7787 ( .A(x[72]), .B(y[187]), .Z(n7056) );
  XNOR U7788 ( .A(n7057), .B(n7056), .Z(n7094) );
  AND U7789 ( .A(x[74]), .B(y[185]), .Z(n7208) );
  NAND U7790 ( .A(x[73]), .B(y[186]), .Z(n7058) );
  XOR U7791 ( .A(n7208), .B(n7058), .Z(n7095) );
  XNOR U7792 ( .A(n7094), .B(n7095), .Z(n7115) );
  XOR U7793 ( .A(n7116), .B(n7115), .Z(n7118) );
  XOR U7794 ( .A(n7117), .B(n7118), .Z(n7155) );
  XOR U7795 ( .A(n7156), .B(n7155), .Z(n7141) );
  XNOR U7796 ( .A(n7142), .B(n7141), .Z(n7143) );
  XOR U7797 ( .A(n7144), .B(n7143), .Z(n7160) );
  XNOR U7798 ( .A(n7159), .B(n7160), .Z(n7162) );
  NANDN U7799 ( .A(n7060), .B(n7059), .Z(n7064) );
  OR U7800 ( .A(n7062), .B(n7061), .Z(n7063) );
  AND U7801 ( .A(n7064), .B(n7063), .Z(n7150) );
  NANDN U7802 ( .A(n7066), .B(n7065), .Z(n7070) );
  NANDN U7803 ( .A(n7068), .B(n7067), .Z(n7069) );
  AND U7804 ( .A(n7070), .B(n7069), .Z(n7080) );
  XNOR U7805 ( .A(n7080), .B(n7079), .Z(n7082) );
  AND U7806 ( .A(y[64]), .B(x[51]), .Z(n7129) );
  AND U7807 ( .A(y[27]), .B(x[40]), .Z(n7127) );
  NAND U7808 ( .A(y[145]), .B(x[66]), .Z(n7126) );
  XNOR U7809 ( .A(n7127), .B(n7126), .Z(n7128) );
  XOR U7810 ( .A(n7129), .B(n7128), .Z(n7107) );
  AND U7811 ( .A(y[67]), .B(x[48]), .Z(n7102) );
  AND U7812 ( .A(y[65]), .B(x[50]), .Z(n7100) );
  NAND U7813 ( .A(y[144]), .B(x[67]), .Z(n7099) );
  XNOR U7814 ( .A(n7100), .B(n7099), .Z(n7101) );
  XOR U7815 ( .A(n7102), .B(n7101), .Z(n7105) );
  AND U7816 ( .A(y[66]), .B(x[49]), .Z(n7106) );
  XOR U7817 ( .A(n7105), .B(n7106), .Z(n7108) );
  XOR U7818 ( .A(n7107), .B(n7108), .Z(n7081) );
  XOR U7819 ( .A(n7082), .B(n7081), .Z(n7148) );
  NAND U7820 ( .A(n7074), .B(n7073), .Z(n7078) );
  NAND U7821 ( .A(n7076), .B(n7075), .Z(n7077) );
  AND U7822 ( .A(n7078), .B(n7077), .Z(n7147) );
  XNOR U7823 ( .A(n7148), .B(n7147), .Z(n7149) );
  XNOR U7824 ( .A(n7150), .B(n7149), .Z(n7161) );
  XOR U7825 ( .A(n7162), .B(n7161), .Z(o[67]) );
  NANDN U7826 ( .A(n7080), .B(n7079), .Z(n7084) );
  NAND U7827 ( .A(n7082), .B(n7081), .Z(n7083) );
  AND U7828 ( .A(n7084), .B(n7083), .Z(n7176) );
  AND U7829 ( .A(y[66]), .B(x[50]), .Z(n7285) );
  AND U7830 ( .A(x[48]), .B(y[68]), .Z(n7086) );
  NAND U7831 ( .A(x[51]), .B(y[65]), .Z(n7085) );
  XOR U7832 ( .A(n7086), .B(n7085), .Z(n7231) );
  XNOR U7833 ( .A(n7285), .B(n7231), .Z(n7241) );
  AND U7834 ( .A(y[67]), .B(x[49]), .Z(n7240) );
  XOR U7835 ( .A(n7241), .B(n7240), .Z(n7243) );
  AND U7836 ( .A(y[144]), .B(x[68]), .Z(n7196) );
  NAND U7837 ( .A(y[27]), .B(x[41]), .Z(n7197) );
  XNOR U7838 ( .A(n7196), .B(n7197), .Z(n7198) );
  NAND U7839 ( .A(y[28]), .B(x[40]), .Z(n7199) );
  XNOR U7840 ( .A(n7198), .B(n7199), .Z(n7242) );
  XOR U7841 ( .A(n7243), .B(n7242), .Z(n7237) );
  NANDN U7842 ( .A(n7088), .B(n7087), .Z(n7092) );
  OR U7843 ( .A(n7090), .B(n7089), .Z(n7091) );
  AND U7844 ( .A(n7092), .B(n7091), .Z(n7235) );
  AND U7845 ( .A(y[187]), .B(x[75]), .Z(n7533) );
  NANDN U7846 ( .A(n7093), .B(n7533), .Z(n7097) );
  NANDN U7847 ( .A(n7095), .B(n7094), .Z(n7096) );
  AND U7848 ( .A(n7097), .B(n7096), .Z(n7234) );
  XNOR U7849 ( .A(n7235), .B(n7234), .Z(n7236) );
  XNOR U7850 ( .A(n7237), .B(n7236), .Z(n7261) );
  NAND U7851 ( .A(y[24]), .B(x[44]), .Z(n7220) );
  NAND U7852 ( .A(y[146]), .B(x[66]), .Z(n7218) );
  NAND U7853 ( .A(y[108]), .B(x[56]), .Z(n7219) );
  XNOR U7854 ( .A(n7218), .B(n7219), .Z(n7221) );
  XOR U7855 ( .A(n7220), .B(n7221), .Z(n7181) );
  AND U7856 ( .A(y[186]), .B(x[74]), .Z(n7134) );
  NAND U7857 ( .A(n7098), .B(n7134), .Z(n7214) );
  NAND U7858 ( .A(y[188]), .B(x[72]), .Z(n7341) );
  NAND U7859 ( .A(y[104]), .B(x[60]), .Z(n7297) );
  XNOR U7860 ( .A(n7341), .B(n7297), .Z(n7215) );
  XOR U7861 ( .A(n7214), .B(n7215), .Z(n7182) );
  XOR U7862 ( .A(n7181), .B(n7182), .Z(n7183) );
  NANDN U7863 ( .A(n7100), .B(n7099), .Z(n7104) );
  NANDN U7864 ( .A(n7102), .B(n7101), .Z(n7103) );
  NAND U7865 ( .A(n7104), .B(n7103), .Z(n7184) );
  XOR U7866 ( .A(n7183), .B(n7184), .Z(n7258) );
  XOR U7867 ( .A(n7258), .B(n7259), .Z(n7260) );
  XNOR U7868 ( .A(n7261), .B(n7260), .Z(n7175) );
  XNOR U7869 ( .A(n7176), .B(n7175), .Z(n7178) );
  NANDN U7870 ( .A(n7110), .B(n7109), .Z(n7114) );
  NANDN U7871 ( .A(n7112), .B(n7111), .Z(n7113) );
  NAND U7872 ( .A(n7114), .B(n7113), .Z(n7250) );
  NANDN U7873 ( .A(n7116), .B(n7115), .Z(n7120) );
  OR U7874 ( .A(n7118), .B(n7117), .Z(n7119) );
  NAND U7875 ( .A(n7120), .B(n7119), .Z(n7251) );
  XOR U7876 ( .A(n7250), .B(n7251), .Z(n7253) );
  AND U7877 ( .A(y[64]), .B(x[52]), .Z(n7202) );
  NAND U7878 ( .A(y[148]), .B(x[64]), .Z(n7203) );
  XNOR U7879 ( .A(n7202), .B(n7203), .Z(n7204) );
  NAND U7880 ( .A(y[147]), .B(x[65]), .Z(n7205) );
  XNOR U7881 ( .A(n7204), .B(n7205), .Z(n7244) );
  AND U7882 ( .A(x[58]), .B(y[106]), .Z(n7125) );
  NAND U7883 ( .A(x[59]), .B(y[105]), .Z(n7124) );
  XNOR U7884 ( .A(n7125), .B(n7124), .Z(n7192) );
  NAND U7885 ( .A(y[107]), .B(x[57]), .Z(n7193) );
  XOR U7886 ( .A(n7192), .B(n7193), .Z(n7245) );
  XNOR U7887 ( .A(n7244), .B(n7245), .Z(n7246) );
  NANDN U7888 ( .A(n7127), .B(n7126), .Z(n7131) );
  NANDN U7889 ( .A(n7129), .B(n7128), .Z(n7130) );
  NAND U7890 ( .A(n7131), .B(n7130), .Z(n7247) );
  XNOR U7891 ( .A(n7246), .B(n7247), .Z(n7255) );
  XOR U7892 ( .A(n7254), .B(n7255), .Z(n7257) );
  NAND U7893 ( .A(y[26]), .B(x[42]), .Z(n7226) );
  NAND U7894 ( .A(y[145]), .B(x[67]), .Z(n7225) );
  NAND U7895 ( .A(y[25]), .B(x[43]), .Z(n7224) );
  XNOR U7896 ( .A(n7225), .B(n7224), .Z(n7227) );
  AND U7897 ( .A(x[76]), .B(y[184]), .Z(n7133) );
  NAND U7898 ( .A(x[73]), .B(y[187]), .Z(n7132) );
  XNOR U7899 ( .A(n7133), .B(n7132), .Z(n7213) );
  AND U7900 ( .A(y[185]), .B(x[75]), .Z(n7303) );
  XOR U7901 ( .A(n7303), .B(n7134), .Z(n7212) );
  XOR U7902 ( .A(n7213), .B(n7212), .Z(n7185) );
  XOR U7903 ( .A(n7186), .B(n7185), .Z(n7187) );
  NANDN U7904 ( .A(n7136), .B(n7135), .Z(n7140) );
  OR U7905 ( .A(n7138), .B(n7137), .Z(n7139) );
  NAND U7906 ( .A(n7140), .B(n7139), .Z(n7188) );
  XNOR U7907 ( .A(n7187), .B(n7188), .Z(n7256) );
  XOR U7908 ( .A(n7257), .B(n7256), .Z(n7252) );
  XOR U7909 ( .A(n7253), .B(n7252), .Z(n7177) );
  XNOR U7910 ( .A(n7178), .B(n7177), .Z(n7168) );
  NANDN U7911 ( .A(n7142), .B(n7141), .Z(n7146) );
  NANDN U7912 ( .A(n7144), .B(n7143), .Z(n7145) );
  AND U7913 ( .A(n7146), .B(n7145), .Z(n7171) );
  NANDN U7914 ( .A(n7148), .B(n7147), .Z(n7152) );
  NAND U7915 ( .A(n7150), .B(n7149), .Z(n7151) );
  NAND U7916 ( .A(n7152), .B(n7151), .Z(n7169) );
  NAND U7917 ( .A(n7154), .B(n7153), .Z(n7158) );
  NAND U7918 ( .A(n7156), .B(n7155), .Z(n7157) );
  AND U7919 ( .A(n7158), .B(n7157), .Z(n7170) );
  XNOR U7920 ( .A(n7169), .B(n7170), .Z(n7172) );
  NANDN U7921 ( .A(n7160), .B(n7159), .Z(n7164) );
  NAND U7922 ( .A(n7162), .B(n7161), .Z(n7163) );
  NAND U7923 ( .A(n7164), .B(n7163), .Z(n7166) );
  XNOR U7924 ( .A(n7167), .B(n7166), .Z(n7165) );
  XNOR U7925 ( .A(n7168), .B(n7165), .Z(o[68]) );
  NAND U7926 ( .A(n7170), .B(n7169), .Z(n7174) );
  NANDN U7927 ( .A(n7172), .B(n7171), .Z(n7173) );
  AND U7928 ( .A(n7174), .B(n7173), .Z(n7379) );
  XNOR U7929 ( .A(n7380), .B(n7379), .Z(n7382) );
  NANDN U7930 ( .A(n7176), .B(n7175), .Z(n7180) );
  NAND U7931 ( .A(n7178), .B(n7177), .Z(n7179) );
  AND U7932 ( .A(n7180), .B(n7179), .Z(n7376) );
  NAND U7933 ( .A(n7186), .B(n7185), .Z(n7190) );
  NANDN U7934 ( .A(n7188), .B(n7187), .Z(n7189) );
  NAND U7935 ( .A(n7190), .B(n7189), .Z(n7312) );
  XOR U7936 ( .A(n7311), .B(n7312), .Z(n7314) );
  AND U7937 ( .A(y[106]), .B(x[59]), .Z(n7299) );
  NAND U7938 ( .A(n7191), .B(n7299), .Z(n7195) );
  NANDN U7939 ( .A(n7193), .B(n7192), .Z(n7194) );
  NAND U7940 ( .A(n7195), .B(n7194), .Z(n7270) );
  NANDN U7941 ( .A(n7197), .B(n7196), .Z(n7201) );
  NANDN U7942 ( .A(n7199), .B(n7198), .Z(n7200) );
  NAND U7943 ( .A(n7201), .B(n7200), .Z(n7278) );
  AND U7944 ( .A(y[64]), .B(x[53]), .Z(n7308) );
  AND U7945 ( .A(y[107]), .B(x[58]), .Z(n7307) );
  XOR U7946 ( .A(n7308), .B(n7307), .Z(n7310) );
  AND U7947 ( .A(y[149]), .B(x[64]), .Z(n7309) );
  XOR U7948 ( .A(n7310), .B(n7309), .Z(n7277) );
  AND U7949 ( .A(y[145]), .B(x[68]), .Z(n7305) );
  AND U7950 ( .A(y[24]), .B(x[45]), .Z(n7304) );
  XOR U7951 ( .A(n7305), .B(n7304), .Z(n7306) );
  AND U7952 ( .A(y[25]), .B(x[44]), .Z(n7538) );
  XOR U7953 ( .A(n7306), .B(n7538), .Z(n7276) );
  XOR U7954 ( .A(n7277), .B(n7276), .Z(n7279) );
  XOR U7955 ( .A(n7278), .B(n7279), .Z(n7271) );
  XOR U7956 ( .A(n7270), .B(n7271), .Z(n7273) );
  NANDN U7957 ( .A(n7203), .B(n7202), .Z(n7207) );
  NANDN U7958 ( .A(n7205), .B(n7204), .Z(n7206) );
  NAND U7959 ( .A(n7207), .B(n7206), .Z(n7373) );
  AND U7960 ( .A(y[186]), .B(x[75]), .Z(n7216) );
  AND U7961 ( .A(n7208), .B(n7216), .Z(n7343) );
  AND U7962 ( .A(x[72]), .B(y[189]), .Z(n7210) );
  AND U7963 ( .A(x[73]), .B(y[188]), .Z(n7209) );
  XOR U7964 ( .A(n7210), .B(n7209), .Z(n7342) );
  XOR U7965 ( .A(n7343), .B(n7342), .Z(n7372) );
  AND U7966 ( .A(y[65]), .B(x[52]), .Z(n7366) );
  AND U7967 ( .A(y[69]), .B(x[48]), .Z(n7364) );
  AND U7968 ( .A(y[28]), .B(x[41]), .Z(n7363) );
  XOR U7969 ( .A(n7364), .B(n7363), .Z(n7365) );
  XOR U7970 ( .A(n7366), .B(n7365), .Z(n7371) );
  XOR U7971 ( .A(n7372), .B(n7371), .Z(n7374) );
  XOR U7972 ( .A(n7373), .B(n7374), .Z(n7272) );
  XOR U7973 ( .A(n7273), .B(n7272), .Z(n7313) );
  XOR U7974 ( .A(n7314), .B(n7313), .Z(n7264) );
  AND U7975 ( .A(y[187]), .B(x[76]), .Z(n7417) );
  XOR U7976 ( .A(n7327), .B(n7328), .Z(n7330) );
  AND U7977 ( .A(y[187]), .B(x[74]), .Z(n7281) );
  AND U7978 ( .A(y[184]), .B(x[77]), .Z(n7280) );
  XOR U7979 ( .A(n7281), .B(n7280), .Z(n7283) );
  AND U7980 ( .A(y[185]), .B(x[76]), .Z(n7412) );
  XOR U7981 ( .A(n7412), .B(n7216), .Z(n7282) );
  XOR U7982 ( .A(n7283), .B(n7282), .Z(n7316) );
  AND U7983 ( .A(y[66]), .B(x[51]), .Z(n7518) );
  NAND U7984 ( .A(x[50]), .B(y[67]), .Z(n7217) );
  XNOR U7985 ( .A(n7518), .B(n7217), .Z(n7287) );
  AND U7986 ( .A(y[68]), .B(x[49]), .Z(n7286) );
  XOR U7987 ( .A(n7287), .B(n7286), .Z(n7315) );
  XOR U7988 ( .A(n7316), .B(n7315), .Z(n7318) );
  XOR U7989 ( .A(n7318), .B(n7317), .Z(n7329) );
  XOR U7990 ( .A(n7330), .B(n7329), .Z(n7338) );
  AND U7991 ( .A(y[105]), .B(x[60]), .Z(n7223) );
  AND U7992 ( .A(x[61]), .B(y[104]), .Z(n7222) );
  XOR U7993 ( .A(n7223), .B(n7222), .Z(n7298) );
  XOR U7994 ( .A(n7299), .B(n7298), .Z(n7358) );
  AND U7995 ( .A(y[144]), .B(x[69]), .Z(n7291) );
  AND U7996 ( .A(y[26]), .B(x[43]), .Z(n7290) );
  XOR U7997 ( .A(n7291), .B(n7290), .Z(n7294) );
  AND U7998 ( .A(y[27]), .B(x[42]), .Z(n7293) );
  XOR U7999 ( .A(n7294), .B(n7293), .Z(n7357) );
  XOR U8000 ( .A(n7358), .B(n7357), .Z(n7360) );
  NAND U8001 ( .A(n7225), .B(n7224), .Z(n7229) );
  NANDN U8002 ( .A(n7227), .B(n7226), .Z(n7228) );
  AND U8003 ( .A(n7229), .B(n7228), .Z(n7359) );
  XOR U8004 ( .A(n7360), .B(n7359), .Z(n7336) );
  AND U8005 ( .A(y[68]), .B(x[51]), .Z(n7510) );
  NAND U8006 ( .A(n7510), .B(n7230), .Z(n7233) );
  NANDN U8007 ( .A(n7231), .B(n7285), .Z(n7232) );
  NAND U8008 ( .A(n7233), .B(n7232), .Z(n7323) );
  AND U8009 ( .A(y[146]), .B(x[67]), .Z(n7352) );
  AND U8010 ( .A(y[108]), .B(x[57]), .Z(n7596) );
  XOR U8011 ( .A(n7352), .B(n7596), .Z(n7354) );
  AND U8012 ( .A(y[109]), .B(x[56]), .Z(n7353) );
  XOR U8013 ( .A(n7354), .B(n7353), .Z(n7322) );
  AND U8014 ( .A(y[29]), .B(x[40]), .Z(n7345) );
  AND U8015 ( .A(y[148]), .B(x[65]), .Z(n7344) );
  XOR U8016 ( .A(n7345), .B(n7344), .Z(n7347) );
  AND U8017 ( .A(y[147]), .B(x[66]), .Z(n7346) );
  XOR U8018 ( .A(n7347), .B(n7346), .Z(n7321) );
  XNOR U8019 ( .A(n7322), .B(n7321), .Z(n7324) );
  XOR U8020 ( .A(n7323), .B(n7324), .Z(n7335) );
  XNOR U8021 ( .A(n7336), .B(n7335), .Z(n7337) );
  XOR U8022 ( .A(n7338), .B(n7337), .Z(n7263) );
  NANDN U8023 ( .A(n7235), .B(n7234), .Z(n7239) );
  NANDN U8024 ( .A(n7237), .B(n7236), .Z(n7238) );
  AND U8025 ( .A(n7239), .B(n7238), .Z(n7334) );
  NANDN U8026 ( .A(n7245), .B(n7244), .Z(n7249) );
  NANDN U8027 ( .A(n7247), .B(n7246), .Z(n7248) );
  NAND U8028 ( .A(n7249), .B(n7248), .Z(n7332) );
  XOR U8029 ( .A(n7331), .B(n7332), .Z(n7333) );
  XOR U8030 ( .A(n7334), .B(n7333), .Z(n7262) );
  XNOR U8031 ( .A(n7263), .B(n7262), .Z(n7265) );
  XNOR U8032 ( .A(n7264), .B(n7265), .Z(n7375) );
  XNOR U8033 ( .A(n7376), .B(n7375), .Z(n7378) );
  XOR U8034 ( .A(n7266), .B(n7267), .Z(n7269) );
  XOR U8035 ( .A(n7268), .B(n7269), .Z(n7377) );
  XOR U8036 ( .A(n7378), .B(n7377), .Z(n7381) );
  XOR U8037 ( .A(n7382), .B(n7381), .Z(o[69]) );
  XNOR U8038 ( .A(n7655), .B(n7656), .Z(n7653) );
  NAND U8039 ( .A(n7271), .B(n7270), .Z(n7275) );
  NAND U8040 ( .A(n7273), .B(n7272), .Z(n7274) );
  AND U8041 ( .A(n7275), .B(n7274), .Z(n7670) );
  AND U8042 ( .A(y[67]), .B(x[51]), .Z(n7284) );
  NAND U8043 ( .A(n7285), .B(n7284), .Z(n7289) );
  NAND U8044 ( .A(n7287), .B(n7286), .Z(n7288) );
  AND U8045 ( .A(n7289), .B(n7288), .Z(n7549) );
  AND U8046 ( .A(y[147]), .B(x[67]), .Z(n7555) );
  NAND U8047 ( .A(y[107]), .B(x[59]), .Z(n7556) );
  XNOR U8048 ( .A(n7555), .B(n7556), .Z(n7553) );
  NAND U8049 ( .A(y[27]), .B(x[43]), .Z(n7554) );
  XNOR U8050 ( .A(n7553), .B(n7554), .Z(n7548) );
  AND U8051 ( .A(y[148]), .B(x[66]), .Z(n7406) );
  NAND U8052 ( .A(y[106]), .B(x[60]), .Z(n7407) );
  XNOR U8053 ( .A(n7406), .B(n7407), .Z(n7404) );
  NAND U8054 ( .A(y[28]), .B(x[42]), .Z(n7405) );
  XNOR U8055 ( .A(n7404), .B(n7405), .Z(n7547) );
  XNOR U8056 ( .A(n7548), .B(n7547), .Z(n7550) );
  XNOR U8057 ( .A(n7549), .B(n7550), .Z(n7399) );
  IV U8058 ( .A(n7290), .Z(n7292) );
  NANDN U8059 ( .A(n7292), .B(n7291), .Z(n7296) );
  NAND U8060 ( .A(n7294), .B(n7293), .Z(n7295) );
  NAND U8061 ( .A(n7296), .B(n7295), .Z(n7398) );
  XNOR U8062 ( .A(n7399), .B(n7398), .Z(n7400) );
  XNOR U8063 ( .A(n7401), .B(n7400), .Z(n7388) );
  XNOR U8064 ( .A(n7389), .B(n7388), .Z(n7386) );
  AND U8065 ( .A(y[105]), .B(x[61]), .Z(n7440) );
  AND U8066 ( .A(x[45]), .B(y[25]), .Z(n7301) );
  NAND U8067 ( .A(x[44]), .B(y[26]), .Z(n7300) );
  XNOR U8068 ( .A(n7301), .B(n7300), .Z(n7539) );
  NAND U8069 ( .A(y[144]), .B(x[70]), .Z(n7540) );
  XNOR U8070 ( .A(n7539), .B(n7540), .Z(n7456) );
  AND U8071 ( .A(y[189]), .B(x[73]), .Z(n7527) );
  AND U8072 ( .A(y[186]), .B(x[76]), .Z(n7302) );
  AND U8073 ( .A(n7303), .B(n7302), .Z(n7525) );
  AND U8074 ( .A(y[188]), .B(x[74]), .Z(n7526) );
  XNOR U8075 ( .A(n7525), .B(n7526), .Z(n7528) );
  XNOR U8076 ( .A(n7527), .B(n7528), .Z(n7455) );
  XNOR U8077 ( .A(n7456), .B(n7455), .Z(n7458) );
  XNOR U8078 ( .A(n7457), .B(n7458), .Z(n7609) );
  IV U8079 ( .A(n7309), .Z(n7436) );
  XNOR U8080 ( .A(n7608), .B(n7607), .Z(n7610) );
  XNOR U8081 ( .A(n7609), .B(n7610), .Z(n7387) );
  XNOR U8082 ( .A(n7386), .B(n7387), .Z(n7640) );
  XNOR U8083 ( .A(n7640), .B(n7639), .Z(n7637) );
  NAND U8084 ( .A(n7316), .B(n7315), .Z(n7320) );
  NAND U8085 ( .A(n7318), .B(n7317), .Z(n7319) );
  AND U8086 ( .A(n7320), .B(n7319), .Z(n7394) );
  NAND U8087 ( .A(n7322), .B(n7321), .Z(n7326) );
  NANDN U8088 ( .A(n7324), .B(n7323), .Z(n7325) );
  AND U8089 ( .A(n7326), .B(n7325), .Z(n7392) );
  XNOR U8090 ( .A(n7392), .B(n7393), .Z(n7395) );
  XNOR U8091 ( .A(n7394), .B(n7395), .Z(n7638) );
  XNOR U8092 ( .A(n7637), .B(n7638), .Z(n7671) );
  XNOR U8093 ( .A(n7670), .B(n7671), .Z(n7668) );
  NANDN U8094 ( .A(n7336), .B(n7335), .Z(n7340) );
  NANDN U8095 ( .A(n7338), .B(n7337), .Z(n7339) );
  AND U8096 ( .A(n7340), .B(n7339), .Z(n7677) );
  NAND U8097 ( .A(n7345), .B(n7344), .Z(n7349) );
  NAND U8098 ( .A(n7347), .B(n7346), .Z(n7348) );
  AND U8099 ( .A(n7349), .B(n7348), .Z(n7450) );
  AND U8100 ( .A(y[29]), .B(x[41]), .Z(n7445) );
  NAND U8101 ( .A(y[64]), .B(x[54]), .Z(n7446) );
  XNOR U8102 ( .A(n7445), .B(n7446), .Z(n7443) );
  NAND U8103 ( .A(y[70]), .B(x[48]), .Z(n7444) );
  XNOR U8104 ( .A(n7443), .B(n7444), .Z(n7452) );
  AND U8105 ( .A(x[77]), .B(y[185]), .Z(n7351) );
  NAND U8106 ( .A(x[76]), .B(y[186]), .Z(n7350) );
  XOR U8107 ( .A(n7351), .B(n7350), .Z(n7531) );
  NAND U8108 ( .A(y[184]), .B(x[78]), .Z(n7532) );
  XOR U8109 ( .A(n7531), .B(n7532), .Z(n7534) );
  XNOR U8110 ( .A(n7533), .B(n7534), .Z(n7451) );
  XNOR U8111 ( .A(n7452), .B(n7451), .Z(n7449) );
  XNOR U8112 ( .A(n7450), .B(n7449), .Z(n7619) );
  XNOR U8113 ( .A(n7620), .B(n7619), .Z(n7621) );
  NAND U8114 ( .A(n7352), .B(n7596), .Z(n7356) );
  NAND U8115 ( .A(n7354), .B(n7353), .Z(n7355) );
  AND U8116 ( .A(n7356), .B(n7355), .Z(n7622) );
  XNOR U8117 ( .A(n7621), .B(n7622), .Z(n7646) );
  AND U8118 ( .A(y[110]), .B(x[56]), .Z(n7591) );
  NAND U8119 ( .A(y[24]), .B(x[46]), .Z(n7592) );
  XNOR U8120 ( .A(n7591), .B(n7592), .Z(n7589) );
  NAND U8121 ( .A(y[145]), .B(x[69]), .Z(n7590) );
  XNOR U8122 ( .A(n7589), .B(n7590), .Z(n7567) );
  AND U8123 ( .A(y[65]), .B(x[53]), .Z(n7424) );
  NAND U8124 ( .A(y[68]), .B(x[50]), .Z(n7425) );
  XNOR U8125 ( .A(n7424), .B(n7425), .Z(n7422) );
  NAND U8126 ( .A(y[69]), .B(x[49]), .Z(n7423) );
  XNOR U8127 ( .A(n7422), .B(n7423), .Z(n7519) );
  AND U8128 ( .A(x[52]), .B(y[66]), .Z(n7362) );
  NAND U8129 ( .A(x[51]), .B(y[67]), .Z(n7361) );
  XNOR U8130 ( .A(n7362), .B(n7361), .Z(n7520) );
  XNOR U8131 ( .A(n7519), .B(n7520), .Z(n7568) );
  XNOR U8132 ( .A(n7567), .B(n7568), .Z(n7565) );
  AND U8133 ( .A(y[190]), .B(x[72]), .Z(n7439) );
  XOR U8134 ( .A(n7440), .B(n7439), .Z(n7441) );
  AND U8135 ( .A(y[104]), .B(x[62]), .Z(n7442) );
  XNOR U8136 ( .A(n7441), .B(n7442), .Z(n7566) );
  XNOR U8137 ( .A(n7565), .B(n7566), .Z(n7628) );
  AND U8138 ( .A(y[146]), .B(x[68]), .Z(n7597) );
  AND U8139 ( .A(x[57]), .B(y[109]), .Z(n7368) );
  AND U8140 ( .A(x[58]), .B(y[108]), .Z(n7367) );
  XNOR U8141 ( .A(n7368), .B(n7367), .Z(n7598) );
  XNOR U8142 ( .A(n7597), .B(n7598), .Z(n7462) );
  AND U8143 ( .A(y[30]), .B(x[40]), .Z(n7437) );
  AND U8144 ( .A(y[150]), .B(x[64]), .Z(n7370) );
  AND U8145 ( .A(x[65]), .B(y[149]), .Z(n7369) );
  XNOR U8146 ( .A(n7370), .B(n7369), .Z(n7438) );
  XNOR U8147 ( .A(n7437), .B(n7438), .Z(n7461) );
  XNOR U8148 ( .A(n7462), .B(n7461), .Z(n7464) );
  XNOR U8149 ( .A(n7463), .B(n7464), .Z(n7627) );
  XNOR U8150 ( .A(n7628), .B(n7627), .Z(n7625) );
  XNOR U8151 ( .A(n7625), .B(n7626), .Z(n7644) );
  XNOR U8152 ( .A(n7643), .B(n7644), .Z(n7645) );
  XNOR U8153 ( .A(n7646), .B(n7645), .Z(n7676) );
  XNOR U8154 ( .A(n7677), .B(n7676), .Z(n7674) );
  XNOR U8155 ( .A(n7675), .B(n7674), .Z(n7669) );
  XNOR U8156 ( .A(n7668), .B(n7669), .Z(n7654) );
  XOR U8157 ( .A(n7653), .B(n7654), .Z(n7659) );
  NANDN U8158 ( .A(n7380), .B(n7379), .Z(n7384) );
  NAND U8159 ( .A(n7382), .B(n7381), .Z(n7383) );
  AND U8160 ( .A(n7384), .B(n7383), .Z(n7660) );
  XNOR U8161 ( .A(n7661), .B(n7660), .Z(n7385) );
  XOR U8162 ( .A(n7659), .B(n7385), .Z(o[70]) );
  NANDN U8163 ( .A(n7387), .B(n7386), .Z(n7391) );
  NANDN U8164 ( .A(n7389), .B(n7388), .Z(n7390) );
  AND U8165 ( .A(n7391), .B(n7390), .Z(n7636) );
  NAND U8166 ( .A(n7393), .B(n7392), .Z(n7397) );
  NANDN U8167 ( .A(n7395), .B(n7394), .Z(n7396) );
  AND U8168 ( .A(n7397), .B(n7396), .Z(n7618) );
  NANDN U8169 ( .A(n7399), .B(n7398), .Z(n7403) );
  NANDN U8170 ( .A(n7401), .B(n7400), .Z(n7402) );
  NAND U8171 ( .A(n7403), .B(n7402), .Z(n7616) );
  NANDN U8172 ( .A(n7405), .B(n7404), .Z(n7409) );
  NANDN U8173 ( .A(n7407), .B(n7406), .Z(n7408) );
  AND U8174 ( .A(n7409), .B(n7408), .Z(n7435) );
  AND U8175 ( .A(x[43]), .B(y[28]), .Z(n7411) );
  NAND U8176 ( .A(x[79]), .B(y[184]), .Z(n7410) );
  XNOR U8177 ( .A(n7411), .B(n7410), .Z(n7421) );
  AND U8178 ( .A(y[186]), .B(x[77]), .Z(n7509) );
  AND U8179 ( .A(n7412), .B(n7509), .Z(n7416) );
  AND U8180 ( .A(x[48]), .B(y[71]), .Z(n7414) );
  NAND U8181 ( .A(x[70]), .B(y[145]), .Z(n7413) );
  XNOR U8182 ( .A(n7414), .B(n7413), .Z(n7415) );
  XOR U8183 ( .A(n7416), .B(n7415), .Z(n7419) );
  AND U8184 ( .A(y[26]), .B(x[45]), .Z(n7537) );
  XNOR U8185 ( .A(n7417), .B(n7537), .Z(n7418) );
  XNOR U8186 ( .A(n7419), .B(n7418), .Z(n7420) );
  XOR U8187 ( .A(n7421), .B(n7420), .Z(n7433) );
  NANDN U8188 ( .A(n7423), .B(n7422), .Z(n7427) );
  NANDN U8189 ( .A(n7425), .B(n7424), .Z(n7426) );
  AND U8190 ( .A(n7427), .B(n7426), .Z(n7431) );
  AND U8191 ( .A(x[42]), .B(y[29]), .Z(n7429) );
  NAND U8192 ( .A(x[54]), .B(y[65]), .Z(n7428) );
  XNOR U8193 ( .A(n7429), .B(n7428), .Z(n7430) );
  XNOR U8194 ( .A(n7431), .B(n7430), .Z(n7432) );
  XNOR U8195 ( .A(n7433), .B(n7432), .Z(n7434) );
  XOR U8196 ( .A(n7435), .B(n7434), .Z(n7448) );
  AND U8197 ( .A(y[150]), .B(x[65]), .Z(n7476) );
  XNOR U8198 ( .A(n7448), .B(n7447), .Z(n7472) );
  NAND U8199 ( .A(n7450), .B(n7449), .Z(n7454) );
  NANDN U8200 ( .A(n7452), .B(n7451), .Z(n7453) );
  NAND U8201 ( .A(n7454), .B(n7453), .Z(n7470) );
  OR U8202 ( .A(n7456), .B(n7455), .Z(n7460) );
  NANDN U8203 ( .A(n7458), .B(n7457), .Z(n7459) );
  AND U8204 ( .A(n7460), .B(n7459), .Z(n7468) );
  OR U8205 ( .A(n7462), .B(n7461), .Z(n7466) );
  NANDN U8206 ( .A(n7464), .B(n7463), .Z(n7465) );
  NAND U8207 ( .A(n7466), .B(n7465), .Z(n7467) );
  XNOR U8208 ( .A(n7468), .B(n7467), .Z(n7469) );
  XNOR U8209 ( .A(n7470), .B(n7469), .Z(n7471) );
  XOR U8210 ( .A(n7472), .B(n7471), .Z(n7606) );
  AND U8211 ( .A(x[55]), .B(y[64]), .Z(n7478) );
  AND U8212 ( .A(x[66]), .B(y[149]), .Z(n7474) );
  NAND U8213 ( .A(x[53]), .B(y[66]), .Z(n7473) );
  XNOR U8214 ( .A(n7474), .B(n7473), .Z(n7475) );
  XNOR U8215 ( .A(n7476), .B(n7475), .Z(n7477) );
  XNOR U8216 ( .A(n7478), .B(n7477), .Z(n7494) );
  AND U8217 ( .A(x[59]), .B(y[108]), .Z(n7480) );
  NAND U8218 ( .A(x[46]), .B(y[25]), .Z(n7479) );
  XNOR U8219 ( .A(n7480), .B(n7479), .Z(n7484) );
  AND U8220 ( .A(x[71]), .B(y[144]), .Z(n7482) );
  NAND U8221 ( .A(x[67]), .B(y[148]), .Z(n7481) );
  XNOR U8222 ( .A(n7482), .B(n7481), .Z(n7483) );
  XOR U8223 ( .A(n7484), .B(n7483), .Z(n7492) );
  AND U8224 ( .A(x[56]), .B(y[111]), .Z(n7486) );
  NAND U8225 ( .A(x[64]), .B(y[151]), .Z(n7485) );
  XNOR U8226 ( .A(n7486), .B(n7485), .Z(n7490) );
  AND U8227 ( .A(x[49]), .B(y[70]), .Z(n7488) );
  NAND U8228 ( .A(x[50]), .B(y[69]), .Z(n7487) );
  XNOR U8229 ( .A(n7488), .B(n7487), .Z(n7489) );
  XNOR U8230 ( .A(n7490), .B(n7489), .Z(n7491) );
  XNOR U8231 ( .A(n7492), .B(n7491), .Z(n7493) );
  XOR U8232 ( .A(n7494), .B(n7493), .Z(n7516) );
  AND U8233 ( .A(x[41]), .B(y[30]), .Z(n7496) );
  NAND U8234 ( .A(x[69]), .B(y[146]), .Z(n7495) );
  XNOR U8235 ( .A(n7496), .B(n7495), .Z(n7500) );
  AND U8236 ( .A(x[78]), .B(y[185]), .Z(n7498) );
  NAND U8237 ( .A(x[61]), .B(y[106]), .Z(n7497) );
  XNOR U8238 ( .A(n7498), .B(n7497), .Z(n7499) );
  XOR U8239 ( .A(n7500), .B(n7499), .Z(n7508) );
  AND U8240 ( .A(x[40]), .B(y[31]), .Z(n7502) );
  NAND U8241 ( .A(x[73]), .B(y[190]), .Z(n7501) );
  XNOR U8242 ( .A(n7502), .B(n7501), .Z(n7506) );
  AND U8243 ( .A(x[72]), .B(y[191]), .Z(n7504) );
  NAND U8244 ( .A(x[63]), .B(y[104]), .Z(n7503) );
  XNOR U8245 ( .A(n7504), .B(n7503), .Z(n7505) );
  XNOR U8246 ( .A(n7506), .B(n7505), .Z(n7507) );
  XNOR U8247 ( .A(n7508), .B(n7507), .Z(n7514) );
  AND U8248 ( .A(y[67]), .B(x[52]), .Z(n7517) );
  AND U8249 ( .A(y[109]), .B(x[58]), .Z(n7595) );
  XOR U8250 ( .A(n7517), .B(n7595), .Z(n7512) );
  XNOR U8251 ( .A(n7510), .B(n7509), .Z(n7511) );
  XNOR U8252 ( .A(n7512), .B(n7511), .Z(n7513) );
  XNOR U8253 ( .A(n7514), .B(n7513), .Z(n7515) );
  XNOR U8254 ( .A(n7516), .B(n7515), .Z(n7524) );
  NAND U8255 ( .A(n7518), .B(n7517), .Z(n7522) );
  NAND U8256 ( .A(n7520), .B(n7519), .Z(n7521) );
  NAND U8257 ( .A(n7522), .B(n7521), .Z(n7523) );
  XNOR U8258 ( .A(n7524), .B(n7523), .Z(n7564) );
  NAND U8259 ( .A(n7526), .B(n7525), .Z(n7530) );
  NANDN U8260 ( .A(n7528), .B(n7527), .Z(n7529) );
  AND U8261 ( .A(n7530), .B(n7529), .Z(n7546) );
  OR U8262 ( .A(n7532), .B(n7531), .Z(n7536) );
  NAND U8263 ( .A(n7534), .B(n7533), .Z(n7535) );
  AND U8264 ( .A(n7536), .B(n7535), .Z(n7544) );
  NAND U8265 ( .A(n7538), .B(n7537), .Z(n7542) );
  NANDN U8266 ( .A(n7540), .B(n7539), .Z(n7541) );
  NAND U8267 ( .A(n7542), .B(n7541), .Z(n7543) );
  XNOR U8268 ( .A(n7544), .B(n7543), .Z(n7545) );
  XOR U8269 ( .A(n7546), .B(n7545), .Z(n7562) );
  OR U8270 ( .A(n7548), .B(n7547), .Z(n7552) );
  NANDN U8271 ( .A(n7550), .B(n7549), .Z(n7551) );
  AND U8272 ( .A(n7552), .B(n7551), .Z(n7560) );
  NANDN U8273 ( .A(n7554), .B(n7553), .Z(n7558) );
  NANDN U8274 ( .A(n7556), .B(n7555), .Z(n7557) );
  AND U8275 ( .A(n7558), .B(n7557), .Z(n7559) );
  XNOR U8276 ( .A(n7560), .B(n7559), .Z(n7561) );
  XNOR U8277 ( .A(n7562), .B(n7561), .Z(n7563) );
  XOR U8278 ( .A(n7564), .B(n7563), .Z(n7588) );
  NANDN U8279 ( .A(n7566), .B(n7565), .Z(n7570) );
  NANDN U8280 ( .A(n7568), .B(n7567), .Z(n7569) );
  AND U8281 ( .A(n7570), .B(n7569), .Z(n7586) );
  AND U8282 ( .A(x[74]), .B(y[189]), .Z(n7572) );
  NAND U8283 ( .A(x[44]), .B(y[27]), .Z(n7571) );
  XNOR U8284 ( .A(n7572), .B(n7571), .Z(n7576) );
  AND U8285 ( .A(x[47]), .B(y[24]), .Z(n7574) );
  NAND U8286 ( .A(x[68]), .B(y[147]), .Z(n7573) );
  XNOR U8287 ( .A(n7574), .B(n7573), .Z(n7575) );
  XOR U8288 ( .A(n7576), .B(n7575), .Z(n7584) );
  AND U8289 ( .A(x[60]), .B(y[107]), .Z(n7578) );
  NAND U8290 ( .A(x[62]), .B(y[105]), .Z(n7577) );
  XNOR U8291 ( .A(n7578), .B(n7577), .Z(n7582) );
  AND U8292 ( .A(x[57]), .B(y[110]), .Z(n7580) );
  NAND U8293 ( .A(x[75]), .B(y[188]), .Z(n7579) );
  XNOR U8294 ( .A(n7580), .B(n7579), .Z(n7581) );
  XNOR U8295 ( .A(n7582), .B(n7581), .Z(n7583) );
  XNOR U8296 ( .A(n7584), .B(n7583), .Z(n7585) );
  XNOR U8297 ( .A(n7586), .B(n7585), .Z(n7587) );
  XNOR U8298 ( .A(n7588), .B(n7587), .Z(n7604) );
  NANDN U8299 ( .A(n7590), .B(n7589), .Z(n7594) );
  NANDN U8300 ( .A(n7592), .B(n7591), .Z(n7593) );
  AND U8301 ( .A(n7594), .B(n7593), .Z(n7602) );
  NAND U8302 ( .A(n7596), .B(n7595), .Z(n7600) );
  NANDN U8303 ( .A(n7598), .B(n7597), .Z(n7599) );
  NAND U8304 ( .A(n7600), .B(n7599), .Z(n7601) );
  XNOR U8305 ( .A(n7602), .B(n7601), .Z(n7603) );
  XNOR U8306 ( .A(n7604), .B(n7603), .Z(n7605) );
  XNOR U8307 ( .A(n7606), .B(n7605), .Z(n7614) );
  OR U8308 ( .A(n7608), .B(n7607), .Z(n7612) );
  OR U8309 ( .A(n7610), .B(n7609), .Z(n7611) );
  NAND U8310 ( .A(n7612), .B(n7611), .Z(n7613) );
  XNOR U8311 ( .A(n7614), .B(n7613), .Z(n7615) );
  XNOR U8312 ( .A(n7616), .B(n7615), .Z(n7617) );
  XOR U8313 ( .A(n7618), .B(n7617), .Z(n7634) );
  NANDN U8314 ( .A(n7620), .B(n7619), .Z(n7624) );
  NANDN U8315 ( .A(n7622), .B(n7621), .Z(n7623) );
  NAND U8316 ( .A(n7624), .B(n7623), .Z(n7632) );
  NAND U8317 ( .A(n7626), .B(n7625), .Z(n7630) );
  NANDN U8318 ( .A(n7628), .B(n7627), .Z(n7629) );
  AND U8319 ( .A(n7630), .B(n7629), .Z(n7631) );
  XOR U8320 ( .A(n7632), .B(n7631), .Z(n7633) );
  XNOR U8321 ( .A(n7634), .B(n7633), .Z(n7635) );
  XOR U8322 ( .A(n7636), .B(n7635), .Z(n7652) );
  NAND U8323 ( .A(n7638), .B(n7637), .Z(n7642) );
  NANDN U8324 ( .A(n7640), .B(n7639), .Z(n7641) );
  AND U8325 ( .A(n7642), .B(n7641), .Z(n7650) );
  NANDN U8326 ( .A(n7644), .B(n7643), .Z(n7648) );
  NANDN U8327 ( .A(n7646), .B(n7645), .Z(n7647) );
  AND U8328 ( .A(n7648), .B(n7647), .Z(n7649) );
  XNOR U8329 ( .A(n7650), .B(n7649), .Z(n7651) );
  XNOR U8330 ( .A(n7652), .B(n7651), .Z(n7667) );
  NAND U8331 ( .A(n7654), .B(n7653), .Z(n7658) );
  NANDN U8332 ( .A(n7656), .B(n7655), .Z(n7657) );
  AND U8333 ( .A(n7658), .B(n7657), .Z(n7665) );
  NAND U8334 ( .A(n7661), .B(n7660), .Z(n7663) );
  AND U8335 ( .A(n7663), .B(n7662), .Z(n7664) );
  XNOR U8336 ( .A(n7665), .B(n7664), .Z(n7666) );
  XOR U8337 ( .A(n7667), .B(n7666), .Z(n7683) );
  NANDN U8338 ( .A(n7669), .B(n7668), .Z(n7673) );
  NANDN U8339 ( .A(n7671), .B(n7670), .Z(n7672) );
  AND U8340 ( .A(n7673), .B(n7672), .Z(n7681) );
  NAND U8341 ( .A(n7675), .B(n7674), .Z(n7679) );
  NANDN U8342 ( .A(n7677), .B(n7676), .Z(n7678) );
  AND U8343 ( .A(n7679), .B(n7678), .Z(n7680) );
  XNOR U8344 ( .A(n7681), .B(n7680), .Z(n7682) );
  XNOR U8345 ( .A(n7683), .B(n7682), .Z(o[71]) );
  NAND U8346 ( .A(y[192]), .B(x[72]), .Z(n7818) );
  NAND U8347 ( .A(y[72]), .B(x[48]), .Z(n7686) );
  XOR U8348 ( .A(n7818), .B(n7686), .Z(n7687) );
  AND U8349 ( .A(y[32]), .B(x[40]), .Z(n7694) );
  AND U8350 ( .A(y[112]), .B(x[56]), .Z(n7691) );
  XOR U8351 ( .A(n7694), .B(n7691), .Z(n7690) );
  AND U8352 ( .A(y[152]), .B(x[64]), .Z(n7689) );
  XNOR U8353 ( .A(n7690), .B(n7689), .Z(n7688) );
  XNOR U8354 ( .A(n7687), .B(n7688), .Z(o[72]) );
  AND U8355 ( .A(x[41]), .B(y[32]), .Z(n7685) );
  NAND U8356 ( .A(x[40]), .B(y[33]), .Z(n7684) );
  XNOR U8357 ( .A(n7685), .B(n7684), .Z(n7695) );
  NAND U8358 ( .A(y[72]), .B(x[49]), .Z(n7696) );
  XOR U8359 ( .A(n7695), .B(n7696), .Z(n7712) );
  AND U8360 ( .A(y[192]), .B(x[73]), .Z(n7919) );
  NAND U8361 ( .A(y[113]), .B(x[56]), .Z(n7699) );
  XNOR U8362 ( .A(n7919), .B(n7699), .Z(n7700) );
  AND U8363 ( .A(y[193]), .B(x[72]), .Z(n7723) );
  NAND U8364 ( .A(y[112]), .B(x[57]), .Z(n7722) );
  XOR U8365 ( .A(n7723), .B(n7722), .Z(n7701) );
  XOR U8366 ( .A(n7700), .B(n7701), .Z(n7711) );
  AND U8367 ( .A(y[73]), .B(x[48]), .Z(n7942) );
  AND U8368 ( .A(y[153]), .B(x[64]), .Z(n7716) );
  XOR U8369 ( .A(n7942), .B(n7716), .Z(n7718) );
  AND U8370 ( .A(y[152]), .B(x[65]), .Z(n7717) );
  XNOR U8371 ( .A(n7718), .B(n7717), .Z(n7710) );
  XOR U8372 ( .A(n7711), .B(n7710), .Z(n7713) );
  XOR U8373 ( .A(n7712), .B(n7713), .Z(n7707) );
  NAND U8374 ( .A(n7690), .B(n7689), .Z(n7693) );
  AND U8375 ( .A(n7694), .B(n7691), .Z(n7692) );
  ANDN U8376 ( .B(n7693), .A(n7692), .Z(n7704) );
  XNOR U8377 ( .A(n7705), .B(n7704), .Z(n7706) );
  XNOR U8378 ( .A(n7707), .B(n7706), .Z(o[73]) );
  AND U8379 ( .A(y[33]), .B(x[41]), .Z(n7754) );
  NAND U8380 ( .A(n7754), .B(n7694), .Z(n7698) );
  NANDN U8381 ( .A(n7696), .B(n7695), .Z(n7697) );
  NAND U8382 ( .A(n7698), .B(n7697), .Z(n7766) );
  NANDN U8383 ( .A(n7699), .B(n7919), .Z(n7703) );
  NANDN U8384 ( .A(n7701), .B(n7700), .Z(n7702) );
  NAND U8385 ( .A(n7703), .B(n7702), .Z(n7764) );
  AND U8386 ( .A(y[154]), .B(x[64]), .Z(n7770) );
  NAND U8387 ( .A(y[34]), .B(x[40]), .Z(n7771) );
  XNOR U8388 ( .A(n7770), .B(n7771), .Z(n7773) );
  AND U8389 ( .A(y[72]), .B(x[50]), .Z(n7772) );
  XOR U8390 ( .A(n7773), .B(n7772), .Z(n7765) );
  XOR U8391 ( .A(n7764), .B(n7765), .Z(n7767) );
  XNOR U8392 ( .A(n7766), .B(n7767), .Z(n7725) );
  NANDN U8393 ( .A(n7705), .B(n7704), .Z(n7709) );
  NAND U8394 ( .A(n7707), .B(n7706), .Z(n7708) );
  NAND U8395 ( .A(n7709), .B(n7708), .Z(n7724) );
  XOR U8396 ( .A(n7725), .B(n7724), .Z(n7727) );
  NAND U8397 ( .A(n7711), .B(n7710), .Z(n7715) );
  NAND U8398 ( .A(n7713), .B(n7712), .Z(n7714) );
  AND U8399 ( .A(n7715), .B(n7714), .Z(n7733) );
  AND U8400 ( .A(y[32]), .B(x[42]), .Z(n7752) );
  AND U8401 ( .A(y[114]), .B(x[56]), .Z(n7751) );
  XOR U8402 ( .A(n7752), .B(n7751), .Z(n7753) );
  XOR U8403 ( .A(n7754), .B(n7753), .Z(n7779) );
  AND U8404 ( .A(y[152]), .B(x[66]), .Z(n7778) );
  XOR U8405 ( .A(n7779), .B(n7778), .Z(n7781) );
  AND U8406 ( .A(y[112]), .B(x[58]), .Z(n7849) );
  AND U8407 ( .A(y[194]), .B(x[72]), .Z(n7742) );
  XOR U8408 ( .A(n7849), .B(n7742), .Z(n7744) );
  AND U8409 ( .A(y[113]), .B(x[57]), .Z(n7743) );
  XOR U8410 ( .A(n7744), .B(n7743), .Z(n7780) );
  XOR U8411 ( .A(n7781), .B(n7780), .Z(n7730) );
  AND U8412 ( .A(n7942), .B(n7716), .Z(n7720) );
  NAND U8413 ( .A(n7718), .B(n7717), .Z(n7719) );
  NANDN U8414 ( .A(n7720), .B(n7719), .Z(n7738) );
  AND U8415 ( .A(x[73]), .B(y[193]), .Z(n7823) );
  NAND U8416 ( .A(x[74]), .B(y[192]), .Z(n7721) );
  XNOR U8417 ( .A(n7823), .B(n7721), .Z(n7777) );
  ANDN U8418 ( .B(n7723), .A(n7722), .Z(n7776) );
  XOR U8419 ( .A(n7777), .B(n7776), .Z(n7737) );
  AND U8420 ( .A(y[153]), .B(x[65]), .Z(n7757) );
  NAND U8421 ( .A(y[73]), .B(x[49]), .Z(n7758) );
  XNOR U8422 ( .A(n7757), .B(n7758), .Z(n7759) );
  NAND U8423 ( .A(y[74]), .B(x[48]), .Z(n7760) );
  XNOR U8424 ( .A(n7759), .B(n7760), .Z(n7736) );
  XOR U8425 ( .A(n7737), .B(n7736), .Z(n7739) );
  XOR U8426 ( .A(n7738), .B(n7739), .Z(n7731) );
  XOR U8427 ( .A(n7730), .B(n7731), .Z(n7732) );
  XNOR U8428 ( .A(n7733), .B(n7732), .Z(n7726) );
  XNOR U8429 ( .A(n7727), .B(n7726), .Z(o[74]) );
  NAND U8430 ( .A(n7725), .B(n7724), .Z(n7729) );
  NAND U8431 ( .A(n7727), .B(n7726), .Z(n7728) );
  AND U8432 ( .A(n7729), .B(n7728), .Z(n7785) );
  NAND U8433 ( .A(n7731), .B(n7730), .Z(n7735) );
  NAND U8434 ( .A(n7733), .B(n7732), .Z(n7734) );
  NAND U8435 ( .A(n7735), .B(n7734), .Z(n7790) );
  NAND U8436 ( .A(n7737), .B(n7736), .Z(n7741) );
  NAND U8437 ( .A(n7739), .B(n7738), .Z(n7740) );
  NAND U8438 ( .A(n7741), .B(n7740), .Z(n7788) );
  AND U8439 ( .A(y[34]), .B(x[41]), .Z(n7814) );
  AND U8440 ( .A(y[33]), .B(x[42]), .Z(n7813) );
  NAND U8441 ( .A(y[154]), .B(x[65]), .Z(n7812) );
  XOR U8442 ( .A(n7813), .B(n7812), .Z(n7815) );
  XOR U8443 ( .A(n7814), .B(n7815), .Z(n7845) );
  NAND U8444 ( .A(n7849), .B(n7742), .Z(n7746) );
  AND U8445 ( .A(n7744), .B(n7743), .Z(n7745) );
  ANDN U8446 ( .B(n7746), .A(n7745), .Z(n7843) );
  AND U8447 ( .A(x[75]), .B(y[192]), .Z(n7748) );
  NAND U8448 ( .A(x[72]), .B(y[195]), .Z(n7747) );
  XNOR U8449 ( .A(n7748), .B(n7747), .Z(n7819) );
  AND U8450 ( .A(x[73]), .B(y[194]), .Z(n7750) );
  NAND U8451 ( .A(x[74]), .B(y[193]), .Z(n7749) );
  XOR U8452 ( .A(n7750), .B(n7749), .Z(n7820) );
  XNOR U8453 ( .A(n7819), .B(n7820), .Z(n7842) );
  XNOR U8454 ( .A(n7843), .B(n7842), .Z(n7844) );
  XNOR U8455 ( .A(n7845), .B(n7844), .Z(n7802) );
  NAND U8456 ( .A(n7752), .B(n7751), .Z(n7756) );
  NAND U8457 ( .A(n7754), .B(n7753), .Z(n7755) );
  NAND U8458 ( .A(n7756), .B(n7755), .Z(n7800) );
  NANDN U8459 ( .A(n7758), .B(n7757), .Z(n7762) );
  NANDN U8460 ( .A(n7760), .B(n7759), .Z(n7761) );
  AND U8461 ( .A(n7762), .B(n7761), .Z(n7838) );
  AND U8462 ( .A(y[155]), .B(x[64]), .Z(n7867) );
  AND U8463 ( .A(y[115]), .B(x[56]), .Z(n7866) );
  NAND U8464 ( .A(y[32]), .B(x[43]), .Z(n7865) );
  XOR U8465 ( .A(n7866), .B(n7865), .Z(n7868) );
  XOR U8466 ( .A(n7867), .B(n7868), .Z(n7837) );
  AND U8467 ( .A(y[113]), .B(x[58]), .Z(n7899) );
  NAND U8468 ( .A(x[59]), .B(y[112]), .Z(n7763) );
  XNOR U8469 ( .A(n7899), .B(n7763), .Z(n7850) );
  NAND U8470 ( .A(y[114]), .B(x[57]), .Z(n7851) );
  XNOR U8471 ( .A(n7850), .B(n7851), .Z(n7836) );
  XOR U8472 ( .A(n7837), .B(n7836), .Z(n7839) );
  XOR U8473 ( .A(n7838), .B(n7839), .Z(n7801) );
  XOR U8474 ( .A(n7800), .B(n7801), .Z(n7803) );
  XOR U8475 ( .A(n7802), .B(n7803), .Z(n7789) );
  XOR U8476 ( .A(n7788), .B(n7789), .Z(n7791) );
  XOR U8477 ( .A(n7790), .B(n7791), .Z(n7784) );
  XOR U8478 ( .A(n7785), .B(n7784), .Z(n7787) );
  NAND U8479 ( .A(n7765), .B(n7764), .Z(n7769) );
  NAND U8480 ( .A(n7767), .B(n7766), .Z(n7768) );
  AND U8481 ( .A(n7769), .B(n7768), .Z(n7797) );
  NANDN U8482 ( .A(n7771), .B(n7770), .Z(n7775) );
  NAND U8483 ( .A(n7773), .B(n7772), .Z(n7774) );
  AND U8484 ( .A(n7775), .B(n7774), .Z(n7807) );
  AND U8485 ( .A(y[193]), .B(x[74]), .Z(n7916) );
  XNOR U8486 ( .A(n7807), .B(n7806), .Z(n7809) );
  NAND U8487 ( .A(y[72]), .B(x[51]), .Z(n7859) );
  NAND U8488 ( .A(y[35]), .B(x[40]), .Z(n7857) );
  NAND U8489 ( .A(y[153]), .B(x[66]), .Z(n7856) );
  XOR U8490 ( .A(n7857), .B(n7856), .Z(n7858) );
  XNOR U8491 ( .A(n7859), .B(n7858), .Z(n7833) );
  NAND U8492 ( .A(y[75]), .B(x[48]), .Z(n7827) );
  NAND U8493 ( .A(y[73]), .B(x[50]), .Z(n7825) );
  NAND U8494 ( .A(y[152]), .B(x[67]), .Z(n7824) );
  XOR U8495 ( .A(n7825), .B(n7824), .Z(n7826) );
  XNOR U8496 ( .A(n7827), .B(n7826), .Z(n7831) );
  AND U8497 ( .A(y[74]), .B(x[49]), .Z(n7830) );
  XOR U8498 ( .A(n7831), .B(n7830), .Z(n7832) );
  XOR U8499 ( .A(n7833), .B(n7832), .Z(n7808) );
  XNOR U8500 ( .A(n7809), .B(n7808), .Z(n7795) );
  NAND U8501 ( .A(n7779), .B(n7778), .Z(n7783) );
  NAND U8502 ( .A(n7781), .B(n7780), .Z(n7782) );
  AND U8503 ( .A(n7783), .B(n7782), .Z(n7794) );
  XOR U8504 ( .A(n7795), .B(n7794), .Z(n7796) );
  XNOR U8505 ( .A(n7797), .B(n7796), .Z(n7786) );
  XOR U8506 ( .A(n7787), .B(n7786), .Z(o[75]) );
  NAND U8507 ( .A(n7789), .B(n7788), .Z(n7793) );
  NAND U8508 ( .A(n7791), .B(n7790), .Z(n7792) );
  AND U8509 ( .A(n7793), .B(n7792), .Z(n7877) );
  NAND U8510 ( .A(n7795), .B(n7794), .Z(n7799) );
  NAND U8511 ( .A(n7797), .B(n7796), .Z(n7798) );
  NAND U8512 ( .A(n7799), .B(n7798), .Z(n7875) );
  NAND U8513 ( .A(n7801), .B(n7800), .Z(n7805) );
  NAND U8514 ( .A(n7803), .B(n7802), .Z(n7804) );
  AND U8515 ( .A(n7805), .B(n7804), .Z(n7876) );
  XOR U8516 ( .A(n7875), .B(n7876), .Z(n7878) );
  XOR U8517 ( .A(n7877), .B(n7878), .Z(n7871) );
  XOR U8518 ( .A(n7872), .B(n7871), .Z(n7874) );
  AND U8519 ( .A(y[74]), .B(x[50]), .Z(n8003) );
  AND U8520 ( .A(x[48]), .B(y[76]), .Z(n7811) );
  NAND U8521 ( .A(x[51]), .B(y[73]), .Z(n7810) );
  XOR U8522 ( .A(n7811), .B(n7810), .Z(n7943) );
  NAND U8523 ( .A(y[75]), .B(x[49]), .Z(n7953) );
  AND U8524 ( .A(y[152]), .B(x[68]), .Z(n7904) );
  NAND U8525 ( .A(y[35]), .B(x[41]), .Z(n7905) );
  NAND U8526 ( .A(y[36]), .B(x[40]), .Z(n7907) );
  XOR U8527 ( .A(n7955), .B(n7954), .Z(n7949) );
  NANDN U8528 ( .A(n7813), .B(n7812), .Z(n7817) );
  OR U8529 ( .A(n7815), .B(n7814), .Z(n7816) );
  AND U8530 ( .A(n7817), .B(n7816), .Z(n7947) );
  AND U8531 ( .A(y[195]), .B(x[75]), .Z(n8222) );
  NANDN U8532 ( .A(n7818), .B(n8222), .Z(n7822) );
  NANDN U8533 ( .A(n7820), .B(n7819), .Z(n7821) );
  AND U8534 ( .A(n7822), .B(n7821), .Z(n7946) );
  NAND U8535 ( .A(y[32]), .B(x[44]), .Z(n7928) );
  NAND U8536 ( .A(y[154]), .B(x[66]), .Z(n7927) );
  NAND U8537 ( .A(y[116]), .B(x[56]), .Z(n7926) );
  XNOR U8538 ( .A(n7927), .B(n7926), .Z(n7929) );
  AND U8539 ( .A(y[194]), .B(x[74]), .Z(n7864) );
  NAND U8540 ( .A(n7864), .B(n7823), .Z(n7924) );
  NAND U8541 ( .A(y[112]), .B(x[60]), .Z(n8024) );
  NAND U8542 ( .A(y[196]), .B(x[72]), .Z(n8068) );
  XNOR U8543 ( .A(n8024), .B(n8068), .Z(n7925) );
  XOR U8544 ( .A(n7924), .B(n7925), .Z(n7887) );
  XOR U8545 ( .A(n7888), .B(n7887), .Z(n7890) );
  NAND U8546 ( .A(n7825), .B(n7824), .Z(n7829) );
  NAND U8547 ( .A(n7827), .B(n7826), .Z(n7828) );
  AND U8548 ( .A(n7829), .B(n7828), .Z(n7889) );
  XOR U8549 ( .A(n7890), .B(n7889), .Z(n7973) );
  NAND U8550 ( .A(n7831), .B(n7830), .Z(n7835) );
  NAND U8551 ( .A(n7833), .B(n7832), .Z(n7834) );
  AND U8552 ( .A(n7835), .B(n7834), .Z(n7972) );
  XNOR U8553 ( .A(n7973), .B(n7972), .Z(n7974) );
  XNOR U8554 ( .A(n7975), .B(n7974), .Z(n7881) );
  XNOR U8555 ( .A(n7882), .B(n7881), .Z(n7884) );
  NANDN U8556 ( .A(n7837), .B(n7836), .Z(n7841) );
  OR U8557 ( .A(n7839), .B(n7838), .Z(n7840) );
  AND U8558 ( .A(n7841), .B(n7840), .Z(n7965) );
  NANDN U8559 ( .A(n7843), .B(n7842), .Z(n7847) );
  NANDN U8560 ( .A(n7845), .B(n7844), .Z(n7846) );
  NAND U8561 ( .A(n7847), .B(n7846), .Z(n7964) );
  XNOR U8562 ( .A(n7965), .B(n7964), .Z(n7967) );
  AND U8563 ( .A(y[113]), .B(x[59]), .Z(n7848) );
  NAND U8564 ( .A(n7849), .B(n7848), .Z(n7853) );
  NANDN U8565 ( .A(n7851), .B(n7850), .Z(n7852) );
  AND U8566 ( .A(n7853), .B(n7852), .Z(n7969) );
  AND U8567 ( .A(y[72]), .B(x[52]), .Z(n7910) );
  NAND U8568 ( .A(y[156]), .B(x[64]), .Z(n7911) );
  NAND U8569 ( .A(y[155]), .B(x[65]), .Z(n7913) );
  AND U8570 ( .A(x[58]), .B(y[114]), .Z(n7855) );
  NAND U8571 ( .A(x[59]), .B(y[113]), .Z(n7854) );
  XNOR U8572 ( .A(n7855), .B(n7854), .Z(n7900) );
  NAND U8573 ( .A(y[115]), .B(x[57]), .Z(n7901) );
  XOR U8574 ( .A(n7959), .B(n7958), .Z(n7960) );
  NAND U8575 ( .A(n7857), .B(n7856), .Z(n7861) );
  NAND U8576 ( .A(n7859), .B(n7858), .Z(n7860) );
  NAND U8577 ( .A(n7861), .B(n7860), .Z(n7961) );
  XNOR U8578 ( .A(n7969), .B(n7968), .Z(n7971) );
  NAND U8579 ( .A(y[34]), .B(x[42]), .Z(n7938) );
  NAND U8580 ( .A(y[153]), .B(x[67]), .Z(n7937) );
  NAND U8581 ( .A(y[33]), .B(x[43]), .Z(n7936) );
  XNOR U8582 ( .A(n7937), .B(n7936), .Z(n7939) );
  AND U8583 ( .A(x[76]), .B(y[192]), .Z(n7863) );
  NAND U8584 ( .A(x[73]), .B(y[195]), .Z(n7862) );
  XNOR U8585 ( .A(n7863), .B(n7862), .Z(n7921) );
  AND U8586 ( .A(y[193]), .B(x[75]), .Z(n8031) );
  XOR U8587 ( .A(n7864), .B(n8031), .Z(n7920) );
  XOR U8588 ( .A(n7921), .B(n7920), .Z(n7894) );
  XOR U8589 ( .A(n7893), .B(n7894), .Z(n7895) );
  NANDN U8590 ( .A(n7866), .B(n7865), .Z(n7870) );
  OR U8591 ( .A(n7868), .B(n7867), .Z(n7869) );
  NAND U8592 ( .A(n7870), .B(n7869), .Z(n7896) );
  XOR U8593 ( .A(n7971), .B(n7970), .Z(n7966) );
  XOR U8594 ( .A(n7967), .B(n7966), .Z(n7883) );
  XNOR U8595 ( .A(n7884), .B(n7883), .Z(n7873) );
  XNOR U8596 ( .A(n7874), .B(n7873), .Z(o[76]) );
  NAND U8597 ( .A(n7876), .B(n7875), .Z(n7880) );
  NAND U8598 ( .A(n7878), .B(n7877), .Z(n7879) );
  NAND U8599 ( .A(n7880), .B(n7879), .Z(n8122) );
  XNOR U8600 ( .A(n8121), .B(n8122), .Z(n8124) );
  NANDN U8601 ( .A(n7882), .B(n7881), .Z(n7886) );
  NAND U8602 ( .A(n7884), .B(n7883), .Z(n7885) );
  AND U8603 ( .A(n7886), .B(n7885), .Z(n7979) );
  NAND U8604 ( .A(n7888), .B(n7887), .Z(n7892) );
  NAND U8605 ( .A(n7890), .B(n7889), .Z(n7891) );
  AND U8606 ( .A(n7892), .B(n7891), .Z(n8033) );
  NAND U8607 ( .A(n7894), .B(n7893), .Z(n7898) );
  NANDN U8608 ( .A(n7896), .B(n7895), .Z(n7897) );
  NAND U8609 ( .A(n7898), .B(n7897), .Z(n8032) );
  AND U8610 ( .A(y[114]), .B(x[59]), .Z(n8025) );
  NAND U8611 ( .A(n7899), .B(n8025), .Z(n7903) );
  NANDN U8612 ( .A(n7901), .B(n7900), .Z(n7902) );
  AND U8613 ( .A(n7903), .B(n7902), .Z(n7985) );
  NANDN U8614 ( .A(n7905), .B(n7904), .Z(n7909) );
  NANDN U8615 ( .A(n7907), .B(n7906), .Z(n7908) );
  NAND U8616 ( .A(n7909), .B(n7908), .Z(n8010) );
  AND U8617 ( .A(y[72]), .B(x[53]), .Z(n8015) );
  AND U8618 ( .A(y[115]), .B(x[58]), .Z(n8014) );
  XOR U8619 ( .A(n8015), .B(n8014), .Z(n8016) );
  AND U8620 ( .A(y[157]), .B(x[64]), .Z(n8181) );
  XOR U8621 ( .A(n8016), .B(n8181), .Z(n8009) );
  AND U8622 ( .A(y[153]), .B(x[68]), .Z(n8020) );
  AND U8623 ( .A(y[32]), .B(x[45]), .Z(n8019) );
  XOR U8624 ( .A(n8020), .B(n8019), .Z(n8021) );
  AND U8625 ( .A(y[33]), .B(x[44]), .Z(n8152) );
  XOR U8626 ( .A(n8021), .B(n8152), .Z(n8008) );
  XOR U8627 ( .A(n8009), .B(n8008), .Z(n8011) );
  XOR U8628 ( .A(n8010), .B(n8011), .Z(n7984) );
  NANDN U8629 ( .A(n7911), .B(n7910), .Z(n7915) );
  NANDN U8630 ( .A(n7913), .B(n7912), .Z(n7914) );
  NAND U8631 ( .A(n7915), .B(n7914), .Z(n8088) );
  AND U8632 ( .A(y[194]), .B(x[75]), .Z(n7933) );
  AND U8633 ( .A(n7916), .B(n7933), .Z(n8070) );
  AND U8634 ( .A(x[72]), .B(y[197]), .Z(n7918) );
  AND U8635 ( .A(x[73]), .B(y[196]), .Z(n7917) );
  XOR U8636 ( .A(n7918), .B(n7917), .Z(n8069) );
  XOR U8637 ( .A(n8070), .B(n8069), .Z(n8087) );
  AND U8638 ( .A(y[77]), .B(x[48]), .Z(n8095) );
  AND U8639 ( .A(y[36]), .B(x[41]), .Z(n8094) );
  XOR U8640 ( .A(n8095), .B(n8094), .Z(n8097) );
  AND U8641 ( .A(y[73]), .B(x[52]), .Z(n8096) );
  XOR U8642 ( .A(n8097), .B(n8096), .Z(n8086) );
  XOR U8643 ( .A(n8087), .B(n8086), .Z(n8089) );
  XOR U8644 ( .A(n8088), .B(n8089), .Z(n7986) );
  XOR U8645 ( .A(n7987), .B(n7986), .Z(n8034) );
  XOR U8646 ( .A(n8035), .B(n8034), .Z(n8119) );
  AND U8647 ( .A(y[195]), .B(x[76]), .Z(n8289) );
  NAND U8648 ( .A(n8289), .B(n7919), .Z(n7923) );
  NAND U8649 ( .A(n7921), .B(n7920), .Z(n7922) );
  AND U8650 ( .A(n7923), .B(n7922), .Z(n8045) );
  NAND U8651 ( .A(n7927), .B(n7926), .Z(n7931) );
  NANDN U8652 ( .A(n7929), .B(n7928), .Z(n7930) );
  AND U8653 ( .A(n7931), .B(n7930), .Z(n8053) );
  AND U8654 ( .A(y[74]), .B(x[51]), .Z(n8212) );
  NAND U8655 ( .A(x[50]), .B(y[75]), .Z(n7932) );
  XNOR U8656 ( .A(n8212), .B(n7932), .Z(n8004) );
  NAND U8657 ( .A(y[76]), .B(x[49]), .Z(n8005) );
  AND U8658 ( .A(y[195]), .B(x[74]), .Z(n7990) );
  NAND U8659 ( .A(y[192]), .B(x[77]), .Z(n7991) );
  NAND U8660 ( .A(y[193]), .B(x[76]), .Z(n8242) );
  XOR U8661 ( .A(n7933), .B(n8242), .Z(n7993) );
  XOR U8662 ( .A(n8051), .B(n8050), .Z(n8052) );
  XOR U8663 ( .A(n8053), .B(n8052), .Z(n8046) );
  XOR U8664 ( .A(n8047), .B(n8046), .Z(n8065) );
  AND U8665 ( .A(x[60]), .B(y[113]), .Z(n7935) );
  NAND U8666 ( .A(x[61]), .B(y[112]), .Z(n7934) );
  XOR U8667 ( .A(n7935), .B(n7934), .Z(n8026) );
  AND U8668 ( .A(y[152]), .B(x[69]), .Z(n7996) );
  NAND U8669 ( .A(y[34]), .B(x[43]), .Z(n7997) );
  AND U8670 ( .A(y[35]), .B(x[42]), .Z(n7998) );
  XOR U8671 ( .A(n7999), .B(n7998), .Z(n8104) );
  XOR U8672 ( .A(n8105), .B(n8104), .Z(n8107) );
  NAND U8673 ( .A(n7937), .B(n7936), .Z(n7941) );
  NANDN U8674 ( .A(n7939), .B(n7938), .Z(n7940) );
  AND U8675 ( .A(n7941), .B(n7940), .Z(n8106) );
  XOR U8676 ( .A(n8107), .B(n8106), .Z(n8063) );
  AND U8677 ( .A(y[76]), .B(x[51]), .Z(n8288) );
  NAND U8678 ( .A(n8288), .B(n7942), .Z(n7945) );
  NANDN U8679 ( .A(n7943), .B(n8003), .Z(n7944) );
  AND U8680 ( .A(n7945), .B(n7944), .Z(n8041) );
  AND U8681 ( .A(y[116]), .B(x[57]), .Z(n8237) );
  AND U8682 ( .A(y[154]), .B(x[67]), .Z(n8081) );
  XOR U8683 ( .A(n8237), .B(n8081), .Z(n8083) );
  AND U8684 ( .A(y[117]), .B(x[56]), .Z(n8082) );
  XOR U8685 ( .A(n8083), .B(n8082), .Z(n8039) );
  AND U8686 ( .A(y[37]), .B(x[40]), .Z(n8074) );
  AND U8687 ( .A(y[156]), .B(x[65]), .Z(n8073) );
  XOR U8688 ( .A(n8074), .B(n8073), .Z(n8076) );
  AND U8689 ( .A(y[155]), .B(x[66]), .Z(n8075) );
  XOR U8690 ( .A(n8076), .B(n8075), .Z(n8038) );
  XOR U8691 ( .A(n8039), .B(n8038), .Z(n8040) );
  XOR U8692 ( .A(n8041), .B(n8040), .Z(n8062) );
  NANDN U8693 ( .A(n7947), .B(n7946), .Z(n7951) );
  NANDN U8694 ( .A(n7949), .B(n7948), .Z(n7950) );
  AND U8695 ( .A(n7951), .B(n7950), .Z(n8059) );
  NANDN U8696 ( .A(n7953), .B(n7952), .Z(n7957) );
  NAND U8697 ( .A(n7955), .B(n7954), .Z(n7956) );
  AND U8698 ( .A(n7957), .B(n7956), .Z(n8057) );
  NAND U8699 ( .A(n7959), .B(n7958), .Z(n7963) );
  NANDN U8700 ( .A(n7961), .B(n7960), .Z(n7962) );
  NAND U8701 ( .A(n7963), .B(n7962), .Z(n8056) );
  XOR U8702 ( .A(n8059), .B(n8058), .Z(n8116) );
  XOR U8703 ( .A(n8117), .B(n8116), .Z(n8118) );
  XOR U8704 ( .A(n8119), .B(n8118), .Z(n7978) );
  XNOR U8705 ( .A(n7979), .B(n7978), .Z(n7980) );
  NANDN U8706 ( .A(n7973), .B(n7972), .Z(n7977) );
  NAND U8707 ( .A(n7975), .B(n7974), .Z(n7976) );
  AND U8708 ( .A(n7977), .B(n7976), .Z(n8110) );
  XNOR U8709 ( .A(n8111), .B(n8110), .Z(n8112) );
  XOR U8710 ( .A(n8113), .B(n8112), .Z(n7981) );
  XNOR U8711 ( .A(n7980), .B(n7981), .Z(n8123) );
  XOR U8712 ( .A(n8124), .B(n8123), .Z(o[77]) );
  NANDN U8713 ( .A(n7979), .B(n7978), .Z(n7983) );
  NANDN U8714 ( .A(n7981), .B(n7980), .Z(n7982) );
  AND U8715 ( .A(n7983), .B(n7982), .Z(n8408) );
  NANDN U8716 ( .A(n7985), .B(n7984), .Z(n7989) );
  NAND U8717 ( .A(n7987), .B(n7986), .Z(n7988) );
  AND U8718 ( .A(n7989), .B(n7988), .Z(n8412) );
  NANDN U8719 ( .A(n7991), .B(n7990), .Z(n7995) );
  NANDN U8720 ( .A(n7993), .B(n7992), .Z(n7994) );
  NAND U8721 ( .A(n7995), .B(n7994), .Z(n8348) );
  NANDN U8722 ( .A(n7997), .B(n7996), .Z(n8001) );
  NAND U8723 ( .A(n7999), .B(n7998), .Z(n8000) );
  NAND U8724 ( .A(n8001), .B(n8000), .Z(n8351) );
  AND U8725 ( .A(y[75]), .B(x[51]), .Z(n8002) );
  NAND U8726 ( .A(n8003), .B(n8002), .Z(n8007) );
  NANDN U8727 ( .A(n8005), .B(n8004), .Z(n8006) );
  AND U8728 ( .A(n8007), .B(n8006), .Z(n8216) );
  AND U8729 ( .A(y[155]), .B(x[67]), .Z(n8187) );
  AND U8730 ( .A(y[115]), .B(x[59]), .Z(n8186) );
  XOR U8731 ( .A(n8187), .B(n8186), .Z(n8185) );
  AND U8732 ( .A(y[35]), .B(x[43]), .Z(n8184) );
  XOR U8733 ( .A(n8185), .B(n8184), .Z(n8218) );
  AND U8734 ( .A(y[156]), .B(x[66]), .Z(n8158) );
  AND U8735 ( .A(y[114]), .B(x[60]), .Z(n8157) );
  XOR U8736 ( .A(n8158), .B(n8157), .Z(n8156) );
  AND U8737 ( .A(y[36]), .B(x[42]), .Z(n8155) );
  XNOR U8738 ( .A(n8156), .B(n8155), .Z(n8217) );
  XNOR U8739 ( .A(n8216), .B(n8215), .Z(n8350) );
  XOR U8740 ( .A(n8351), .B(n8350), .Z(n8349) );
  XOR U8741 ( .A(n8348), .B(n8349), .Z(n8137) );
  NAND U8742 ( .A(n8009), .B(n8008), .Z(n8013) );
  NAND U8743 ( .A(n8011), .B(n8010), .Z(n8012) );
  NAND U8744 ( .A(n8013), .B(n8012), .Z(n8136) );
  XOR U8745 ( .A(n8137), .B(n8136), .Z(n8135) );
  NAND U8746 ( .A(n8015), .B(n8014), .Z(n8018) );
  NAND U8747 ( .A(n8016), .B(n8181), .Z(n8017) );
  NAND U8748 ( .A(n8018), .B(n8017), .Z(n8335) );
  NAND U8749 ( .A(n8020), .B(n8019), .Z(n8023) );
  NAND U8750 ( .A(n8021), .B(n8152), .Z(n8022) );
  NAND U8751 ( .A(n8023), .B(n8022), .Z(n8334) );
  XOR U8752 ( .A(n8335), .B(n8334), .Z(n8333) );
  AND U8753 ( .A(y[113]), .B(x[61]), .Z(n8166) );
  NANDN U8754 ( .A(n8024), .B(n8166), .Z(n8028) );
  NANDN U8755 ( .A(n8026), .B(n8025), .Z(n8027) );
  AND U8756 ( .A(n8028), .B(n8027), .Z(n8361) );
  AND U8757 ( .A(x[45]), .B(y[33]), .Z(n8030) );
  NAND U8758 ( .A(x[44]), .B(y[34]), .Z(n8029) );
  XNOR U8759 ( .A(n8030), .B(n8029), .Z(n8151) );
  AND U8760 ( .A(y[152]), .B(x[70]), .Z(n8150) );
  XOR U8761 ( .A(n8151), .B(n8150), .Z(n8363) );
  AND U8762 ( .A(y[197]), .B(x[73]), .Z(n8230) );
  AND U8763 ( .A(y[194]), .B(x[76]), .Z(n8080) );
  AND U8764 ( .A(n8031), .B(n8080), .Z(n8228) );
  AND U8765 ( .A(y[196]), .B(x[74]), .Z(n8227) );
  XOR U8766 ( .A(n8228), .B(n8227), .Z(n8229) );
  XNOR U8767 ( .A(n8230), .B(n8229), .Z(n8362) );
  XNOR U8768 ( .A(n8361), .B(n8360), .Z(n8332) );
  XOR U8769 ( .A(n8333), .B(n8332), .Z(n8134) );
  XOR U8770 ( .A(n8135), .B(n8134), .Z(n8133) );
  NANDN U8771 ( .A(n8033), .B(n8032), .Z(n8037) );
  NAND U8772 ( .A(n8035), .B(n8034), .Z(n8036) );
  AND U8773 ( .A(n8037), .B(n8036), .Z(n8132) );
  NAND U8774 ( .A(n8039), .B(n8038), .Z(n8043) );
  NANDN U8775 ( .A(n8041), .B(n8040), .Z(n8042) );
  AND U8776 ( .A(n8043), .B(n8042), .Z(n8377) );
  NANDN U8777 ( .A(n8045), .B(n8044), .Z(n8049) );
  NAND U8778 ( .A(n8047), .B(n8046), .Z(n8048) );
  AND U8779 ( .A(n8049), .B(n8048), .Z(n8376) );
  XOR U8780 ( .A(n8377), .B(n8376), .Z(n8375) );
  NAND U8781 ( .A(n8051), .B(n8050), .Z(n8055) );
  NAND U8782 ( .A(n8053), .B(n8052), .Z(n8054) );
  AND U8783 ( .A(n8055), .B(n8054), .Z(n8374) );
  XOR U8784 ( .A(n8375), .B(n8374), .Z(n8130) );
  XOR U8785 ( .A(n8131), .B(n8130), .Z(n8411) );
  XOR U8786 ( .A(n8412), .B(n8411), .Z(n8414) );
  NANDN U8787 ( .A(n8057), .B(n8056), .Z(n8061) );
  NAND U8788 ( .A(n8059), .B(n8058), .Z(n8060) );
  AND U8789 ( .A(n8061), .B(n8060), .Z(n8391) );
  NANDN U8790 ( .A(n8063), .B(n8062), .Z(n8067) );
  NANDN U8791 ( .A(n8065), .B(n8064), .Z(n8066) );
  NAND U8792 ( .A(n8067), .B(n8066), .Z(n8392) );
  NANDN U8793 ( .A(n8068), .B(n8230), .Z(n8072) );
  NAND U8794 ( .A(n8070), .B(n8069), .Z(n8071) );
  NAND U8795 ( .A(n8072), .B(n8071), .Z(n8329) );
  NAND U8796 ( .A(n8074), .B(n8073), .Z(n8078) );
  NAND U8797 ( .A(n8076), .B(n8075), .Z(n8077) );
  AND U8798 ( .A(n8078), .B(n8077), .Z(n8355) );
  AND U8799 ( .A(y[37]), .B(x[41]), .Z(n8172) );
  AND U8800 ( .A(y[72]), .B(x[54]), .Z(n8171) );
  XOR U8801 ( .A(n8172), .B(n8171), .Z(n8170) );
  AND U8802 ( .A(y[78]), .B(x[48]), .Z(n8169) );
  XOR U8803 ( .A(n8170), .B(n8169), .Z(n8357) );
  NAND U8804 ( .A(x[77]), .B(y[193]), .Z(n8079) );
  XNOR U8805 ( .A(n8080), .B(n8079), .Z(n8224) );
  AND U8806 ( .A(y[192]), .B(x[78]), .Z(n8223) );
  XOR U8807 ( .A(n8224), .B(n8223), .Z(n8221) );
  XNOR U8808 ( .A(n8222), .B(n8221), .Z(n8356) );
  XNOR U8809 ( .A(n8355), .B(n8354), .Z(n8328) );
  XOR U8810 ( .A(n8329), .B(n8328), .Z(n8327) );
  AND U8811 ( .A(n8237), .B(n8081), .Z(n8085) );
  NAND U8812 ( .A(n8083), .B(n8082), .Z(n8084) );
  NANDN U8813 ( .A(n8085), .B(n8084), .Z(n8326) );
  XOR U8814 ( .A(n8327), .B(n8326), .Z(n8399) );
  NAND U8815 ( .A(n8087), .B(n8086), .Z(n8091) );
  NAND U8816 ( .A(n8089), .B(n8088), .Z(n8090) );
  AND U8817 ( .A(n8091), .B(n8090), .Z(n8138) );
  AND U8818 ( .A(y[118]), .B(x[56]), .Z(n8201) );
  AND U8819 ( .A(y[32]), .B(x[46]), .Z(n8200) );
  XOR U8820 ( .A(n8201), .B(n8200), .Z(n8199) );
  AND U8821 ( .A(y[153]), .B(x[69]), .Z(n8198) );
  XOR U8822 ( .A(n8199), .B(n8198), .Z(n8371) );
  AND U8823 ( .A(y[73]), .B(x[53]), .Z(n8195) );
  AND U8824 ( .A(y[76]), .B(x[50]), .Z(n8194) );
  XOR U8825 ( .A(n8195), .B(n8194), .Z(n8193) );
  AND U8826 ( .A(y[77]), .B(x[49]), .Z(n8192) );
  XOR U8827 ( .A(n8193), .B(n8192), .Z(n8211) );
  AND U8828 ( .A(x[52]), .B(y[74]), .Z(n8093) );
  NAND U8829 ( .A(x[51]), .B(y[75]), .Z(n8092) );
  XNOR U8830 ( .A(n8093), .B(n8092), .Z(n8210) );
  XOR U8831 ( .A(n8211), .B(n8210), .Z(n8370) );
  XOR U8832 ( .A(n8371), .B(n8370), .Z(n8369) );
  AND U8833 ( .A(y[198]), .B(x[72]), .Z(n8165) );
  XOR U8834 ( .A(n8166), .B(n8165), .Z(n8164) );
  AND U8835 ( .A(y[112]), .B(x[62]), .Z(n8163) );
  XOR U8836 ( .A(n8164), .B(n8163), .Z(n8368) );
  XOR U8837 ( .A(n8369), .B(n8368), .Z(n8141) );
  NAND U8838 ( .A(n8095), .B(n8094), .Z(n8099) );
  NAND U8839 ( .A(n8097), .B(n8096), .Z(n8098) );
  AND U8840 ( .A(n8099), .B(n8098), .Z(n8145) );
  AND U8841 ( .A(y[154]), .B(x[68]), .Z(n8236) );
  AND U8842 ( .A(x[57]), .B(y[117]), .Z(n8101) );
  AND U8843 ( .A(x[58]), .B(y[116]), .Z(n8100) );
  XOR U8844 ( .A(n8101), .B(n8100), .Z(n8235) );
  XOR U8845 ( .A(n8236), .B(n8235), .Z(n8147) );
  AND U8846 ( .A(y[38]), .B(x[40]), .Z(n8180) );
  AND U8847 ( .A(x[64]), .B(y[158]), .Z(n8103) );
  NAND U8848 ( .A(x[65]), .B(y[157]), .Z(n8102) );
  XNOR U8849 ( .A(n8103), .B(n8102), .Z(n8179) );
  XNOR U8850 ( .A(n8180), .B(n8179), .Z(n8146) );
  XOR U8851 ( .A(n8145), .B(n8144), .Z(n8140) );
  XNOR U8852 ( .A(n8138), .B(n8139), .Z(n8398) );
  NAND U8853 ( .A(n8105), .B(n8104), .Z(n8109) );
  NAND U8854 ( .A(n8107), .B(n8106), .Z(n8108) );
  AND U8855 ( .A(n8109), .B(n8108), .Z(n8396) );
  XOR U8856 ( .A(n8397), .B(n8396), .Z(n8393) );
  XOR U8857 ( .A(n8392), .B(n8393), .Z(n8390) );
  XOR U8858 ( .A(n8391), .B(n8390), .Z(n8413) );
  XOR U8859 ( .A(n8414), .B(n8413), .Z(n8129) );
  NANDN U8860 ( .A(n8111), .B(n8110), .Z(n8115) );
  NANDN U8861 ( .A(n8113), .B(n8112), .Z(n8114) );
  AND U8862 ( .A(n8115), .B(n8114), .Z(n8128) );
  XOR U8863 ( .A(n8128), .B(n8127), .Z(n8120) );
  XOR U8864 ( .A(n8129), .B(n8120), .Z(n8407) );
  NANDN U8865 ( .A(n8122), .B(n8121), .Z(n8126) );
  NAND U8866 ( .A(n8124), .B(n8123), .Z(n8125) );
  NAND U8867 ( .A(n8126), .B(n8125), .Z(n8405) );
  XOR U8868 ( .A(n8406), .B(n8405), .Z(o[78]) );
  NANDN U8869 ( .A(n8139), .B(n8138), .Z(n8143) );
  NANDN U8870 ( .A(n8141), .B(n8140), .Z(n8142) );
  AND U8871 ( .A(n8143), .B(n8142), .Z(n8389) );
  NAND U8872 ( .A(n8145), .B(n8144), .Z(n8149) );
  NANDN U8873 ( .A(n8147), .B(n8146), .Z(n8148) );
  AND U8874 ( .A(n8149), .B(n8148), .Z(n8347) );
  NAND U8875 ( .A(n8151), .B(n8150), .Z(n8154) );
  AND U8876 ( .A(y[34]), .B(x[45]), .Z(n8287) );
  NAND U8877 ( .A(n8152), .B(n8287), .Z(n8153) );
  AND U8878 ( .A(n8154), .B(n8153), .Z(n8162) );
  NAND U8879 ( .A(n8156), .B(n8155), .Z(n8160) );
  NAND U8880 ( .A(n8158), .B(n8157), .Z(n8159) );
  NAND U8881 ( .A(n8160), .B(n8159), .Z(n8161) );
  XNOR U8882 ( .A(n8162), .B(n8161), .Z(n8178) );
  NAND U8883 ( .A(n8164), .B(n8163), .Z(n8168) );
  NAND U8884 ( .A(n8166), .B(n8165), .Z(n8167) );
  AND U8885 ( .A(n8168), .B(n8167), .Z(n8176) );
  NAND U8886 ( .A(n8170), .B(n8169), .Z(n8174) );
  NAND U8887 ( .A(n8172), .B(n8171), .Z(n8173) );
  NAND U8888 ( .A(n8174), .B(n8173), .Z(n8175) );
  XNOR U8889 ( .A(n8176), .B(n8175), .Z(n8177) );
  XOR U8890 ( .A(n8178), .B(n8177), .Z(n8209) );
  NAND U8891 ( .A(n8180), .B(n8179), .Z(n8183) );
  AND U8892 ( .A(y[158]), .B(x[65]), .Z(n8292) );
  NAND U8893 ( .A(n8181), .B(n8292), .Z(n8182) );
  AND U8894 ( .A(n8183), .B(n8182), .Z(n8191) );
  NAND U8895 ( .A(n8185), .B(n8184), .Z(n8189) );
  NAND U8896 ( .A(n8187), .B(n8186), .Z(n8188) );
  NAND U8897 ( .A(n8189), .B(n8188), .Z(n8190) );
  XNOR U8898 ( .A(n8191), .B(n8190), .Z(n8207) );
  NAND U8899 ( .A(n8193), .B(n8192), .Z(n8197) );
  NAND U8900 ( .A(n8195), .B(n8194), .Z(n8196) );
  AND U8901 ( .A(n8197), .B(n8196), .Z(n8205) );
  NAND U8902 ( .A(n8199), .B(n8198), .Z(n8203) );
  NAND U8903 ( .A(n8201), .B(n8200), .Z(n8202) );
  NAND U8904 ( .A(n8203), .B(n8202), .Z(n8204) );
  XNOR U8905 ( .A(n8205), .B(n8204), .Z(n8206) );
  XNOR U8906 ( .A(n8207), .B(n8206), .Z(n8208) );
  XNOR U8907 ( .A(n8209), .B(n8208), .Z(n8345) );
  NAND U8908 ( .A(n8211), .B(n8210), .Z(n8214) );
  AND U8909 ( .A(y[75]), .B(x[52]), .Z(n8286) );
  NAND U8910 ( .A(n8212), .B(n8286), .Z(n8213) );
  AND U8911 ( .A(n8214), .B(n8213), .Z(n8343) );
  NAND U8912 ( .A(n8216), .B(n8215), .Z(n8220) );
  NANDN U8913 ( .A(n8218), .B(n8217), .Z(n8219) );
  AND U8914 ( .A(n8220), .B(n8219), .Z(n8325) );
  NAND U8915 ( .A(n8222), .B(n8221), .Z(n8226) );
  AND U8916 ( .A(n8224), .B(n8223), .Z(n8225) );
  ANDN U8917 ( .B(n8226), .A(n8225), .Z(n8234) );
  AND U8918 ( .A(n8228), .B(n8227), .Z(n8232) );
  AND U8919 ( .A(n8230), .B(n8229), .Z(n8231) );
  OR U8920 ( .A(n8232), .B(n8231), .Z(n8233) );
  XNOR U8921 ( .A(n8234), .B(n8233), .Z(n8323) );
  NAND U8922 ( .A(n8236), .B(n8235), .Z(n8239) );
  AND U8923 ( .A(y[117]), .B(x[58]), .Z(n8293) );
  NAND U8924 ( .A(n8237), .B(n8293), .Z(n8238) );
  AND U8925 ( .A(n8239), .B(n8238), .Z(n8321) );
  AND U8926 ( .A(x[49]), .B(y[78]), .Z(n8241) );
  NAND U8927 ( .A(x[55]), .B(y[72]), .Z(n8240) );
  XNOR U8928 ( .A(n8241), .B(n8240), .Z(n8247) );
  AND U8929 ( .A(x[64]), .B(y[159]), .Z(n8245) );
  AND U8930 ( .A(x[77]), .B(n8242), .Z(n8243) );
  NAND U8931 ( .A(n8243), .B(y[194]), .Z(n8244) );
  XNOR U8932 ( .A(n8245), .B(n8244), .Z(n8246) );
  XOR U8933 ( .A(n8247), .B(n8246), .Z(n8255) );
  AND U8934 ( .A(x[73]), .B(y[198]), .Z(n8249) );
  NAND U8935 ( .A(x[53]), .B(y[74]), .Z(n8248) );
  XNOR U8936 ( .A(n8249), .B(n8248), .Z(n8253) );
  AND U8937 ( .A(x[50]), .B(y[77]), .Z(n8251) );
  NAND U8938 ( .A(x[66]), .B(y[157]), .Z(n8250) );
  XNOR U8939 ( .A(n8251), .B(n8250), .Z(n8252) );
  XNOR U8940 ( .A(n8253), .B(n8252), .Z(n8254) );
  XNOR U8941 ( .A(n8255), .B(n8254), .Z(n8319) );
  AND U8942 ( .A(x[40]), .B(y[39]), .Z(n8257) );
  NAND U8943 ( .A(x[63]), .B(y[112]), .Z(n8256) );
  XNOR U8944 ( .A(n8257), .B(n8256), .Z(n8261) );
  AND U8945 ( .A(x[72]), .B(y[199]), .Z(n8259) );
  NAND U8946 ( .A(x[69]), .B(y[154]), .Z(n8258) );
  XNOR U8947 ( .A(n8259), .B(n8258), .Z(n8260) );
  XOR U8948 ( .A(n8261), .B(n8260), .Z(n8269) );
  AND U8949 ( .A(x[41]), .B(y[38]), .Z(n8263) );
  NAND U8950 ( .A(x[61]), .B(y[114]), .Z(n8262) );
  XNOR U8951 ( .A(n8263), .B(n8262), .Z(n8267) );
  AND U8952 ( .A(x[42]), .B(y[37]), .Z(n8265) );
  NAND U8953 ( .A(x[70]), .B(y[153]), .Z(n8264) );
  XNOR U8954 ( .A(n8265), .B(n8264), .Z(n8266) );
  XNOR U8955 ( .A(n8267), .B(n8266), .Z(n8268) );
  XNOR U8956 ( .A(n8269), .B(n8268), .Z(n8285) );
  AND U8957 ( .A(x[43]), .B(y[36]), .Z(n8271) );
  NAND U8958 ( .A(x[54]), .B(y[73]), .Z(n8270) );
  XNOR U8959 ( .A(n8271), .B(n8270), .Z(n8275) );
  AND U8960 ( .A(x[57]), .B(y[118]), .Z(n8273) );
  NAND U8961 ( .A(x[60]), .B(y[115]), .Z(n8272) );
  XNOR U8962 ( .A(n8273), .B(n8272), .Z(n8274) );
  XOR U8963 ( .A(n8275), .B(n8274), .Z(n8283) );
  AND U8964 ( .A(x[59]), .B(y[116]), .Z(n8277) );
  NAND U8965 ( .A(x[78]), .B(y[193]), .Z(n8276) );
  XNOR U8966 ( .A(n8277), .B(n8276), .Z(n8281) );
  AND U8967 ( .A(x[79]), .B(y[192]), .Z(n8279) );
  NAND U8968 ( .A(x[62]), .B(y[113]), .Z(n8278) );
  XNOR U8969 ( .A(n8279), .B(n8278), .Z(n8280) );
  XNOR U8970 ( .A(n8281), .B(n8280), .Z(n8282) );
  XNOR U8971 ( .A(n8283), .B(n8282), .Z(n8284) );
  XOR U8972 ( .A(n8285), .B(n8284), .Z(n8317) );
  XOR U8973 ( .A(n8287), .B(n8286), .Z(n8291) );
  XNOR U8974 ( .A(n8289), .B(n8288), .Z(n8290) );
  XNOR U8975 ( .A(n8291), .B(n8290), .Z(n8315) );
  AND U8976 ( .A(x[71]), .B(y[152]), .Z(n8313) );
  AND U8977 ( .A(x[56]), .B(y[119]), .Z(n8295) );
  XNOR U8978 ( .A(n8293), .B(n8292), .Z(n8294) );
  XNOR U8979 ( .A(n8295), .B(n8294), .Z(n8311) );
  AND U8980 ( .A(x[47]), .B(y[32]), .Z(n8297) );
  NAND U8981 ( .A(x[46]), .B(y[33]), .Z(n8296) );
  XNOR U8982 ( .A(n8297), .B(n8296), .Z(n8301) );
  AND U8983 ( .A(x[75]), .B(y[196]), .Z(n8299) );
  NAND U8984 ( .A(x[68]), .B(y[155]), .Z(n8298) );
  XNOR U8985 ( .A(n8299), .B(n8298), .Z(n8300) );
  XOR U8986 ( .A(n8301), .B(n8300), .Z(n8309) );
  AND U8987 ( .A(x[74]), .B(y[197]), .Z(n8303) );
  NAND U8988 ( .A(x[44]), .B(y[35]), .Z(n8302) );
  XNOR U8989 ( .A(n8303), .B(n8302), .Z(n8307) );
  AND U8990 ( .A(x[48]), .B(y[79]), .Z(n8305) );
  NAND U8991 ( .A(x[67]), .B(y[156]), .Z(n8304) );
  XNOR U8992 ( .A(n8305), .B(n8304), .Z(n8306) );
  XNOR U8993 ( .A(n8307), .B(n8306), .Z(n8308) );
  XNOR U8994 ( .A(n8309), .B(n8308), .Z(n8310) );
  XNOR U8995 ( .A(n8311), .B(n8310), .Z(n8312) );
  XNOR U8996 ( .A(n8313), .B(n8312), .Z(n8314) );
  XNOR U8997 ( .A(n8315), .B(n8314), .Z(n8316) );
  XNOR U8998 ( .A(n8317), .B(n8316), .Z(n8318) );
  XNOR U8999 ( .A(n8319), .B(n8318), .Z(n8320) );
  XNOR U9000 ( .A(n8321), .B(n8320), .Z(n8322) );
  XNOR U9001 ( .A(n8323), .B(n8322), .Z(n8324) );
  XNOR U9002 ( .A(n8325), .B(n8324), .Z(n8341) );
  NAND U9003 ( .A(n8327), .B(n8326), .Z(n8331) );
  NAND U9004 ( .A(n8329), .B(n8328), .Z(n8330) );
  AND U9005 ( .A(n8331), .B(n8330), .Z(n8339) );
  NAND U9006 ( .A(n8333), .B(n8332), .Z(n8337) );
  NAND U9007 ( .A(n8335), .B(n8334), .Z(n8336) );
  NAND U9008 ( .A(n8337), .B(n8336), .Z(n8338) );
  XNOR U9009 ( .A(n8339), .B(n8338), .Z(n8340) );
  XNOR U9010 ( .A(n8341), .B(n8340), .Z(n8342) );
  XNOR U9011 ( .A(n8343), .B(n8342), .Z(n8344) );
  XNOR U9012 ( .A(n8345), .B(n8344), .Z(n8346) );
  XNOR U9013 ( .A(n8347), .B(n8346), .Z(n8387) );
  NAND U9014 ( .A(n8349), .B(n8348), .Z(n8353) );
  NAND U9015 ( .A(n8351), .B(n8350), .Z(n8352) );
  AND U9016 ( .A(n8353), .B(n8352), .Z(n8385) );
  NAND U9017 ( .A(n8355), .B(n8354), .Z(n8359) );
  NANDN U9018 ( .A(n8357), .B(n8356), .Z(n8358) );
  AND U9019 ( .A(n8359), .B(n8358), .Z(n8367) );
  NAND U9020 ( .A(n8361), .B(n8360), .Z(n8365) );
  NANDN U9021 ( .A(n8363), .B(n8362), .Z(n8364) );
  NAND U9022 ( .A(n8365), .B(n8364), .Z(n8366) );
  XNOR U9023 ( .A(n8367), .B(n8366), .Z(n8383) );
  NAND U9024 ( .A(n8369), .B(n8368), .Z(n8373) );
  NAND U9025 ( .A(n8371), .B(n8370), .Z(n8372) );
  AND U9026 ( .A(n8373), .B(n8372), .Z(n8381) );
  NAND U9027 ( .A(n8375), .B(n8374), .Z(n8379) );
  NAND U9028 ( .A(n8377), .B(n8376), .Z(n8378) );
  NAND U9029 ( .A(n8379), .B(n8378), .Z(n8380) );
  XNOR U9030 ( .A(n8381), .B(n8380), .Z(n8382) );
  XNOR U9031 ( .A(n8383), .B(n8382), .Z(n8384) );
  XNOR U9032 ( .A(n8385), .B(n8384), .Z(n8386) );
  XNOR U9033 ( .A(n8387), .B(n8386), .Z(n8388) );
  NAND U9034 ( .A(n8391), .B(n8390), .Z(n8395) );
  NAND U9035 ( .A(n8393), .B(n8392), .Z(n8394) );
  AND U9036 ( .A(n8395), .B(n8394), .Z(n8403) );
  NAND U9037 ( .A(n8397), .B(n8396), .Z(n8401) );
  NANDN U9038 ( .A(n8399), .B(n8398), .Z(n8400) );
  NAND U9039 ( .A(n8401), .B(n8400), .Z(n8402) );
  XNOR U9040 ( .A(n8403), .B(n8402), .Z(n8404) );
  NAND U9041 ( .A(n8406), .B(n8405), .Z(n8410) );
  NANDN U9042 ( .A(n8408), .B(n8407), .Z(n8409) );
  AND U9043 ( .A(n8412), .B(n8411), .Z(n8416) );
  AND U9044 ( .A(n8414), .B(n8413), .Z(n8415) );
  NAND U9045 ( .A(y[160]), .B(x[112]), .Z(n8555) );
  NAND U9046 ( .A(y[40]), .B(x[88]), .Z(n8419) );
  XOR U9047 ( .A(n8555), .B(n8419), .Z(n8420) );
  AND U9048 ( .A(y[0]), .B(x[80]), .Z(n8427) );
  AND U9049 ( .A(y[80]), .B(x[96]), .Z(n8424) );
  XOR U9050 ( .A(n8427), .B(n8424), .Z(n8423) );
  AND U9051 ( .A(y[120]), .B(x[104]), .Z(n8422) );
  XNOR U9052 ( .A(n8423), .B(n8422), .Z(n8421) );
  XNOR U9053 ( .A(n8420), .B(n8421), .Z(o[80]) );
  AND U9054 ( .A(x[80]), .B(y[1]), .Z(n8418) );
  NAND U9055 ( .A(x[81]), .B(y[0]), .Z(n8417) );
  XNOR U9056 ( .A(n8418), .B(n8417), .Z(n8429) );
  AND U9057 ( .A(y[40]), .B(x[89]), .Z(n8428) );
  XOR U9058 ( .A(n8429), .B(n8428), .Z(n8446) );
  AND U9059 ( .A(y[160]), .B(x[113]), .Z(n8658) );
  NAND U9060 ( .A(y[81]), .B(x[96]), .Z(n8432) );
  XNOR U9061 ( .A(n8658), .B(n8432), .Z(n8434) );
  AND U9062 ( .A(y[161]), .B(x[112]), .Z(n8456) );
  NAND U9063 ( .A(y[80]), .B(x[97]), .Z(n8455) );
  XNOR U9064 ( .A(n8456), .B(n8455), .Z(n8433) );
  XOR U9065 ( .A(n8434), .B(n8433), .Z(n8444) );
  AND U9066 ( .A(y[41]), .B(x[88]), .Z(n8682) );
  AND U9067 ( .A(y[121]), .B(x[104]), .Z(n8449) );
  XOR U9068 ( .A(n8682), .B(n8449), .Z(n8451) );
  AND U9069 ( .A(y[120]), .B(x[105]), .Z(n8450) );
  XNOR U9070 ( .A(n8451), .B(n8450), .Z(n8443) );
  XNOR U9071 ( .A(n8444), .B(n8443), .Z(n8445) );
  XNOR U9072 ( .A(n8446), .B(n8445), .Z(n8440) );
  NAND U9073 ( .A(n8423), .B(n8422), .Z(n8426) );
  AND U9074 ( .A(n8427), .B(n8424), .Z(n8425) );
  ANDN U9075 ( .B(n8426), .A(n8425), .Z(n8437) );
  XNOR U9076 ( .A(n8438), .B(n8437), .Z(n8439) );
  XNOR U9077 ( .A(n8440), .B(n8439), .Z(o[81]) );
  NAND U9078 ( .A(y[1]), .B(x[81]), .Z(n8478) );
  NANDN U9079 ( .A(n8478), .B(n8427), .Z(n8431) );
  NAND U9080 ( .A(n8429), .B(n8428), .Z(n8430) );
  AND U9081 ( .A(n8431), .B(n8430), .Z(n8513) );
  NANDN U9082 ( .A(n8432), .B(n8658), .Z(n8436) );
  NAND U9083 ( .A(n8434), .B(n8433), .Z(n8435) );
  AND U9084 ( .A(n8436), .B(n8435), .Z(n8512) );
  AND U9085 ( .A(y[122]), .B(x[104]), .Z(n8497) );
  NAND U9086 ( .A(y[2]), .B(x[80]), .Z(n8498) );
  XNOR U9087 ( .A(n8497), .B(n8498), .Z(n8499) );
  NAND U9088 ( .A(y[40]), .B(x[90]), .Z(n8500) );
  XNOR U9089 ( .A(n8499), .B(n8500), .Z(n8511) );
  XOR U9090 ( .A(n8512), .B(n8511), .Z(n8514) );
  XOR U9091 ( .A(n8513), .B(n8514), .Z(n8458) );
  NANDN U9092 ( .A(n8438), .B(n8437), .Z(n8442) );
  NAND U9093 ( .A(n8440), .B(n8439), .Z(n8441) );
  NAND U9094 ( .A(n8442), .B(n8441), .Z(n8457) );
  XNOR U9095 ( .A(n8458), .B(n8457), .Z(n8460) );
  NANDN U9096 ( .A(n8444), .B(n8443), .Z(n8448) );
  NANDN U9097 ( .A(n8446), .B(n8445), .Z(n8447) );
  AND U9098 ( .A(n8448), .B(n8447), .Z(n8466) );
  AND U9099 ( .A(y[0]), .B(x[82]), .Z(n8475) );
  NAND U9100 ( .A(y[82]), .B(x[96]), .Z(n8476) );
  XNOR U9101 ( .A(n8475), .B(n8476), .Z(n8477) );
  NAND U9102 ( .A(y[120]), .B(x[106]), .Z(n8506) );
  XNOR U9103 ( .A(n8505), .B(n8506), .Z(n8507) );
  AND U9104 ( .A(y[80]), .B(x[98]), .Z(n8585) );
  AND U9105 ( .A(y[162]), .B(x[112]), .Z(n8488) );
  XOR U9106 ( .A(n8585), .B(n8488), .Z(n8490) );
  NAND U9107 ( .A(y[81]), .B(x[97]), .Z(n8489) );
  XOR U9108 ( .A(n8490), .B(n8489), .Z(n8508) );
  XNOR U9109 ( .A(n8507), .B(n8508), .Z(n8463) );
  NAND U9110 ( .A(n8682), .B(n8449), .Z(n8453) );
  AND U9111 ( .A(n8451), .B(n8450), .Z(n8452) );
  ANDN U9112 ( .B(n8453), .A(n8452), .Z(n8472) );
  AND U9113 ( .A(x[113]), .B(y[161]), .Z(n8560) );
  NAND U9114 ( .A(x[114]), .B(y[160]), .Z(n8454) );
  XNOR U9115 ( .A(n8560), .B(n8454), .Z(n8504) );
  ANDN U9116 ( .B(n8456), .A(n8455), .Z(n8503) );
  XOR U9117 ( .A(n8504), .B(n8503), .Z(n8469) );
  AND U9118 ( .A(y[121]), .B(x[105]), .Z(n8481) );
  NAND U9119 ( .A(y[41]), .B(x[89]), .Z(n8482) );
  XNOR U9120 ( .A(n8481), .B(n8482), .Z(n8483) );
  NAND U9121 ( .A(y[42]), .B(x[88]), .Z(n8484) );
  XOR U9122 ( .A(n8483), .B(n8484), .Z(n8470) );
  XNOR U9123 ( .A(n8469), .B(n8470), .Z(n8471) );
  XOR U9124 ( .A(n8472), .B(n8471), .Z(n8464) );
  XNOR U9125 ( .A(n8463), .B(n8464), .Z(n8465) );
  XNOR U9126 ( .A(n8466), .B(n8465), .Z(n8459) );
  XNOR U9127 ( .A(n8460), .B(n8459), .Z(o[82]) );
  NANDN U9128 ( .A(n8458), .B(n8457), .Z(n8462) );
  NAND U9129 ( .A(n8460), .B(n8459), .Z(n8461) );
  AND U9130 ( .A(n8462), .B(n8461), .Z(n8535) );
  NANDN U9131 ( .A(n8464), .B(n8463), .Z(n8468) );
  NAND U9132 ( .A(n8466), .B(n8465), .Z(n8467) );
  AND U9133 ( .A(n8468), .B(n8467), .Z(n8532) );
  NANDN U9134 ( .A(n8470), .B(n8469), .Z(n8474) );
  NANDN U9135 ( .A(n8472), .B(n8471), .Z(n8473) );
  AND U9136 ( .A(n8474), .B(n8473), .Z(n8530) );
  NANDN U9137 ( .A(n8476), .B(n8475), .Z(n8480) );
  NANDN U9138 ( .A(n8478), .B(n8477), .Z(n8479) );
  AND U9139 ( .A(n8480), .B(n8479), .Z(n8524) );
  NANDN U9140 ( .A(n8482), .B(n8481), .Z(n8486) );
  NANDN U9141 ( .A(n8484), .B(n8483), .Z(n8485) );
  AND U9142 ( .A(n8486), .B(n8485), .Z(n8576) );
  AND U9143 ( .A(y[123]), .B(x[104]), .Z(n8604) );
  AND U9144 ( .A(y[83]), .B(x[96]), .Z(n8603) );
  NAND U9145 ( .A(y[0]), .B(x[83]), .Z(n8602) );
  XOR U9146 ( .A(n8603), .B(n8602), .Z(n8605) );
  XOR U9147 ( .A(n8604), .B(n8605), .Z(n8574) );
  AND U9148 ( .A(x[98]), .B(y[81]), .Z(n8638) );
  NAND U9149 ( .A(x[99]), .B(y[80]), .Z(n8487) );
  XNOR U9150 ( .A(n8638), .B(n8487), .Z(n8587) );
  NAND U9151 ( .A(y[82]), .B(x[97]), .Z(n8588) );
  XNOR U9152 ( .A(n8574), .B(n8573), .Z(n8575) );
  XNOR U9153 ( .A(n8576), .B(n8575), .Z(n8523) );
  XNOR U9154 ( .A(n8524), .B(n8523), .Z(n8525) );
  NAND U9155 ( .A(n8585), .B(n8488), .Z(n8492) );
  ANDN U9156 ( .B(n8490), .A(n8489), .Z(n8491) );
  ANDN U9157 ( .B(n8492), .A(n8491), .Z(n8582) );
  AND U9158 ( .A(y[2]), .B(x[81]), .Z(n8551) );
  AND U9159 ( .A(y[1]), .B(x[82]), .Z(n8550) );
  NAND U9160 ( .A(y[122]), .B(x[105]), .Z(n8549) );
  XOR U9161 ( .A(n8550), .B(n8549), .Z(n8552) );
  XOR U9162 ( .A(n8551), .B(n8552), .Z(n8580) );
  AND U9163 ( .A(x[115]), .B(y[160]), .Z(n8494) );
  NAND U9164 ( .A(x[112]), .B(y[163]), .Z(n8493) );
  XNOR U9165 ( .A(n8494), .B(n8493), .Z(n8556) );
  AND U9166 ( .A(x[113]), .B(y[162]), .Z(n8496) );
  NAND U9167 ( .A(x[114]), .B(y[161]), .Z(n8495) );
  XOR U9168 ( .A(n8496), .B(n8495), .Z(n8557) );
  XNOR U9169 ( .A(n8556), .B(n8557), .Z(n8579) );
  XNOR U9170 ( .A(n8580), .B(n8579), .Z(n8581) );
  XOR U9171 ( .A(n8582), .B(n8581), .Z(n8526) );
  XNOR U9172 ( .A(n8525), .B(n8526), .Z(n8529) );
  XNOR U9173 ( .A(n8530), .B(n8529), .Z(n8531) );
  XOR U9174 ( .A(n8532), .B(n8531), .Z(n8536) );
  XNOR U9175 ( .A(n8535), .B(n8536), .Z(n8538) );
  NANDN U9176 ( .A(n8498), .B(n8497), .Z(n8502) );
  NANDN U9177 ( .A(n8500), .B(n8499), .Z(n8501) );
  AND U9178 ( .A(n8502), .B(n8501), .Z(n8542) );
  AND U9179 ( .A(y[161]), .B(x[114]), .Z(n8655) );
  XNOR U9180 ( .A(n8542), .B(n8541), .Z(n8544) );
  AND U9181 ( .A(y[40]), .B(x[91]), .Z(n8595) );
  AND U9182 ( .A(y[3]), .B(x[80]), .Z(n8594) );
  NAND U9183 ( .A(y[121]), .B(x[106]), .Z(n8593) );
  XOR U9184 ( .A(n8594), .B(n8593), .Z(n8596) );
  XOR U9185 ( .A(n8595), .B(n8596), .Z(n8570) );
  AND U9186 ( .A(y[43]), .B(x[88]), .Z(n8563) );
  AND U9187 ( .A(y[41]), .B(x[90]), .Z(n8562) );
  NAND U9188 ( .A(y[120]), .B(x[107]), .Z(n8561) );
  XOR U9189 ( .A(n8562), .B(n8561), .Z(n8564) );
  XOR U9190 ( .A(n8563), .B(n8564), .Z(n8568) );
  AND U9191 ( .A(y[42]), .B(x[89]), .Z(n8567) );
  XOR U9192 ( .A(n8544), .B(n8543), .Z(n8518) );
  NANDN U9193 ( .A(n8506), .B(n8505), .Z(n8510) );
  NANDN U9194 ( .A(n8508), .B(n8507), .Z(n8509) );
  AND U9195 ( .A(n8510), .B(n8509), .Z(n8517) );
  XNOR U9196 ( .A(n8518), .B(n8517), .Z(n8520) );
  NANDN U9197 ( .A(n8512), .B(n8511), .Z(n8516) );
  OR U9198 ( .A(n8514), .B(n8513), .Z(n8515) );
  AND U9199 ( .A(n8516), .B(n8515), .Z(n8519) );
  XNOR U9200 ( .A(n8520), .B(n8519), .Z(n8537) );
  XOR U9201 ( .A(n8538), .B(n8537), .Z(o[83]) );
  NANDN U9202 ( .A(n8518), .B(n8517), .Z(n8522) );
  NAND U9203 ( .A(n8520), .B(n8519), .Z(n8521) );
  AND U9204 ( .A(n8522), .B(n8521), .Z(n8609) );
  NANDN U9205 ( .A(n8524), .B(n8523), .Z(n8528) );
  NANDN U9206 ( .A(n8526), .B(n8525), .Z(n8527) );
  AND U9207 ( .A(n8528), .B(n8527), .Z(n8608) );
  XNOR U9208 ( .A(n8609), .B(n8608), .Z(n8610) );
  NANDN U9209 ( .A(n8530), .B(n8529), .Z(n8534) );
  NANDN U9210 ( .A(n8532), .B(n8531), .Z(n8533) );
  NAND U9211 ( .A(n8534), .B(n8533), .Z(n8611) );
  XNOR U9212 ( .A(n8610), .B(n8611), .Z(n8614) );
  NANDN U9213 ( .A(n8536), .B(n8535), .Z(n8540) );
  NAND U9214 ( .A(n8538), .B(n8537), .Z(n8539) );
  NAND U9215 ( .A(n8540), .B(n8539), .Z(n8615) );
  XNOR U9216 ( .A(n8614), .B(n8615), .Z(n8617) );
  NANDN U9217 ( .A(n8542), .B(n8541), .Z(n8546) );
  NAND U9218 ( .A(n8544), .B(n8543), .Z(n8545) );
  AND U9219 ( .A(n8546), .B(n8545), .Z(n8621) );
  AND U9220 ( .A(y[42]), .B(x[90]), .Z(n8760) );
  AND U9221 ( .A(x[91]), .B(y[41]), .Z(n8548) );
  NAND U9222 ( .A(x[88]), .B(y[44]), .Z(n8547) );
  XOR U9223 ( .A(n8548), .B(n8547), .Z(n8683) );
  XNOR U9224 ( .A(n8760), .B(n8683), .Z(n8692) );
  NAND U9225 ( .A(y[43]), .B(x[89]), .Z(n8693) );
  XNOR U9226 ( .A(n8692), .B(n8693), .Z(n8695) );
  AND U9227 ( .A(y[120]), .B(x[108]), .Z(n8643) );
  NAND U9228 ( .A(y[3]), .B(x[81]), .Z(n8644) );
  XNOR U9229 ( .A(n8643), .B(n8644), .Z(n8645) );
  NAND U9230 ( .A(y[4]), .B(x[80]), .Z(n8646) );
  XNOR U9231 ( .A(n8645), .B(n8646), .Z(n8694) );
  XOR U9232 ( .A(n8695), .B(n8694), .Z(n8689) );
  NANDN U9233 ( .A(n8550), .B(n8549), .Z(n8554) );
  OR U9234 ( .A(n8552), .B(n8551), .Z(n8553) );
  AND U9235 ( .A(n8554), .B(n8553), .Z(n8687) );
  AND U9236 ( .A(y[163]), .B(x[115]), .Z(n8946) );
  NANDN U9237 ( .A(n8555), .B(n8946), .Z(n8559) );
  NANDN U9238 ( .A(n8557), .B(n8556), .Z(n8558) );
  AND U9239 ( .A(n8559), .B(n8558), .Z(n8686) );
  XNOR U9240 ( .A(n8687), .B(n8686), .Z(n8688) );
  XNOR U9241 ( .A(n8689), .B(n8688), .Z(n8719) );
  NAND U9242 ( .A(y[0]), .B(x[84]), .Z(n8670) );
  NAND U9243 ( .A(y[122]), .B(x[106]), .Z(n8669) );
  NAND U9244 ( .A(y[84]), .B(x[96]), .Z(n8668) );
  XOR U9245 ( .A(n8669), .B(n8668), .Z(n8671) );
  XNOR U9246 ( .A(n8670), .B(n8671), .Z(n8627) );
  AND U9247 ( .A(y[162]), .B(x[114]), .Z(n8601) );
  NAND U9248 ( .A(n8560), .B(n8601), .Z(n8663) );
  NAND U9249 ( .A(y[164]), .B(x[112]), .Z(n8815) );
  NAND U9250 ( .A(y[80]), .B(x[100]), .Z(n8775) );
  XNOR U9251 ( .A(n8815), .B(n8775), .Z(n8664) );
  XOR U9252 ( .A(n8663), .B(n8664), .Z(n8626) );
  XOR U9253 ( .A(n8627), .B(n8626), .Z(n8629) );
  NANDN U9254 ( .A(n8562), .B(n8561), .Z(n8566) );
  OR U9255 ( .A(n8564), .B(n8563), .Z(n8565) );
  AND U9256 ( .A(n8566), .B(n8565), .Z(n8628) );
  XOR U9257 ( .A(n8629), .B(n8628), .Z(n8717) );
  NANDN U9258 ( .A(n8568), .B(n8567), .Z(n8572) );
  NANDN U9259 ( .A(n8570), .B(n8569), .Z(n8571) );
  AND U9260 ( .A(n8572), .B(n8571), .Z(n8716) );
  XNOR U9261 ( .A(n8719), .B(n8718), .Z(n8620) );
  XNOR U9262 ( .A(n8621), .B(n8620), .Z(n8623) );
  NANDN U9263 ( .A(n8574), .B(n8573), .Z(n8578) );
  NANDN U9264 ( .A(n8576), .B(n8575), .Z(n8577) );
  AND U9265 ( .A(n8578), .B(n8577), .Z(n8705) );
  NANDN U9266 ( .A(n8580), .B(n8579), .Z(n8584) );
  NANDN U9267 ( .A(n8582), .B(n8581), .Z(n8583) );
  NAND U9268 ( .A(n8584), .B(n8583), .Z(n8704) );
  AND U9269 ( .A(y[81]), .B(x[99]), .Z(n8586) );
  NAND U9270 ( .A(n8586), .B(n8585), .Z(n8590) );
  NANDN U9271 ( .A(n8588), .B(n8587), .Z(n8589) );
  AND U9272 ( .A(n8590), .B(n8589), .Z(n8711) );
  AND U9273 ( .A(y[40]), .B(x[92]), .Z(n8649) );
  NAND U9274 ( .A(y[124]), .B(x[104]), .Z(n8650) );
  XNOR U9275 ( .A(n8649), .B(n8650), .Z(n8651) );
  NAND U9276 ( .A(y[123]), .B(x[105]), .Z(n8652) );
  XNOR U9277 ( .A(n8651), .B(n8652), .Z(n8698) );
  AND U9278 ( .A(x[98]), .B(y[82]), .Z(n8592) );
  NAND U9279 ( .A(x[99]), .B(y[81]), .Z(n8591) );
  XNOR U9280 ( .A(n8592), .B(n8591), .Z(n8639) );
  NAND U9281 ( .A(y[83]), .B(x[97]), .Z(n8640) );
  XOR U9282 ( .A(n8639), .B(n8640), .Z(n8699) );
  XNOR U9283 ( .A(n8698), .B(n8699), .Z(n8700) );
  NANDN U9284 ( .A(n8594), .B(n8593), .Z(n8598) );
  OR U9285 ( .A(n8596), .B(n8595), .Z(n8597) );
  NAND U9286 ( .A(n8598), .B(n8597), .Z(n8701) );
  XNOR U9287 ( .A(n8700), .B(n8701), .Z(n8710) );
  NAND U9288 ( .A(y[2]), .B(x[82]), .Z(n8678) );
  NAND U9289 ( .A(y[121]), .B(x[107]), .Z(n8677) );
  NAND U9290 ( .A(y[1]), .B(x[83]), .Z(n8676) );
  XNOR U9291 ( .A(n8677), .B(n8676), .Z(n8679) );
  AND U9292 ( .A(x[116]), .B(y[160]), .Z(n8600) );
  NAND U9293 ( .A(x[113]), .B(y[163]), .Z(n8599) );
  XNOR U9294 ( .A(n8600), .B(n8599), .Z(n8660) );
  AND U9295 ( .A(y[161]), .B(x[115]), .Z(n8782) );
  XOR U9296 ( .A(n8601), .B(n8782), .Z(n8659) );
  XOR U9297 ( .A(n8660), .B(n8659), .Z(n8632) );
  XOR U9298 ( .A(n8633), .B(n8632), .Z(n8634) );
  NANDN U9299 ( .A(n8603), .B(n8602), .Z(n8607) );
  OR U9300 ( .A(n8605), .B(n8604), .Z(n8606) );
  NAND U9301 ( .A(n8607), .B(n8606), .Z(n8635) );
  XOR U9302 ( .A(n8634), .B(n8635), .Z(n8713) );
  XOR U9303 ( .A(n8707), .B(n8706), .Z(n8622) );
  XNOR U9304 ( .A(n8623), .B(n8622), .Z(n8616) );
  XNOR U9305 ( .A(n8617), .B(n8616), .Z(o[84]) );
  NANDN U9306 ( .A(n8609), .B(n8608), .Z(n8613) );
  NANDN U9307 ( .A(n8611), .B(n8610), .Z(n8612) );
  AND U9308 ( .A(n8613), .B(n8612), .Z(n8857) );
  NANDN U9309 ( .A(n8615), .B(n8614), .Z(n8619) );
  NAND U9310 ( .A(n8617), .B(n8616), .Z(n8618) );
  NAND U9311 ( .A(n8619), .B(n8618), .Z(n8858) );
  XNOR U9312 ( .A(n8857), .B(n8858), .Z(n8860) );
  NANDN U9313 ( .A(n8621), .B(n8620), .Z(n8625) );
  NAND U9314 ( .A(n8623), .B(n8622), .Z(n8624) );
  AND U9315 ( .A(n8625), .B(n8624), .Z(n8723) );
  NAND U9316 ( .A(n8627), .B(n8626), .Z(n8631) );
  NAND U9317 ( .A(n8629), .B(n8628), .Z(n8630) );
  AND U9318 ( .A(n8631), .B(n8630), .Z(n8784) );
  NAND U9319 ( .A(n8633), .B(n8632), .Z(n8637) );
  NANDN U9320 ( .A(n8635), .B(n8634), .Z(n8636) );
  NAND U9321 ( .A(n8637), .B(n8636), .Z(n8783) );
  XNOR U9322 ( .A(n8784), .B(n8783), .Z(n8786) );
  AND U9323 ( .A(y[82]), .B(x[99]), .Z(n8776) );
  NAND U9324 ( .A(n8638), .B(n8776), .Z(n8642) );
  NANDN U9325 ( .A(n8640), .B(n8639), .Z(n8641) );
  AND U9326 ( .A(n8642), .B(n8641), .Z(n8739) );
  NANDN U9327 ( .A(n8644), .B(n8643), .Z(n8648) );
  NANDN U9328 ( .A(n8646), .B(n8645), .Z(n8647) );
  NAND U9329 ( .A(n8648), .B(n8647), .Z(n8746) );
  AND U9330 ( .A(y[125]), .B(x[104]), .Z(n8883) );
  AND U9331 ( .A(y[40]), .B(x[93]), .Z(n8766) );
  AND U9332 ( .A(y[83]), .B(x[98]), .Z(n8765) );
  XOR U9333 ( .A(n8766), .B(n8765), .Z(n8767) );
  XOR U9334 ( .A(n8883), .B(n8767), .Z(n8745) );
  AND U9335 ( .A(y[1]), .B(x[84]), .Z(n8888) );
  AND U9336 ( .A(y[121]), .B(x[108]), .Z(n8771) );
  AND U9337 ( .A(y[0]), .B(x[85]), .Z(n8770) );
  XOR U9338 ( .A(n8771), .B(n8770), .Z(n8772) );
  XOR U9339 ( .A(n8888), .B(n8772), .Z(n8744) );
  XOR U9340 ( .A(n8745), .B(n8744), .Z(n8747) );
  XOR U9341 ( .A(n8746), .B(n8747), .Z(n8738) );
  NANDN U9342 ( .A(n8650), .B(n8649), .Z(n8654) );
  NANDN U9343 ( .A(n8652), .B(n8651), .Z(n8653) );
  NAND U9344 ( .A(n8654), .B(n8653), .Z(n8853) );
  AND U9345 ( .A(y[162]), .B(x[115]), .Z(n8665) );
  AND U9346 ( .A(n8665), .B(n8655), .Z(n8817) );
  AND U9347 ( .A(x[112]), .B(y[165]), .Z(n8657) );
  AND U9348 ( .A(x[113]), .B(y[164]), .Z(n8656) );
  XOR U9349 ( .A(n8657), .B(n8656), .Z(n8816) );
  XOR U9350 ( .A(n8817), .B(n8816), .Z(n8852) );
  AND U9351 ( .A(y[45]), .B(x[88]), .Z(n8842) );
  AND U9352 ( .A(y[4]), .B(x[81]), .Z(n8841) );
  XOR U9353 ( .A(n8842), .B(n8841), .Z(n8844) );
  AND U9354 ( .A(y[41]), .B(x[92]), .Z(n8843) );
  XOR U9355 ( .A(n8844), .B(n8843), .Z(n8851) );
  XOR U9356 ( .A(n8852), .B(n8851), .Z(n8854) );
  XOR U9357 ( .A(n8853), .B(n8854), .Z(n8740) );
  XOR U9358 ( .A(n8741), .B(n8740), .Z(n8785) );
  XOR U9359 ( .A(n8786), .B(n8785), .Z(n8729) );
  AND U9360 ( .A(y[163]), .B(x[116]), .Z(n9013) );
  NAND U9361 ( .A(n9013), .B(n8658), .Z(n8662) );
  NAND U9362 ( .A(n8660), .B(n8659), .Z(n8661) );
  AND U9363 ( .A(n8662), .B(n8661), .Z(n8798) );
  XNOR U9364 ( .A(n8798), .B(n8797), .Z(n8800) );
  AND U9365 ( .A(y[163]), .B(x[114]), .Z(n8748) );
  NAND U9366 ( .A(y[160]), .B(x[117]), .Z(n8749) );
  XNOR U9367 ( .A(n8748), .B(n8749), .Z(n8750) );
  NAND U9368 ( .A(y[161]), .B(x[116]), .Z(n8967) );
  XOR U9369 ( .A(n8665), .B(n8967), .Z(n8751) );
  XNOR U9370 ( .A(n8750), .B(n8751), .Z(n8787) );
  AND U9371 ( .A(x[90]), .B(y[43]), .Z(n8667) );
  NAND U9372 ( .A(x[91]), .B(y[42]), .Z(n8666) );
  XNOR U9373 ( .A(n8667), .B(n8666), .Z(n8761) );
  NAND U9374 ( .A(y[44]), .B(x[89]), .Z(n8762) );
  XOR U9375 ( .A(n8761), .B(n8762), .Z(n8788) );
  XNOR U9376 ( .A(n8787), .B(n8788), .Z(n8789) );
  NAND U9377 ( .A(n8669), .B(n8668), .Z(n8673) );
  NAND U9378 ( .A(n8671), .B(n8670), .Z(n8672) );
  NAND U9379 ( .A(n8673), .B(n8672), .Z(n8790) );
  XNOR U9380 ( .A(n8789), .B(n8790), .Z(n8799) );
  XOR U9381 ( .A(n8800), .B(n8799), .Z(n8811) );
  AND U9382 ( .A(x[100]), .B(y[81]), .Z(n8675) );
  NAND U9383 ( .A(x[101]), .B(y[80]), .Z(n8674) );
  XOR U9384 ( .A(n8675), .B(n8674), .Z(n8777) );
  XNOR U9385 ( .A(n8776), .B(n8777), .Z(n8834) );
  AND U9386 ( .A(y[120]), .B(x[109]), .Z(n8754) );
  NAND U9387 ( .A(y[2]), .B(x[83]), .Z(n8755) );
  XNOR U9388 ( .A(n8754), .B(n8755), .Z(n8757) );
  AND U9389 ( .A(y[3]), .B(x[82]), .Z(n8756) );
  XOR U9390 ( .A(n8757), .B(n8756), .Z(n8833) );
  XOR U9391 ( .A(n8834), .B(n8833), .Z(n8836) );
  NAND U9392 ( .A(n8677), .B(n8676), .Z(n8681) );
  NANDN U9393 ( .A(n8679), .B(n8678), .Z(n8680) );
  AND U9394 ( .A(n8681), .B(n8680), .Z(n8835) );
  XOR U9395 ( .A(n8836), .B(n8835), .Z(n8810) );
  AND U9396 ( .A(y[44]), .B(x[91]), .Z(n9012) );
  NAND U9397 ( .A(n9012), .B(n8682), .Z(n8685) );
  NANDN U9398 ( .A(n8683), .B(n8760), .Z(n8684) );
  AND U9399 ( .A(n8685), .B(n8684), .Z(n8796) );
  AND U9400 ( .A(y[122]), .B(x[107]), .Z(n8828) );
  AND U9401 ( .A(y[84]), .B(x[97]), .Z(n8895) );
  XOR U9402 ( .A(n8828), .B(n8895), .Z(n8830) );
  AND U9403 ( .A(y[85]), .B(x[96]), .Z(n8829) );
  XOR U9404 ( .A(n8830), .B(n8829), .Z(n8794) );
  AND U9405 ( .A(y[5]), .B(x[80]), .Z(n8821) );
  AND U9406 ( .A(y[124]), .B(x[105]), .Z(n8820) );
  XOR U9407 ( .A(n8821), .B(n8820), .Z(n8823) );
  AND U9408 ( .A(y[123]), .B(x[106]), .Z(n8822) );
  XOR U9409 ( .A(n8823), .B(n8822), .Z(n8793) );
  XOR U9410 ( .A(n8794), .B(n8793), .Z(n8795) );
  XOR U9411 ( .A(n8796), .B(n8795), .Z(n8809) );
  XOR U9412 ( .A(n8810), .B(n8809), .Z(n8812) );
  XOR U9413 ( .A(n8811), .B(n8812), .Z(n8727) );
  NANDN U9414 ( .A(n8687), .B(n8686), .Z(n8691) );
  NANDN U9415 ( .A(n8689), .B(n8688), .Z(n8690) );
  AND U9416 ( .A(n8691), .B(n8690), .Z(n8805) );
  NANDN U9417 ( .A(n8693), .B(n8692), .Z(n8697) );
  NAND U9418 ( .A(n8695), .B(n8694), .Z(n8696) );
  AND U9419 ( .A(n8697), .B(n8696), .Z(n8804) );
  NANDN U9420 ( .A(n8699), .B(n8698), .Z(n8703) );
  NANDN U9421 ( .A(n8701), .B(n8700), .Z(n8702) );
  NAND U9422 ( .A(n8703), .B(n8702), .Z(n8803) );
  XOR U9423 ( .A(n8804), .B(n8803), .Z(n8806) );
  XNOR U9424 ( .A(n8805), .B(n8806), .Z(n8726) );
  XOR U9425 ( .A(n8729), .B(n8728), .Z(n8722) );
  XNOR U9426 ( .A(n8723), .B(n8722), .Z(n8725) );
  NANDN U9427 ( .A(n8705), .B(n8704), .Z(n8709) );
  NAND U9428 ( .A(n8707), .B(n8706), .Z(n8708) );
  AND U9429 ( .A(n8709), .B(n8708), .Z(n8735) );
  NANDN U9430 ( .A(n8711), .B(n8710), .Z(n8715) );
  NANDN U9431 ( .A(n8713), .B(n8712), .Z(n8714) );
  AND U9432 ( .A(n8715), .B(n8714), .Z(n8733) );
  NANDN U9433 ( .A(n8717), .B(n8716), .Z(n8721) );
  NAND U9434 ( .A(n8719), .B(n8718), .Z(n8720) );
  AND U9435 ( .A(n8721), .B(n8720), .Z(n8732) );
  XOR U9436 ( .A(n8725), .B(n8724), .Z(n8859) );
  XOR U9437 ( .A(n8860), .B(n8859), .Z(o[85]) );
  NANDN U9438 ( .A(n8727), .B(n8726), .Z(n8731) );
  NAND U9439 ( .A(n8729), .B(n8728), .Z(n8730) );
  AND U9440 ( .A(n8731), .B(n8730), .Z(n9131) );
  NANDN U9441 ( .A(n8733), .B(n8732), .Z(n8737) );
  NANDN U9442 ( .A(n8735), .B(n8734), .Z(n8736) );
  NAND U9443 ( .A(n8737), .B(n8736), .Z(n9132) );
  NANDN U9444 ( .A(n8739), .B(n8738), .Z(n8743) );
  NAND U9445 ( .A(n8741), .B(n8740), .Z(n8742) );
  AND U9446 ( .A(n8743), .B(n8742), .Z(n9138) );
  NANDN U9447 ( .A(n8749), .B(n8748), .Z(n8753) );
  NANDN U9448 ( .A(n8751), .B(n8750), .Z(n8752) );
  NAND U9449 ( .A(n8753), .B(n8752), .Z(n9093) );
  NANDN U9450 ( .A(n8755), .B(n8754), .Z(n8759) );
  NAND U9451 ( .A(n8757), .B(n8756), .Z(n8758) );
  NAND U9452 ( .A(n8759), .B(n8758), .Z(n9096) );
  AND U9453 ( .A(x[91]), .B(y[43]), .Z(n8840) );
  NAND U9454 ( .A(n8760), .B(n8840), .Z(n8764) );
  NANDN U9455 ( .A(n8762), .B(n8761), .Z(n8763) );
  AND U9456 ( .A(n8764), .B(n8763), .Z(n8935) );
  AND U9457 ( .A(y[123]), .B(x[107]), .Z(n8917) );
  AND U9458 ( .A(y[83]), .B(x[99]), .Z(n8916) );
  XOR U9459 ( .A(n8917), .B(n8916), .Z(n8915) );
  AND U9460 ( .A(y[3]), .B(x[83]), .Z(n8914) );
  XOR U9461 ( .A(n8915), .B(n8914), .Z(n8937) );
  AND U9462 ( .A(y[124]), .B(x[106]), .Z(n8929) );
  AND U9463 ( .A(y[82]), .B(x[100]), .Z(n8928) );
  XOR U9464 ( .A(n8929), .B(n8928), .Z(n8927) );
  AND U9465 ( .A(y[4]), .B(x[82]), .Z(n8926) );
  XNOR U9466 ( .A(n8927), .B(n8926), .Z(n8936) );
  XNOR U9467 ( .A(n8935), .B(n8934), .Z(n9095) );
  XOR U9468 ( .A(n9096), .B(n9095), .Z(n9094) );
  XOR U9469 ( .A(n9093), .B(n9094), .Z(n8870) );
  XOR U9470 ( .A(n8869), .B(n8870), .Z(n8868) );
  NAND U9471 ( .A(n8766), .B(n8765), .Z(n8769) );
  NAND U9472 ( .A(n8883), .B(n8767), .Z(n8768) );
  NAND U9473 ( .A(n8769), .B(n8768), .Z(n9056) );
  NAND U9474 ( .A(n8771), .B(n8770), .Z(n8774) );
  NAND U9475 ( .A(n8888), .B(n8772), .Z(n8773) );
  NAND U9476 ( .A(n8774), .B(n8773), .Z(n9055) );
  XOR U9477 ( .A(n9056), .B(n9055), .Z(n9058) );
  AND U9478 ( .A(y[81]), .B(x[101]), .Z(n8901) );
  NANDN U9479 ( .A(n8775), .B(n8901), .Z(n8779) );
  NANDN U9480 ( .A(n8777), .B(n8776), .Z(n8778) );
  AND U9481 ( .A(n8779), .B(n8778), .Z(n9080) );
  AND U9482 ( .A(x[85]), .B(y[1]), .Z(n8781) );
  NAND U9483 ( .A(x[84]), .B(y[2]), .Z(n8780) );
  XNOR U9484 ( .A(n8781), .B(n8780), .Z(n8887) );
  AND U9485 ( .A(y[120]), .B(x[110]), .Z(n8886) );
  XOR U9486 ( .A(n8887), .B(n8886), .Z(n9082) );
  AND U9487 ( .A(y[165]), .B(x[113]), .Z(n8954) );
  AND U9488 ( .A(y[162]), .B(x[116]), .Z(n8827) );
  AND U9489 ( .A(n8827), .B(n8782), .Z(n8952) );
  AND U9490 ( .A(y[164]), .B(x[114]), .Z(n8951) );
  XOR U9491 ( .A(n8952), .B(n8951), .Z(n8953) );
  XNOR U9492 ( .A(n8954), .B(n8953), .Z(n9081) );
  XNOR U9493 ( .A(n9080), .B(n9079), .Z(n9057) );
  XOR U9494 ( .A(n9058), .B(n9057), .Z(n8867) );
  XOR U9495 ( .A(n8868), .B(n8867), .Z(n8866) );
  NANDN U9496 ( .A(n8788), .B(n8787), .Z(n8792) );
  NANDN U9497 ( .A(n8790), .B(n8789), .Z(n8791) );
  AND U9498 ( .A(n8792), .B(n8791), .Z(n9068) );
  NANDN U9499 ( .A(n8798), .B(n8797), .Z(n8802) );
  NAND U9500 ( .A(n8800), .B(n8799), .Z(n8801) );
  AND U9501 ( .A(n8802), .B(n8801), .Z(n9069) );
  XOR U9502 ( .A(n9070), .B(n9069), .Z(n9067) );
  XOR U9503 ( .A(n9068), .B(n9067), .Z(n8863) );
  XOR U9504 ( .A(n8864), .B(n8863), .Z(n9137) );
  XOR U9505 ( .A(n9138), .B(n9137), .Z(n9135) );
  NANDN U9506 ( .A(n8804), .B(n8803), .Z(n8808) );
  NANDN U9507 ( .A(n8806), .B(n8805), .Z(n8807) );
  AND U9508 ( .A(n8808), .B(n8807), .Z(n9109) );
  NANDN U9509 ( .A(n8810), .B(n8809), .Z(n8814) );
  OR U9510 ( .A(n8812), .B(n8811), .Z(n8813) );
  NAND U9511 ( .A(n8814), .B(n8813), .Z(n9112) );
  NANDN U9512 ( .A(n8815), .B(n8954), .Z(n8819) );
  NAND U9513 ( .A(n8817), .B(n8816), .Z(n8818) );
  NAND U9514 ( .A(n8819), .B(n8818), .Z(n9054) );
  NAND U9515 ( .A(n8821), .B(n8820), .Z(n8825) );
  NAND U9516 ( .A(n8823), .B(n8822), .Z(n8824) );
  AND U9517 ( .A(n8825), .B(n8824), .Z(n9074) );
  AND U9518 ( .A(y[5]), .B(x[81]), .Z(n8925) );
  AND U9519 ( .A(y[40]), .B(x[94]), .Z(n8924) );
  XOR U9520 ( .A(n8925), .B(n8924), .Z(n8923) );
  AND U9521 ( .A(y[46]), .B(x[88]), .Z(n8922) );
  XOR U9522 ( .A(n8923), .B(n8922), .Z(n9076) );
  NAND U9523 ( .A(x[117]), .B(y[161]), .Z(n8826) );
  XNOR U9524 ( .A(n8827), .B(n8826), .Z(n8948) );
  AND U9525 ( .A(y[160]), .B(x[118]), .Z(n8947) );
  XOR U9526 ( .A(n8948), .B(n8947), .Z(n8945) );
  XNOR U9527 ( .A(n8946), .B(n8945), .Z(n9075) );
  XNOR U9528 ( .A(n9074), .B(n9073), .Z(n9053) );
  XOR U9529 ( .A(n9054), .B(n9053), .Z(n9052) );
  NAND U9530 ( .A(n8828), .B(n8895), .Z(n8832) );
  NAND U9531 ( .A(n8830), .B(n8829), .Z(n8831) );
  NAND U9532 ( .A(n8832), .B(n8831), .Z(n9051) );
  XOR U9533 ( .A(n9052), .B(n9051), .Z(n9117) );
  NAND U9534 ( .A(n8834), .B(n8833), .Z(n8838) );
  NAND U9535 ( .A(n8836), .B(n8835), .Z(n8837) );
  AND U9536 ( .A(n8838), .B(n8837), .Z(n9116) );
  AND U9537 ( .A(y[166]), .B(x[112]), .Z(n8900) );
  XOR U9538 ( .A(n8901), .B(n8900), .Z(n8899) );
  AND U9539 ( .A(y[80]), .B(x[102]), .Z(n8898) );
  XOR U9540 ( .A(n8899), .B(n8898), .Z(n9088) );
  AND U9541 ( .A(y[86]), .B(x[96]), .Z(n8911) );
  AND U9542 ( .A(y[0]), .B(x[86]), .Z(n8910) );
  XOR U9543 ( .A(n8911), .B(n8910), .Z(n8909) );
  AND U9544 ( .A(y[121]), .B(x[109]), .Z(n8908) );
  XOR U9545 ( .A(n8909), .B(n8908), .Z(n9090) );
  AND U9546 ( .A(y[41]), .B(x[93]), .Z(n8962) );
  AND U9547 ( .A(y[44]), .B(x[90]), .Z(n8961) );
  XOR U9548 ( .A(n8962), .B(n8961), .Z(n8960) );
  AND U9549 ( .A(y[45]), .B(x[89]), .Z(n8959) );
  XOR U9550 ( .A(n8960), .B(n8959), .Z(n8941) );
  AND U9551 ( .A(x[92]), .B(y[42]), .Z(n8839) );
  XOR U9552 ( .A(n8840), .B(n8839), .Z(n8940) );
  XOR U9553 ( .A(n8941), .B(n8940), .Z(n9089) );
  XOR U9554 ( .A(n9090), .B(n9089), .Z(n9087) );
  XOR U9555 ( .A(n9088), .B(n9087), .Z(n8874) );
  NAND U9556 ( .A(n8842), .B(n8841), .Z(n8846) );
  NAND U9557 ( .A(n8844), .B(n8843), .Z(n8845) );
  AND U9558 ( .A(n8846), .B(n8845), .Z(n8875) );
  AND U9559 ( .A(y[122]), .B(x[108]), .Z(n8894) );
  AND U9560 ( .A(x[97]), .B(y[85]), .Z(n8848) );
  AND U9561 ( .A(x[98]), .B(y[84]), .Z(n8847) );
  XOR U9562 ( .A(n8848), .B(n8847), .Z(n8893) );
  XOR U9563 ( .A(n8894), .B(n8893), .Z(n8878) );
  AND U9564 ( .A(y[6]), .B(x[80]), .Z(n8882) );
  AND U9565 ( .A(y[126]), .B(x[104]), .Z(n8850) );
  AND U9566 ( .A(x[105]), .B(y[125]), .Z(n8849) );
  XOR U9567 ( .A(n8850), .B(n8849), .Z(n8881) );
  XNOR U9568 ( .A(n8882), .B(n8881), .Z(n8877) );
  XNOR U9569 ( .A(n8875), .B(n8876), .Z(n8873) );
  NAND U9570 ( .A(n8852), .B(n8851), .Z(n8856) );
  NAND U9571 ( .A(n8854), .B(n8853), .Z(n8855) );
  AND U9572 ( .A(n8856), .B(n8855), .Z(n8871) );
  XOR U9573 ( .A(n8872), .B(n8871), .Z(n9115) );
  XOR U9574 ( .A(n9116), .B(n9115), .Z(n9118) );
  XOR U9575 ( .A(n9112), .B(n9111), .Z(n9110) );
  XOR U9576 ( .A(n9109), .B(n9110), .Z(n9136) );
  XNOR U9577 ( .A(n9130), .B(n9129), .Z(n9125) );
  NANDN U9578 ( .A(n8858), .B(n8857), .Z(n8862) );
  NAND U9579 ( .A(n8860), .B(n8859), .Z(n8861) );
  NAND U9580 ( .A(n8862), .B(n8861), .Z(n9123) );
  XOR U9581 ( .A(n9124), .B(n9123), .Z(o[86]) );
  NANDN U9582 ( .A(n8876), .B(n8875), .Z(n8880) );
  NANDN U9583 ( .A(n8878), .B(n8877), .Z(n8879) );
  AND U9584 ( .A(n8880), .B(n8879), .Z(n9066) );
  NAND U9585 ( .A(n8882), .B(n8881), .Z(n8885) );
  AND U9586 ( .A(y[126]), .B(x[105]), .Z(n9017) );
  NAND U9587 ( .A(n8883), .B(n9017), .Z(n8884) );
  AND U9588 ( .A(n8885), .B(n8884), .Z(n8892) );
  NAND U9589 ( .A(n8887), .B(n8886), .Z(n8890) );
  AND U9590 ( .A(y[2]), .B(x[85]), .Z(n9014) );
  NAND U9591 ( .A(n8888), .B(n9014), .Z(n8889) );
  NAND U9592 ( .A(n8890), .B(n8889), .Z(n8891) );
  XNOR U9593 ( .A(n8892), .B(n8891), .Z(n8907) );
  NAND U9594 ( .A(n8894), .B(n8893), .Z(n8897) );
  AND U9595 ( .A(y[85]), .B(x[98]), .Z(n9018) );
  NAND U9596 ( .A(n8895), .B(n9018), .Z(n8896) );
  AND U9597 ( .A(n8897), .B(n8896), .Z(n8905) );
  NAND U9598 ( .A(n8899), .B(n8898), .Z(n8903) );
  NAND U9599 ( .A(n8901), .B(n8900), .Z(n8902) );
  NAND U9600 ( .A(n8903), .B(n8902), .Z(n8904) );
  XNOR U9601 ( .A(n8905), .B(n8904), .Z(n8906) );
  XOR U9602 ( .A(n8907), .B(n8906), .Z(n8933) );
  NAND U9603 ( .A(n8909), .B(n8908), .Z(n8913) );
  NAND U9604 ( .A(n8911), .B(n8910), .Z(n8912) );
  AND U9605 ( .A(n8913), .B(n8912), .Z(n8921) );
  NAND U9606 ( .A(n8915), .B(n8914), .Z(n8919) );
  NAND U9607 ( .A(n8917), .B(n8916), .Z(n8918) );
  NAND U9608 ( .A(n8919), .B(n8918), .Z(n8920) );
  XNOR U9609 ( .A(n8921), .B(n8920), .Z(n8931) );
  XNOR U9610 ( .A(n8931), .B(n8930), .Z(n8932) );
  XNOR U9611 ( .A(n8933), .B(n8932), .Z(n9064) );
  NAND U9612 ( .A(n8935), .B(n8934), .Z(n8939) );
  NANDN U9613 ( .A(n8937), .B(n8936), .Z(n8938) );
  AND U9614 ( .A(n8939), .B(n8938), .Z(n9062) );
  NAND U9615 ( .A(n8941), .B(n8940), .Z(n8944) );
  AND U9616 ( .A(y[42]), .B(x[91]), .Z(n8942) );
  AND U9617 ( .A(y[43]), .B(x[92]), .Z(n9011) );
  NAND U9618 ( .A(n8942), .B(n9011), .Z(n8943) );
  AND U9619 ( .A(n8944), .B(n8943), .Z(n9050) );
  NAND U9620 ( .A(n8946), .B(n8945), .Z(n8950) );
  AND U9621 ( .A(n8948), .B(n8947), .Z(n8949) );
  ANDN U9622 ( .B(n8950), .A(n8949), .Z(n8958) );
  AND U9623 ( .A(n8952), .B(n8951), .Z(n8956) );
  AND U9624 ( .A(n8954), .B(n8953), .Z(n8955) );
  OR U9625 ( .A(n8956), .B(n8955), .Z(n8957) );
  XNOR U9626 ( .A(n8958), .B(n8957), .Z(n9048) );
  NAND U9627 ( .A(n8960), .B(n8959), .Z(n8964) );
  NAND U9628 ( .A(n8962), .B(n8961), .Z(n8963) );
  AND U9629 ( .A(n8964), .B(n8963), .Z(n9046) );
  AND U9630 ( .A(x[84]), .B(y[3]), .Z(n8966) );
  NAND U9631 ( .A(x[101]), .B(y[82]), .Z(n8965) );
  XNOR U9632 ( .A(n8966), .B(n8965), .Z(n8972) );
  AND U9633 ( .A(x[81]), .B(y[6]), .Z(n8970) );
  AND U9634 ( .A(x[117]), .B(n8967), .Z(n8968) );
  NAND U9635 ( .A(n8968), .B(y[162]), .Z(n8969) );
  XNOR U9636 ( .A(n8970), .B(n8969), .Z(n8971) );
  XOR U9637 ( .A(n8972), .B(n8971), .Z(n8980) );
  AND U9638 ( .A(x[97]), .B(y[86]), .Z(n8974) );
  NAND U9639 ( .A(x[109]), .B(y[122]), .Z(n8973) );
  XNOR U9640 ( .A(n8974), .B(n8973), .Z(n8978) );
  AND U9641 ( .A(x[114]), .B(y[165]), .Z(n8976) );
  NAND U9642 ( .A(x[115]), .B(y[164]), .Z(n8975) );
  XNOR U9643 ( .A(n8976), .B(n8975), .Z(n8977) );
  XNOR U9644 ( .A(n8978), .B(n8977), .Z(n8979) );
  XNOR U9645 ( .A(n8980), .B(n8979), .Z(n9044) );
  AND U9646 ( .A(x[82]), .B(y[5]), .Z(n8982) );
  NAND U9647 ( .A(x[99]), .B(y[84]), .Z(n8981) );
  XNOR U9648 ( .A(n8982), .B(n8981), .Z(n8986) );
  AND U9649 ( .A(x[83]), .B(y[4]), .Z(n8984) );
  NAND U9650 ( .A(x[110]), .B(y[121]), .Z(n8983) );
  XNOR U9651 ( .A(n8984), .B(n8983), .Z(n8985) );
  XOR U9652 ( .A(n8986), .B(n8985), .Z(n8994) );
  AND U9653 ( .A(x[100]), .B(y[83]), .Z(n8988) );
  NAND U9654 ( .A(x[94]), .B(y[41]), .Z(n8987) );
  XNOR U9655 ( .A(n8988), .B(n8987), .Z(n8992) );
  AND U9656 ( .A(x[118]), .B(y[161]), .Z(n8990) );
  NAND U9657 ( .A(x[119]), .B(y[160]), .Z(n8989) );
  XNOR U9658 ( .A(n8990), .B(n8989), .Z(n8991) );
  XNOR U9659 ( .A(n8992), .B(n8991), .Z(n8993) );
  XNOR U9660 ( .A(n8994), .B(n8993), .Z(n9010) );
  AND U9661 ( .A(x[112]), .B(y[167]), .Z(n8996) );
  NAND U9662 ( .A(x[103]), .B(y[80]), .Z(n8995) );
  XNOR U9663 ( .A(n8996), .B(n8995), .Z(n9000) );
  AND U9664 ( .A(x[80]), .B(y[7]), .Z(n8998) );
  NAND U9665 ( .A(x[113]), .B(y[166]), .Z(n8997) );
  XNOR U9666 ( .A(n8998), .B(n8997), .Z(n8999) );
  XOR U9667 ( .A(n9000), .B(n8999), .Z(n9008) );
  AND U9668 ( .A(x[108]), .B(y[123]), .Z(n9002) );
  NAND U9669 ( .A(x[87]), .B(y[0]), .Z(n9001) );
  XNOR U9670 ( .A(n9002), .B(n9001), .Z(n9006) );
  AND U9671 ( .A(x[88]), .B(y[47]), .Z(n9004) );
  NAND U9672 ( .A(x[111]), .B(y[120]), .Z(n9003) );
  XNOR U9673 ( .A(n9004), .B(n9003), .Z(n9005) );
  XNOR U9674 ( .A(n9006), .B(n9005), .Z(n9007) );
  XNOR U9675 ( .A(n9008), .B(n9007), .Z(n9009) );
  XOR U9676 ( .A(n9010), .B(n9009), .Z(n9042) );
  XOR U9677 ( .A(n9012), .B(n9011), .Z(n9016) );
  XNOR U9678 ( .A(n9014), .B(n9013), .Z(n9015) );
  XNOR U9679 ( .A(n9016), .B(n9015), .Z(n9040) );
  AND U9680 ( .A(x[89]), .B(y[46]), .Z(n9038) );
  AND U9681 ( .A(x[104]), .B(y[127]), .Z(n9020) );
  XNOR U9682 ( .A(n9018), .B(n9017), .Z(n9019) );
  XNOR U9683 ( .A(n9020), .B(n9019), .Z(n9036) );
  AND U9684 ( .A(x[86]), .B(y[1]), .Z(n9022) );
  NAND U9685 ( .A(x[102]), .B(y[81]), .Z(n9021) );
  XNOR U9686 ( .A(n9022), .B(n9021), .Z(n9026) );
  AND U9687 ( .A(x[96]), .B(y[87]), .Z(n9024) );
  NAND U9688 ( .A(x[107]), .B(y[124]), .Z(n9023) );
  XNOR U9689 ( .A(n9024), .B(n9023), .Z(n9025) );
  XOR U9690 ( .A(n9026), .B(n9025), .Z(n9034) );
  AND U9691 ( .A(x[106]), .B(y[125]), .Z(n9028) );
  NAND U9692 ( .A(x[95]), .B(y[40]), .Z(n9027) );
  XNOR U9693 ( .A(n9028), .B(n9027), .Z(n9032) );
  AND U9694 ( .A(x[90]), .B(y[45]), .Z(n9030) );
  NAND U9695 ( .A(x[93]), .B(y[42]), .Z(n9029) );
  XNOR U9696 ( .A(n9030), .B(n9029), .Z(n9031) );
  XNOR U9697 ( .A(n9032), .B(n9031), .Z(n9033) );
  XNOR U9698 ( .A(n9034), .B(n9033), .Z(n9035) );
  XNOR U9699 ( .A(n9036), .B(n9035), .Z(n9037) );
  XNOR U9700 ( .A(n9038), .B(n9037), .Z(n9039) );
  XNOR U9701 ( .A(n9040), .B(n9039), .Z(n9041) );
  XNOR U9702 ( .A(n9042), .B(n9041), .Z(n9043) );
  XNOR U9703 ( .A(n9044), .B(n9043), .Z(n9045) );
  XNOR U9704 ( .A(n9046), .B(n9045), .Z(n9047) );
  XNOR U9705 ( .A(n9048), .B(n9047), .Z(n9049) );
  XNOR U9706 ( .A(n9050), .B(n9049), .Z(n9060) );
  XNOR U9707 ( .A(n9060), .B(n9059), .Z(n9061) );
  XNOR U9708 ( .A(n9062), .B(n9061), .Z(n9063) );
  XNOR U9709 ( .A(n9064), .B(n9063), .Z(n9065) );
  XNOR U9710 ( .A(n9066), .B(n9065), .Z(n9106) );
  NAND U9711 ( .A(n9068), .B(n9067), .Z(n9072) );
  NAND U9712 ( .A(n9070), .B(n9069), .Z(n9071) );
  AND U9713 ( .A(n9072), .B(n9071), .Z(n9104) );
  NAND U9714 ( .A(n9074), .B(n9073), .Z(n9078) );
  NANDN U9715 ( .A(n9076), .B(n9075), .Z(n9077) );
  AND U9716 ( .A(n9078), .B(n9077), .Z(n9086) );
  NAND U9717 ( .A(n9080), .B(n9079), .Z(n9084) );
  NANDN U9718 ( .A(n9082), .B(n9081), .Z(n9083) );
  NAND U9719 ( .A(n9084), .B(n9083), .Z(n9085) );
  XNOR U9720 ( .A(n9086), .B(n9085), .Z(n9102) );
  NAND U9721 ( .A(n9088), .B(n9087), .Z(n9092) );
  NAND U9722 ( .A(n9090), .B(n9089), .Z(n9091) );
  AND U9723 ( .A(n9092), .B(n9091), .Z(n9100) );
  NAND U9724 ( .A(n9094), .B(n9093), .Z(n9098) );
  NAND U9725 ( .A(n9096), .B(n9095), .Z(n9097) );
  NAND U9726 ( .A(n9098), .B(n9097), .Z(n9099) );
  XNOR U9727 ( .A(n9100), .B(n9099), .Z(n9101) );
  XNOR U9728 ( .A(n9102), .B(n9101), .Z(n9103) );
  XNOR U9729 ( .A(n9104), .B(n9103), .Z(n9105) );
  XNOR U9730 ( .A(n9106), .B(n9105), .Z(n9107) );
  NANDN U9731 ( .A(n9110), .B(n9109), .Z(n9114) );
  ANDN U9732 ( .B(n9112), .A(n9111), .Z(n9113) );
  ANDN U9733 ( .B(n9114), .A(n9113), .Z(n9122) );
  AND U9734 ( .A(n9116), .B(n9115), .Z(n9120) );
  ANDN U9735 ( .B(n9118), .A(n9117), .Z(n9119) );
  OR U9736 ( .A(n9120), .B(n9119), .Z(n9121) );
  NAND U9737 ( .A(n9124), .B(n9123), .Z(n9128) );
  NANDN U9738 ( .A(n9126), .B(n9125), .Z(n9127) );
  NAND U9739 ( .A(n9130), .B(n9129), .Z(n9134) );
  NANDN U9740 ( .A(n9132), .B(n9131), .Z(n9133) );
  NAND U9741 ( .A(y[168]), .B(x[112]), .Z(n9272) );
  NAND U9742 ( .A(y[48]), .B(x[88]), .Z(n9141) );
  XOR U9743 ( .A(n9272), .B(n9141), .Z(n9142) );
  AND U9744 ( .A(y[8]), .B(x[80]), .Z(n9149) );
  AND U9745 ( .A(y[88]), .B(x[96]), .Z(n9146) );
  XOR U9746 ( .A(n9149), .B(n9146), .Z(n9145) );
  AND U9747 ( .A(y[128]), .B(x[104]), .Z(n9144) );
  XNOR U9748 ( .A(n9145), .B(n9144), .Z(n9143) );
  XNOR U9749 ( .A(n9142), .B(n9143), .Z(o[88]) );
  AND U9750 ( .A(x[80]), .B(y[9]), .Z(n9140) );
  NAND U9751 ( .A(x[81]), .B(y[8]), .Z(n9139) );
  XNOR U9752 ( .A(n9140), .B(n9139), .Z(n9150) );
  NAND U9753 ( .A(y[48]), .B(x[89]), .Z(n9151) );
  XOR U9754 ( .A(n9150), .B(n9151), .Z(n9167) );
  AND U9755 ( .A(y[168]), .B(x[113]), .Z(n9368) );
  NAND U9756 ( .A(y[89]), .B(x[96]), .Z(n9154) );
  XNOR U9757 ( .A(n9368), .B(n9154), .Z(n9155) );
  AND U9758 ( .A(y[169]), .B(x[112]), .Z(n9178) );
  NAND U9759 ( .A(y[88]), .B(x[97]), .Z(n9177) );
  XOR U9760 ( .A(n9178), .B(n9177), .Z(n9156) );
  XOR U9761 ( .A(n9155), .B(n9156), .Z(n9166) );
  AND U9762 ( .A(y[49]), .B(x[88]), .Z(n9397) );
  AND U9763 ( .A(y[129]), .B(x[104]), .Z(n9171) );
  XOR U9764 ( .A(n9397), .B(n9171), .Z(n9173) );
  AND U9765 ( .A(y[128]), .B(x[105]), .Z(n9172) );
  XNOR U9766 ( .A(n9173), .B(n9172), .Z(n9165) );
  XOR U9767 ( .A(n9166), .B(n9165), .Z(n9168) );
  XOR U9768 ( .A(n9167), .B(n9168), .Z(n9162) );
  NAND U9769 ( .A(n9145), .B(n9144), .Z(n9148) );
  AND U9770 ( .A(n9149), .B(n9146), .Z(n9147) );
  ANDN U9771 ( .B(n9148), .A(n9147), .Z(n9159) );
  XNOR U9772 ( .A(n9160), .B(n9159), .Z(n9161) );
  XNOR U9773 ( .A(n9162), .B(n9161), .Z(o[89]) );
  AND U9774 ( .A(y[9]), .B(x[81]), .Z(n9200) );
  NAND U9775 ( .A(n9200), .B(n9149), .Z(n9153) );
  NANDN U9776 ( .A(n9151), .B(n9150), .Z(n9152) );
  NAND U9777 ( .A(n9153), .B(n9152), .Z(n9220) );
  NANDN U9778 ( .A(n9154), .B(n9368), .Z(n9158) );
  NANDN U9779 ( .A(n9156), .B(n9155), .Z(n9157) );
  NAND U9780 ( .A(n9158), .B(n9157), .Z(n9218) );
  AND U9781 ( .A(y[130]), .B(x[104]), .Z(n9224) );
  NAND U9782 ( .A(y[10]), .B(x[80]), .Z(n9225) );
  XNOR U9783 ( .A(n9224), .B(n9225), .Z(n9227) );
  AND U9784 ( .A(y[48]), .B(x[90]), .Z(n9226) );
  XOR U9785 ( .A(n9227), .B(n9226), .Z(n9219) );
  XOR U9786 ( .A(n9218), .B(n9219), .Z(n9221) );
  XNOR U9787 ( .A(n9220), .B(n9221), .Z(n9180) );
  NANDN U9788 ( .A(n9160), .B(n9159), .Z(n9164) );
  NAND U9789 ( .A(n9162), .B(n9161), .Z(n9163) );
  NAND U9790 ( .A(n9164), .B(n9163), .Z(n9179) );
  XOR U9791 ( .A(n9180), .B(n9179), .Z(n9182) );
  NAND U9792 ( .A(n9166), .B(n9165), .Z(n9170) );
  NAND U9793 ( .A(n9168), .B(n9167), .Z(n9169) );
  AND U9794 ( .A(n9170), .B(n9169), .Z(n9188) );
  AND U9795 ( .A(y[8]), .B(x[82]), .Z(n9198) );
  AND U9796 ( .A(y[90]), .B(x[96]), .Z(n9197) );
  XOR U9797 ( .A(n9198), .B(n9197), .Z(n9199) );
  XOR U9798 ( .A(n9200), .B(n9199), .Z(n9233) );
  AND U9799 ( .A(y[128]), .B(x[106]), .Z(n9232) );
  XOR U9800 ( .A(n9233), .B(n9232), .Z(n9235) );
  AND U9801 ( .A(y[88]), .B(x[98]), .Z(n9303) );
  AND U9802 ( .A(y[170]), .B(x[112]), .Z(n9210) );
  XOR U9803 ( .A(n9303), .B(n9210), .Z(n9212) );
  AND U9804 ( .A(y[89]), .B(x[97]), .Z(n9211) );
  XOR U9805 ( .A(n9212), .B(n9211), .Z(n9234) );
  XOR U9806 ( .A(n9235), .B(n9234), .Z(n9185) );
  AND U9807 ( .A(n9397), .B(n9171), .Z(n9175) );
  NAND U9808 ( .A(n9173), .B(n9172), .Z(n9174) );
  NANDN U9809 ( .A(n9175), .B(n9174), .Z(n9193) );
  AND U9810 ( .A(x[113]), .B(y[169]), .Z(n9277) );
  NAND U9811 ( .A(x[114]), .B(y[168]), .Z(n9176) );
  XNOR U9812 ( .A(n9277), .B(n9176), .Z(n9231) );
  ANDN U9813 ( .B(n9178), .A(n9177), .Z(n9230) );
  XOR U9814 ( .A(n9231), .B(n9230), .Z(n9192) );
  AND U9815 ( .A(y[129]), .B(x[105]), .Z(n9203) );
  NAND U9816 ( .A(y[49]), .B(x[89]), .Z(n9204) );
  XNOR U9817 ( .A(n9203), .B(n9204), .Z(n9205) );
  NAND U9818 ( .A(y[50]), .B(x[88]), .Z(n9206) );
  XNOR U9819 ( .A(n9205), .B(n9206), .Z(n9191) );
  XOR U9820 ( .A(n9192), .B(n9191), .Z(n9194) );
  XOR U9821 ( .A(n9193), .B(n9194), .Z(n9186) );
  XOR U9822 ( .A(n9185), .B(n9186), .Z(n9187) );
  XNOR U9823 ( .A(n9188), .B(n9187), .Z(n9181) );
  XNOR U9824 ( .A(n9182), .B(n9181), .Z(o[90]) );
  NAND U9825 ( .A(n9180), .B(n9179), .Z(n9184) );
  NAND U9826 ( .A(n9182), .B(n9181), .Z(n9183) );
  AND U9827 ( .A(n9184), .B(n9183), .Z(n9239) );
  NAND U9828 ( .A(n9186), .B(n9185), .Z(n9190) );
  NAND U9829 ( .A(n9188), .B(n9187), .Z(n9189) );
  NAND U9830 ( .A(n9190), .B(n9189), .Z(n9244) );
  NAND U9831 ( .A(n9192), .B(n9191), .Z(n9196) );
  NAND U9832 ( .A(n9194), .B(n9193), .Z(n9195) );
  NAND U9833 ( .A(n9196), .B(n9195), .Z(n9242) );
  NAND U9834 ( .A(n9198), .B(n9197), .Z(n9202) );
  NAND U9835 ( .A(n9200), .B(n9199), .Z(n9201) );
  NAND U9836 ( .A(n9202), .B(n9201), .Z(n9254) );
  NANDN U9837 ( .A(n9204), .B(n9203), .Z(n9208) );
  NANDN U9838 ( .A(n9206), .B(n9205), .Z(n9207) );
  AND U9839 ( .A(n9208), .B(n9207), .Z(n9294) );
  AND U9840 ( .A(y[131]), .B(x[104]), .Z(n9321) );
  AND U9841 ( .A(y[91]), .B(x[96]), .Z(n9320) );
  NAND U9842 ( .A(y[8]), .B(x[83]), .Z(n9319) );
  XOR U9843 ( .A(n9320), .B(n9319), .Z(n9322) );
  XOR U9844 ( .A(n9321), .B(n9322), .Z(n9292) );
  AND U9845 ( .A(x[98]), .B(y[89]), .Z(n9341) );
  NAND U9846 ( .A(x[99]), .B(y[88]), .Z(n9209) );
  XNOR U9847 ( .A(n9341), .B(n9209), .Z(n9304) );
  NAND U9848 ( .A(y[90]), .B(x[97]), .Z(n9305) );
  XNOR U9849 ( .A(n9292), .B(n9291), .Z(n9293) );
  XNOR U9850 ( .A(n9294), .B(n9293), .Z(n9255) );
  XOR U9851 ( .A(n9254), .B(n9255), .Z(n9257) );
  NAND U9852 ( .A(n9303), .B(n9210), .Z(n9214) );
  AND U9853 ( .A(n9212), .B(n9211), .Z(n9213) );
  ANDN U9854 ( .B(n9214), .A(n9213), .Z(n9299) );
  AND U9855 ( .A(y[10]), .B(x[81]), .Z(n9268) );
  AND U9856 ( .A(y[9]), .B(x[82]), .Z(n9267) );
  NAND U9857 ( .A(y[130]), .B(x[105]), .Z(n9266) );
  XOR U9858 ( .A(n9267), .B(n9266), .Z(n9269) );
  XOR U9859 ( .A(n9268), .B(n9269), .Z(n9298) );
  AND U9860 ( .A(x[115]), .B(y[168]), .Z(n9216) );
  NAND U9861 ( .A(x[112]), .B(y[171]), .Z(n9215) );
  XNOR U9862 ( .A(n9216), .B(n9215), .Z(n9273) );
  AND U9863 ( .A(x[114]), .B(y[169]), .Z(n9353) );
  NAND U9864 ( .A(x[113]), .B(y[170]), .Z(n9217) );
  XOR U9865 ( .A(n9353), .B(n9217), .Z(n9274) );
  XNOR U9866 ( .A(n9273), .B(n9274), .Z(n9297) );
  XOR U9867 ( .A(n9298), .B(n9297), .Z(n9300) );
  XOR U9868 ( .A(n9299), .B(n9300), .Z(n9256) );
  XOR U9869 ( .A(n9257), .B(n9256), .Z(n9243) );
  XOR U9870 ( .A(n9242), .B(n9243), .Z(n9245) );
  XOR U9871 ( .A(n9244), .B(n9245), .Z(n9238) );
  XOR U9872 ( .A(n9239), .B(n9238), .Z(n9241) );
  NAND U9873 ( .A(n9219), .B(n9218), .Z(n9223) );
  NAND U9874 ( .A(n9221), .B(n9220), .Z(n9222) );
  AND U9875 ( .A(n9223), .B(n9222), .Z(n9251) );
  NANDN U9876 ( .A(n9225), .B(n9224), .Z(n9229) );
  NAND U9877 ( .A(n9227), .B(n9226), .Z(n9228) );
  AND U9878 ( .A(n9229), .B(n9228), .Z(n9261) );
  XNOR U9879 ( .A(n9261), .B(n9260), .Z(n9263) );
  AND U9880 ( .A(y[48]), .B(x[91]), .Z(n9312) );
  AND U9881 ( .A(y[11]), .B(x[80]), .Z(n9311) );
  NAND U9882 ( .A(y[129]), .B(x[106]), .Z(n9310) );
  XOR U9883 ( .A(n9311), .B(n9310), .Z(n9313) );
  XOR U9884 ( .A(n9312), .B(n9313), .Z(n9288) );
  AND U9885 ( .A(y[51]), .B(x[88]), .Z(n9281) );
  AND U9886 ( .A(y[49]), .B(x[90]), .Z(n9280) );
  NAND U9887 ( .A(y[128]), .B(x[107]), .Z(n9279) );
  XOR U9888 ( .A(n9280), .B(n9279), .Z(n9282) );
  XOR U9889 ( .A(n9281), .B(n9282), .Z(n9286) );
  AND U9890 ( .A(y[50]), .B(x[89]), .Z(n9285) );
  XNOR U9891 ( .A(n9263), .B(n9262), .Z(n9249) );
  NAND U9892 ( .A(n9233), .B(n9232), .Z(n9237) );
  NAND U9893 ( .A(n9235), .B(n9234), .Z(n9236) );
  AND U9894 ( .A(n9237), .B(n9236), .Z(n9248) );
  XOR U9895 ( .A(n9249), .B(n9248), .Z(n9250) );
  XNOR U9896 ( .A(n9251), .B(n9250), .Z(n9240) );
  XOR U9897 ( .A(n9241), .B(n9240), .Z(o[91]) );
  NAND U9898 ( .A(n9243), .B(n9242), .Z(n9247) );
  NAND U9899 ( .A(n9245), .B(n9244), .Z(n9246) );
  AND U9900 ( .A(n9247), .B(n9246), .Z(n9331) );
  NAND U9901 ( .A(n9249), .B(n9248), .Z(n9253) );
  NAND U9902 ( .A(n9251), .B(n9250), .Z(n9252) );
  NAND U9903 ( .A(n9253), .B(n9252), .Z(n9329) );
  NAND U9904 ( .A(n9255), .B(n9254), .Z(n9259) );
  NAND U9905 ( .A(n9257), .B(n9256), .Z(n9258) );
  AND U9906 ( .A(n9259), .B(n9258), .Z(n9330) );
  XOR U9907 ( .A(n9329), .B(n9330), .Z(n9332) );
  XOR U9908 ( .A(n9331), .B(n9332), .Z(n9325) );
  XOR U9909 ( .A(n9326), .B(n9325), .Z(n9328) );
  AND U9910 ( .A(y[50]), .B(x[90]), .Z(n9461) );
  AND U9911 ( .A(x[91]), .B(y[49]), .Z(n9265) );
  AND U9912 ( .A(x[88]), .B(y[52]), .Z(n9264) );
  XOR U9913 ( .A(n9265), .B(n9264), .Z(n9398) );
  XOR U9914 ( .A(n9461), .B(n9398), .Z(n9406) );
  AND U9915 ( .A(y[51]), .B(x[89]), .Z(n9405) );
  XOR U9916 ( .A(n9406), .B(n9405), .Z(n9408) );
  AND U9917 ( .A(y[128]), .B(x[108]), .Z(n9345) );
  AND U9918 ( .A(y[11]), .B(x[81]), .Z(n9344) );
  XOR U9919 ( .A(n9345), .B(n9344), .Z(n9347) );
  AND U9920 ( .A(y[12]), .B(x[80]), .Z(n9346) );
  XOR U9921 ( .A(n9347), .B(n9346), .Z(n9407) );
  XOR U9922 ( .A(n9408), .B(n9407), .Z(n9402) );
  NANDN U9923 ( .A(n9267), .B(n9266), .Z(n9271) );
  OR U9924 ( .A(n9269), .B(n9268), .Z(n9270) );
  AND U9925 ( .A(n9271), .B(n9270), .Z(n9400) );
  AND U9926 ( .A(y[171]), .B(x[115]), .Z(n9603) );
  NANDN U9927 ( .A(n9272), .B(n9603), .Z(n9276) );
  NANDN U9928 ( .A(n9274), .B(n9273), .Z(n9275) );
  AND U9929 ( .A(n9276), .B(n9275), .Z(n9399) );
  XNOR U9930 ( .A(n9400), .B(n9399), .Z(n9401) );
  XNOR U9931 ( .A(n9402), .B(n9401), .Z(n9428) );
  AND U9932 ( .A(y[8]), .B(x[84]), .Z(n9382) );
  AND U9933 ( .A(y[130]), .B(x[106]), .Z(n9380) );
  NAND U9934 ( .A(y[92]), .B(x[96]), .Z(n9379) );
  AND U9935 ( .A(y[170]), .B(x[114]), .Z(n9278) );
  AND U9936 ( .A(n9278), .B(n9277), .Z(n9376) );
  AND U9937 ( .A(y[172]), .B(x[112]), .Z(n9374) );
  IV U9938 ( .A(n9374), .Z(n9547) );
  AND U9939 ( .A(y[88]), .B(x[100]), .Z(n9373) );
  XNOR U9940 ( .A(n9547), .B(n9373), .Z(n9375) );
  XOR U9941 ( .A(n9376), .B(n9375), .Z(n9356) );
  XOR U9942 ( .A(n9357), .B(n9356), .Z(n9359) );
  NANDN U9943 ( .A(n9280), .B(n9279), .Z(n9284) );
  OR U9944 ( .A(n9282), .B(n9281), .Z(n9283) );
  AND U9945 ( .A(n9284), .B(n9283), .Z(n9358) );
  XOR U9946 ( .A(n9359), .B(n9358), .Z(n9426) );
  NANDN U9947 ( .A(n9286), .B(n9285), .Z(n9290) );
  NANDN U9948 ( .A(n9288), .B(n9287), .Z(n9289) );
  AND U9949 ( .A(n9290), .B(n9289), .Z(n9425) );
  XNOR U9950 ( .A(n9428), .B(n9427), .Z(n9335) );
  XNOR U9951 ( .A(n9336), .B(n9335), .Z(n9338) );
  NANDN U9952 ( .A(n9292), .B(n9291), .Z(n9296) );
  NANDN U9953 ( .A(n9294), .B(n9293), .Z(n9295) );
  AND U9954 ( .A(n9296), .B(n9295), .Z(n9414) );
  NANDN U9955 ( .A(n9298), .B(n9297), .Z(n9302) );
  OR U9956 ( .A(n9300), .B(n9299), .Z(n9301) );
  NAND U9957 ( .A(n9302), .B(n9301), .Z(n9413) );
  AND U9958 ( .A(y[89]), .B(x[99]), .Z(n9309) );
  NAND U9959 ( .A(n9309), .B(n9303), .Z(n9307) );
  NANDN U9960 ( .A(n9305), .B(n9304), .Z(n9306) );
  AND U9961 ( .A(n9307), .B(n9306), .Z(n9420) );
  AND U9962 ( .A(y[48]), .B(x[92]), .Z(n9349) );
  AND U9963 ( .A(y[132]), .B(x[104]), .Z(n9348) );
  XOR U9964 ( .A(n9349), .B(n9348), .Z(n9351) );
  AND U9965 ( .A(y[131]), .B(x[105]), .Z(n9350) );
  XOR U9966 ( .A(n9351), .B(n9350), .Z(n9410) );
  NAND U9967 ( .A(x[98]), .B(y[90]), .Z(n9308) );
  XNOR U9968 ( .A(n9309), .B(n9308), .Z(n9343) );
  AND U9969 ( .A(y[91]), .B(x[97]), .Z(n9342) );
  XOR U9970 ( .A(n9343), .B(n9342), .Z(n9409) );
  XOR U9971 ( .A(n9410), .B(n9409), .Z(n9411) );
  NANDN U9972 ( .A(n9311), .B(n9310), .Z(n9315) );
  OR U9973 ( .A(n9313), .B(n9312), .Z(n9314) );
  NAND U9974 ( .A(n9315), .B(n9314), .Z(n9412) );
  XNOR U9975 ( .A(n9411), .B(n9412), .Z(n9419) );
  AND U9976 ( .A(y[10]), .B(x[82]), .Z(n9394) );
  AND U9977 ( .A(y[129]), .B(x[107]), .Z(n9392) );
  NAND U9978 ( .A(y[9]), .B(x[83]), .Z(n9391) );
  AND U9979 ( .A(x[116]), .B(y[168]), .Z(n9317) );
  NAND U9980 ( .A(x[113]), .B(y[171]), .Z(n9316) );
  XNOR U9981 ( .A(n9317), .B(n9316), .Z(n9369) );
  AND U9982 ( .A(x[115]), .B(y[169]), .Z(n9486) );
  NAND U9983 ( .A(x[114]), .B(y[170]), .Z(n9318) );
  XOR U9984 ( .A(n9486), .B(n9318), .Z(n9370) );
  XOR U9985 ( .A(n9363), .B(n9362), .Z(n9364) );
  NANDN U9986 ( .A(n9320), .B(n9319), .Z(n9324) );
  OR U9987 ( .A(n9322), .B(n9321), .Z(n9323) );
  NAND U9988 ( .A(n9324), .B(n9323), .Z(n9365) );
  XOR U9989 ( .A(n9364), .B(n9365), .Z(n9422) );
  XOR U9990 ( .A(n9416), .B(n9415), .Z(n9337) );
  XNOR U9991 ( .A(n9338), .B(n9337), .Z(n9327) );
  XNOR U9992 ( .A(n9328), .B(n9327), .Z(o[92]) );
  NAND U9993 ( .A(n9330), .B(n9329), .Z(n9334) );
  NAND U9994 ( .A(n9332), .B(n9331), .Z(n9333) );
  NAND U9995 ( .A(n9334), .B(n9333), .Z(n9561) );
  XNOR U9996 ( .A(n9560), .B(n9561), .Z(n9563) );
  NANDN U9997 ( .A(n9336), .B(n9335), .Z(n9340) );
  NAND U9998 ( .A(n9338), .B(n9337), .Z(n9339) );
  AND U9999 ( .A(n9340), .B(n9339), .Z(n9432) );
  AND U10000 ( .A(y[90]), .B(x[99]), .Z(n9390) );
  IV U10001 ( .A(n9390), .Z(n9480) );
  AND U10002 ( .A(y[133]), .B(x[104]), .Z(n9690) );
  AND U10003 ( .A(y[48]), .B(x[93]), .Z(n9469) );
  AND U10004 ( .A(y[91]), .B(x[98]), .Z(n9468) );
  XOR U10005 ( .A(n9469), .B(n9468), .Z(n9470) );
  XOR U10006 ( .A(n9690), .B(n9470), .Z(n9465) );
  AND U10007 ( .A(y[129]), .B(x[108]), .Z(n9474) );
  AND U10008 ( .A(y[8]), .B(x[85]), .Z(n9473) );
  XOR U10009 ( .A(n9474), .B(n9473), .Z(n9475) );
  AND U10010 ( .A(y[9]), .B(x[84]), .Z(n9768) );
  XOR U10011 ( .A(n9475), .B(n9768), .Z(n9464) );
  XOR U10012 ( .A(n9465), .B(n9464), .Z(n9467) );
  XOR U10013 ( .A(n9466), .B(n9467), .Z(n9448) );
  XOR U10014 ( .A(n9447), .B(n9448), .Z(n9449) );
  AND U10015 ( .A(y[170]), .B(x[115]), .Z(n9352) );
  AND U10016 ( .A(n9353), .B(n9352), .Z(n9549) );
  AND U10017 ( .A(x[112]), .B(y[173]), .Z(n9355) );
  AND U10018 ( .A(x[113]), .B(y[172]), .Z(n9354) );
  XOR U10019 ( .A(n9355), .B(n9354), .Z(n9548) );
  XOR U10020 ( .A(n9549), .B(n9548), .Z(n9537) );
  AND U10021 ( .A(y[49]), .B(x[92]), .Z(n9529) );
  AND U10022 ( .A(y[53]), .B(x[88]), .Z(n9527) );
  AND U10023 ( .A(y[12]), .B(x[81]), .Z(n9526) );
  XOR U10024 ( .A(n9527), .B(n9526), .Z(n9528) );
  XOR U10025 ( .A(n9529), .B(n9528), .Z(n9536) );
  XOR U10026 ( .A(n9537), .B(n9536), .Z(n9539) );
  XNOR U10027 ( .A(n9538), .B(n9539), .Z(n9450) );
  NAND U10028 ( .A(n9357), .B(n9356), .Z(n9361) );
  NAND U10029 ( .A(n9359), .B(n9358), .Z(n9360) );
  NAND U10030 ( .A(n9361), .B(n9360), .Z(n9487) );
  NAND U10031 ( .A(n9363), .B(n9362), .Z(n9367) );
  NANDN U10032 ( .A(n9365), .B(n9364), .Z(n9366) );
  NAND U10033 ( .A(n9367), .B(n9366), .Z(n9488) );
  XNOR U10034 ( .A(n9487), .B(n9488), .Z(n9491) );
  XNOR U10035 ( .A(n9490), .B(n9491), .Z(n9438) );
  AND U10036 ( .A(y[171]), .B(x[116]), .Z(n9754) );
  NAND U10037 ( .A(n9754), .B(n9368), .Z(n9372) );
  NANDN U10038 ( .A(n9370), .B(n9369), .Z(n9371) );
  NAND U10039 ( .A(n9372), .B(n9371), .Z(n9498) );
  IV U10040 ( .A(n9373), .Z(n9478) );
  NANDN U10041 ( .A(n9374), .B(n9478), .Z(n9378) );
  NANDN U10042 ( .A(n9376), .B(n9375), .Z(n9377) );
  AND U10043 ( .A(n9378), .B(n9377), .Z(n9499) );
  XOR U10044 ( .A(n9498), .B(n9499), .Z(n9501) );
  NANDN U10045 ( .A(n9380), .B(n9379), .Z(n9384) );
  NANDN U10046 ( .A(n9382), .B(n9381), .Z(n9383) );
  AND U10047 ( .A(n9384), .B(n9383), .Z(n9505) );
  AND U10048 ( .A(x[90]), .B(y[51]), .Z(n9386) );
  NAND U10049 ( .A(x[91]), .B(y[50]), .Z(n9385) );
  XNOR U10050 ( .A(n9386), .B(n9385), .Z(n9463) );
  AND U10051 ( .A(y[52]), .B(x[89]), .Z(n9462) );
  XOR U10052 ( .A(n9463), .B(n9462), .Z(n9503) );
  AND U10053 ( .A(y[171]), .B(x[114]), .Z(n9454) );
  AND U10054 ( .A(y[168]), .B(x[117]), .Z(n9453) );
  XOR U10055 ( .A(n9454), .B(n9453), .Z(n9456) );
  AND U10056 ( .A(y[169]), .B(x[116]), .Z(n9736) );
  NAND U10057 ( .A(x[115]), .B(y[170]), .Z(n9387) );
  XNOR U10058 ( .A(n9736), .B(n9387), .Z(n9455) );
  XOR U10059 ( .A(n9456), .B(n9455), .Z(n9502) );
  XOR U10060 ( .A(n9503), .B(n9502), .Z(n9504) );
  XOR U10061 ( .A(n9505), .B(n9504), .Z(n9500) );
  XOR U10062 ( .A(n9501), .B(n9500), .Z(n9515) );
  AND U10063 ( .A(x[100]), .B(y[89]), .Z(n9389) );
  NAND U10064 ( .A(x[101]), .B(y[88]), .Z(n9388) );
  XNOR U10065 ( .A(n9389), .B(n9388), .Z(n9479) );
  XOR U10066 ( .A(n9479), .B(n9390), .Z(n9519) );
  AND U10067 ( .A(y[128]), .B(x[109]), .Z(n9458) );
  AND U10068 ( .A(y[10]), .B(x[83]), .Z(n9457) );
  XOR U10069 ( .A(n9458), .B(n9457), .Z(n9460) );
  AND U10070 ( .A(y[11]), .B(x[82]), .Z(n9459) );
  XOR U10071 ( .A(n9460), .B(n9459), .Z(n9518) );
  XOR U10072 ( .A(n9519), .B(n9518), .Z(n9521) );
  NANDN U10073 ( .A(n9392), .B(n9391), .Z(n9396) );
  NANDN U10074 ( .A(n9394), .B(n9393), .Z(n9395) );
  AND U10075 ( .A(n9396), .B(n9395), .Z(n9520) );
  XOR U10076 ( .A(n9521), .B(n9520), .Z(n9513) );
  AND U10077 ( .A(y[52]), .B(x[91]), .Z(n9753) );
  AND U10078 ( .A(y[130]), .B(x[107]), .Z(n9542) );
  AND U10079 ( .A(y[92]), .B(x[97]), .Z(n9676) );
  XOR U10080 ( .A(n9542), .B(n9676), .Z(n9544) );
  AND U10081 ( .A(y[93]), .B(x[96]), .Z(n9543) );
  XOR U10082 ( .A(n9544), .B(n9543), .Z(n9495) );
  AND U10083 ( .A(y[13]), .B(x[80]), .Z(n9553) );
  AND U10084 ( .A(y[132]), .B(x[105]), .Z(n9552) );
  XOR U10085 ( .A(n9553), .B(n9552), .Z(n9555) );
  AND U10086 ( .A(y[131]), .B(x[106]), .Z(n9554) );
  XOR U10087 ( .A(n9555), .B(n9554), .Z(n9494) );
  XOR U10088 ( .A(n9495), .B(n9494), .Z(n9497) );
  XOR U10089 ( .A(n9496), .B(n9497), .Z(n9512) );
  XOR U10090 ( .A(n9513), .B(n9512), .Z(n9514) );
  XOR U10091 ( .A(n9515), .B(n9514), .Z(n9435) );
  NANDN U10092 ( .A(n9400), .B(n9399), .Z(n9404) );
  NANDN U10093 ( .A(n9402), .B(n9401), .Z(n9403) );
  AND U10094 ( .A(n9404), .B(n9403), .Z(n9510) );
  XNOR U10095 ( .A(n9508), .B(n9509), .Z(n9511) );
  XNOR U10096 ( .A(n9510), .B(n9511), .Z(n9436) );
  XOR U10097 ( .A(n9435), .B(n9436), .Z(n9437) );
  XOR U10098 ( .A(n9438), .B(n9437), .Z(n9431) );
  XNOR U10099 ( .A(n9432), .B(n9431), .Z(n9434) );
  NANDN U10100 ( .A(n9414), .B(n9413), .Z(n9418) );
  NAND U10101 ( .A(n9416), .B(n9415), .Z(n9417) );
  AND U10102 ( .A(n9418), .B(n9417), .Z(n9444) );
  NANDN U10103 ( .A(n9420), .B(n9419), .Z(n9424) );
  NANDN U10104 ( .A(n9422), .B(n9421), .Z(n9423) );
  AND U10105 ( .A(n9424), .B(n9423), .Z(n9442) );
  NANDN U10106 ( .A(n9426), .B(n9425), .Z(n9430) );
  NAND U10107 ( .A(n9428), .B(n9427), .Z(n9429) );
  AND U10108 ( .A(n9430), .B(n9429), .Z(n9441) );
  XOR U10109 ( .A(n9434), .B(n9433), .Z(n9562) );
  XOR U10110 ( .A(n9563), .B(n9562), .Z(o[93]) );
  NAND U10111 ( .A(n9436), .B(n9435), .Z(n9440) );
  NAND U10112 ( .A(n9438), .B(n9437), .Z(n9439) );
  AND U10113 ( .A(n9440), .B(n9439), .Z(n9851) );
  NANDN U10114 ( .A(n9442), .B(n9441), .Z(n9446) );
  NANDN U10115 ( .A(n9444), .B(n9443), .Z(n9445) );
  NAND U10116 ( .A(n9446), .B(n9445), .Z(n9852) );
  NAND U10117 ( .A(n9448), .B(n9447), .Z(n9452) );
  NANDN U10118 ( .A(n9450), .B(n9449), .Z(n9451) );
  AND U10119 ( .A(n9452), .B(n9451), .Z(n9840) );
  AND U10120 ( .A(x[91]), .B(y[51]), .Z(n9525) );
  AND U10121 ( .A(y[131]), .B(x[107]), .Z(n9782) );
  AND U10122 ( .A(y[91]), .B(x[99]), .Z(n9781) );
  XOR U10123 ( .A(n9782), .B(n9781), .Z(n9780) );
  AND U10124 ( .A(y[11]), .B(x[83]), .Z(n9779) );
  XOR U10125 ( .A(n9780), .B(n9779), .Z(n9804) );
  AND U10126 ( .A(y[132]), .B(x[106]), .Z(n9740) );
  AND U10127 ( .A(y[90]), .B(x[100]), .Z(n9739) );
  XOR U10128 ( .A(n9740), .B(n9739), .Z(n9738) );
  AND U10129 ( .A(y[12]), .B(x[82]), .Z(n9737) );
  XNOR U10130 ( .A(n9738), .B(n9737), .Z(n9803) );
  XNOR U10131 ( .A(n9802), .B(n9801), .Z(n9594) );
  XOR U10132 ( .A(n9595), .B(n9594), .Z(n9593) );
  XOR U10133 ( .A(n9592), .B(n9593), .Z(n9575) );
  XOR U10134 ( .A(n9575), .B(n9574), .Z(n9573) );
  NAND U10135 ( .A(n9469), .B(n9468), .Z(n9472) );
  NAND U10136 ( .A(n9690), .B(n9470), .Z(n9471) );
  NAND U10137 ( .A(n9472), .B(n9471), .Z(n9710) );
  NAND U10138 ( .A(n9474), .B(n9473), .Z(n9477) );
  NAND U10139 ( .A(n9475), .B(n9768), .Z(n9476) );
  NAND U10140 ( .A(n9477), .B(n9476), .Z(n9709) );
  XOR U10141 ( .A(n9710), .B(n9709), .Z(n9708) );
  AND U10142 ( .A(y[89]), .B(x[101]), .Z(n9762) );
  NANDN U10143 ( .A(n9478), .B(n9762), .Z(n9482) );
  NANDN U10144 ( .A(n9480), .B(n9479), .Z(n9481) );
  AND U10145 ( .A(n9482), .B(n9481), .Z(n9714) );
  AND U10146 ( .A(x[85]), .B(y[9]), .Z(n9484) );
  NAND U10147 ( .A(x[84]), .B(y[10]), .Z(n9483) );
  XNOR U10148 ( .A(n9484), .B(n9483), .Z(n9766) );
  AND U10149 ( .A(y[128]), .B(x[110]), .Z(n9765) );
  XOR U10150 ( .A(n9766), .B(n9765), .Z(n9716) );
  AND U10151 ( .A(y[173]), .B(x[113]), .Z(n9682) );
  AND U10152 ( .A(y[170]), .B(x[116]), .Z(n9485) );
  AND U10153 ( .A(n9486), .B(n9485), .Z(n9680) );
  AND U10154 ( .A(y[172]), .B(x[114]), .Z(n9679) );
  XOR U10155 ( .A(n9680), .B(n9679), .Z(n9681) );
  XNOR U10156 ( .A(n9682), .B(n9681), .Z(n9715) );
  XNOR U10157 ( .A(n9714), .B(n9713), .Z(n9707) );
  XOR U10158 ( .A(n9708), .B(n9707), .Z(n9572) );
  XOR U10159 ( .A(n9573), .B(n9572), .Z(n9569) );
  IV U10160 ( .A(n9487), .Z(n9489) );
  NANDN U10161 ( .A(n9489), .B(n9488), .Z(n9493) );
  NANDN U10162 ( .A(n9491), .B(n9490), .Z(n9492) );
  AND U10163 ( .A(n9493), .B(n9492), .Z(n9568) );
  XOR U10164 ( .A(n9581), .B(n9580), .Z(n9579) );
  NAND U10165 ( .A(n9503), .B(n9502), .Z(n9507) );
  NAND U10166 ( .A(n9505), .B(n9504), .Z(n9506) );
  AND U10167 ( .A(n9507), .B(n9506), .Z(n9578) );
  XOR U10168 ( .A(n9579), .B(n9578), .Z(n9566) );
  XOR U10169 ( .A(n9567), .B(n9566), .Z(n9839) );
  XOR U10170 ( .A(n9840), .B(n9839), .Z(n9838) );
  OR U10171 ( .A(n9513), .B(n9512), .Z(n9517) );
  NANDN U10172 ( .A(n9515), .B(n9514), .Z(n9516) );
  NAND U10173 ( .A(n9517), .B(n9516), .Z(n9815) );
  NAND U10174 ( .A(n9519), .B(n9518), .Z(n9523) );
  NAND U10175 ( .A(n9521), .B(n9520), .Z(n9522) );
  AND U10176 ( .A(n9523), .B(n9522), .Z(n9820) );
  AND U10177 ( .A(y[94]), .B(x[96]), .Z(n9776) );
  AND U10178 ( .A(y[8]), .B(x[86]), .Z(n9775) );
  XOR U10179 ( .A(n9776), .B(n9775), .Z(n9774) );
  AND U10180 ( .A(y[129]), .B(x[109]), .Z(n9773) );
  XOR U10181 ( .A(n9774), .B(n9773), .Z(n9798) );
  AND U10182 ( .A(y[49]), .B(x[93]), .Z(n9728) );
  AND U10183 ( .A(y[52]), .B(x[90]), .Z(n9727) );
  XOR U10184 ( .A(n9728), .B(n9727), .Z(n9726) );
  AND U10185 ( .A(y[53]), .B(x[89]), .Z(n9725) );
  XOR U10186 ( .A(n9726), .B(n9725), .Z(n9694) );
  NAND U10187 ( .A(x[92]), .B(y[50]), .Z(n9524) );
  XNOR U10188 ( .A(n9525), .B(n9524), .Z(n9693) );
  XOR U10189 ( .A(n9694), .B(n9693), .Z(n9797) );
  XOR U10190 ( .A(n9798), .B(n9797), .Z(n9796) );
  AND U10191 ( .A(y[174]), .B(x[112]), .Z(n9761) );
  XOR U10192 ( .A(n9762), .B(n9761), .Z(n9760) );
  AND U10193 ( .A(y[88]), .B(x[102]), .Z(n9759) );
  XOR U10194 ( .A(n9760), .B(n9759), .Z(n9795) );
  XOR U10195 ( .A(n9796), .B(n9795), .Z(n9588) );
  NAND U10196 ( .A(n9527), .B(n9526), .Z(n9531) );
  NAND U10197 ( .A(n9529), .B(n9528), .Z(n9530) );
  AND U10198 ( .A(n9531), .B(n9530), .Z(n9596) );
  AND U10199 ( .A(y[130]), .B(x[108]), .Z(n9674) );
  AND U10200 ( .A(x[97]), .B(y[93]), .Z(n9533) );
  AND U10201 ( .A(x[98]), .B(y[92]), .Z(n9532) );
  XOR U10202 ( .A(n9533), .B(n9532), .Z(n9673) );
  XOR U10203 ( .A(n9674), .B(n9673), .Z(n9599) );
  AND U10204 ( .A(y[14]), .B(x[80]), .Z(n9688) );
  AND U10205 ( .A(y[134]), .B(x[104]), .Z(n9535) );
  AND U10206 ( .A(x[105]), .B(y[133]), .Z(n9534) );
  XOR U10207 ( .A(n9535), .B(n9534), .Z(n9687) );
  XNOR U10208 ( .A(n9688), .B(n9687), .Z(n9598) );
  XNOR U10209 ( .A(n9596), .B(n9597), .Z(n9589) );
  XNOR U10210 ( .A(n9588), .B(n9589), .Z(n9591) );
  NAND U10211 ( .A(n9537), .B(n9536), .Z(n9541) );
  NAND U10212 ( .A(n9539), .B(n9538), .Z(n9540) );
  AND U10213 ( .A(n9541), .B(n9540), .Z(n9590) );
  XOR U10214 ( .A(n9591), .B(n9590), .Z(n9819) );
  XOR U10215 ( .A(n9820), .B(n9819), .Z(n9822) );
  NAND U10216 ( .A(n9542), .B(n9676), .Z(n9546) );
  NAND U10217 ( .A(n9544), .B(n9543), .Z(n9545) );
  NAND U10218 ( .A(n9546), .B(n9545), .Z(n9584) );
  NANDN U10219 ( .A(n9547), .B(n9682), .Z(n9551) );
  NAND U10220 ( .A(n9549), .B(n9548), .Z(n9550) );
  NAND U10221 ( .A(n9551), .B(n9550), .Z(n9587) );
  NAND U10222 ( .A(n9553), .B(n9552), .Z(n9557) );
  NAND U10223 ( .A(n9555), .B(n9554), .Z(n9556) );
  AND U10224 ( .A(n9557), .B(n9556), .Z(n9668) );
  AND U10225 ( .A(y[13]), .B(x[81]), .Z(n9722) );
  AND U10226 ( .A(y[48]), .B(x[94]), .Z(n9721) );
  XOR U10227 ( .A(n9722), .B(n9721), .Z(n9720) );
  AND U10228 ( .A(y[54]), .B(x[88]), .Z(n9719) );
  XOR U10229 ( .A(n9720), .B(n9719), .Z(n9669) );
  AND U10230 ( .A(x[117]), .B(y[169]), .Z(n9559) );
  NAND U10231 ( .A(x[116]), .B(y[170]), .Z(n9558) );
  XNOR U10232 ( .A(n9559), .B(n9558), .Z(n9605) );
  AND U10233 ( .A(y[168]), .B(x[118]), .Z(n9604) );
  XOR U10234 ( .A(n9605), .B(n9604), .Z(n9602) );
  XNOR U10235 ( .A(n9603), .B(n9602), .Z(n9670) );
  XNOR U10236 ( .A(n9668), .B(n9667), .Z(n9586) );
  XOR U10237 ( .A(n9587), .B(n9586), .Z(n9585) );
  XOR U10238 ( .A(n9584), .B(n9585), .Z(n9821) );
  XOR U10239 ( .A(n9815), .B(n9816), .Z(n9813) );
  XOR U10240 ( .A(n9814), .B(n9813), .Z(n9837) );
  XOR U10241 ( .A(n9838), .B(n9837), .Z(n9849) );
  XNOR U10242 ( .A(n9850), .B(n9849), .Z(n9833) );
  NANDN U10243 ( .A(n9561), .B(n9560), .Z(n9565) );
  NAND U10244 ( .A(n9563), .B(n9562), .Z(n9564) );
  NAND U10245 ( .A(n9565), .B(n9564), .Z(n9831) );
  XOR U10246 ( .A(n9832), .B(n9831), .Z(o[94]) );
  NAND U10247 ( .A(n9567), .B(n9566), .Z(n9571) );
  NANDN U10248 ( .A(n9569), .B(n9568), .Z(n9570) );
  AND U10249 ( .A(n9571), .B(n9570), .Z(n9848) );
  NAND U10250 ( .A(n9573), .B(n9572), .Z(n9577) );
  NAND U10251 ( .A(n9575), .B(n9574), .Z(n9576) );
  AND U10252 ( .A(n9577), .B(n9576), .Z(n9830) );
  NAND U10253 ( .A(n9579), .B(n9578), .Z(n9583) );
  NAND U10254 ( .A(n9581), .B(n9580), .Z(n9582) );
  AND U10255 ( .A(n9583), .B(n9582), .Z(n9812) );
  NANDN U10256 ( .A(n9597), .B(n9596), .Z(n9601) );
  NANDN U10257 ( .A(n9599), .B(n9598), .Z(n9600) );
  NAND U10258 ( .A(n9603), .B(n9602), .Z(n9607) );
  NAND U10259 ( .A(n9605), .B(n9604), .Z(n9606) );
  AND U10260 ( .A(n9607), .B(n9606), .Z(n9666) );
  AND U10261 ( .A(x[86]), .B(y[9]), .Z(n9609) );
  NAND U10262 ( .A(x[102]), .B(y[89]), .Z(n9608) );
  XNOR U10263 ( .A(n9609), .B(n9608), .Z(n9613) );
  AND U10264 ( .A(x[118]), .B(y[169]), .Z(n9611) );
  NAND U10265 ( .A(x[119]), .B(y[168]), .Z(n9610) );
  XNOR U10266 ( .A(n9611), .B(n9610), .Z(n9612) );
  XOR U10267 ( .A(n9613), .B(n9612), .Z(n9621) );
  AND U10268 ( .A(x[100]), .B(y[91]), .Z(n9615) );
  NAND U10269 ( .A(x[99]), .B(y[92]), .Z(n9614) );
  XNOR U10270 ( .A(n9615), .B(n9614), .Z(n9619) );
  AND U10271 ( .A(x[108]), .B(y[131]), .Z(n9617) );
  NAND U10272 ( .A(x[87]), .B(y[8]), .Z(n9616) );
  XNOR U10273 ( .A(n9617), .B(n9616), .Z(n9618) );
  XNOR U10274 ( .A(n9619), .B(n9618), .Z(n9620) );
  XNOR U10275 ( .A(n9621), .B(n9620), .Z(n9664) );
  AND U10276 ( .A(x[93]), .B(y[50]), .Z(n9626) );
  AND U10277 ( .A(y[170]), .B(x[117]), .Z(n9735) );
  AND U10278 ( .A(x[106]), .B(y[133]), .Z(n9623) );
  NAND U10279 ( .A(x[95]), .B(y[48]), .Z(n9622) );
  XNOR U10280 ( .A(n9623), .B(n9622), .Z(n9624) );
  XNOR U10281 ( .A(n9735), .B(n9624), .Z(n9625) );
  XNOR U10282 ( .A(n9626), .B(n9625), .Z(n9642) );
  AND U10283 ( .A(x[96]), .B(y[95]), .Z(n9628) );
  NAND U10284 ( .A(x[97]), .B(y[94]), .Z(n9627) );
  XNOR U10285 ( .A(n9628), .B(n9627), .Z(n9632) );
  AND U10286 ( .A(x[88]), .B(y[55]), .Z(n9630) );
  NAND U10287 ( .A(x[107]), .B(y[132]), .Z(n9629) );
  XNOR U10288 ( .A(n9630), .B(n9629), .Z(n9631) );
  XOR U10289 ( .A(n9632), .B(n9631), .Z(n9640) );
  AND U10290 ( .A(x[104]), .B(y[135]), .Z(n9634) );
  NAND U10291 ( .A(x[111]), .B(y[128]), .Z(n9633) );
  XNOR U10292 ( .A(n9634), .B(n9633), .Z(n9638) );
  AND U10293 ( .A(x[89]), .B(y[54]), .Z(n9636) );
  NAND U10294 ( .A(x[90]), .B(y[53]), .Z(n9635) );
  XNOR U10295 ( .A(n9636), .B(n9635), .Z(n9637) );
  XNOR U10296 ( .A(n9638), .B(n9637), .Z(n9639) );
  XNOR U10297 ( .A(n9640), .B(n9639), .Z(n9641) );
  XOR U10298 ( .A(n9642), .B(n9641), .Z(n9662) );
  AND U10299 ( .A(x[113]), .B(y[174]), .Z(n9644) );
  NAND U10300 ( .A(x[103]), .B(y[88]), .Z(n9643) );
  XNOR U10301 ( .A(n9644), .B(n9643), .Z(n9648) );
  AND U10302 ( .A(x[82]), .B(y[13]), .Z(n9646) );
  NAND U10303 ( .A(x[110]), .B(y[129]), .Z(n9645) );
  XNOR U10304 ( .A(n9646), .B(n9645), .Z(n9647) );
  XOR U10305 ( .A(n9648), .B(n9647), .Z(n9656) );
  AND U10306 ( .A(x[114]), .B(y[173]), .Z(n9650) );
  NAND U10307 ( .A(x[115]), .B(y[172]), .Z(n9649) );
  XNOR U10308 ( .A(n9650), .B(n9649), .Z(n9654) );
  AND U10309 ( .A(x[80]), .B(y[15]), .Z(n9652) );
  NAND U10310 ( .A(x[84]), .B(y[11]), .Z(n9651) );
  XNOR U10311 ( .A(n9652), .B(n9651), .Z(n9653) );
  XNOR U10312 ( .A(n9654), .B(n9653), .Z(n9655) );
  XNOR U10313 ( .A(n9656), .B(n9655), .Z(n9660) );
  AND U10314 ( .A(y[93]), .B(x[98]), .Z(n9675) );
  AND U10315 ( .A(y[134]), .B(x[105]), .Z(n9689) );
  XOR U10316 ( .A(n9675), .B(n9689), .Z(n9658) );
  AND U10317 ( .A(y[10]), .B(x[85]), .Z(n9767) );
  AND U10318 ( .A(y[51]), .B(x[92]), .Z(n9695) );
  XNOR U10319 ( .A(n9767), .B(n9695), .Z(n9657) );
  XNOR U10320 ( .A(n9658), .B(n9657), .Z(n9659) );
  XNOR U10321 ( .A(n9660), .B(n9659), .Z(n9661) );
  XNOR U10322 ( .A(n9662), .B(n9661), .Z(n9663) );
  XNOR U10323 ( .A(n9664), .B(n9663), .Z(n9665) );
  XNOR U10324 ( .A(n9666), .B(n9665), .Z(n9706) );
  NAND U10325 ( .A(n9668), .B(n9667), .Z(n9672) );
  ANDN U10326 ( .B(n9670), .A(n9669), .Z(n9671) );
  ANDN U10327 ( .B(n9672), .A(n9671), .Z(n9704) );
  NAND U10328 ( .A(n9674), .B(n9673), .Z(n9678) );
  AND U10329 ( .A(n9676), .B(n9675), .Z(n9677) );
  ANDN U10330 ( .B(n9678), .A(n9677), .Z(n9686) );
  AND U10331 ( .A(n9680), .B(n9679), .Z(n9684) );
  AND U10332 ( .A(n9682), .B(n9681), .Z(n9683) );
  OR U10333 ( .A(n9684), .B(n9683), .Z(n9685) );
  XNOR U10334 ( .A(n9686), .B(n9685), .Z(n9702) );
  NAND U10335 ( .A(n9688), .B(n9687), .Z(n9692) );
  NAND U10336 ( .A(n9690), .B(n9689), .Z(n9691) );
  AND U10337 ( .A(n9692), .B(n9691), .Z(n9700) );
  NAND U10338 ( .A(n9694), .B(n9693), .Z(n9698) );
  AND U10339 ( .A(y[50]), .B(x[91]), .Z(n9696) );
  NAND U10340 ( .A(n9696), .B(n9695), .Z(n9697) );
  NAND U10341 ( .A(n9698), .B(n9697), .Z(n9699) );
  XNOR U10342 ( .A(n9700), .B(n9699), .Z(n9701) );
  XNOR U10343 ( .A(n9702), .B(n9701), .Z(n9703) );
  XNOR U10344 ( .A(n9704), .B(n9703), .Z(n9705) );
  NAND U10345 ( .A(n9708), .B(n9707), .Z(n9712) );
  NAND U10346 ( .A(n9710), .B(n9709), .Z(n9711) );
  NAND U10347 ( .A(n9714), .B(n9713), .Z(n9718) );
  NANDN U10348 ( .A(n9716), .B(n9715), .Z(n9717) );
  AND U10349 ( .A(n9718), .B(n9717), .Z(n9794) );
  NAND U10350 ( .A(n9720), .B(n9719), .Z(n9724) );
  NAND U10351 ( .A(n9722), .B(n9721), .Z(n9723) );
  AND U10352 ( .A(n9724), .B(n9723), .Z(n9732) );
  NAND U10353 ( .A(n9726), .B(n9725), .Z(n9730) );
  NAND U10354 ( .A(n9728), .B(n9727), .Z(n9729) );
  NAND U10355 ( .A(n9730), .B(n9729), .Z(n9731) );
  XNOR U10356 ( .A(n9732), .B(n9731), .Z(n9792) );
  AND U10357 ( .A(x[101]), .B(y[90]), .Z(n9734) );
  NAND U10358 ( .A(x[109]), .B(y[130]), .Z(n9733) );
  XNOR U10359 ( .A(n9734), .B(n9733), .Z(n9758) );
  AND U10360 ( .A(n9736), .B(n9735), .Z(n9752) );
  NAND U10361 ( .A(n9738), .B(n9737), .Z(n9742) );
  NAND U10362 ( .A(n9740), .B(n9739), .Z(n9741) );
  AND U10363 ( .A(n9742), .B(n9741), .Z(n9750) );
  AND U10364 ( .A(x[81]), .B(y[14]), .Z(n9744) );
  NAND U10365 ( .A(x[94]), .B(y[49]), .Z(n9743) );
  XNOR U10366 ( .A(n9744), .B(n9743), .Z(n9748) );
  AND U10367 ( .A(x[112]), .B(y[175]), .Z(n9746) );
  NAND U10368 ( .A(x[83]), .B(y[12]), .Z(n9745) );
  XNOR U10369 ( .A(n9746), .B(n9745), .Z(n9747) );
  XNOR U10370 ( .A(n9748), .B(n9747), .Z(n9749) );
  XNOR U10371 ( .A(n9750), .B(n9749), .Z(n9751) );
  XOR U10372 ( .A(n9752), .B(n9751), .Z(n9756) );
  XNOR U10373 ( .A(n9754), .B(n9753), .Z(n9755) );
  XNOR U10374 ( .A(n9756), .B(n9755), .Z(n9757) );
  XOR U10375 ( .A(n9758), .B(n9757), .Z(n9790) );
  NAND U10376 ( .A(n9760), .B(n9759), .Z(n9764) );
  NAND U10377 ( .A(n9762), .B(n9761), .Z(n9763) );
  AND U10378 ( .A(n9764), .B(n9763), .Z(n9772) );
  NAND U10379 ( .A(n9766), .B(n9765), .Z(n9770) );
  NAND U10380 ( .A(n9768), .B(n9767), .Z(n9769) );
  NAND U10381 ( .A(n9770), .B(n9769), .Z(n9771) );
  XNOR U10382 ( .A(n9772), .B(n9771), .Z(n9788) );
  NAND U10383 ( .A(n9774), .B(n9773), .Z(n9778) );
  NAND U10384 ( .A(n9776), .B(n9775), .Z(n9777) );
  AND U10385 ( .A(n9778), .B(n9777), .Z(n9786) );
  NAND U10386 ( .A(n9780), .B(n9779), .Z(n9784) );
  NAND U10387 ( .A(n9782), .B(n9781), .Z(n9783) );
  NAND U10388 ( .A(n9784), .B(n9783), .Z(n9785) );
  XNOR U10389 ( .A(n9786), .B(n9785), .Z(n9787) );
  XNOR U10390 ( .A(n9788), .B(n9787), .Z(n9789) );
  XNOR U10391 ( .A(n9790), .B(n9789), .Z(n9791) );
  XNOR U10392 ( .A(n9792), .B(n9791), .Z(n9793) );
  XNOR U10393 ( .A(n9794), .B(n9793), .Z(n9810) );
  NAND U10394 ( .A(n9796), .B(n9795), .Z(n9800) );
  NAND U10395 ( .A(n9798), .B(n9797), .Z(n9799) );
  AND U10396 ( .A(n9800), .B(n9799), .Z(n9808) );
  NAND U10397 ( .A(n9802), .B(n9801), .Z(n9806) );
  NANDN U10398 ( .A(n9804), .B(n9803), .Z(n9805) );
  NAND U10399 ( .A(n9806), .B(n9805), .Z(n9807) );
  XNOR U10400 ( .A(n9808), .B(n9807), .Z(n9809) );
  XNOR U10401 ( .A(n9812), .B(n9811), .Z(n9828) );
  NAND U10402 ( .A(n9814), .B(n9813), .Z(n9818) );
  AND U10403 ( .A(n9816), .B(n9815), .Z(n9817) );
  ANDN U10404 ( .B(n9818), .A(n9817), .Z(n9826) );
  AND U10405 ( .A(n9820), .B(n9819), .Z(n9824) );
  ANDN U10406 ( .B(n9822), .A(n9821), .Z(n9823) );
  OR U10407 ( .A(n9824), .B(n9823), .Z(n9825) );
  XNOR U10408 ( .A(n9826), .B(n9825), .Z(n9827) );
  XNOR U10409 ( .A(n9828), .B(n9827), .Z(n9829) );
  XNOR U10410 ( .A(n9830), .B(n9829), .Z(n9846) );
  NAND U10411 ( .A(n9832), .B(n9831), .Z(n9836) );
  NANDN U10412 ( .A(n9834), .B(n9833), .Z(n9835) );
  AND U10413 ( .A(n9836), .B(n9835), .Z(n9844) );
  NAND U10414 ( .A(n9838), .B(n9837), .Z(n9842) );
  NAND U10415 ( .A(n9840), .B(n9839), .Z(n9841) );
  NAND U10416 ( .A(n9842), .B(n9841), .Z(n9843) );
  XNOR U10417 ( .A(n9844), .B(n9843), .Z(n9845) );
  XNOR U10418 ( .A(n9846), .B(n9845), .Z(n9847) );
  XNOR U10419 ( .A(n9848), .B(n9847), .Z(n9856) );
  NAND U10420 ( .A(n9850), .B(n9849), .Z(n9854) );
  NANDN U10421 ( .A(n9852), .B(n9851), .Z(n9853) );
  NAND U10422 ( .A(n9854), .B(n9853), .Z(n9855) );
  XNOR U10423 ( .A(n9856), .B(n9855), .Z(o[95]) );
  NAND U10424 ( .A(y[176]), .B(x[112]), .Z(n9992) );
  NAND U10425 ( .A(y[56]), .B(x[88]), .Z(n9859) );
  XOR U10426 ( .A(n9992), .B(n9859), .Z(n9860) );
  AND U10427 ( .A(y[16]), .B(x[80]), .Z(n9867) );
  AND U10428 ( .A(y[96]), .B(x[96]), .Z(n9864) );
  XOR U10429 ( .A(n9867), .B(n9864), .Z(n9863) );
  AND U10430 ( .A(y[136]), .B(x[104]), .Z(n9862) );
  XNOR U10431 ( .A(n9863), .B(n9862), .Z(n9861) );
  XNOR U10432 ( .A(n9860), .B(n9861), .Z(o[96]) );
  AND U10433 ( .A(x[81]), .B(y[16]), .Z(n9858) );
  NAND U10434 ( .A(x[80]), .B(y[17]), .Z(n9857) );
  XNOR U10435 ( .A(n9858), .B(n9857), .Z(n9868) );
  NAND U10436 ( .A(y[56]), .B(x[89]), .Z(n9869) );
  XOR U10437 ( .A(n9868), .B(n9869), .Z(n9885) );
  AND U10438 ( .A(y[176]), .B(x[113]), .Z(n10087) );
  NAND U10439 ( .A(y[97]), .B(x[96]), .Z(n9872) );
  XNOR U10440 ( .A(n10087), .B(n9872), .Z(n9873) );
  AND U10441 ( .A(y[177]), .B(x[112]), .Z(n9897) );
  NAND U10442 ( .A(y[96]), .B(x[97]), .Z(n9896) );
  XOR U10443 ( .A(n9897), .B(n9896), .Z(n9874) );
  XOR U10444 ( .A(n9873), .B(n9874), .Z(n9884) );
  AND U10445 ( .A(y[57]), .B(x[88]), .Z(n10115) );
  AND U10446 ( .A(y[137]), .B(x[104]), .Z(n9889) );
  XOR U10447 ( .A(n10115), .B(n9889), .Z(n9891) );
  AND U10448 ( .A(y[136]), .B(x[105]), .Z(n9890) );
  XNOR U10449 ( .A(n9891), .B(n9890), .Z(n9883) );
  XOR U10450 ( .A(n9884), .B(n9883), .Z(n9886) );
  XOR U10451 ( .A(n9885), .B(n9886), .Z(n9880) );
  NAND U10452 ( .A(n9863), .B(n9862), .Z(n9866) );
  AND U10453 ( .A(n9867), .B(n9864), .Z(n9865) );
  ANDN U10454 ( .B(n9866), .A(n9865), .Z(n9877) );
  XNOR U10455 ( .A(n9878), .B(n9877), .Z(n9879) );
  XNOR U10456 ( .A(n9880), .B(n9879), .Z(o[97]) );
  AND U10457 ( .A(y[17]), .B(x[81]), .Z(n9919) );
  NAND U10458 ( .A(n9919), .B(n9867), .Z(n9871) );
  NANDN U10459 ( .A(n9869), .B(n9868), .Z(n9870) );
  NAND U10460 ( .A(n9871), .B(n9870), .Z(n9940) );
  NANDN U10461 ( .A(n9872), .B(n10087), .Z(n9876) );
  NANDN U10462 ( .A(n9874), .B(n9873), .Z(n9875) );
  NAND U10463 ( .A(n9876), .B(n9875), .Z(n9938) );
  AND U10464 ( .A(y[138]), .B(x[104]), .Z(n9944) );
  NAND U10465 ( .A(y[18]), .B(x[80]), .Z(n9945) );
  XNOR U10466 ( .A(n9944), .B(n9945), .Z(n9947) );
  AND U10467 ( .A(y[56]), .B(x[90]), .Z(n9946) );
  XOR U10468 ( .A(n9947), .B(n9946), .Z(n9939) );
  XOR U10469 ( .A(n9938), .B(n9939), .Z(n9941) );
  XNOR U10470 ( .A(n9940), .B(n9941), .Z(n9899) );
  NANDN U10471 ( .A(n9878), .B(n9877), .Z(n9882) );
  NAND U10472 ( .A(n9880), .B(n9879), .Z(n9881) );
  NAND U10473 ( .A(n9882), .B(n9881), .Z(n9898) );
  XOR U10474 ( .A(n9899), .B(n9898), .Z(n9901) );
  NAND U10475 ( .A(n9884), .B(n9883), .Z(n9888) );
  NAND U10476 ( .A(n9886), .B(n9885), .Z(n9887) );
  AND U10477 ( .A(n9888), .B(n9887), .Z(n9907) );
  AND U10478 ( .A(y[16]), .B(x[82]), .Z(n9917) );
  AND U10479 ( .A(y[98]), .B(x[96]), .Z(n9916) );
  XOR U10480 ( .A(n9917), .B(n9916), .Z(n9918) );
  XOR U10481 ( .A(n9919), .B(n9918), .Z(n9953) );
  AND U10482 ( .A(y[136]), .B(x[106]), .Z(n9952) );
  XOR U10483 ( .A(n9953), .B(n9952), .Z(n9955) );
  AND U10484 ( .A(y[96]), .B(x[98]), .Z(n10023) );
  AND U10485 ( .A(y[178]), .B(x[112]), .Z(n9930) );
  XOR U10486 ( .A(n10023), .B(n9930), .Z(n9932) );
  AND U10487 ( .A(y[97]), .B(x[97]), .Z(n9931) );
  XOR U10488 ( .A(n9932), .B(n9931), .Z(n9954) );
  XOR U10489 ( .A(n9955), .B(n9954), .Z(n9904) );
  AND U10490 ( .A(n10115), .B(n9889), .Z(n9893) );
  NAND U10491 ( .A(n9891), .B(n9890), .Z(n9892) );
  NANDN U10492 ( .A(n9893), .B(n9892), .Z(n9912) );
  AND U10493 ( .A(x[114]), .B(y[176]), .Z(n9895) );
  NAND U10494 ( .A(x[113]), .B(y[177]), .Z(n9894) );
  XNOR U10495 ( .A(n9895), .B(n9894), .Z(n9951) );
  ANDN U10496 ( .B(n9897), .A(n9896), .Z(n9950) );
  XOR U10497 ( .A(n9951), .B(n9950), .Z(n9911) );
  AND U10498 ( .A(y[137]), .B(x[105]), .Z(n9922) );
  NAND U10499 ( .A(y[57]), .B(x[89]), .Z(n9923) );
  XNOR U10500 ( .A(n9922), .B(n9923), .Z(n9924) );
  NAND U10501 ( .A(y[58]), .B(x[88]), .Z(n9925) );
  XNOR U10502 ( .A(n9924), .B(n9925), .Z(n9910) );
  XOR U10503 ( .A(n9911), .B(n9910), .Z(n9913) );
  XOR U10504 ( .A(n9912), .B(n9913), .Z(n9905) );
  XOR U10505 ( .A(n9904), .B(n9905), .Z(n9906) );
  XNOR U10506 ( .A(n9907), .B(n9906), .Z(n9900) );
  XNOR U10507 ( .A(n9901), .B(n9900), .Z(o[98]) );
  NAND U10508 ( .A(n9899), .B(n9898), .Z(n9903) );
  NAND U10509 ( .A(n9901), .B(n9900), .Z(n9902) );
  AND U10510 ( .A(n9903), .B(n9902), .Z(n9959) );
  NAND U10511 ( .A(n9905), .B(n9904), .Z(n9909) );
  NAND U10512 ( .A(n9907), .B(n9906), .Z(n9908) );
  NAND U10513 ( .A(n9909), .B(n9908), .Z(n9964) );
  NAND U10514 ( .A(n9911), .B(n9910), .Z(n9915) );
  NAND U10515 ( .A(n9913), .B(n9912), .Z(n9914) );
  NAND U10516 ( .A(n9915), .B(n9914), .Z(n9962) );
  NAND U10517 ( .A(n9917), .B(n9916), .Z(n9921) );
  NAND U10518 ( .A(n9919), .B(n9918), .Z(n9920) );
  NAND U10519 ( .A(n9921), .B(n9920), .Z(n9974) );
  NANDN U10520 ( .A(n9923), .B(n9922), .Z(n9927) );
  NANDN U10521 ( .A(n9925), .B(n9924), .Z(n9926) );
  AND U10522 ( .A(n9927), .B(n9926), .Z(n10014) );
  AND U10523 ( .A(y[139]), .B(x[104]), .Z(n10041) );
  AND U10524 ( .A(y[99]), .B(x[96]), .Z(n10040) );
  NAND U10525 ( .A(y[16]), .B(x[83]), .Z(n10039) );
  XOR U10526 ( .A(n10040), .B(n10039), .Z(n10042) );
  XOR U10527 ( .A(n10041), .B(n10042), .Z(n10012) );
  AND U10528 ( .A(x[99]), .B(y[96]), .Z(n9929) );
  NAND U10529 ( .A(x[98]), .B(y[97]), .Z(n9928) );
  XNOR U10530 ( .A(n9929), .B(n9928), .Z(n10024) );
  NAND U10531 ( .A(y[98]), .B(x[97]), .Z(n10025) );
  XNOR U10532 ( .A(n10012), .B(n10011), .Z(n10013) );
  XNOR U10533 ( .A(n10014), .B(n10013), .Z(n9975) );
  XOR U10534 ( .A(n9974), .B(n9975), .Z(n9977) );
  NAND U10535 ( .A(n10023), .B(n9930), .Z(n9934) );
  AND U10536 ( .A(n9932), .B(n9931), .Z(n9933) );
  ANDN U10537 ( .B(n9934), .A(n9933), .Z(n10019) );
  AND U10538 ( .A(y[18]), .B(x[81]), .Z(n9988) );
  AND U10539 ( .A(y[17]), .B(x[82]), .Z(n9987) );
  NAND U10540 ( .A(y[138]), .B(x[105]), .Z(n9986) );
  XOR U10541 ( .A(n9987), .B(n9986), .Z(n9989) );
  XOR U10542 ( .A(n9988), .B(n9989), .Z(n10018) );
  AND U10543 ( .A(x[115]), .B(y[176]), .Z(n9936) );
  NAND U10544 ( .A(x[112]), .B(y[179]), .Z(n9935) );
  XNOR U10545 ( .A(n9936), .B(n9935), .Z(n9993) );
  AND U10546 ( .A(x[114]), .B(y[177]), .Z(n10084) );
  NAND U10547 ( .A(x[113]), .B(y[178]), .Z(n9937) );
  XOR U10548 ( .A(n10084), .B(n9937), .Z(n9994) );
  XNOR U10549 ( .A(n9993), .B(n9994), .Z(n10017) );
  XOR U10550 ( .A(n10018), .B(n10017), .Z(n10020) );
  XOR U10551 ( .A(n10019), .B(n10020), .Z(n9976) );
  XOR U10552 ( .A(n9977), .B(n9976), .Z(n9963) );
  XOR U10553 ( .A(n9962), .B(n9963), .Z(n9965) );
  XOR U10554 ( .A(n9964), .B(n9965), .Z(n9958) );
  XOR U10555 ( .A(n9959), .B(n9958), .Z(n9961) );
  NAND U10556 ( .A(n9939), .B(n9938), .Z(n9943) );
  NAND U10557 ( .A(n9941), .B(n9940), .Z(n9942) );
  AND U10558 ( .A(n9943), .B(n9942), .Z(n9971) );
  NANDN U10559 ( .A(n9945), .B(n9944), .Z(n9949) );
  NAND U10560 ( .A(n9947), .B(n9946), .Z(n9948) );
  AND U10561 ( .A(n9949), .B(n9948), .Z(n9981) );
  XNOR U10562 ( .A(n9981), .B(n9980), .Z(n9983) );
  AND U10563 ( .A(y[56]), .B(x[91]), .Z(n10032) );
  AND U10564 ( .A(y[19]), .B(x[80]), .Z(n10031) );
  NAND U10565 ( .A(y[137]), .B(x[106]), .Z(n10030) );
  XOR U10566 ( .A(n10031), .B(n10030), .Z(n10033) );
  XOR U10567 ( .A(n10032), .B(n10033), .Z(n10008) );
  AND U10568 ( .A(y[59]), .B(x[88]), .Z(n10001) );
  AND U10569 ( .A(y[57]), .B(x[90]), .Z(n10000) );
  NAND U10570 ( .A(y[136]), .B(x[107]), .Z(n9999) );
  XOR U10571 ( .A(n10000), .B(n9999), .Z(n10002) );
  XOR U10572 ( .A(n10001), .B(n10002), .Z(n10006) );
  AND U10573 ( .A(y[58]), .B(x[89]), .Z(n10005) );
  XNOR U10574 ( .A(n9983), .B(n9982), .Z(n9969) );
  NAND U10575 ( .A(n9953), .B(n9952), .Z(n9957) );
  NAND U10576 ( .A(n9955), .B(n9954), .Z(n9956) );
  AND U10577 ( .A(n9957), .B(n9956), .Z(n9968) );
  XOR U10578 ( .A(n9969), .B(n9968), .Z(n9970) );
  XNOR U10579 ( .A(n9971), .B(n9970), .Z(n9960) );
  XOR U10580 ( .A(n9961), .B(n9960), .Z(o[99]) );
  NAND U10581 ( .A(n9963), .B(n9962), .Z(n9967) );
  NAND U10582 ( .A(n9965), .B(n9964), .Z(n9966) );
  AND U10583 ( .A(n9967), .B(n9966), .Z(n10051) );
  NAND U10584 ( .A(n9969), .B(n9968), .Z(n9973) );
  NAND U10585 ( .A(n9971), .B(n9970), .Z(n9972) );
  NAND U10586 ( .A(n9973), .B(n9972), .Z(n10049) );
  NAND U10587 ( .A(n9975), .B(n9974), .Z(n9979) );
  NAND U10588 ( .A(n9977), .B(n9976), .Z(n9978) );
  AND U10589 ( .A(n9979), .B(n9978), .Z(n10050) );
  XOR U10590 ( .A(n10049), .B(n10050), .Z(n10052) );
  XOR U10591 ( .A(n10051), .B(n10052), .Z(n10045) );
  XOR U10592 ( .A(n10046), .B(n10045), .Z(n10048) );
  AND U10593 ( .A(y[58]), .B(x[90]), .Z(n10179) );
  AND U10594 ( .A(y[60]), .B(x[88]), .Z(n9985) );
  AND U10595 ( .A(x[91]), .B(y[57]), .Z(n9984) );
  XOR U10596 ( .A(n9985), .B(n9984), .Z(n10116) );
  XOR U10597 ( .A(n10179), .B(n10116), .Z(n10124) );
  AND U10598 ( .A(y[59]), .B(x[89]), .Z(n10123) );
  XOR U10599 ( .A(n10124), .B(n10123), .Z(n10126) );
  AND U10600 ( .A(y[136]), .B(x[108]), .Z(n10076) );
  AND U10601 ( .A(y[19]), .B(x[81]), .Z(n10075) );
  XOR U10602 ( .A(n10076), .B(n10075), .Z(n10078) );
  AND U10603 ( .A(y[20]), .B(x[80]), .Z(n10077) );
  XOR U10604 ( .A(n10078), .B(n10077), .Z(n10125) );
  XOR U10605 ( .A(n10126), .B(n10125), .Z(n10120) );
  NANDN U10606 ( .A(n9987), .B(n9986), .Z(n9991) );
  OR U10607 ( .A(n9989), .B(n9988), .Z(n9990) );
  AND U10608 ( .A(n9991), .B(n9990), .Z(n10118) );
  AND U10609 ( .A(y[179]), .B(x[115]), .Z(n10322) );
  NANDN U10610 ( .A(n9992), .B(n10322), .Z(n9996) );
  NANDN U10611 ( .A(n9994), .B(n9993), .Z(n9995) );
  AND U10612 ( .A(n9996), .B(n9995), .Z(n10117) );
  XNOR U10613 ( .A(n10118), .B(n10117), .Z(n10119) );
  XNOR U10614 ( .A(n10120), .B(n10119), .Z(n10146) );
  AND U10615 ( .A(y[16]), .B(x[84]), .Z(n10101) );
  AND U10616 ( .A(y[138]), .B(x[106]), .Z(n10099) );
  NAND U10617 ( .A(y[100]), .B(x[96]), .Z(n10098) );
  AND U10618 ( .A(y[178]), .B(x[114]), .Z(n9998) );
  AND U10619 ( .A(y[177]), .B(x[113]), .Z(n9997) );
  AND U10620 ( .A(n9998), .B(n9997), .Z(n10095) );
  AND U10621 ( .A(y[180]), .B(x[112]), .Z(n10093) );
  IV U10622 ( .A(n10093), .Z(n10242) );
  AND U10623 ( .A(y[96]), .B(x[100]), .Z(n10092) );
  XNOR U10624 ( .A(n10242), .B(n10092), .Z(n10094) );
  XOR U10625 ( .A(n10095), .B(n10094), .Z(n10061) );
  XOR U10626 ( .A(n10062), .B(n10061), .Z(n10064) );
  NANDN U10627 ( .A(n10000), .B(n9999), .Z(n10004) );
  OR U10628 ( .A(n10002), .B(n10001), .Z(n10003) );
  AND U10629 ( .A(n10004), .B(n10003), .Z(n10063) );
  XOR U10630 ( .A(n10064), .B(n10063), .Z(n10144) );
  NANDN U10631 ( .A(n10006), .B(n10005), .Z(n10010) );
  NANDN U10632 ( .A(n10008), .B(n10007), .Z(n10009) );
  AND U10633 ( .A(n10010), .B(n10009), .Z(n10143) );
  XNOR U10634 ( .A(n10146), .B(n10145), .Z(n10055) );
  XNOR U10635 ( .A(n10056), .B(n10055), .Z(n10058) );
  NANDN U10636 ( .A(n10012), .B(n10011), .Z(n10016) );
  NANDN U10637 ( .A(n10014), .B(n10013), .Z(n10015) );
  AND U10638 ( .A(n10016), .B(n10015), .Z(n10132) );
  NANDN U10639 ( .A(n10018), .B(n10017), .Z(n10022) );
  OR U10640 ( .A(n10020), .B(n10019), .Z(n10021) );
  NAND U10641 ( .A(n10022), .B(n10021), .Z(n10131) );
  AND U10642 ( .A(y[97]), .B(x[99]), .Z(n10029) );
  NAND U10643 ( .A(n10029), .B(n10023), .Z(n10027) );
  NANDN U10644 ( .A(n10025), .B(n10024), .Z(n10026) );
  AND U10645 ( .A(n10027), .B(n10026), .Z(n10138) );
  AND U10646 ( .A(y[56]), .B(x[92]), .Z(n10080) );
  AND U10647 ( .A(y[140]), .B(x[104]), .Z(n10079) );
  XOR U10648 ( .A(n10080), .B(n10079), .Z(n10082) );
  AND U10649 ( .A(y[139]), .B(x[105]), .Z(n10081) );
  XOR U10650 ( .A(n10082), .B(n10081), .Z(n10128) );
  NAND U10651 ( .A(x[98]), .B(y[98]), .Z(n10028) );
  XNOR U10652 ( .A(n10029), .B(n10028), .Z(n10074) );
  AND U10653 ( .A(y[99]), .B(x[97]), .Z(n10073) );
  XOR U10654 ( .A(n10074), .B(n10073), .Z(n10127) );
  XOR U10655 ( .A(n10128), .B(n10127), .Z(n10129) );
  NANDN U10656 ( .A(n10031), .B(n10030), .Z(n10035) );
  OR U10657 ( .A(n10033), .B(n10032), .Z(n10034) );
  NAND U10658 ( .A(n10035), .B(n10034), .Z(n10130) );
  XNOR U10659 ( .A(n10129), .B(n10130), .Z(n10137) );
  AND U10660 ( .A(y[18]), .B(x[82]), .Z(n10112) );
  AND U10661 ( .A(y[137]), .B(x[107]), .Z(n10110) );
  NAND U10662 ( .A(y[17]), .B(x[83]), .Z(n10109) );
  AND U10663 ( .A(x[116]), .B(y[176]), .Z(n10037) );
  NAND U10664 ( .A(x[113]), .B(y[179]), .Z(n10036) );
  XNOR U10665 ( .A(n10037), .B(n10036), .Z(n10088) );
  AND U10666 ( .A(x[115]), .B(y[177]), .Z(n10204) );
  NAND U10667 ( .A(x[114]), .B(y[178]), .Z(n10038) );
  XOR U10668 ( .A(n10204), .B(n10038), .Z(n10089) );
  XOR U10669 ( .A(n10068), .B(n10067), .Z(n10069) );
  NANDN U10670 ( .A(n10040), .B(n10039), .Z(n10044) );
  OR U10671 ( .A(n10042), .B(n10041), .Z(n10043) );
  NAND U10672 ( .A(n10044), .B(n10043), .Z(n10070) );
  XOR U10673 ( .A(n10069), .B(n10070), .Z(n10140) );
  XOR U10674 ( .A(n10134), .B(n10133), .Z(n10057) );
  XNOR U10675 ( .A(n10058), .B(n10057), .Z(n10047) );
  XNOR U10676 ( .A(n10048), .B(n10047), .Z(o[100]) );
  NAND U10677 ( .A(n10050), .B(n10049), .Z(n10054) );
  NAND U10678 ( .A(n10052), .B(n10051), .Z(n10053) );
  NAND U10679 ( .A(n10054), .B(n10053), .Z(n10280) );
  XNOR U10680 ( .A(n10279), .B(n10280), .Z(n10282) );
  NANDN U10681 ( .A(n10056), .B(n10055), .Z(n10060) );
  NAND U10682 ( .A(n10058), .B(n10057), .Z(n10059) );
  AND U10683 ( .A(n10060), .B(n10059), .Z(n10150) );
  NAND U10684 ( .A(n10062), .B(n10061), .Z(n10066) );
  NAND U10685 ( .A(n10064), .B(n10063), .Z(n10065) );
  NAND U10686 ( .A(n10066), .B(n10065), .Z(n10205) );
  NAND U10687 ( .A(n10068), .B(n10067), .Z(n10072) );
  NANDN U10688 ( .A(n10070), .B(n10069), .Z(n10071) );
  NAND U10689 ( .A(n10072), .B(n10071), .Z(n10206) );
  XOR U10690 ( .A(n10205), .B(n10206), .Z(n10209) );
  AND U10691 ( .A(y[98]), .B(x[99]), .Z(n10108) );
  IV U10692 ( .A(n10108), .Z(n10198) );
  AND U10693 ( .A(y[141]), .B(x[104]), .Z(n10495) );
  AND U10694 ( .A(y[56]), .B(x[93]), .Z(n10187) );
  AND U10695 ( .A(y[99]), .B(x[98]), .Z(n10186) );
  XOR U10696 ( .A(n10187), .B(n10186), .Z(n10188) );
  XOR U10697 ( .A(n10495), .B(n10188), .Z(n10183) );
  AND U10698 ( .A(y[137]), .B(x[108]), .Z(n10192) );
  AND U10699 ( .A(y[16]), .B(x[85]), .Z(n10191) );
  XOR U10700 ( .A(n10192), .B(n10191), .Z(n10193) );
  AND U10701 ( .A(y[17]), .B(x[84]), .Z(n10447) );
  XOR U10702 ( .A(n10193), .B(n10447), .Z(n10182) );
  XOR U10703 ( .A(n10183), .B(n10182), .Z(n10185) );
  XOR U10704 ( .A(n10184), .B(n10185), .Z(n10166) );
  XOR U10705 ( .A(n10165), .B(n10166), .Z(n10168) );
  AND U10706 ( .A(y[178]), .B(x[115]), .Z(n10083) );
  AND U10707 ( .A(n10084), .B(n10083), .Z(n10244) );
  AND U10708 ( .A(x[112]), .B(y[181]), .Z(n10086) );
  AND U10709 ( .A(x[113]), .B(y[180]), .Z(n10085) );
  XOR U10710 ( .A(n10086), .B(n10085), .Z(n10243) );
  XOR U10711 ( .A(n10244), .B(n10243), .Z(n10262) );
  AND U10712 ( .A(y[61]), .B(x[88]), .Z(n10270) );
  AND U10713 ( .A(y[20]), .B(x[81]), .Z(n10269) );
  XOR U10714 ( .A(n10270), .B(n10269), .Z(n10272) );
  AND U10715 ( .A(y[57]), .B(x[92]), .Z(n10271) );
  XOR U10716 ( .A(n10272), .B(n10271), .Z(n10261) );
  XOR U10717 ( .A(n10262), .B(n10261), .Z(n10264) );
  XOR U10718 ( .A(n10263), .B(n10264), .Z(n10167) );
  XOR U10719 ( .A(n10168), .B(n10167), .Z(n10208) );
  XOR U10720 ( .A(n10209), .B(n10208), .Z(n10156) );
  AND U10721 ( .A(y[179]), .B(x[116]), .Z(n10473) );
  NAND U10722 ( .A(n10473), .B(n10087), .Z(n10091) );
  NANDN U10723 ( .A(n10089), .B(n10088), .Z(n10090) );
  NAND U10724 ( .A(n10091), .B(n10090), .Z(n10217) );
  IV U10725 ( .A(n10092), .Z(n10196) );
  NANDN U10726 ( .A(n10093), .B(n10196), .Z(n10097) );
  NANDN U10727 ( .A(n10095), .B(n10094), .Z(n10096) );
  AND U10728 ( .A(n10097), .B(n10096), .Z(n10218) );
  XOR U10729 ( .A(n10217), .B(n10218), .Z(n10220) );
  NANDN U10730 ( .A(n10099), .B(n10098), .Z(n10103) );
  NANDN U10731 ( .A(n10101), .B(n10100), .Z(n10102) );
  AND U10732 ( .A(n10103), .B(n10102), .Z(n10224) );
  AND U10733 ( .A(y[58]), .B(x[91]), .Z(n10395) );
  NAND U10734 ( .A(x[90]), .B(y[59]), .Z(n10104) );
  XNOR U10735 ( .A(n10395), .B(n10104), .Z(n10181) );
  AND U10736 ( .A(y[60]), .B(x[89]), .Z(n10180) );
  XOR U10737 ( .A(n10181), .B(n10180), .Z(n10222) );
  AND U10738 ( .A(y[179]), .B(x[114]), .Z(n10172) );
  AND U10739 ( .A(y[176]), .B(x[117]), .Z(n10171) );
  XOR U10740 ( .A(n10172), .B(n10171), .Z(n10174) );
  AND U10741 ( .A(y[177]), .B(x[116]), .Z(n10455) );
  NAND U10742 ( .A(x[115]), .B(y[178]), .Z(n10105) );
  XNOR U10743 ( .A(n10455), .B(n10105), .Z(n10173) );
  XOR U10744 ( .A(n10174), .B(n10173), .Z(n10221) );
  XOR U10745 ( .A(n10222), .B(n10221), .Z(n10223) );
  XOR U10746 ( .A(n10224), .B(n10223), .Z(n10219) );
  XOR U10747 ( .A(n10220), .B(n10219), .Z(n10234) );
  AND U10748 ( .A(x[101]), .B(y[96]), .Z(n10107) );
  NAND U10749 ( .A(x[100]), .B(y[97]), .Z(n10106) );
  XNOR U10750 ( .A(n10107), .B(n10106), .Z(n10197) );
  XOR U10751 ( .A(n10197), .B(n10108), .Z(n10256) );
  AND U10752 ( .A(y[136]), .B(x[109]), .Z(n10176) );
  AND U10753 ( .A(y[18]), .B(x[83]), .Z(n10175) );
  XOR U10754 ( .A(n10176), .B(n10175), .Z(n10178) );
  AND U10755 ( .A(y[19]), .B(x[82]), .Z(n10177) );
  XOR U10756 ( .A(n10178), .B(n10177), .Z(n10255) );
  XOR U10757 ( .A(n10256), .B(n10255), .Z(n10258) );
  NANDN U10758 ( .A(n10110), .B(n10109), .Z(n10114) );
  NANDN U10759 ( .A(n10112), .B(n10111), .Z(n10113) );
  AND U10760 ( .A(n10114), .B(n10113), .Z(n10257) );
  XOR U10761 ( .A(n10258), .B(n10257), .Z(n10232) );
  AND U10762 ( .A(y[60]), .B(x[91]), .Z(n10472) );
  AND U10763 ( .A(y[100]), .B(x[97]), .Z(n10501) );
  AND U10764 ( .A(y[138]), .B(x[107]), .Z(n10237) );
  XOR U10765 ( .A(n10501), .B(n10237), .Z(n10239) );
  AND U10766 ( .A(y[101]), .B(x[96]), .Z(n10238) );
  XOR U10767 ( .A(n10239), .B(n10238), .Z(n10214) );
  AND U10768 ( .A(y[21]), .B(x[80]), .Z(n10248) );
  AND U10769 ( .A(y[140]), .B(x[105]), .Z(n10247) );
  XOR U10770 ( .A(n10248), .B(n10247), .Z(n10250) );
  AND U10771 ( .A(y[139]), .B(x[106]), .Z(n10249) );
  XOR U10772 ( .A(n10250), .B(n10249), .Z(n10213) );
  XOR U10773 ( .A(n10214), .B(n10213), .Z(n10216) );
  XOR U10774 ( .A(n10215), .B(n10216), .Z(n10231) );
  XOR U10775 ( .A(n10232), .B(n10231), .Z(n10233) );
  XOR U10776 ( .A(n10234), .B(n10233), .Z(n10153) );
  NANDN U10777 ( .A(n10118), .B(n10117), .Z(n10122) );
  NANDN U10778 ( .A(n10120), .B(n10119), .Z(n10121) );
  AND U10779 ( .A(n10122), .B(n10121), .Z(n10229) );
  XNOR U10780 ( .A(n10227), .B(n10228), .Z(n10230) );
  XNOR U10781 ( .A(n10229), .B(n10230), .Z(n10154) );
  XOR U10782 ( .A(n10153), .B(n10154), .Z(n10155) );
  XOR U10783 ( .A(n10156), .B(n10155), .Z(n10149) );
  XNOR U10784 ( .A(n10150), .B(n10149), .Z(n10152) );
  NANDN U10785 ( .A(n10132), .B(n10131), .Z(n10136) );
  NAND U10786 ( .A(n10134), .B(n10133), .Z(n10135) );
  AND U10787 ( .A(n10136), .B(n10135), .Z(n10162) );
  NANDN U10788 ( .A(n10138), .B(n10137), .Z(n10142) );
  NANDN U10789 ( .A(n10140), .B(n10139), .Z(n10141) );
  AND U10790 ( .A(n10142), .B(n10141), .Z(n10160) );
  NANDN U10791 ( .A(n10144), .B(n10143), .Z(n10148) );
  NAND U10792 ( .A(n10146), .B(n10145), .Z(n10147) );
  AND U10793 ( .A(n10148), .B(n10147), .Z(n10159) );
  XOR U10794 ( .A(n10152), .B(n10151), .Z(n10281) );
  XOR U10795 ( .A(n10282), .B(n10281), .Z(o[101]) );
  NAND U10796 ( .A(n10154), .B(n10153), .Z(n10158) );
  NAND U10797 ( .A(n10156), .B(n10155), .Z(n10157) );
  AND U10798 ( .A(n10158), .B(n10157), .Z(n10571) );
  NANDN U10799 ( .A(n10160), .B(n10159), .Z(n10164) );
  NANDN U10800 ( .A(n10162), .B(n10161), .Z(n10163) );
  NAND U10801 ( .A(n10164), .B(n10163), .Z(n10572) );
  NAND U10802 ( .A(n10166), .B(n10165), .Z(n10170) );
  NAND U10803 ( .A(n10168), .B(n10167), .Z(n10169) );
  AND U10804 ( .A(n10170), .B(n10169), .Z(n10560) );
  AND U10805 ( .A(y[139]), .B(x[107]), .Z(n10415) );
  AND U10806 ( .A(y[99]), .B(x[99]), .Z(n10414) );
  XOR U10807 ( .A(n10415), .B(n10414), .Z(n10413) );
  AND U10808 ( .A(y[19]), .B(x[83]), .Z(n10412) );
  XOR U10809 ( .A(n10413), .B(n10412), .Z(n10523) );
  AND U10810 ( .A(y[140]), .B(x[106]), .Z(n10487) );
  AND U10811 ( .A(y[98]), .B(x[100]), .Z(n10486) );
  XOR U10812 ( .A(n10487), .B(n10486), .Z(n10485) );
  AND U10813 ( .A(y[20]), .B(x[82]), .Z(n10484) );
  XNOR U10814 ( .A(n10485), .B(n10484), .Z(n10522) );
  XNOR U10815 ( .A(n10521), .B(n10520), .Z(n10313) );
  XOR U10816 ( .A(n10314), .B(n10313), .Z(n10312) );
  XOR U10817 ( .A(n10311), .B(n10312), .Z(n10294) );
  XOR U10818 ( .A(n10294), .B(n10293), .Z(n10292) );
  NAND U10819 ( .A(n10187), .B(n10186), .Z(n10190) );
  NAND U10820 ( .A(n10495), .B(n10188), .Z(n10189) );
  NAND U10821 ( .A(n10190), .B(n10189), .Z(n10429) );
  NAND U10822 ( .A(n10192), .B(n10191), .Z(n10195) );
  NAND U10823 ( .A(n10193), .B(n10447), .Z(n10194) );
  NAND U10824 ( .A(n10195), .B(n10194), .Z(n10428) );
  XOR U10825 ( .A(n10429), .B(n10428), .Z(n10427) );
  AND U10826 ( .A(y[97]), .B(x[101]), .Z(n10459) );
  NANDN U10827 ( .A(n10196), .B(n10459), .Z(n10200) );
  NANDN U10828 ( .A(n10198), .B(n10197), .Z(n10199) );
  AND U10829 ( .A(n10200), .B(n10199), .Z(n10515) );
  AND U10830 ( .A(x[84]), .B(y[18]), .Z(n10202) );
  NAND U10831 ( .A(x[85]), .B(y[17]), .Z(n10201) );
  XNOR U10832 ( .A(n10202), .B(n10201), .Z(n10445) );
  AND U10833 ( .A(y[136]), .B(x[110]), .Z(n10444) );
  XOR U10834 ( .A(n10445), .B(n10444), .Z(n10517) );
  AND U10835 ( .A(y[181]), .B(x[113]), .Z(n10399) );
  AND U10836 ( .A(y[178]), .B(x[116]), .Z(n10203) );
  AND U10837 ( .A(n10204), .B(n10203), .Z(n10401) );
  AND U10838 ( .A(y[180]), .B(x[114]), .Z(n10400) );
  XOR U10839 ( .A(n10401), .B(n10400), .Z(n10398) );
  XNOR U10840 ( .A(n10399), .B(n10398), .Z(n10516) );
  XNOR U10841 ( .A(n10515), .B(n10514), .Z(n10426) );
  XOR U10842 ( .A(n10427), .B(n10426), .Z(n10291) );
  XOR U10843 ( .A(n10292), .B(n10291), .Z(n10288) );
  IV U10844 ( .A(n10205), .Z(n10207) );
  NANDN U10845 ( .A(n10207), .B(n10206), .Z(n10212) );
  IV U10846 ( .A(n10208), .Z(n10210) );
  NANDN U10847 ( .A(n10210), .B(n10209), .Z(n10211) );
  AND U10848 ( .A(n10212), .B(n10211), .Z(n10287) );
  XOR U10849 ( .A(n10300), .B(n10299), .Z(n10298) );
  NAND U10850 ( .A(n10222), .B(n10221), .Z(n10226) );
  NAND U10851 ( .A(n10224), .B(n10223), .Z(n10225) );
  AND U10852 ( .A(n10226), .B(n10225), .Z(n10297) );
  XOR U10853 ( .A(n10298), .B(n10297), .Z(n10285) );
  XOR U10854 ( .A(n10286), .B(n10285), .Z(n10559) );
  XOR U10855 ( .A(n10560), .B(n10559), .Z(n10558) );
  OR U10856 ( .A(n10232), .B(n10231), .Z(n10236) );
  NANDN U10857 ( .A(n10234), .B(n10233), .Z(n10235) );
  NAND U10858 ( .A(n10236), .B(n10235), .Z(n10535) );
  AND U10859 ( .A(n10501), .B(n10237), .Z(n10241) );
  NAND U10860 ( .A(n10239), .B(n10238), .Z(n10240) );
  NANDN U10861 ( .A(n10241), .B(n10240), .Z(n10309) );
  NANDN U10862 ( .A(n10242), .B(n10399), .Z(n10246) );
  NAND U10863 ( .A(n10244), .B(n10243), .Z(n10245) );
  NAND U10864 ( .A(n10246), .B(n10245), .Z(n10307) );
  NAND U10865 ( .A(n10248), .B(n10247), .Z(n10252) );
  NAND U10866 ( .A(n10250), .B(n10249), .Z(n10251) );
  AND U10867 ( .A(n10252), .B(n10251), .Z(n10316) );
  AND U10868 ( .A(y[21]), .B(x[81]), .Z(n10481) );
  AND U10869 ( .A(y[56]), .B(x[94]), .Z(n10480) );
  XOR U10870 ( .A(n10481), .B(n10480), .Z(n10479) );
  AND U10871 ( .A(y[62]), .B(x[88]), .Z(n10478) );
  XOR U10872 ( .A(n10479), .B(n10478), .Z(n10318) );
  AND U10873 ( .A(x[117]), .B(y[177]), .Z(n10254) );
  NAND U10874 ( .A(x[116]), .B(y[178]), .Z(n10253) );
  XNOR U10875 ( .A(n10254), .B(n10253), .Z(n10324) );
  AND U10876 ( .A(y[176]), .B(x[118]), .Z(n10323) );
  XOR U10877 ( .A(n10324), .B(n10323), .Z(n10321) );
  XNOR U10878 ( .A(n10322), .B(n10321), .Z(n10317) );
  XNOR U10879 ( .A(n10316), .B(n10315), .Z(n10308) );
  XOR U10880 ( .A(n10307), .B(n10308), .Z(n10310) );
  XOR U10881 ( .A(n10309), .B(n10310), .Z(n10539) );
  NAND U10882 ( .A(n10256), .B(n10255), .Z(n10260) );
  NAND U10883 ( .A(n10258), .B(n10257), .Z(n10259) );
  AND U10884 ( .A(n10260), .B(n10259), .Z(n10540) );
  NAND U10885 ( .A(n10262), .B(n10261), .Z(n10266) );
  NAND U10886 ( .A(n10264), .B(n10263), .Z(n10265) );
  AND U10887 ( .A(n10266), .B(n10265), .Z(n10304) );
  AND U10888 ( .A(y[102]), .B(x[96]), .Z(n10409) );
  AND U10889 ( .A(y[16]), .B(x[86]), .Z(n10408) );
  XOR U10890 ( .A(n10409), .B(n10408), .Z(n10407) );
  AND U10891 ( .A(y[137]), .B(x[109]), .Z(n10406) );
  XOR U10892 ( .A(n10407), .B(n10406), .Z(n10435) );
  AND U10893 ( .A(y[57]), .B(x[93]), .Z(n10441) );
  AND U10894 ( .A(y[60]), .B(x[90]), .Z(n10440) );
  XOR U10895 ( .A(n10441), .B(n10440), .Z(n10439) );
  AND U10896 ( .A(y[61]), .B(x[89]), .Z(n10438) );
  XOR U10897 ( .A(n10439), .B(n10438), .Z(n10393) );
  AND U10898 ( .A(x[92]), .B(y[58]), .Z(n10268) );
  NAND U10899 ( .A(x[91]), .B(y[59]), .Z(n10267) );
  XNOR U10900 ( .A(n10268), .B(n10267), .Z(n10392) );
  XOR U10901 ( .A(n10393), .B(n10392), .Z(n10434) );
  XOR U10902 ( .A(n10435), .B(n10434), .Z(n10433) );
  AND U10903 ( .A(y[182]), .B(x[112]), .Z(n10458) );
  XOR U10904 ( .A(n10459), .B(n10458), .Z(n10457) );
  AND U10905 ( .A(y[96]), .B(x[102]), .Z(n10456) );
  XOR U10906 ( .A(n10457), .B(n10456), .Z(n10432) );
  XOR U10907 ( .A(n10433), .B(n10432), .Z(n10306) );
  NAND U10908 ( .A(n10270), .B(n10269), .Z(n10274) );
  NAND U10909 ( .A(n10272), .B(n10271), .Z(n10273) );
  AND U10910 ( .A(n10274), .B(n10273), .Z(n10386) );
  AND U10911 ( .A(y[138]), .B(x[108]), .Z(n10499) );
  AND U10912 ( .A(x[97]), .B(y[101]), .Z(n10276) );
  AND U10913 ( .A(x[98]), .B(y[100]), .Z(n10275) );
  XOR U10914 ( .A(n10276), .B(n10275), .Z(n10498) );
  XOR U10915 ( .A(n10499), .B(n10498), .Z(n10389) );
  AND U10916 ( .A(y[22]), .B(x[80]), .Z(n10493) );
  AND U10917 ( .A(y[142]), .B(x[104]), .Z(n10278) );
  AND U10918 ( .A(x[105]), .B(y[141]), .Z(n10277) );
  XOR U10919 ( .A(n10278), .B(n10277), .Z(n10492) );
  XNOR U10920 ( .A(n10493), .B(n10492), .Z(n10388) );
  XNOR U10921 ( .A(n10386), .B(n10387), .Z(n10305) );
  XOR U10922 ( .A(n10304), .B(n10303), .Z(n10541) );
  XOR U10923 ( .A(n10542), .B(n10541), .Z(n10536) );
  XOR U10924 ( .A(n10535), .B(n10536), .Z(n10533) );
  XOR U10925 ( .A(n10534), .B(n10533), .Z(n10557) );
  XOR U10926 ( .A(n10558), .B(n10557), .Z(n10569) );
  XNOR U10927 ( .A(n10570), .B(n10569), .Z(n10553) );
  NANDN U10928 ( .A(n10280), .B(n10279), .Z(n10284) );
  NAND U10929 ( .A(n10282), .B(n10281), .Z(n10283) );
  NAND U10930 ( .A(n10284), .B(n10283), .Z(n10551) );
  XOR U10931 ( .A(n10552), .B(n10551), .Z(o[102]) );
  NAND U10932 ( .A(n10286), .B(n10285), .Z(n10290) );
  NANDN U10933 ( .A(n10288), .B(n10287), .Z(n10289) );
  AND U10934 ( .A(n10290), .B(n10289), .Z(n10568) );
  NAND U10935 ( .A(n10292), .B(n10291), .Z(n10296) );
  NAND U10936 ( .A(n10294), .B(n10293), .Z(n10295) );
  AND U10937 ( .A(n10296), .B(n10295), .Z(n10550) );
  NAND U10938 ( .A(n10298), .B(n10297), .Z(n10302) );
  NAND U10939 ( .A(n10300), .B(n10299), .Z(n10301) );
  AND U10940 ( .A(n10302), .B(n10301), .Z(n10532) );
  NAND U10941 ( .A(n10316), .B(n10315), .Z(n10320) );
  NANDN U10942 ( .A(n10318), .B(n10317), .Z(n10319) );
  NAND U10943 ( .A(n10322), .B(n10321), .Z(n10326) );
  NAND U10944 ( .A(n10324), .B(n10323), .Z(n10325) );
  AND U10945 ( .A(n10326), .B(n10325), .Z(n10385) );
  AND U10946 ( .A(x[94]), .B(y[57]), .Z(n10328) );
  NAND U10947 ( .A(x[100]), .B(y[99]), .Z(n10327) );
  XNOR U10948 ( .A(n10328), .B(n10327), .Z(n10332) );
  AND U10949 ( .A(x[112]), .B(y[183]), .Z(n10330) );
  NAND U10950 ( .A(x[99]), .B(y[100]), .Z(n10329) );
  XNOR U10951 ( .A(n10330), .B(n10329), .Z(n10331) );
  XOR U10952 ( .A(n10332), .B(n10331), .Z(n10340) );
  AND U10953 ( .A(x[118]), .B(y[177]), .Z(n10334) );
  NAND U10954 ( .A(x[101]), .B(y[98]), .Z(n10333) );
  XNOR U10955 ( .A(n10334), .B(n10333), .Z(n10338) );
  AND U10956 ( .A(x[109]), .B(y[138]), .Z(n10336) );
  NAND U10957 ( .A(x[83]), .B(y[20]), .Z(n10335) );
  XNOR U10958 ( .A(n10336), .B(n10335), .Z(n10337) );
  XNOR U10959 ( .A(n10338), .B(n10337), .Z(n10339) );
  XNOR U10960 ( .A(n10340), .B(n10339), .Z(n10383) );
  AND U10961 ( .A(x[115]), .B(y[180]), .Z(n10345) );
  AND U10962 ( .A(y[142]), .B(x[105]), .Z(n10494) );
  AND U10963 ( .A(x[81]), .B(y[22]), .Z(n10342) );
  NAND U10964 ( .A(x[114]), .B(y[181]), .Z(n10341) );
  XNOR U10965 ( .A(n10342), .B(n10341), .Z(n10343) );
  XNOR U10966 ( .A(n10494), .B(n10343), .Z(n10344) );
  XNOR U10967 ( .A(n10345), .B(n10344), .Z(n10361) );
  AND U10968 ( .A(x[119]), .B(y[176]), .Z(n10347) );
  NAND U10969 ( .A(x[110]), .B(y[137]), .Z(n10346) );
  XNOR U10970 ( .A(n10347), .B(n10346), .Z(n10351) );
  AND U10971 ( .A(x[96]), .B(y[103]), .Z(n10349) );
  NAND U10972 ( .A(x[82]), .B(y[21]), .Z(n10348) );
  XNOR U10973 ( .A(n10349), .B(n10348), .Z(n10350) );
  XOR U10974 ( .A(n10351), .B(n10350), .Z(n10359) );
  AND U10975 ( .A(x[88]), .B(y[63]), .Z(n10353) );
  NAND U10976 ( .A(x[107]), .B(y[140]), .Z(n10352) );
  XNOR U10977 ( .A(n10353), .B(n10352), .Z(n10357) );
  AND U10978 ( .A(x[84]), .B(y[19]), .Z(n10355) );
  NAND U10979 ( .A(x[111]), .B(y[136]), .Z(n10354) );
  XNOR U10980 ( .A(n10355), .B(n10354), .Z(n10356) );
  XNOR U10981 ( .A(n10357), .B(n10356), .Z(n10358) );
  XNOR U10982 ( .A(n10359), .B(n10358), .Z(n10360) );
  XOR U10983 ( .A(n10361), .B(n10360), .Z(n10381) );
  AND U10984 ( .A(x[80]), .B(y[23]), .Z(n10363) );
  NAND U10985 ( .A(x[87]), .B(y[16]), .Z(n10362) );
  XNOR U10986 ( .A(n10363), .B(n10362), .Z(n10367) );
  AND U10987 ( .A(x[113]), .B(y[182]), .Z(n10365) );
  NAND U10988 ( .A(x[97]), .B(y[102]), .Z(n10364) );
  XNOR U10989 ( .A(n10365), .B(n10364), .Z(n10366) );
  XOR U10990 ( .A(n10367), .B(n10366), .Z(n10375) );
  AND U10991 ( .A(x[103]), .B(y[96]), .Z(n10369) );
  NAND U10992 ( .A(x[86]), .B(y[17]), .Z(n10368) );
  XNOR U10993 ( .A(n10369), .B(n10368), .Z(n10373) );
  AND U10994 ( .A(x[108]), .B(y[139]), .Z(n10371) );
  NAND U10995 ( .A(x[102]), .B(y[97]), .Z(n10370) );
  XNOR U10996 ( .A(n10371), .B(n10370), .Z(n10372) );
  XNOR U10997 ( .A(n10373), .B(n10372), .Z(n10374) );
  XNOR U10998 ( .A(n10375), .B(n10374), .Z(n10379) );
  AND U10999 ( .A(y[59]), .B(x[92]), .Z(n10394) );
  AND U11000 ( .A(y[101]), .B(x[98]), .Z(n10500) );
  XOR U11001 ( .A(n10394), .B(n10500), .Z(n10377) );
  AND U11002 ( .A(y[18]), .B(x[85]), .Z(n10446) );
  AND U11003 ( .A(y[178]), .B(x[117]), .Z(n10454) );
  XNOR U11004 ( .A(n10446), .B(n10454), .Z(n10376) );
  XNOR U11005 ( .A(n10377), .B(n10376), .Z(n10378) );
  XNOR U11006 ( .A(n10379), .B(n10378), .Z(n10380) );
  XNOR U11007 ( .A(n10381), .B(n10380), .Z(n10382) );
  XNOR U11008 ( .A(n10383), .B(n10382), .Z(n10384) );
  XNOR U11009 ( .A(n10385), .B(n10384), .Z(n10425) );
  NANDN U11010 ( .A(n10387), .B(n10386), .Z(n10391) );
  NANDN U11011 ( .A(n10389), .B(n10388), .Z(n10390) );
  AND U11012 ( .A(n10391), .B(n10390), .Z(n10423) );
  NAND U11013 ( .A(n10393), .B(n10392), .Z(n10397) );
  NAND U11014 ( .A(n10395), .B(n10394), .Z(n10396) );
  AND U11015 ( .A(n10397), .B(n10396), .Z(n10405) );
  NAND U11016 ( .A(n10399), .B(n10398), .Z(n10403) );
  NAND U11017 ( .A(n10401), .B(n10400), .Z(n10402) );
  NAND U11018 ( .A(n10403), .B(n10402), .Z(n10404) );
  XNOR U11019 ( .A(n10405), .B(n10404), .Z(n10421) );
  NAND U11020 ( .A(n10407), .B(n10406), .Z(n10411) );
  NAND U11021 ( .A(n10409), .B(n10408), .Z(n10410) );
  AND U11022 ( .A(n10411), .B(n10410), .Z(n10419) );
  NAND U11023 ( .A(n10413), .B(n10412), .Z(n10417) );
  NAND U11024 ( .A(n10415), .B(n10414), .Z(n10416) );
  NAND U11025 ( .A(n10417), .B(n10416), .Z(n10418) );
  XNOR U11026 ( .A(n10419), .B(n10418), .Z(n10420) );
  XNOR U11027 ( .A(n10421), .B(n10420), .Z(n10422) );
  XNOR U11028 ( .A(n10423), .B(n10422), .Z(n10424) );
  NAND U11029 ( .A(n10427), .B(n10426), .Z(n10431) );
  NAND U11030 ( .A(n10429), .B(n10428), .Z(n10430) );
  NAND U11031 ( .A(n10433), .B(n10432), .Z(n10437) );
  NAND U11032 ( .A(n10435), .B(n10434), .Z(n10436) );
  AND U11033 ( .A(n10437), .B(n10436), .Z(n10513) );
  NAND U11034 ( .A(n10439), .B(n10438), .Z(n10443) );
  NAND U11035 ( .A(n10441), .B(n10440), .Z(n10442) );
  AND U11036 ( .A(n10443), .B(n10442), .Z(n10451) );
  NAND U11037 ( .A(n10445), .B(n10444), .Z(n10449) );
  NAND U11038 ( .A(n10447), .B(n10446), .Z(n10448) );
  NAND U11039 ( .A(n10449), .B(n10448), .Z(n10450) );
  XNOR U11040 ( .A(n10451), .B(n10450), .Z(n10511) );
  AND U11041 ( .A(x[104]), .B(y[143]), .Z(n10453) );
  NAND U11042 ( .A(x[89]), .B(y[62]), .Z(n10452) );
  XNOR U11043 ( .A(n10453), .B(n10452), .Z(n10477) );
  AND U11044 ( .A(n10455), .B(n10454), .Z(n10471) );
  NAND U11045 ( .A(n10457), .B(n10456), .Z(n10461) );
  NAND U11046 ( .A(n10459), .B(n10458), .Z(n10460) );
  AND U11047 ( .A(n10461), .B(n10460), .Z(n10469) );
  AND U11048 ( .A(x[93]), .B(y[58]), .Z(n10463) );
  NAND U11049 ( .A(x[90]), .B(y[61]), .Z(n10462) );
  XNOR U11050 ( .A(n10463), .B(n10462), .Z(n10467) );
  AND U11051 ( .A(x[95]), .B(y[56]), .Z(n10465) );
  NAND U11052 ( .A(x[106]), .B(y[141]), .Z(n10464) );
  XNOR U11053 ( .A(n10465), .B(n10464), .Z(n10466) );
  XNOR U11054 ( .A(n10467), .B(n10466), .Z(n10468) );
  XNOR U11055 ( .A(n10469), .B(n10468), .Z(n10470) );
  XOR U11056 ( .A(n10471), .B(n10470), .Z(n10475) );
  XNOR U11057 ( .A(n10473), .B(n10472), .Z(n10474) );
  XNOR U11058 ( .A(n10475), .B(n10474), .Z(n10476) );
  XOR U11059 ( .A(n10477), .B(n10476), .Z(n10509) );
  NAND U11060 ( .A(n10479), .B(n10478), .Z(n10483) );
  NAND U11061 ( .A(n10481), .B(n10480), .Z(n10482) );
  AND U11062 ( .A(n10483), .B(n10482), .Z(n10491) );
  NAND U11063 ( .A(n10485), .B(n10484), .Z(n10489) );
  NAND U11064 ( .A(n10487), .B(n10486), .Z(n10488) );
  NAND U11065 ( .A(n10489), .B(n10488), .Z(n10490) );
  XNOR U11066 ( .A(n10491), .B(n10490), .Z(n10507) );
  NAND U11067 ( .A(n10493), .B(n10492), .Z(n10497) );
  NAND U11068 ( .A(n10495), .B(n10494), .Z(n10496) );
  AND U11069 ( .A(n10497), .B(n10496), .Z(n10505) );
  NAND U11070 ( .A(n10499), .B(n10498), .Z(n10503) );
  NAND U11071 ( .A(n10501), .B(n10500), .Z(n10502) );
  NAND U11072 ( .A(n10503), .B(n10502), .Z(n10504) );
  XNOR U11073 ( .A(n10505), .B(n10504), .Z(n10506) );
  XNOR U11074 ( .A(n10507), .B(n10506), .Z(n10508) );
  XNOR U11075 ( .A(n10509), .B(n10508), .Z(n10510) );
  XNOR U11076 ( .A(n10511), .B(n10510), .Z(n10512) );
  XNOR U11077 ( .A(n10513), .B(n10512), .Z(n10529) );
  NAND U11078 ( .A(n10515), .B(n10514), .Z(n10519) );
  NANDN U11079 ( .A(n10517), .B(n10516), .Z(n10518) );
  AND U11080 ( .A(n10519), .B(n10518), .Z(n10527) );
  NAND U11081 ( .A(n10521), .B(n10520), .Z(n10525) );
  NANDN U11082 ( .A(n10523), .B(n10522), .Z(n10524) );
  NAND U11083 ( .A(n10525), .B(n10524), .Z(n10526) );
  XNOR U11084 ( .A(n10527), .B(n10526), .Z(n10528) );
  XNOR U11085 ( .A(n10529), .B(n10528), .Z(n10530) );
  XNOR U11086 ( .A(n10532), .B(n10531), .Z(n10548) );
  NAND U11087 ( .A(n10534), .B(n10533), .Z(n10538) );
  AND U11088 ( .A(n10536), .B(n10535), .Z(n10537) );
  ANDN U11089 ( .B(n10538), .A(n10537), .Z(n10546) );
  ANDN U11090 ( .B(n10540), .A(n10539), .Z(n10544) );
  AND U11091 ( .A(n10542), .B(n10541), .Z(n10543) );
  OR U11092 ( .A(n10544), .B(n10543), .Z(n10545) );
  XNOR U11093 ( .A(n10546), .B(n10545), .Z(n10547) );
  XNOR U11094 ( .A(n10548), .B(n10547), .Z(n10549) );
  XNOR U11095 ( .A(n10550), .B(n10549), .Z(n10566) );
  NAND U11096 ( .A(n10552), .B(n10551), .Z(n10556) );
  NANDN U11097 ( .A(n10554), .B(n10553), .Z(n10555) );
  AND U11098 ( .A(n10556), .B(n10555), .Z(n10564) );
  NAND U11099 ( .A(n10558), .B(n10557), .Z(n10562) );
  NAND U11100 ( .A(n10560), .B(n10559), .Z(n10561) );
  NAND U11101 ( .A(n10562), .B(n10561), .Z(n10563) );
  XNOR U11102 ( .A(n10564), .B(n10563), .Z(n10565) );
  XNOR U11103 ( .A(n10566), .B(n10565), .Z(n10567) );
  XNOR U11104 ( .A(n10568), .B(n10567), .Z(n10576) );
  NAND U11105 ( .A(n10570), .B(n10569), .Z(n10574) );
  NANDN U11106 ( .A(n10572), .B(n10571), .Z(n10573) );
  NAND U11107 ( .A(n10574), .B(n10573), .Z(n10575) );
  XNOR U11108 ( .A(n10576), .B(n10575), .Z(o[103]) );
  AND U11109 ( .A(y[184]), .B(x[112]), .Z(n10580) );
  IV U11110 ( .A(n10580), .Z(n10689) );
  NAND U11111 ( .A(y[64]), .B(x[88]), .Z(n10579) );
  XOR U11112 ( .A(n10689), .B(n10579), .Z(n10581) );
  AND U11113 ( .A(y[24]), .B(x[80]), .Z(n10596) );
  AND U11114 ( .A(y[104]), .B(x[96]), .Z(n10587) );
  XOR U11115 ( .A(n10596), .B(n10587), .Z(n10586) );
  AND U11116 ( .A(y[144]), .B(x[104]), .Z(n10585) );
  XNOR U11117 ( .A(n10586), .B(n10585), .Z(n10582) );
  XNOR U11118 ( .A(n10581), .B(n10582), .Z(o[104]) );
  AND U11119 ( .A(x[81]), .B(y[24]), .Z(n10578) );
  NAND U11120 ( .A(x[80]), .B(y[25]), .Z(n10577) );
  XNOR U11121 ( .A(n10578), .B(n10577), .Z(n10598) );
  AND U11122 ( .A(y[64]), .B(x[89]), .Z(n10597) );
  XOR U11123 ( .A(n10598), .B(n10597), .Z(n10609) );
  AND U11124 ( .A(y[184]), .B(x[113]), .Z(n10798) );
  AND U11125 ( .A(y[105]), .B(x[96]), .Z(n10601) );
  XOR U11126 ( .A(n10798), .B(n10601), .Z(n10603) );
  AND U11127 ( .A(y[185]), .B(x[112]), .Z(n10618) );
  NAND U11128 ( .A(y[104]), .B(x[97]), .Z(n10617) );
  XNOR U11129 ( .A(n10618), .B(n10617), .Z(n10602) );
  XOR U11130 ( .A(n10603), .B(n10602), .Z(n10607) );
  AND U11131 ( .A(y[65]), .B(x[88]), .Z(n10823) );
  AND U11132 ( .A(y[145]), .B(x[104]), .Z(n10612) );
  XOR U11133 ( .A(n10823), .B(n10612), .Z(n10614) );
  AND U11134 ( .A(y[144]), .B(x[105]), .Z(n10613) );
  XNOR U11135 ( .A(n10614), .B(n10613), .Z(n10606) );
  XNOR U11136 ( .A(n10607), .B(n10606), .Z(n10608) );
  XNOR U11137 ( .A(n10609), .B(n10608), .Z(n10593) );
  NANDN U11138 ( .A(n10580), .B(n10579), .Z(n10584) );
  NAND U11139 ( .A(n10582), .B(n10581), .Z(n10583) );
  AND U11140 ( .A(n10584), .B(n10583), .Z(n10591) );
  NAND U11141 ( .A(n10586), .B(n10585), .Z(n10589) );
  AND U11142 ( .A(n10596), .B(n10587), .Z(n10588) );
  ANDN U11143 ( .B(n10589), .A(n10588), .Z(n10590) );
  XNOR U11144 ( .A(n10591), .B(n10590), .Z(n10592) );
  XNOR U11145 ( .A(n10593), .B(n10592), .Z(o[105]) );
  NANDN U11146 ( .A(n10591), .B(n10590), .Z(n10595) );
  NAND U11147 ( .A(n10593), .B(n10592), .Z(n10594) );
  AND U11148 ( .A(n10595), .B(n10594), .Z(n10621) );
  AND U11149 ( .A(y[25]), .B(x[81]), .Z(n10639) );
  NAND U11150 ( .A(n10596), .B(n10639), .Z(n10600) );
  NAND U11151 ( .A(n10598), .B(n10597), .Z(n10599) );
  NAND U11152 ( .A(n10600), .B(n10599), .Z(n10673) );
  NAND U11153 ( .A(n10798), .B(n10601), .Z(n10605) );
  NAND U11154 ( .A(n10603), .B(n10602), .Z(n10604) );
  NAND U11155 ( .A(n10605), .B(n10604), .Z(n10671) );
  AND U11156 ( .A(y[146]), .B(x[104]), .Z(n10656) );
  AND U11157 ( .A(y[26]), .B(x[80]), .Z(n10655) );
  XOR U11158 ( .A(n10656), .B(n10655), .Z(n10658) );
  AND U11159 ( .A(y[64]), .B(x[90]), .Z(n10657) );
  XOR U11160 ( .A(n10658), .B(n10657), .Z(n10672) );
  XOR U11161 ( .A(n10671), .B(n10672), .Z(n10674) );
  XOR U11162 ( .A(n10673), .B(n10674), .Z(n10620) );
  XOR U11163 ( .A(n10621), .B(n10620), .Z(n10623) );
  NANDN U11164 ( .A(n10607), .B(n10606), .Z(n10611) );
  NANDN U11165 ( .A(n10609), .B(n10608), .Z(n10610) );
  AND U11166 ( .A(n10611), .B(n10610), .Z(n10626) );
  AND U11167 ( .A(y[24]), .B(x[82]), .Z(n10637) );
  AND U11168 ( .A(y[106]), .B(x[96]), .Z(n10636) );
  XOR U11169 ( .A(n10637), .B(n10636), .Z(n10638) );
  XOR U11170 ( .A(n10639), .B(n10638), .Z(n10666) );
  AND U11171 ( .A(y[144]), .B(x[106]), .Z(n10665) );
  XOR U11172 ( .A(n10666), .B(n10665), .Z(n10668) );
  AND U11173 ( .A(y[104]), .B(x[98]), .Z(n10715) );
  AND U11174 ( .A(y[186]), .B(x[112]), .Z(n10647) );
  XOR U11175 ( .A(n10715), .B(n10647), .Z(n10649) );
  AND U11176 ( .A(y[105]), .B(x[97]), .Z(n10648) );
  XOR U11177 ( .A(n10649), .B(n10648), .Z(n10667) );
  XOR U11178 ( .A(n10668), .B(n10667), .Z(n10624) );
  AND U11179 ( .A(n10823), .B(n10612), .Z(n10616) );
  NAND U11180 ( .A(n10614), .B(n10613), .Z(n10615) );
  NANDN U11181 ( .A(n10616), .B(n10615), .Z(n10632) );
  ANDN U11182 ( .B(n10618), .A(n10617), .Z(n10662) );
  AND U11183 ( .A(x[113]), .B(y[185]), .Z(n10694) );
  AND U11184 ( .A(x[114]), .B(y[184]), .Z(n10619) );
  XOR U11185 ( .A(n10694), .B(n10619), .Z(n10661) );
  XOR U11186 ( .A(n10662), .B(n10661), .Z(n10631) );
  AND U11187 ( .A(y[145]), .B(x[105]), .Z(n10643) );
  AND U11188 ( .A(y[65]), .B(x[89]), .Z(n10642) );
  XOR U11189 ( .A(n10643), .B(n10642), .Z(n10645) );
  AND U11190 ( .A(y[66]), .B(x[88]), .Z(n10644) );
  XOR U11191 ( .A(n10645), .B(n10644), .Z(n10630) );
  XOR U11192 ( .A(n10631), .B(n10630), .Z(n10633) );
  XNOR U11193 ( .A(n10632), .B(n10633), .Z(n10625) );
  XOR U11194 ( .A(n10624), .B(n10625), .Z(n10627) );
  XNOR U11195 ( .A(n10626), .B(n10627), .Z(n10622) );
  XOR U11196 ( .A(n10623), .B(n10622), .Z(o[106]) );
  NANDN U11197 ( .A(n10625), .B(n10624), .Z(n10629) );
  NANDN U11198 ( .A(n10627), .B(n10626), .Z(n10628) );
  NAND U11199 ( .A(n10629), .B(n10628), .Z(n10739) );
  NAND U11200 ( .A(n10631), .B(n10630), .Z(n10635) );
  NAND U11201 ( .A(n10633), .B(n10632), .Z(n10634) );
  NAND U11202 ( .A(n10635), .B(n10634), .Z(n10737) );
  NAND U11203 ( .A(n10637), .B(n10636), .Z(n10641) );
  NAND U11204 ( .A(n10639), .B(n10638), .Z(n10640) );
  NAND U11205 ( .A(n10641), .B(n10640), .Z(n10749) );
  NAND U11206 ( .A(y[147]), .B(x[104]), .Z(n10729) );
  NAND U11207 ( .A(y[107]), .B(x[96]), .Z(n10727) );
  NAND U11208 ( .A(y[24]), .B(x[83]), .Z(n10728) );
  XOR U11209 ( .A(n10727), .B(n10728), .Z(n10730) );
  XOR U11210 ( .A(n10729), .B(n10730), .Z(n10706) );
  AND U11211 ( .A(x[98]), .B(y[105]), .Z(n10771) );
  NAND U11212 ( .A(x[99]), .B(y[104]), .Z(n10646) );
  XNOR U11213 ( .A(n10771), .B(n10646), .Z(n10717) );
  AND U11214 ( .A(y[106]), .B(x[97]), .Z(n10716) );
  XOR U11215 ( .A(n10717), .B(n10716), .Z(n10705) );
  XNOR U11216 ( .A(n10706), .B(n10705), .Z(n10708) );
  XOR U11217 ( .A(n10707), .B(n10708), .Z(n10750) );
  XOR U11218 ( .A(n10749), .B(n10750), .Z(n10751) );
  AND U11219 ( .A(n10715), .B(n10647), .Z(n10651) );
  NAND U11220 ( .A(n10649), .B(n10648), .Z(n10650) );
  NANDN U11221 ( .A(n10651), .B(n10650), .Z(n10711) );
  NAND U11222 ( .A(y[26]), .B(x[81]), .Z(n10687) );
  NAND U11223 ( .A(y[25]), .B(x[82]), .Z(n10685) );
  NAND U11224 ( .A(y[146]), .B(x[105]), .Z(n10686) );
  XOR U11225 ( .A(n10685), .B(n10686), .Z(n10688) );
  XOR U11226 ( .A(n10687), .B(n10688), .Z(n10710) );
  AND U11227 ( .A(x[115]), .B(y[184]), .Z(n10653) );
  NAND U11228 ( .A(x[112]), .B(y[187]), .Z(n10652) );
  XNOR U11229 ( .A(n10653), .B(n10652), .Z(n10691) );
  AND U11230 ( .A(x[114]), .B(y[185]), .Z(n10780) );
  NAND U11231 ( .A(x[113]), .B(y[186]), .Z(n10654) );
  XNOR U11232 ( .A(n10780), .B(n10654), .Z(n10690) );
  XOR U11233 ( .A(n10691), .B(n10690), .Z(n10709) );
  XOR U11234 ( .A(n10710), .B(n10709), .Z(n10712) );
  XOR U11235 ( .A(n10711), .B(n10712), .Z(n10752) );
  XOR U11236 ( .A(n10737), .B(n10738), .Z(n10740) );
  XOR U11237 ( .A(n10739), .B(n10740), .Z(n10731) );
  XNOR U11238 ( .A(n10732), .B(n10731), .Z(n10734) );
  NAND U11239 ( .A(n10656), .B(n10655), .Z(n10660) );
  NAND U11240 ( .A(n10658), .B(n10657), .Z(n10659) );
  NAND U11241 ( .A(n10660), .B(n10659), .Z(n10678) );
  AND U11242 ( .A(n10662), .B(n10661), .Z(n10664) );
  NAND U11243 ( .A(n10798), .B(n10780), .Z(n10663) );
  NANDN U11244 ( .A(n10664), .B(n10663), .Z(n10677) );
  XOR U11245 ( .A(n10678), .B(n10677), .Z(n10680) );
  NAND U11246 ( .A(y[64]), .B(x[91]), .Z(n10722) );
  NAND U11247 ( .A(y[27]), .B(x[80]), .Z(n10720) );
  NAND U11248 ( .A(y[145]), .B(x[106]), .Z(n10721) );
  XOR U11249 ( .A(n10720), .B(n10721), .Z(n10723) );
  XOR U11250 ( .A(n10722), .B(n10723), .Z(n10701) );
  NAND U11251 ( .A(y[67]), .B(x[88]), .Z(n10697) );
  NAND U11252 ( .A(y[65]), .B(x[90]), .Z(n10695) );
  NAND U11253 ( .A(y[144]), .B(x[107]), .Z(n10696) );
  XOR U11254 ( .A(n10695), .B(n10696), .Z(n10698) );
  XOR U11255 ( .A(n10697), .B(n10698), .Z(n10700) );
  AND U11256 ( .A(y[66]), .B(x[89]), .Z(n10699) );
  XOR U11257 ( .A(n10700), .B(n10699), .Z(n10702) );
  XOR U11258 ( .A(n10701), .B(n10702), .Z(n10679) );
  XOR U11259 ( .A(n10680), .B(n10679), .Z(n10744) );
  NAND U11260 ( .A(n10666), .B(n10665), .Z(n10670) );
  NAND U11261 ( .A(n10668), .B(n10667), .Z(n10669) );
  AND U11262 ( .A(n10670), .B(n10669), .Z(n10743) );
  NAND U11263 ( .A(n10672), .B(n10671), .Z(n10676) );
  NAND U11264 ( .A(n10674), .B(n10673), .Z(n10675) );
  AND U11265 ( .A(n10676), .B(n10675), .Z(n10745) );
  XNOR U11266 ( .A(n10746), .B(n10745), .Z(n10733) );
  XOR U11267 ( .A(n10734), .B(n10733), .Z(o[107]) );
  NAND U11268 ( .A(n10678), .B(n10677), .Z(n10682) );
  NAND U11269 ( .A(n10680), .B(n10679), .Z(n10681) );
  NAND U11270 ( .A(n10682), .B(n10681), .Z(n10766) );
  AND U11271 ( .A(x[88]), .B(y[68]), .Z(n10684) );
  NAND U11272 ( .A(x[91]), .B(y[65]), .Z(n10683) );
  XNOR U11273 ( .A(n10684), .B(n10683), .Z(n10825) );
  AND U11274 ( .A(y[66]), .B(x[90]), .Z(n10824) );
  XOR U11275 ( .A(n10825), .B(n10824), .Z(n10829) );
  AND U11276 ( .A(y[67]), .B(x[89]), .Z(n10828) );
  XOR U11277 ( .A(n10829), .B(n10828), .Z(n10831) );
  AND U11278 ( .A(y[144]), .B(x[108]), .Z(n10777) );
  AND U11279 ( .A(y[27]), .B(x[81]), .Z(n10776) );
  XOR U11280 ( .A(n10777), .B(n10776), .Z(n10779) );
  AND U11281 ( .A(y[28]), .B(x[80]), .Z(n10778) );
  XOR U11282 ( .A(n10779), .B(n10778), .Z(n10830) );
  XOR U11283 ( .A(n10831), .B(n10830), .Z(n10843) );
  AND U11284 ( .A(y[187]), .B(x[115]), .Z(n11117) );
  NANDN U11285 ( .A(n10689), .B(n11117), .Z(n10693) );
  NAND U11286 ( .A(n10691), .B(n10690), .Z(n10692) );
  AND U11287 ( .A(n10693), .B(n10692), .Z(n10841) );
  XOR U11288 ( .A(n10840), .B(n10841), .Z(n10842) );
  XNOR U11289 ( .A(n10843), .B(n10842), .Z(n10855) );
  NAND U11290 ( .A(y[24]), .B(x[84]), .Z(n10809) );
  NAND U11291 ( .A(y[146]), .B(x[106]), .Z(n10808) );
  NAND U11292 ( .A(y[108]), .B(x[96]), .Z(n10807) );
  XOR U11293 ( .A(n10808), .B(n10807), .Z(n10810) );
  XOR U11294 ( .A(n10809), .B(n10810), .Z(n10791) );
  AND U11295 ( .A(x[114]), .B(y[186]), .Z(n10726) );
  NAND U11296 ( .A(n10726), .B(n10694), .Z(n10803) );
  NAND U11297 ( .A(y[104]), .B(x[100]), .Z(n10907) );
  NAND U11298 ( .A(y[188]), .B(x[112]), .Z(n10977) );
  XNOR U11299 ( .A(n10907), .B(n10977), .Z(n10804) );
  XOR U11300 ( .A(n10803), .B(n10804), .Z(n10790) );
  XNOR U11301 ( .A(n10791), .B(n10790), .Z(n10793) );
  XOR U11302 ( .A(n10793), .B(n10792), .Z(n10853) );
  NANDN U11303 ( .A(n10700), .B(n10699), .Z(n10704) );
  OR U11304 ( .A(n10702), .B(n10701), .Z(n10703) );
  AND U11305 ( .A(n10704), .B(n10703), .Z(n10852) );
  XNOR U11306 ( .A(n10853), .B(n10852), .Z(n10854) );
  XNOR U11307 ( .A(n10855), .B(n10854), .Z(n10765) );
  XOR U11308 ( .A(n10766), .B(n10765), .Z(n10768) );
  NANDN U11309 ( .A(n10710), .B(n10709), .Z(n10714) );
  NANDN U11310 ( .A(n10712), .B(n10711), .Z(n10713) );
  NAND U11311 ( .A(n10714), .B(n10713), .Z(n10845) );
  XOR U11312 ( .A(n10844), .B(n10845), .Z(n10847) );
  AND U11313 ( .A(y[64]), .B(x[92]), .Z(n10784) );
  NAND U11314 ( .A(y[148]), .B(x[104]), .Z(n10785) );
  XNOR U11315 ( .A(n10784), .B(n10785), .Z(n10786) );
  NAND U11316 ( .A(y[147]), .B(x[105]), .Z(n10787) );
  XNOR U11317 ( .A(n10786), .B(n10787), .Z(n10833) );
  AND U11318 ( .A(x[98]), .B(y[106]), .Z(n10719) );
  NAND U11319 ( .A(x[99]), .B(y[105]), .Z(n10718) );
  XNOR U11320 ( .A(n10719), .B(n10718), .Z(n10773) );
  AND U11321 ( .A(y[107]), .B(x[97]), .Z(n10772) );
  XOR U11322 ( .A(n10773), .B(n10772), .Z(n10832) );
  XOR U11323 ( .A(n10833), .B(n10832), .Z(n10836) );
  XOR U11324 ( .A(n10836), .B(n10835), .Z(n10849) );
  XOR U11325 ( .A(n10848), .B(n10849), .Z(n10851) );
  AND U11326 ( .A(y[26]), .B(x[82]), .Z(n10820) );
  AND U11327 ( .A(y[145]), .B(x[107]), .Z(n10818) );
  NAND U11328 ( .A(y[25]), .B(x[83]), .Z(n10817) );
  XNOR U11329 ( .A(n10818), .B(n10817), .Z(n10819) );
  XOR U11330 ( .A(n10820), .B(n10819), .Z(n10794) );
  AND U11331 ( .A(x[116]), .B(y[184]), .Z(n10725) );
  NAND U11332 ( .A(x[113]), .B(y[187]), .Z(n10724) );
  XNOR U11333 ( .A(n10725), .B(n10724), .Z(n10800) );
  AND U11334 ( .A(y[185]), .B(x[115]), .Z(n10915) );
  XOR U11335 ( .A(n10915), .B(n10726), .Z(n10799) );
  XOR U11336 ( .A(n10800), .B(n10799), .Z(n10795) );
  XOR U11337 ( .A(n10794), .B(n10795), .Z(n10797) );
  XOR U11338 ( .A(n10797), .B(n10796), .Z(n10850) );
  XOR U11339 ( .A(n10851), .B(n10850), .Z(n10846) );
  XOR U11340 ( .A(n10847), .B(n10846), .Z(n10767) );
  XNOR U11341 ( .A(n10768), .B(n10767), .Z(n10758) );
  NANDN U11342 ( .A(n10732), .B(n10731), .Z(n10736) );
  NAND U11343 ( .A(n10734), .B(n10733), .Z(n10735) );
  NAND U11344 ( .A(n10736), .B(n10735), .Z(n10756) );
  NAND U11345 ( .A(n10738), .B(n10737), .Z(n10742) );
  NAND U11346 ( .A(n10740), .B(n10739), .Z(n10741) );
  AND U11347 ( .A(n10742), .B(n10741), .Z(n10761) );
  NANDN U11348 ( .A(n10744), .B(n10743), .Z(n10748) );
  NAND U11349 ( .A(n10746), .B(n10745), .Z(n10747) );
  NAND U11350 ( .A(n10748), .B(n10747), .Z(n10759) );
  NAND U11351 ( .A(n10750), .B(n10749), .Z(n10754) );
  NANDN U11352 ( .A(n10752), .B(n10751), .Z(n10753) );
  AND U11353 ( .A(n10754), .B(n10753), .Z(n10760) );
  XOR U11354 ( .A(n10759), .B(n10760), .Z(n10762) );
  XNOR U11355 ( .A(n10761), .B(n10762), .Z(n10757) );
  XOR U11356 ( .A(n10756), .B(n10757), .Z(n10755) );
  XNOR U11357 ( .A(n10758), .B(n10755), .Z(o[108]) );
  NAND U11358 ( .A(n10760), .B(n10759), .Z(n10764) );
  NAND U11359 ( .A(n10762), .B(n10761), .Z(n10763) );
  AND U11360 ( .A(n10764), .B(n10763), .Z(n10864) );
  XNOR U11361 ( .A(n10865), .B(n10864), .Z(n10867) );
  NAND U11362 ( .A(n10766), .B(n10765), .Z(n10770) );
  NAND U11363 ( .A(n10768), .B(n10767), .Z(n10769) );
  NAND U11364 ( .A(n10770), .B(n10769), .Z(n10858) );
  AND U11365 ( .A(y[106]), .B(x[99]), .Z(n10909) );
  NAND U11366 ( .A(n10771), .B(n10909), .Z(n10775) );
  NAND U11367 ( .A(n10773), .B(n10772), .Z(n10774) );
  NAND U11368 ( .A(n10775), .B(n10774), .Z(n10870) );
  AND U11369 ( .A(y[64]), .B(x[93]), .Z(n10898) );
  AND U11370 ( .A(y[107]), .B(x[98]), .Z(n10897) );
  XOR U11371 ( .A(n10898), .B(n10897), .Z(n10899) );
  AND U11372 ( .A(y[149]), .B(x[104]), .Z(n11167) );
  XOR U11373 ( .A(n10899), .B(n11167), .Z(n10892) );
  AND U11374 ( .A(y[145]), .B(x[108]), .Z(n10903) );
  AND U11375 ( .A(y[24]), .B(x[85]), .Z(n10902) );
  XOR U11376 ( .A(n10903), .B(n10902), .Z(n10904) );
  AND U11377 ( .A(y[25]), .B(x[84]), .Z(n11213) );
  XOR U11378 ( .A(n10904), .B(n11213), .Z(n10891) );
  XOR U11379 ( .A(n10892), .B(n10891), .Z(n10894) );
  XOR U11380 ( .A(n10893), .B(n10894), .Z(n10871) );
  XOR U11381 ( .A(n10870), .B(n10871), .Z(n10874) );
  AND U11382 ( .A(y[186]), .B(x[115]), .Z(n10781) );
  AND U11383 ( .A(n10781), .B(n10780), .Z(n10979) );
  AND U11384 ( .A(x[112]), .B(y[189]), .Z(n10783) );
  AND U11385 ( .A(x[113]), .B(y[188]), .Z(n10782) );
  XOR U11386 ( .A(n10783), .B(n10782), .Z(n10978) );
  XOR U11387 ( .A(n10979), .B(n10978), .Z(n10966) );
  AND U11388 ( .A(y[65]), .B(x[92]), .Z(n10958) );
  AND U11389 ( .A(y[69]), .B(x[88]), .Z(n10956) );
  NAND U11390 ( .A(y[28]), .B(x[81]), .Z(n10957) );
  XOR U11391 ( .A(n10956), .B(n10957), .Z(n10959) );
  XOR U11392 ( .A(n10958), .B(n10959), .Z(n10967) );
  XNOR U11393 ( .A(n10966), .B(n10967), .Z(n10969) );
  NANDN U11394 ( .A(n10785), .B(n10784), .Z(n10789) );
  NANDN U11395 ( .A(n10787), .B(n10786), .Z(n10788) );
  NAND U11396 ( .A(n10789), .B(n10788), .Z(n10968) );
  XOR U11397 ( .A(n10969), .B(n10968), .Z(n10873) );
  XOR U11398 ( .A(n10874), .B(n10873), .Z(n10919) );
  XNOR U11399 ( .A(n10916), .B(n10917), .Z(n10920) );
  XNOR U11400 ( .A(n10919), .B(n10920), .Z(n10996) );
  AND U11401 ( .A(y[187]), .B(x[116]), .Z(n11199) );
  NAND U11402 ( .A(n11199), .B(n10798), .Z(n10802) );
  NAND U11403 ( .A(n10800), .B(n10799), .Z(n10801) );
  NAND U11404 ( .A(n10802), .B(n10801), .Z(n10929) );
  NAND U11405 ( .A(n10907), .B(n10977), .Z(n10806) );
  NANDN U11406 ( .A(n10804), .B(n10803), .Z(n10805) );
  AND U11407 ( .A(n10806), .B(n10805), .Z(n10930) );
  XOR U11408 ( .A(n10929), .B(n10930), .Z(n10932) );
  NAND U11409 ( .A(n10808), .B(n10807), .Z(n10812) );
  NAND U11410 ( .A(n10810), .B(n10809), .Z(n10811) );
  AND U11411 ( .A(n10812), .B(n10811), .Z(n10936) );
  AND U11412 ( .A(y[68]), .B(x[89]), .Z(n10890) );
  AND U11413 ( .A(y[66]), .B(x[91]), .Z(n11047) );
  AND U11414 ( .A(x[90]), .B(y[67]), .Z(n10813) );
  XOR U11415 ( .A(n11047), .B(n10813), .Z(n10889) );
  XOR U11416 ( .A(n10890), .B(n10889), .Z(n10934) );
  AND U11417 ( .A(y[185]), .B(x[116]), .Z(n11181) );
  NAND U11418 ( .A(x[115]), .B(y[186]), .Z(n10814) );
  XNOR U11419 ( .A(n11181), .B(n10814), .Z(n10881) );
  AND U11420 ( .A(y[184]), .B(x[117]), .Z(n10879) );
  AND U11421 ( .A(y[187]), .B(x[114]), .Z(n10878) );
  XOR U11422 ( .A(n10879), .B(n10878), .Z(n10880) );
  XOR U11423 ( .A(n10881), .B(n10880), .Z(n10933) );
  XOR U11424 ( .A(n10934), .B(n10933), .Z(n10935) );
  XOR U11425 ( .A(n10936), .B(n10935), .Z(n10931) );
  XOR U11426 ( .A(n10932), .B(n10931), .Z(n10946) );
  AND U11427 ( .A(y[105]), .B(x[100]), .Z(n10816) );
  AND U11428 ( .A(x[101]), .B(y[104]), .Z(n10815) );
  XOR U11429 ( .A(n10816), .B(n10815), .Z(n10908) );
  XOR U11430 ( .A(n10909), .B(n10908), .Z(n10948) );
  AND U11431 ( .A(y[144]), .B(x[109]), .Z(n10883) );
  AND U11432 ( .A(y[26]), .B(x[83]), .Z(n10882) );
  XOR U11433 ( .A(n10883), .B(n10882), .Z(n10885) );
  AND U11434 ( .A(y[27]), .B(x[82]), .Z(n10884) );
  XOR U11435 ( .A(n10885), .B(n10884), .Z(n10947) );
  XOR U11436 ( .A(n10948), .B(n10947), .Z(n10950) );
  NANDN U11437 ( .A(n10818), .B(n10817), .Z(n10822) );
  NANDN U11438 ( .A(n10820), .B(n10819), .Z(n10821) );
  NAND U11439 ( .A(n10822), .B(n10821), .Z(n10951) );
  XOR U11440 ( .A(n10950), .B(n10951), .Z(n10943) );
  AND U11441 ( .A(y[68]), .B(x[91]), .Z(n11198) );
  NAND U11442 ( .A(n11198), .B(n10823), .Z(n10827) );
  IV U11443 ( .A(n10824), .Z(n10888) );
  NANDN U11444 ( .A(n10888), .B(n10825), .Z(n10826) );
  NAND U11445 ( .A(n10827), .B(n10826), .Z(n10925) );
  AND U11446 ( .A(y[108]), .B(x[97]), .Z(n11221) );
  AND U11447 ( .A(y[146]), .B(x[107]), .Z(n10972) );
  XOR U11448 ( .A(n11221), .B(n10972), .Z(n10973) );
  NAND U11449 ( .A(y[109]), .B(x[96]), .Z(n10974) );
  XNOR U11450 ( .A(n10973), .B(n10974), .Z(n10924) );
  AND U11451 ( .A(y[29]), .B(x[80]), .Z(n10982) );
  NAND U11452 ( .A(y[148]), .B(x[105]), .Z(n10983) );
  XNOR U11453 ( .A(n10982), .B(n10983), .Z(n10984) );
  NAND U11454 ( .A(y[147]), .B(x[106]), .Z(n10985) );
  XNOR U11455 ( .A(n10984), .B(n10985), .Z(n10923) );
  XNOR U11456 ( .A(n10924), .B(n10923), .Z(n10926) );
  XOR U11457 ( .A(n10925), .B(n10926), .Z(n10944) );
  XOR U11458 ( .A(n10943), .B(n10944), .Z(n10945) );
  XOR U11459 ( .A(n10946), .B(n10945), .Z(n10995) );
  IV U11460 ( .A(n10832), .Z(n10834) );
  NANDN U11461 ( .A(n10834), .B(n10833), .Z(n10839) );
  IV U11462 ( .A(n10835), .Z(n10837) );
  NANDN U11463 ( .A(n10837), .B(n10836), .Z(n10838) );
  NAND U11464 ( .A(n10839), .B(n10838), .Z(n10940) );
  XOR U11465 ( .A(n10939), .B(n10940), .Z(n10942) );
  XOR U11466 ( .A(n10942), .B(n10941), .Z(n10994) );
  XNOR U11467 ( .A(n10995), .B(n10994), .Z(n10997) );
  XNOR U11468 ( .A(n10996), .B(n10997), .Z(n10859) );
  XOR U11469 ( .A(n10858), .B(n10859), .Z(n10860) );
  NANDN U11470 ( .A(n10853), .B(n10852), .Z(n10857) );
  NAND U11471 ( .A(n10855), .B(n10854), .Z(n10856) );
  AND U11472 ( .A(n10857), .B(n10856), .Z(n10990) );
  XNOR U11473 ( .A(n10991), .B(n10990), .Z(n10993) );
  XOR U11474 ( .A(n10992), .B(n10993), .Z(n10861) );
  XOR U11475 ( .A(n10867), .B(n10866), .Z(o[109]) );
  NAND U11476 ( .A(n10859), .B(n10858), .Z(n10863) );
  NANDN U11477 ( .A(n10861), .B(n10860), .Z(n10862) );
  AND U11478 ( .A(n10863), .B(n10862), .Z(n11005) );
  NANDN U11479 ( .A(n10865), .B(n10864), .Z(n10869) );
  NAND U11480 ( .A(n10867), .B(n10866), .Z(n10868) );
  NAND U11481 ( .A(n10869), .B(n10868), .Z(n11003) );
  IV U11482 ( .A(n10870), .Z(n10872) );
  NANDN U11483 ( .A(n10872), .B(n10871), .Z(n10877) );
  IV U11484 ( .A(n10873), .Z(n10875) );
  NANDN U11485 ( .A(n10875), .B(n10874), .Z(n10876) );
  AND U11486 ( .A(n10877), .B(n10876), .Z(n11285) );
  NAND U11487 ( .A(n10883), .B(n10882), .Z(n10887) );
  NAND U11488 ( .A(n10885), .B(n10884), .Z(n10886) );
  NAND U11489 ( .A(n10887), .B(n10886), .Z(n11036) );
  AND U11490 ( .A(y[147]), .B(x[107]), .Z(n11185) );
  AND U11491 ( .A(y[107]), .B(x[99]), .Z(n11184) );
  XOR U11492 ( .A(n11185), .B(n11184), .Z(n11183) );
  AND U11493 ( .A(y[27]), .B(x[83]), .Z(n11182) );
  XOR U11494 ( .A(n11183), .B(n11182), .Z(n11042) );
  AND U11495 ( .A(y[148]), .B(x[106]), .Z(n11173) );
  AND U11496 ( .A(y[106]), .B(x[100]), .Z(n11172) );
  XOR U11497 ( .A(n11173), .B(n11172), .Z(n11171) );
  AND U11498 ( .A(y[28]), .B(x[82]), .Z(n11170) );
  XNOR U11499 ( .A(n11171), .B(n11170), .Z(n11041) );
  XNOR U11500 ( .A(n11040), .B(n11039), .Z(n11035) );
  XOR U11501 ( .A(n11036), .B(n11035), .Z(n11034) );
  XOR U11502 ( .A(n11033), .B(n11034), .Z(n11010) );
  NAND U11503 ( .A(n10892), .B(n10891), .Z(n10896) );
  NAND U11504 ( .A(n10894), .B(n10893), .Z(n10895) );
  NAND U11505 ( .A(n10896), .B(n10895), .Z(n11009) );
  XOR U11506 ( .A(n11010), .B(n11009), .Z(n11008) );
  NAND U11507 ( .A(n10898), .B(n10897), .Z(n10901) );
  NAND U11508 ( .A(n10899), .B(n11167), .Z(n10900) );
  NAND U11509 ( .A(n10901), .B(n10900), .Z(n11155) );
  NAND U11510 ( .A(n10903), .B(n10902), .Z(n10906) );
  NAND U11511 ( .A(n10904), .B(n11213), .Z(n10905) );
  NAND U11512 ( .A(n10906), .B(n10905), .Z(n11154) );
  XOR U11513 ( .A(n11155), .B(n11154), .Z(n11153) );
  AND U11514 ( .A(y[105]), .B(x[101]), .Z(n11207) );
  NANDN U11515 ( .A(n10907), .B(n11207), .Z(n10911) );
  NAND U11516 ( .A(n10909), .B(n10908), .Z(n10910) );
  AND U11517 ( .A(n10911), .B(n10910), .Z(n11249) );
  AND U11518 ( .A(x[85]), .B(y[25]), .Z(n10913) );
  NAND U11519 ( .A(x[84]), .B(y[26]), .Z(n10912) );
  XNOR U11520 ( .A(n10913), .B(n10912), .Z(n11211) );
  AND U11521 ( .A(y[144]), .B(x[110]), .Z(n11210) );
  XOR U11522 ( .A(n11211), .B(n11210), .Z(n11246) );
  AND U11523 ( .A(y[189]), .B(x[113]), .Z(n11125) );
  AND U11524 ( .A(y[186]), .B(x[116]), .Z(n10914) );
  AND U11525 ( .A(n10915), .B(n10914), .Z(n11123) );
  AND U11526 ( .A(y[188]), .B(x[114]), .Z(n11122) );
  XOR U11527 ( .A(n11123), .B(n11122), .Z(n11124) );
  XNOR U11528 ( .A(n11125), .B(n11124), .Z(n11247) );
  XNOR U11529 ( .A(n11249), .B(n11248), .Z(n11152) );
  XOR U11530 ( .A(n11153), .B(n11152), .Z(n11007) );
  XOR U11531 ( .A(n11008), .B(n11007), .Z(n11275) );
  IV U11532 ( .A(n10916), .Z(n10918) );
  NANDN U11533 ( .A(n10918), .B(n10917), .Z(n10922) );
  NANDN U11534 ( .A(n10920), .B(n10919), .Z(n10921) );
  AND U11535 ( .A(n10922), .B(n10921), .Z(n11274) );
  NAND U11536 ( .A(n10924), .B(n10923), .Z(n10928) );
  NANDN U11537 ( .A(n10926), .B(n10925), .Z(n10927) );
  AND U11538 ( .A(n10928), .B(n10927), .Z(n11016) );
  XOR U11539 ( .A(n11016), .B(n11015), .Z(n11014) );
  NAND U11540 ( .A(n10934), .B(n10933), .Z(n10938) );
  NAND U11541 ( .A(n10936), .B(n10935), .Z(n10937) );
  AND U11542 ( .A(n10938), .B(n10937), .Z(n11013) );
  XOR U11543 ( .A(n11014), .B(n11013), .Z(n11272) );
  XOR U11544 ( .A(n11273), .B(n11272), .Z(n11284) );
  XOR U11545 ( .A(n11285), .B(n11284), .Z(n11283) );
  IV U11546 ( .A(n10947), .Z(n10949) );
  NANDN U11547 ( .A(n10949), .B(n10948), .Z(n10953) );
  NANDN U11548 ( .A(n10951), .B(n10950), .Z(n10952) );
  AND U11549 ( .A(n10953), .B(n10952), .Z(n11002) );
  AND U11550 ( .A(y[110]), .B(x[96]), .Z(n11227) );
  AND U11551 ( .A(y[24]), .B(x[86]), .Z(n11226) );
  XOR U11552 ( .A(n11227), .B(n11226), .Z(n11225) );
  AND U11553 ( .A(y[145]), .B(x[109]), .Z(n11224) );
  XOR U11554 ( .A(n11225), .B(n11224), .Z(n11113) );
  AND U11555 ( .A(y[65]), .B(x[93]), .Z(n11139) );
  AND U11556 ( .A(y[68]), .B(x[90]), .Z(n11138) );
  XOR U11557 ( .A(n11139), .B(n11138), .Z(n11137) );
  AND U11558 ( .A(y[69]), .B(x[89]), .Z(n11136) );
  XOR U11559 ( .A(n11137), .B(n11136), .Z(n11046) );
  AND U11560 ( .A(x[92]), .B(y[66]), .Z(n10955) );
  NAND U11561 ( .A(x[91]), .B(y[67]), .Z(n10954) );
  XNOR U11562 ( .A(n10955), .B(n10954), .Z(n11045) );
  XOR U11563 ( .A(n11046), .B(n11045), .Z(n11112) );
  XOR U11564 ( .A(n11113), .B(n11112), .Z(n11111) );
  AND U11565 ( .A(y[190]), .B(x[112]), .Z(n11206) );
  XOR U11566 ( .A(n11207), .B(n11206), .Z(n11205) );
  AND U11567 ( .A(y[104]), .B(x[102]), .Z(n11204) );
  XOR U11568 ( .A(n11205), .B(n11204), .Z(n11110) );
  XOR U11569 ( .A(n11111), .B(n11110), .Z(n11025) );
  NANDN U11570 ( .A(n10957), .B(n10956), .Z(n10961) );
  NANDN U11571 ( .A(n10959), .B(n10958), .Z(n10960) );
  AND U11572 ( .A(n10961), .B(n10960), .Z(n11158) );
  AND U11573 ( .A(y[146]), .B(x[108]), .Z(n11219) );
  AND U11574 ( .A(x[97]), .B(y[109]), .Z(n10963) );
  AND U11575 ( .A(x[98]), .B(y[108]), .Z(n10962) );
  XOR U11576 ( .A(n10963), .B(n10962), .Z(n11218) );
  XOR U11577 ( .A(n11219), .B(n11218), .Z(n11161) );
  AND U11578 ( .A(y[30]), .B(x[80]), .Z(n11165) );
  AND U11579 ( .A(y[150]), .B(x[104]), .Z(n10965) );
  AND U11580 ( .A(x[105]), .B(y[149]), .Z(n10964) );
  XOR U11581 ( .A(n10965), .B(n10964), .Z(n11164) );
  XNOR U11582 ( .A(n11165), .B(n11164), .Z(n11160) );
  XNOR U11583 ( .A(n11158), .B(n11159), .Z(n11026) );
  NANDN U11584 ( .A(n10967), .B(n10966), .Z(n10971) );
  NAND U11585 ( .A(n10969), .B(n10968), .Z(n10970) );
  AND U11586 ( .A(n10971), .B(n10970), .Z(n11027) );
  XOR U11587 ( .A(n11028), .B(n11027), .Z(n11001) );
  XOR U11588 ( .A(n11002), .B(n11001), .Z(n10999) );
  AND U11589 ( .A(n11221), .B(n10972), .Z(n10976) );
  NANDN U11590 ( .A(n10974), .B(n10973), .Z(n10975) );
  NANDN U11591 ( .A(n10976), .B(n10975), .Z(n11019) );
  NANDN U11592 ( .A(n10977), .B(n11125), .Z(n10981) );
  NAND U11593 ( .A(n10979), .B(n10978), .Z(n10980) );
  NAND U11594 ( .A(n10981), .B(n10980), .Z(n11022) );
  NANDN U11595 ( .A(n10983), .B(n10982), .Z(n10987) );
  NANDN U11596 ( .A(n10985), .B(n10984), .Z(n10986) );
  AND U11597 ( .A(n10987), .B(n10986), .Z(n11240) );
  AND U11598 ( .A(y[29]), .B(x[81]), .Z(n11133) );
  AND U11599 ( .A(y[64]), .B(x[94]), .Z(n11132) );
  XOR U11600 ( .A(n11133), .B(n11132), .Z(n11131) );
  AND U11601 ( .A(y[70]), .B(x[88]), .Z(n11130) );
  XNOR U11602 ( .A(n11131), .B(n11130), .Z(n11243) );
  AND U11603 ( .A(x[117]), .B(y[185]), .Z(n10989) );
  NAND U11604 ( .A(x[116]), .B(y[186]), .Z(n10988) );
  XNOR U11605 ( .A(n10989), .B(n10988), .Z(n11119) );
  AND U11606 ( .A(y[184]), .B(x[118]), .Z(n11118) );
  XOR U11607 ( .A(n11119), .B(n11118), .Z(n11116) );
  XOR U11608 ( .A(n11117), .B(n11116), .Z(n11242) );
  XNOR U11609 ( .A(n11240), .B(n11241), .Z(n11021) );
  XOR U11610 ( .A(n11019), .B(n11020), .Z(n11000) );
  XOR U11611 ( .A(n10999), .B(n11000), .Z(n11269) );
  XOR U11612 ( .A(n11268), .B(n11269), .Z(n11266) );
  XOR U11613 ( .A(n11267), .B(n11266), .Z(n11282) );
  XNOR U11614 ( .A(n11283), .B(n11282), .Z(n11286) );
  XNOR U11615 ( .A(n11289), .B(n11288), .Z(n11287) );
  XOR U11616 ( .A(n11003), .B(n11004), .Z(n10998) );
  XNOR U11617 ( .A(n11005), .B(n10998), .Z(o[110]) );
  NAND U11618 ( .A(n11008), .B(n11007), .Z(n11012) );
  NAND U11619 ( .A(n11010), .B(n11009), .Z(n11011) );
  NAND U11620 ( .A(n11014), .B(n11013), .Z(n11018) );
  NAND U11621 ( .A(n11016), .B(n11015), .Z(n11017) );
  AND U11622 ( .A(n11018), .B(n11017), .Z(n11265) );
  NANDN U11623 ( .A(n11020), .B(n11019), .Z(n11024) );
  ANDN U11624 ( .B(n11022), .A(n11021), .Z(n11023) );
  ANDN U11625 ( .B(n11024), .A(n11023), .Z(n11032) );
  ANDN U11626 ( .B(n11026), .A(n11025), .Z(n11030) );
  AND U11627 ( .A(n11028), .B(n11027), .Z(n11029) );
  OR U11628 ( .A(n11030), .B(n11029), .Z(n11031) );
  XNOR U11629 ( .A(n11032), .B(n11031), .Z(n11263) );
  NAND U11630 ( .A(n11034), .B(n11033), .Z(n11038) );
  NAND U11631 ( .A(n11036), .B(n11035), .Z(n11037) );
  AND U11632 ( .A(n11038), .B(n11037), .Z(n11261) );
  NAND U11633 ( .A(n11040), .B(n11039), .Z(n11044) );
  NANDN U11634 ( .A(n11042), .B(n11041), .Z(n11043) );
  AND U11635 ( .A(n11044), .B(n11043), .Z(n11151) );
  NAND U11636 ( .A(n11046), .B(n11045), .Z(n11049) );
  AND U11637 ( .A(y[67]), .B(x[92]), .Z(n11099) );
  NAND U11638 ( .A(n11047), .B(n11099), .Z(n11048) );
  AND U11639 ( .A(n11049), .B(n11048), .Z(n11109) );
  AND U11640 ( .A(x[88]), .B(y[71]), .Z(n11051) );
  NAND U11641 ( .A(x[111]), .B(y[144]), .Z(n11050) );
  XNOR U11642 ( .A(n11051), .B(n11050), .Z(n11055) );
  AND U11643 ( .A(x[81]), .B(y[30]), .Z(n11053) );
  NAND U11644 ( .A(x[101]), .B(y[106]), .Z(n11052) );
  XNOR U11645 ( .A(n11053), .B(n11052), .Z(n11054) );
  XOR U11646 ( .A(n11055), .B(n11054), .Z(n11063) );
  AND U11647 ( .A(x[82]), .B(y[29]), .Z(n11057) );
  NAND U11648 ( .A(x[110]), .B(y[145]), .Z(n11056) );
  XNOR U11649 ( .A(n11057), .B(n11056), .Z(n11061) );
  AND U11650 ( .A(x[83]), .B(y[28]), .Z(n11059) );
  NAND U11651 ( .A(x[94]), .B(y[65]), .Z(n11058) );
  XNOR U11652 ( .A(n11059), .B(n11058), .Z(n11060) );
  XNOR U11653 ( .A(n11061), .B(n11060), .Z(n11062) );
  XNOR U11654 ( .A(n11063), .B(n11062), .Z(n11107) );
  AND U11655 ( .A(x[93]), .B(y[66]), .Z(n11068) );
  AND U11656 ( .A(y[186]), .B(x[117]), .Z(n11180) );
  AND U11657 ( .A(x[104]), .B(y[151]), .Z(n11065) );
  NAND U11658 ( .A(x[89]), .B(y[70]), .Z(n11064) );
  XNOR U11659 ( .A(n11065), .B(n11064), .Z(n11066) );
  XNOR U11660 ( .A(n11180), .B(n11066), .Z(n11067) );
  XNOR U11661 ( .A(n11068), .B(n11067), .Z(n11084) );
  AND U11662 ( .A(x[118]), .B(y[185]), .Z(n11070) );
  NAND U11663 ( .A(x[119]), .B(y[184]), .Z(n11069) );
  XNOR U11664 ( .A(n11070), .B(n11069), .Z(n11074) );
  AND U11665 ( .A(x[97]), .B(y[110]), .Z(n11072) );
  NAND U11666 ( .A(x[99]), .B(y[108]), .Z(n11071) );
  XNOR U11667 ( .A(n11072), .B(n11071), .Z(n11073) );
  XOR U11668 ( .A(n11074), .B(n11073), .Z(n11082) );
  AND U11669 ( .A(x[100]), .B(y[107]), .Z(n11076) );
  NAND U11670 ( .A(x[95]), .B(y[64]), .Z(n11075) );
  XNOR U11671 ( .A(n11076), .B(n11075), .Z(n11080) );
  AND U11672 ( .A(x[90]), .B(y[69]), .Z(n11078) );
  NAND U11673 ( .A(x[106]), .B(y[149]), .Z(n11077) );
  XNOR U11674 ( .A(n11078), .B(n11077), .Z(n11079) );
  XNOR U11675 ( .A(n11080), .B(n11079), .Z(n11081) );
  XNOR U11676 ( .A(n11082), .B(n11081), .Z(n11083) );
  XOR U11677 ( .A(n11084), .B(n11083), .Z(n11105) );
  AND U11678 ( .A(x[102]), .B(y[105]), .Z(n11086) );
  NAND U11679 ( .A(x[103]), .B(y[104]), .Z(n11085) );
  XNOR U11680 ( .A(n11086), .B(n11085), .Z(n11090) );
  AND U11681 ( .A(x[112]), .B(y[191]), .Z(n11088) );
  NAND U11682 ( .A(x[80]), .B(y[31]), .Z(n11087) );
  XNOR U11683 ( .A(n11088), .B(n11087), .Z(n11089) );
  XOR U11684 ( .A(n11090), .B(n11089), .Z(n11098) );
  AND U11685 ( .A(x[109]), .B(y[146]), .Z(n11092) );
  NAND U11686 ( .A(x[108]), .B(y[147]), .Z(n11091) );
  XNOR U11687 ( .A(n11092), .B(n11091), .Z(n11096) );
  AND U11688 ( .A(x[87]), .B(y[24]), .Z(n11094) );
  NAND U11689 ( .A(x[86]), .B(y[25]), .Z(n11093) );
  XNOR U11690 ( .A(n11094), .B(n11093), .Z(n11095) );
  XNOR U11691 ( .A(n11096), .B(n11095), .Z(n11097) );
  XNOR U11692 ( .A(n11098), .B(n11097), .Z(n11103) );
  AND U11693 ( .A(y[109]), .B(x[98]), .Z(n11220) );
  AND U11694 ( .A(y[150]), .B(x[105]), .Z(n11166) );
  XOR U11695 ( .A(n11220), .B(n11166), .Z(n11101) );
  AND U11696 ( .A(y[26]), .B(x[85]), .Z(n11212) );
  XNOR U11697 ( .A(n11212), .B(n11099), .Z(n11100) );
  XNOR U11698 ( .A(n11101), .B(n11100), .Z(n11102) );
  XNOR U11699 ( .A(n11103), .B(n11102), .Z(n11104) );
  XNOR U11700 ( .A(n11105), .B(n11104), .Z(n11106) );
  XNOR U11701 ( .A(n11107), .B(n11106), .Z(n11108) );
  XNOR U11702 ( .A(n11109), .B(n11108), .Z(n11149) );
  NAND U11703 ( .A(n11111), .B(n11110), .Z(n11115) );
  NAND U11704 ( .A(n11113), .B(n11112), .Z(n11114) );
  AND U11705 ( .A(n11115), .B(n11114), .Z(n11147) );
  NAND U11706 ( .A(n11117), .B(n11116), .Z(n11121) );
  AND U11707 ( .A(n11119), .B(n11118), .Z(n11120) );
  ANDN U11708 ( .B(n11121), .A(n11120), .Z(n11129) );
  AND U11709 ( .A(n11123), .B(n11122), .Z(n11127) );
  AND U11710 ( .A(n11125), .B(n11124), .Z(n11126) );
  OR U11711 ( .A(n11127), .B(n11126), .Z(n11128) );
  XNOR U11712 ( .A(n11129), .B(n11128), .Z(n11145) );
  NAND U11713 ( .A(n11131), .B(n11130), .Z(n11135) );
  NAND U11714 ( .A(n11133), .B(n11132), .Z(n11134) );
  AND U11715 ( .A(n11135), .B(n11134), .Z(n11143) );
  NAND U11716 ( .A(n11137), .B(n11136), .Z(n11141) );
  NAND U11717 ( .A(n11139), .B(n11138), .Z(n11140) );
  NAND U11718 ( .A(n11141), .B(n11140), .Z(n11142) );
  XNOR U11719 ( .A(n11143), .B(n11142), .Z(n11144) );
  XNOR U11720 ( .A(n11145), .B(n11144), .Z(n11146) );
  XNOR U11721 ( .A(n11147), .B(n11146), .Z(n11148) );
  XNOR U11722 ( .A(n11149), .B(n11148), .Z(n11150) );
  XNOR U11723 ( .A(n11151), .B(n11150), .Z(n11259) );
  NAND U11724 ( .A(n11153), .B(n11152), .Z(n11157) );
  NAND U11725 ( .A(n11155), .B(n11154), .Z(n11156) );
  AND U11726 ( .A(n11157), .B(n11156), .Z(n11257) );
  NANDN U11727 ( .A(n11159), .B(n11158), .Z(n11163) );
  NANDN U11728 ( .A(n11161), .B(n11160), .Z(n11162) );
  AND U11729 ( .A(n11163), .B(n11162), .Z(n11239) );
  NAND U11730 ( .A(n11165), .B(n11164), .Z(n11169) );
  NAND U11731 ( .A(n11167), .B(n11166), .Z(n11168) );
  AND U11732 ( .A(n11169), .B(n11168), .Z(n11177) );
  NAND U11733 ( .A(n11171), .B(n11170), .Z(n11175) );
  NAND U11734 ( .A(n11173), .B(n11172), .Z(n11174) );
  NAND U11735 ( .A(n11175), .B(n11174), .Z(n11176) );
  XNOR U11736 ( .A(n11177), .B(n11176), .Z(n11237) );
  AND U11737 ( .A(x[115]), .B(y[188]), .Z(n11179) );
  NAND U11738 ( .A(x[84]), .B(y[27]), .Z(n11178) );
  XNOR U11739 ( .A(n11179), .B(n11178), .Z(n11203) );
  AND U11740 ( .A(n11181), .B(n11180), .Z(n11197) );
  NAND U11741 ( .A(n11183), .B(n11182), .Z(n11187) );
  NAND U11742 ( .A(n11185), .B(n11184), .Z(n11186) );
  AND U11743 ( .A(n11187), .B(n11186), .Z(n11195) );
  AND U11744 ( .A(x[113]), .B(y[190]), .Z(n11189) );
  NAND U11745 ( .A(x[114]), .B(y[189]), .Z(n11188) );
  XNOR U11746 ( .A(n11189), .B(n11188), .Z(n11193) );
  AND U11747 ( .A(x[96]), .B(y[111]), .Z(n11191) );
  NAND U11748 ( .A(x[107]), .B(y[148]), .Z(n11190) );
  XNOR U11749 ( .A(n11191), .B(n11190), .Z(n11192) );
  XNOR U11750 ( .A(n11193), .B(n11192), .Z(n11194) );
  XNOR U11751 ( .A(n11195), .B(n11194), .Z(n11196) );
  XOR U11752 ( .A(n11197), .B(n11196), .Z(n11201) );
  XNOR U11753 ( .A(n11199), .B(n11198), .Z(n11200) );
  XNOR U11754 ( .A(n11201), .B(n11200), .Z(n11202) );
  XOR U11755 ( .A(n11203), .B(n11202), .Z(n11235) );
  NAND U11756 ( .A(n11205), .B(n11204), .Z(n11209) );
  NAND U11757 ( .A(n11207), .B(n11206), .Z(n11208) );
  AND U11758 ( .A(n11209), .B(n11208), .Z(n11217) );
  NAND U11759 ( .A(n11211), .B(n11210), .Z(n11215) );
  NAND U11760 ( .A(n11213), .B(n11212), .Z(n11214) );
  NAND U11761 ( .A(n11215), .B(n11214), .Z(n11216) );
  XNOR U11762 ( .A(n11217), .B(n11216), .Z(n11233) );
  NAND U11763 ( .A(n11219), .B(n11218), .Z(n11223) );
  NAND U11764 ( .A(n11221), .B(n11220), .Z(n11222) );
  AND U11765 ( .A(n11223), .B(n11222), .Z(n11231) );
  NAND U11766 ( .A(n11225), .B(n11224), .Z(n11229) );
  NAND U11767 ( .A(n11227), .B(n11226), .Z(n11228) );
  NAND U11768 ( .A(n11229), .B(n11228), .Z(n11230) );
  XNOR U11769 ( .A(n11231), .B(n11230), .Z(n11232) );
  XNOR U11770 ( .A(n11233), .B(n11232), .Z(n11234) );
  XNOR U11771 ( .A(n11235), .B(n11234), .Z(n11236) );
  XNOR U11772 ( .A(n11237), .B(n11236), .Z(n11238) );
  XNOR U11773 ( .A(n11239), .B(n11238), .Z(n11255) );
  NANDN U11774 ( .A(n11241), .B(n11240), .Z(n11245) );
  ANDN U11775 ( .B(n11243), .A(n11242), .Z(n11244) );
  ANDN U11776 ( .B(n11245), .A(n11244), .Z(n11253) );
  ANDN U11777 ( .B(n11247), .A(n11246), .Z(n11251) );
  AND U11778 ( .A(n11249), .B(n11248), .Z(n11250) );
  OR U11779 ( .A(n11251), .B(n11250), .Z(n11252) );
  XNOR U11780 ( .A(n11253), .B(n11252), .Z(n11254) );
  XNOR U11781 ( .A(n11255), .B(n11254), .Z(n11256) );
  XNOR U11782 ( .A(n11257), .B(n11256), .Z(n11258) );
  XNOR U11783 ( .A(n11259), .B(n11258), .Z(n11260) );
  XNOR U11784 ( .A(n11261), .B(n11260), .Z(n11262) );
  XNOR U11785 ( .A(n11263), .B(n11262), .Z(n11264) );
  XNOR U11786 ( .A(n11265), .B(n11264), .Z(n11281) );
  NAND U11787 ( .A(n11267), .B(n11266), .Z(n11271) );
  NAND U11788 ( .A(n11269), .B(n11268), .Z(n11270) );
  AND U11789 ( .A(n11271), .B(n11270), .Z(n11279) );
  NAND U11790 ( .A(n11273), .B(n11272), .Z(n11277) );
  NANDN U11791 ( .A(n11275), .B(n11274), .Z(n11276) );
  NAND U11792 ( .A(n11277), .B(n11276), .Z(n11278) );
  XNOR U11793 ( .A(n11279), .B(n11278), .Z(n11280) );
  NAND U11794 ( .A(y[192]), .B(x[112]), .Z(n11428) );
  NAND U11795 ( .A(y[72]), .B(x[88]), .Z(n11292) );
  XOR U11796 ( .A(n11428), .B(n11292), .Z(n11293) );
  AND U11797 ( .A(y[32]), .B(x[80]), .Z(n11300) );
  AND U11798 ( .A(y[112]), .B(x[96]), .Z(n11297) );
  XOR U11799 ( .A(n11300), .B(n11297), .Z(n11296) );
  AND U11800 ( .A(y[152]), .B(x[104]), .Z(n11295) );
  XNOR U11801 ( .A(n11296), .B(n11295), .Z(n11294) );
  XNOR U11802 ( .A(n11293), .B(n11294), .Z(o[112]) );
  AND U11803 ( .A(x[81]), .B(y[32]), .Z(n11291) );
  NAND U11804 ( .A(x[80]), .B(y[33]), .Z(n11290) );
  XNOR U11805 ( .A(n11291), .B(n11290), .Z(n11302) );
  AND U11806 ( .A(y[72]), .B(x[89]), .Z(n11301) );
  XOR U11807 ( .A(n11302), .B(n11301), .Z(n11319) );
  AND U11808 ( .A(y[192]), .B(x[113]), .Z(n11531) );
  AND U11809 ( .A(y[113]), .B(x[96]), .Z(n11305) );
  XOR U11810 ( .A(n11531), .B(n11305), .Z(n11307) );
  AND U11811 ( .A(y[193]), .B(x[112]), .Z(n11329) );
  NAND U11812 ( .A(y[112]), .B(x[97]), .Z(n11328) );
  XNOR U11813 ( .A(n11329), .B(n11328), .Z(n11306) );
  XOR U11814 ( .A(n11307), .B(n11306), .Z(n11317) );
  AND U11815 ( .A(y[73]), .B(x[88]), .Z(n11555) );
  AND U11816 ( .A(y[153]), .B(x[104]), .Z(n11322) );
  XOR U11817 ( .A(n11555), .B(n11322), .Z(n11324) );
  AND U11818 ( .A(y[152]), .B(x[105]), .Z(n11323) );
  XNOR U11819 ( .A(n11324), .B(n11323), .Z(n11316) );
  XNOR U11820 ( .A(n11317), .B(n11316), .Z(n11318) );
  XNOR U11821 ( .A(n11319), .B(n11318), .Z(n11313) );
  NAND U11822 ( .A(n11296), .B(n11295), .Z(n11299) );
  AND U11823 ( .A(n11300), .B(n11297), .Z(n11298) );
  ANDN U11824 ( .B(n11299), .A(n11298), .Z(n11310) );
  XNOR U11825 ( .A(n11311), .B(n11310), .Z(n11312) );
  XNOR U11826 ( .A(n11313), .B(n11312), .Z(o[113]) );
  NAND U11827 ( .A(y[33]), .B(x[81]), .Z(n11351) );
  NANDN U11828 ( .A(n11351), .B(n11300), .Z(n11304) );
  NAND U11829 ( .A(n11302), .B(n11301), .Z(n11303) );
  AND U11830 ( .A(n11304), .B(n11303), .Z(n11386) );
  NAND U11831 ( .A(n11531), .B(n11305), .Z(n11309) );
  NAND U11832 ( .A(n11307), .B(n11306), .Z(n11308) );
  AND U11833 ( .A(n11309), .B(n11308), .Z(n11385) );
  AND U11834 ( .A(y[154]), .B(x[104]), .Z(n11370) );
  NAND U11835 ( .A(y[34]), .B(x[80]), .Z(n11371) );
  XNOR U11836 ( .A(n11370), .B(n11371), .Z(n11372) );
  NAND U11837 ( .A(y[72]), .B(x[90]), .Z(n11373) );
  XNOR U11838 ( .A(n11372), .B(n11373), .Z(n11384) );
  XOR U11839 ( .A(n11385), .B(n11384), .Z(n11387) );
  XOR U11840 ( .A(n11386), .B(n11387), .Z(n11331) );
  NANDN U11841 ( .A(n11311), .B(n11310), .Z(n11315) );
  NAND U11842 ( .A(n11313), .B(n11312), .Z(n11314) );
  NAND U11843 ( .A(n11315), .B(n11314), .Z(n11330) );
  XNOR U11844 ( .A(n11331), .B(n11330), .Z(n11333) );
  NANDN U11845 ( .A(n11317), .B(n11316), .Z(n11321) );
  NANDN U11846 ( .A(n11319), .B(n11318), .Z(n11320) );
  AND U11847 ( .A(n11321), .B(n11320), .Z(n11339) );
  AND U11848 ( .A(y[32]), .B(x[82]), .Z(n11348) );
  NAND U11849 ( .A(y[114]), .B(x[96]), .Z(n11349) );
  XNOR U11850 ( .A(n11348), .B(n11349), .Z(n11350) );
  AND U11851 ( .A(y[152]), .B(x[106]), .Z(n11378) );
  XOR U11852 ( .A(n11379), .B(n11378), .Z(n11381) );
  AND U11853 ( .A(y[112]), .B(x[98]), .Z(n11458) );
  AND U11854 ( .A(y[194]), .B(x[112]), .Z(n11361) );
  XOR U11855 ( .A(n11458), .B(n11361), .Z(n11363) );
  AND U11856 ( .A(y[113]), .B(x[97]), .Z(n11362) );
  XOR U11857 ( .A(n11363), .B(n11362), .Z(n11380) );
  XOR U11858 ( .A(n11381), .B(n11380), .Z(n11336) );
  NAND U11859 ( .A(n11555), .B(n11322), .Z(n11326) );
  AND U11860 ( .A(n11324), .B(n11323), .Z(n11325) );
  ANDN U11861 ( .B(n11326), .A(n11325), .Z(n11345) );
  AND U11862 ( .A(x[113]), .B(y[193]), .Z(n11433) );
  NAND U11863 ( .A(x[114]), .B(y[192]), .Z(n11327) );
  XNOR U11864 ( .A(n11433), .B(n11327), .Z(n11377) );
  ANDN U11865 ( .B(n11329), .A(n11328), .Z(n11376) );
  XOR U11866 ( .A(n11377), .B(n11376), .Z(n11342) );
  AND U11867 ( .A(y[153]), .B(x[105]), .Z(n11354) );
  NAND U11868 ( .A(y[73]), .B(x[89]), .Z(n11355) );
  XNOR U11869 ( .A(n11354), .B(n11355), .Z(n11356) );
  NAND U11870 ( .A(y[74]), .B(x[88]), .Z(n11357) );
  XOR U11871 ( .A(n11356), .B(n11357), .Z(n11343) );
  XNOR U11872 ( .A(n11342), .B(n11343), .Z(n11344) );
  XOR U11873 ( .A(n11345), .B(n11344), .Z(n11337) );
  XNOR U11874 ( .A(n11336), .B(n11337), .Z(n11338) );
  XNOR U11875 ( .A(n11339), .B(n11338), .Z(n11332) );
  XNOR U11876 ( .A(n11333), .B(n11332), .Z(o[114]) );
  NANDN U11877 ( .A(n11331), .B(n11330), .Z(n11335) );
  NAND U11878 ( .A(n11333), .B(n11332), .Z(n11334) );
  AND U11879 ( .A(n11335), .B(n11334), .Z(n11408) );
  NANDN U11880 ( .A(n11337), .B(n11336), .Z(n11341) );
  NAND U11881 ( .A(n11339), .B(n11338), .Z(n11340) );
  AND U11882 ( .A(n11341), .B(n11340), .Z(n11393) );
  NANDN U11883 ( .A(n11343), .B(n11342), .Z(n11347) );
  NANDN U11884 ( .A(n11345), .B(n11344), .Z(n11346) );
  AND U11885 ( .A(n11347), .B(n11346), .Z(n11391) );
  NANDN U11886 ( .A(n11349), .B(n11348), .Z(n11353) );
  NANDN U11887 ( .A(n11351), .B(n11350), .Z(n11352) );
  NAND U11888 ( .A(n11353), .B(n11352), .Z(n11402) );
  NANDN U11889 ( .A(n11355), .B(n11354), .Z(n11359) );
  NANDN U11890 ( .A(n11357), .B(n11356), .Z(n11358) );
  AND U11891 ( .A(n11359), .B(n11358), .Z(n11449) );
  AND U11892 ( .A(y[155]), .B(x[104]), .Z(n11477) );
  AND U11893 ( .A(y[115]), .B(x[96]), .Z(n11476) );
  NAND U11894 ( .A(y[32]), .B(x[83]), .Z(n11475) );
  XOR U11895 ( .A(n11476), .B(n11475), .Z(n11478) );
  XOR U11896 ( .A(n11477), .B(n11478), .Z(n11447) );
  AND U11897 ( .A(x[98]), .B(y[113]), .Z(n11511) );
  NAND U11898 ( .A(x[99]), .B(y[112]), .Z(n11360) );
  XNOR U11899 ( .A(n11511), .B(n11360), .Z(n11460) );
  NAND U11900 ( .A(y[114]), .B(x[97]), .Z(n11461) );
  XNOR U11901 ( .A(n11460), .B(n11461), .Z(n11446) );
  XNOR U11902 ( .A(n11447), .B(n11446), .Z(n11448) );
  XNOR U11903 ( .A(n11449), .B(n11448), .Z(n11403) );
  XOR U11904 ( .A(n11402), .B(n11403), .Z(n11405) );
  NAND U11905 ( .A(n11458), .B(n11361), .Z(n11365) );
  AND U11906 ( .A(n11363), .B(n11362), .Z(n11364) );
  ANDN U11907 ( .B(n11365), .A(n11364), .Z(n11454) );
  AND U11908 ( .A(y[34]), .B(x[81]), .Z(n11424) );
  AND U11909 ( .A(y[33]), .B(x[82]), .Z(n11423) );
  NAND U11910 ( .A(y[154]), .B(x[105]), .Z(n11422) );
  XOR U11911 ( .A(n11423), .B(n11422), .Z(n11425) );
  XOR U11912 ( .A(n11424), .B(n11425), .Z(n11453) );
  AND U11913 ( .A(x[115]), .B(y[192]), .Z(n11367) );
  NAND U11914 ( .A(x[112]), .B(y[195]), .Z(n11366) );
  XNOR U11915 ( .A(n11367), .B(n11366), .Z(n11429) );
  AND U11916 ( .A(x[113]), .B(y[194]), .Z(n11369) );
  NAND U11917 ( .A(x[114]), .B(y[193]), .Z(n11368) );
  XOR U11918 ( .A(n11369), .B(n11368), .Z(n11430) );
  XNOR U11919 ( .A(n11429), .B(n11430), .Z(n11452) );
  XOR U11920 ( .A(n11453), .B(n11452), .Z(n11455) );
  XOR U11921 ( .A(n11454), .B(n11455), .Z(n11404) );
  XOR U11922 ( .A(n11405), .B(n11404), .Z(n11390) );
  XNOR U11923 ( .A(n11391), .B(n11390), .Z(n11392) );
  XOR U11924 ( .A(n11393), .B(n11392), .Z(n11409) );
  XNOR U11925 ( .A(n11408), .B(n11409), .Z(n11411) );
  NANDN U11926 ( .A(n11371), .B(n11370), .Z(n11375) );
  NANDN U11927 ( .A(n11373), .B(n11372), .Z(n11374) );
  AND U11928 ( .A(n11375), .B(n11374), .Z(n11415) );
  AND U11929 ( .A(y[193]), .B(x[114]), .Z(n11530) );
  XNOR U11930 ( .A(n11415), .B(n11414), .Z(n11417) );
  AND U11931 ( .A(y[72]), .B(x[91]), .Z(n11468) );
  AND U11932 ( .A(y[35]), .B(x[80]), .Z(n11467) );
  NAND U11933 ( .A(y[153]), .B(x[106]), .Z(n11466) );
  XOR U11934 ( .A(n11467), .B(n11466), .Z(n11469) );
  XOR U11935 ( .A(n11468), .B(n11469), .Z(n11443) );
  AND U11936 ( .A(y[75]), .B(x[88]), .Z(n11436) );
  AND U11937 ( .A(y[73]), .B(x[90]), .Z(n11435) );
  NAND U11938 ( .A(y[152]), .B(x[107]), .Z(n11434) );
  XOR U11939 ( .A(n11435), .B(n11434), .Z(n11437) );
  XOR U11940 ( .A(n11436), .B(n11437), .Z(n11441) );
  AND U11941 ( .A(y[74]), .B(x[89]), .Z(n11440) );
  XNOR U11942 ( .A(n11441), .B(n11440), .Z(n11442) );
  XNOR U11943 ( .A(n11443), .B(n11442), .Z(n11416) );
  XOR U11944 ( .A(n11417), .B(n11416), .Z(n11397) );
  NAND U11945 ( .A(n11379), .B(n11378), .Z(n11383) );
  NAND U11946 ( .A(n11381), .B(n11380), .Z(n11382) );
  AND U11947 ( .A(n11383), .B(n11382), .Z(n11396) );
  XNOR U11948 ( .A(n11397), .B(n11396), .Z(n11399) );
  NANDN U11949 ( .A(n11385), .B(n11384), .Z(n11389) );
  OR U11950 ( .A(n11387), .B(n11386), .Z(n11388) );
  AND U11951 ( .A(n11389), .B(n11388), .Z(n11398) );
  XNOR U11952 ( .A(n11399), .B(n11398), .Z(n11410) );
  XOR U11953 ( .A(n11411), .B(n11410), .Z(o[115]) );
  NANDN U11954 ( .A(n11391), .B(n11390), .Z(n11395) );
  NANDN U11955 ( .A(n11393), .B(n11392), .Z(n11394) );
  AND U11956 ( .A(n11395), .B(n11394), .Z(n11489) );
  NANDN U11957 ( .A(n11397), .B(n11396), .Z(n11401) );
  NAND U11958 ( .A(n11399), .B(n11398), .Z(n11400) );
  NAND U11959 ( .A(n11401), .B(n11400), .Z(n11487) );
  NAND U11960 ( .A(n11403), .B(n11402), .Z(n11407) );
  NAND U11961 ( .A(n11405), .B(n11404), .Z(n11406) );
  AND U11962 ( .A(n11407), .B(n11406), .Z(n11488) );
  XOR U11963 ( .A(n11487), .B(n11488), .Z(n11490) );
  XOR U11964 ( .A(n11489), .B(n11490), .Z(n11481) );
  NANDN U11965 ( .A(n11409), .B(n11408), .Z(n11413) );
  NAND U11966 ( .A(n11411), .B(n11410), .Z(n11412) );
  NAND U11967 ( .A(n11413), .B(n11412), .Z(n11482) );
  XNOR U11968 ( .A(n11481), .B(n11482), .Z(n11484) );
  NANDN U11969 ( .A(n11415), .B(n11414), .Z(n11419) );
  NAND U11970 ( .A(n11417), .B(n11416), .Z(n11418) );
  AND U11971 ( .A(n11419), .B(n11418), .Z(n11494) );
  AND U11972 ( .A(y[74]), .B(x[90]), .Z(n11618) );
  AND U11973 ( .A(x[88]), .B(y[76]), .Z(n11421) );
  NAND U11974 ( .A(x[91]), .B(y[73]), .Z(n11420) );
  XOR U11975 ( .A(n11421), .B(n11420), .Z(n11556) );
  XNOR U11976 ( .A(n11618), .B(n11556), .Z(n11565) );
  NAND U11977 ( .A(y[75]), .B(x[89]), .Z(n11566) );
  XNOR U11978 ( .A(n11565), .B(n11566), .Z(n11568) );
  AND U11979 ( .A(y[152]), .B(x[108]), .Z(n11516) );
  NAND U11980 ( .A(y[35]), .B(x[81]), .Z(n11517) );
  XNOR U11981 ( .A(n11516), .B(n11517), .Z(n11518) );
  NAND U11982 ( .A(y[36]), .B(x[80]), .Z(n11519) );
  XNOR U11983 ( .A(n11518), .B(n11519), .Z(n11567) );
  XOR U11984 ( .A(n11568), .B(n11567), .Z(n11562) );
  NANDN U11985 ( .A(n11423), .B(n11422), .Z(n11427) );
  OR U11986 ( .A(n11425), .B(n11424), .Z(n11426) );
  AND U11987 ( .A(n11427), .B(n11426), .Z(n11560) );
  AND U11988 ( .A(y[195]), .B(x[115]), .Z(n11879) );
  NANDN U11989 ( .A(n11428), .B(n11879), .Z(n11432) );
  NANDN U11990 ( .A(n11430), .B(n11429), .Z(n11431) );
  AND U11991 ( .A(n11432), .B(n11431), .Z(n11559) );
  XNOR U11992 ( .A(n11560), .B(n11559), .Z(n11561) );
  XNOR U11993 ( .A(n11562), .B(n11561), .Z(n11592) );
  NAND U11994 ( .A(y[32]), .B(x[84]), .Z(n11540) );
  NAND U11995 ( .A(y[154]), .B(x[106]), .Z(n11539) );
  NAND U11996 ( .A(y[116]), .B(x[96]), .Z(n11538) );
  XNOR U11997 ( .A(n11539), .B(n11538), .Z(n11541) );
  AND U11998 ( .A(x[114]), .B(y[194]), .Z(n11474) );
  NAND U11999 ( .A(n11433), .B(n11474), .Z(n11536) );
  NAND U12000 ( .A(y[196]), .B(x[112]), .Z(n11716) );
  NAND U12001 ( .A(y[112]), .B(x[100]), .Z(n11639) );
  XNOR U12002 ( .A(n11716), .B(n11639), .Z(n11537) );
  XOR U12003 ( .A(n11536), .B(n11537), .Z(n11499) );
  XOR U12004 ( .A(n11500), .B(n11499), .Z(n11502) );
  NANDN U12005 ( .A(n11435), .B(n11434), .Z(n11439) );
  OR U12006 ( .A(n11437), .B(n11436), .Z(n11438) );
  AND U12007 ( .A(n11439), .B(n11438), .Z(n11501) );
  XOR U12008 ( .A(n11502), .B(n11501), .Z(n11590) );
  NANDN U12009 ( .A(n11441), .B(n11440), .Z(n11445) );
  NANDN U12010 ( .A(n11443), .B(n11442), .Z(n11444) );
  AND U12011 ( .A(n11445), .B(n11444), .Z(n11589) );
  XNOR U12012 ( .A(n11590), .B(n11589), .Z(n11591) );
  XNOR U12013 ( .A(n11592), .B(n11591), .Z(n11493) );
  XNOR U12014 ( .A(n11494), .B(n11493), .Z(n11496) );
  NANDN U12015 ( .A(n11447), .B(n11446), .Z(n11451) );
  NANDN U12016 ( .A(n11449), .B(n11448), .Z(n11450) );
  AND U12017 ( .A(n11451), .B(n11450), .Z(n11578) );
  NANDN U12018 ( .A(n11453), .B(n11452), .Z(n11457) );
  OR U12019 ( .A(n11455), .B(n11454), .Z(n11456) );
  NAND U12020 ( .A(n11457), .B(n11456), .Z(n11577) );
  XNOR U12021 ( .A(n11578), .B(n11577), .Z(n11579) );
  AND U12022 ( .A(y[113]), .B(x[99]), .Z(n11459) );
  NAND U12023 ( .A(n11459), .B(n11458), .Z(n11463) );
  NANDN U12024 ( .A(n11461), .B(n11460), .Z(n11462) );
  AND U12025 ( .A(n11463), .B(n11462), .Z(n11584) );
  AND U12026 ( .A(y[72]), .B(x[92]), .Z(n11522) );
  NAND U12027 ( .A(y[156]), .B(x[104]), .Z(n11523) );
  XNOR U12028 ( .A(n11522), .B(n11523), .Z(n11524) );
  NAND U12029 ( .A(y[155]), .B(x[105]), .Z(n11525) );
  XNOR U12030 ( .A(n11524), .B(n11525), .Z(n11571) );
  AND U12031 ( .A(x[98]), .B(y[114]), .Z(n11465) );
  NAND U12032 ( .A(x[99]), .B(y[113]), .Z(n11464) );
  XNOR U12033 ( .A(n11465), .B(n11464), .Z(n11512) );
  NAND U12034 ( .A(y[115]), .B(x[97]), .Z(n11513) );
  XOR U12035 ( .A(n11512), .B(n11513), .Z(n11572) );
  XNOR U12036 ( .A(n11571), .B(n11572), .Z(n11573) );
  NANDN U12037 ( .A(n11467), .B(n11466), .Z(n11471) );
  OR U12038 ( .A(n11469), .B(n11468), .Z(n11470) );
  NAND U12039 ( .A(n11471), .B(n11470), .Z(n11574) );
  XNOR U12040 ( .A(n11573), .B(n11574), .Z(n11583) );
  XNOR U12041 ( .A(n11584), .B(n11583), .Z(n11585) );
  NAND U12042 ( .A(y[34]), .B(x[82]), .Z(n11551) );
  NAND U12043 ( .A(y[153]), .B(x[107]), .Z(n11550) );
  NAND U12044 ( .A(y[33]), .B(x[83]), .Z(n11549) );
  XNOR U12045 ( .A(n11550), .B(n11549), .Z(n11552) );
  AND U12046 ( .A(x[116]), .B(y[192]), .Z(n11473) );
  NAND U12047 ( .A(x[113]), .B(y[195]), .Z(n11472) );
  XNOR U12048 ( .A(n11473), .B(n11472), .Z(n11533) );
  AND U12049 ( .A(x[115]), .B(y[193]), .Z(n11646) );
  XOR U12050 ( .A(n11474), .B(n11646), .Z(n11532) );
  XOR U12051 ( .A(n11533), .B(n11532), .Z(n11505) );
  XOR U12052 ( .A(n11506), .B(n11505), .Z(n11507) );
  NANDN U12053 ( .A(n11476), .B(n11475), .Z(n11480) );
  OR U12054 ( .A(n11478), .B(n11477), .Z(n11479) );
  NAND U12055 ( .A(n11480), .B(n11479), .Z(n11508) );
  XOR U12056 ( .A(n11507), .B(n11508), .Z(n11586) );
  XOR U12057 ( .A(n11585), .B(n11586), .Z(n11580) );
  XNOR U12058 ( .A(n11579), .B(n11580), .Z(n11495) );
  XNOR U12059 ( .A(n11496), .B(n11495), .Z(n11483) );
  XNOR U12060 ( .A(n11484), .B(n11483), .Z(o[116]) );
  NANDN U12061 ( .A(n11482), .B(n11481), .Z(n11486) );
  NAND U12062 ( .A(n11484), .B(n11483), .Z(n11485) );
  AND U12063 ( .A(n11486), .B(n11485), .Z(n11734) );
  NAND U12064 ( .A(n11488), .B(n11487), .Z(n11492) );
  NAND U12065 ( .A(n11490), .B(n11489), .Z(n11491) );
  NAND U12066 ( .A(n11492), .B(n11491), .Z(n11735) );
  XNOR U12067 ( .A(n11734), .B(n11735), .Z(n11737) );
  NANDN U12068 ( .A(n11494), .B(n11493), .Z(n11498) );
  NAND U12069 ( .A(n11496), .B(n11495), .Z(n11497) );
  AND U12070 ( .A(n11498), .B(n11497), .Z(n11596) );
  NAND U12071 ( .A(n11500), .B(n11499), .Z(n11504) );
  NAND U12072 ( .A(n11502), .B(n11501), .Z(n11503) );
  AND U12073 ( .A(n11504), .B(n11503), .Z(n11648) );
  NAND U12074 ( .A(n11506), .B(n11505), .Z(n11510) );
  NANDN U12075 ( .A(n11508), .B(n11507), .Z(n11509) );
  NAND U12076 ( .A(n11510), .B(n11509), .Z(n11647) );
  XNOR U12077 ( .A(n11648), .B(n11647), .Z(n11650) );
  AND U12078 ( .A(y[114]), .B(x[99]), .Z(n11640) );
  NAND U12079 ( .A(n11640), .B(n11511), .Z(n11515) );
  NANDN U12080 ( .A(n11513), .B(n11512), .Z(n11514) );
  AND U12081 ( .A(n11515), .B(n11514), .Z(n11602) );
  NANDN U12082 ( .A(n11517), .B(n11516), .Z(n11521) );
  NANDN U12083 ( .A(n11519), .B(n11518), .Z(n11520) );
  NAND U12084 ( .A(n11521), .B(n11520), .Z(n11609) );
  AND U12085 ( .A(y[157]), .B(x[104]), .Z(n11784) );
  AND U12086 ( .A(y[72]), .B(x[93]), .Z(n11630) );
  AND U12087 ( .A(y[115]), .B(x[98]), .Z(n11629) );
  XOR U12088 ( .A(n11630), .B(n11629), .Z(n11631) );
  XOR U12089 ( .A(n11784), .B(n11631), .Z(n11608) );
  AND U12090 ( .A(y[153]), .B(x[108]), .Z(n11635) );
  AND U12091 ( .A(y[32]), .B(x[85]), .Z(n11634) );
  XOR U12092 ( .A(n11635), .B(n11634), .Z(n11636) );
  AND U12093 ( .A(y[33]), .B(x[84]), .Z(n11841) );
  XOR U12094 ( .A(n11636), .B(n11841), .Z(n11607) );
  XOR U12095 ( .A(n11608), .B(n11607), .Z(n11610) );
  XOR U12096 ( .A(n11609), .B(n11610), .Z(n11601) );
  NANDN U12097 ( .A(n11523), .B(n11522), .Z(n11527) );
  NANDN U12098 ( .A(n11525), .B(n11524), .Z(n11526) );
  NAND U12099 ( .A(n11527), .B(n11526), .Z(n11699) );
  AND U12100 ( .A(x[112]), .B(y[197]), .Z(n11529) );
  NAND U12101 ( .A(x[113]), .B(y[196]), .Z(n11528) );
  XNOR U12102 ( .A(n11529), .B(n11528), .Z(n11718) );
  AND U12103 ( .A(y[194]), .B(x[115]), .Z(n11546) );
  AND U12104 ( .A(n11530), .B(n11546), .Z(n11717) );
  XOR U12105 ( .A(n11718), .B(n11717), .Z(n11698) );
  AND U12106 ( .A(y[77]), .B(x[88]), .Z(n11688) );
  AND U12107 ( .A(y[36]), .B(x[81]), .Z(n11687) );
  XOR U12108 ( .A(n11688), .B(n11687), .Z(n11690) );
  AND U12109 ( .A(y[73]), .B(x[92]), .Z(n11689) );
  XOR U12110 ( .A(n11690), .B(n11689), .Z(n11697) );
  XOR U12111 ( .A(n11698), .B(n11697), .Z(n11700) );
  XOR U12112 ( .A(n11699), .B(n11700), .Z(n11603) );
  XOR U12113 ( .A(n11604), .B(n11603), .Z(n11649) );
  XOR U12114 ( .A(n11650), .B(n11649), .Z(n11723) );
  AND U12115 ( .A(y[195]), .B(x[116]), .Z(n11814) );
  NAND U12116 ( .A(n11814), .B(n11531), .Z(n11535) );
  NAND U12117 ( .A(n11533), .B(n11532), .Z(n11534) );
  AND U12118 ( .A(n11535), .B(n11534), .Z(n11656) );
  XNOR U12119 ( .A(n11656), .B(n11655), .Z(n11658) );
  NAND U12120 ( .A(n11539), .B(n11538), .Z(n11543) );
  NANDN U12121 ( .A(n11541), .B(n11540), .Z(n11542) );
  AND U12122 ( .A(n11543), .B(n11542), .Z(n11664) );
  AND U12123 ( .A(y[74]), .B(x[91]), .Z(n11970) );
  NAND U12124 ( .A(x[90]), .B(y[75]), .Z(n11544) );
  XNOR U12125 ( .A(n11970), .B(n11544), .Z(n11619) );
  NAND U12126 ( .A(y[76]), .B(x[89]), .Z(n11620) );
  XNOR U12127 ( .A(n11619), .B(n11620), .Z(n11662) );
  AND U12128 ( .A(y[195]), .B(x[114]), .Z(n11611) );
  NAND U12129 ( .A(y[192]), .B(x[117]), .Z(n11612) );
  XNOR U12130 ( .A(n11611), .B(n11612), .Z(n11613) );
  NAND U12131 ( .A(x[116]), .B(y[193]), .Z(n11545) );
  XOR U12132 ( .A(n11546), .B(n11545), .Z(n11614) );
  XNOR U12133 ( .A(n11613), .B(n11614), .Z(n11661) );
  XOR U12134 ( .A(n11662), .B(n11661), .Z(n11663) );
  XOR U12135 ( .A(n11664), .B(n11663), .Z(n11657) );
  XOR U12136 ( .A(n11658), .B(n11657), .Z(n11675) );
  AND U12137 ( .A(x[100]), .B(y[113]), .Z(n11548) );
  NAND U12138 ( .A(x[101]), .B(y[112]), .Z(n11547) );
  XOR U12139 ( .A(n11548), .B(n11547), .Z(n11641) );
  XNOR U12140 ( .A(n11640), .B(n11641), .Z(n11680) );
  AND U12141 ( .A(y[152]), .B(x[109]), .Z(n11623) );
  NAND U12142 ( .A(y[34]), .B(x[83]), .Z(n11624) );
  XNOR U12143 ( .A(n11623), .B(n11624), .Z(n11626) );
  AND U12144 ( .A(y[35]), .B(x[82]), .Z(n11625) );
  XOR U12145 ( .A(n11626), .B(n11625), .Z(n11679) );
  XOR U12146 ( .A(n11680), .B(n11679), .Z(n11682) );
  NAND U12147 ( .A(n11550), .B(n11549), .Z(n11554) );
  NANDN U12148 ( .A(n11552), .B(n11551), .Z(n11553) );
  AND U12149 ( .A(n11554), .B(n11553), .Z(n11681) );
  XOR U12150 ( .A(n11682), .B(n11681), .Z(n11674) );
  AND U12151 ( .A(y[76]), .B(x[91]), .Z(n11936) );
  NAND U12152 ( .A(n11936), .B(n11555), .Z(n11558) );
  NANDN U12153 ( .A(n11556), .B(n11618), .Z(n11557) );
  AND U12154 ( .A(n11558), .B(n11557), .Z(n11654) );
  AND U12155 ( .A(y[154]), .B(x[107]), .Z(n11703) );
  AND U12156 ( .A(y[116]), .B(x[97]), .Z(n11835) );
  XOR U12157 ( .A(n11703), .B(n11835), .Z(n11705) );
  AND U12158 ( .A(y[117]), .B(x[96]), .Z(n11704) );
  XOR U12159 ( .A(n11705), .B(n11704), .Z(n11652) );
  AND U12160 ( .A(y[37]), .B(x[80]), .Z(n11709) );
  AND U12161 ( .A(y[156]), .B(x[105]), .Z(n11708) );
  XOR U12162 ( .A(n11709), .B(n11708), .Z(n11711) );
  AND U12163 ( .A(y[155]), .B(x[106]), .Z(n11710) );
  XOR U12164 ( .A(n11711), .B(n11710), .Z(n11651) );
  XOR U12165 ( .A(n11652), .B(n11651), .Z(n11653) );
  XOR U12166 ( .A(n11654), .B(n11653), .Z(n11673) );
  XOR U12167 ( .A(n11674), .B(n11673), .Z(n11676) );
  XOR U12168 ( .A(n11675), .B(n11676), .Z(n11722) );
  NANDN U12169 ( .A(n11560), .B(n11559), .Z(n11564) );
  NANDN U12170 ( .A(n11562), .B(n11561), .Z(n11563) );
  AND U12171 ( .A(n11564), .B(n11563), .Z(n11669) );
  NANDN U12172 ( .A(n11566), .B(n11565), .Z(n11570) );
  NAND U12173 ( .A(n11568), .B(n11567), .Z(n11569) );
  AND U12174 ( .A(n11570), .B(n11569), .Z(n11668) );
  NANDN U12175 ( .A(n11572), .B(n11571), .Z(n11576) );
  NANDN U12176 ( .A(n11574), .B(n11573), .Z(n11575) );
  NAND U12177 ( .A(n11576), .B(n11575), .Z(n11667) );
  XOR U12178 ( .A(n11668), .B(n11667), .Z(n11670) );
  XNOR U12179 ( .A(n11669), .B(n11670), .Z(n11721) );
  XOR U12180 ( .A(n11722), .B(n11721), .Z(n11724) );
  XNOR U12181 ( .A(n11723), .B(n11724), .Z(n11595) );
  XNOR U12182 ( .A(n11596), .B(n11595), .Z(n11597) );
  NANDN U12183 ( .A(n11578), .B(n11577), .Z(n11582) );
  NANDN U12184 ( .A(n11580), .B(n11579), .Z(n11581) );
  AND U12185 ( .A(n11582), .B(n11581), .Z(n11730) );
  NANDN U12186 ( .A(n11584), .B(n11583), .Z(n11588) );
  NANDN U12187 ( .A(n11586), .B(n11585), .Z(n11587) );
  AND U12188 ( .A(n11588), .B(n11587), .Z(n11728) );
  NANDN U12189 ( .A(n11590), .B(n11589), .Z(n11594) );
  NAND U12190 ( .A(n11592), .B(n11591), .Z(n11593) );
  AND U12191 ( .A(n11594), .B(n11593), .Z(n11727) );
  XNOR U12192 ( .A(n11728), .B(n11727), .Z(n11729) );
  XOR U12193 ( .A(n11730), .B(n11729), .Z(n11598) );
  XNOR U12194 ( .A(n11597), .B(n11598), .Z(n11736) );
  XOR U12195 ( .A(n11737), .B(n11736), .Z(o[117]) );
  NANDN U12196 ( .A(n11596), .B(n11595), .Z(n11600) );
  NANDN U12197 ( .A(n11598), .B(n11597), .Z(n11599) );
  AND U12198 ( .A(n11600), .B(n11599), .Z(n12022) );
  NANDN U12199 ( .A(n11602), .B(n11601), .Z(n11606) );
  NAND U12200 ( .A(n11604), .B(n11603), .Z(n11605) );
  AND U12201 ( .A(n11606), .B(n11605), .Z(n12027) );
  NANDN U12202 ( .A(n11612), .B(n11611), .Z(n11616) );
  NANDN U12203 ( .A(n11614), .B(n11613), .Z(n11615) );
  NAND U12204 ( .A(n11616), .B(n11615), .Z(n11770) );
  AND U12205 ( .A(y[75]), .B(x[91]), .Z(n11617) );
  NAND U12206 ( .A(n11618), .B(n11617), .Z(n11622) );
  NANDN U12207 ( .A(n11620), .B(n11619), .Z(n11621) );
  AND U12208 ( .A(n11622), .B(n11621), .Z(n11985) );
  AND U12209 ( .A(y[155]), .B(x[107]), .Z(n11976) );
  AND U12210 ( .A(y[115]), .B(x[99]), .Z(n11975) );
  XOR U12211 ( .A(n11976), .B(n11975), .Z(n11974) );
  AND U12212 ( .A(y[35]), .B(x[83]), .Z(n11973) );
  XOR U12213 ( .A(n11974), .B(n11973), .Z(n11988) );
  AND U12214 ( .A(y[156]), .B(x[106]), .Z(n11828) );
  AND U12215 ( .A(y[114]), .B(x[100]), .Z(n11827) );
  XOR U12216 ( .A(n11828), .B(n11827), .Z(n11826) );
  AND U12217 ( .A(y[36]), .B(x[82]), .Z(n11825) );
  XNOR U12218 ( .A(n11826), .B(n11825), .Z(n11987) );
  XNOR U12219 ( .A(n11985), .B(n11986), .Z(n11773) );
  NANDN U12220 ( .A(n11624), .B(n11623), .Z(n11628) );
  NAND U12221 ( .A(n11626), .B(n11625), .Z(n11627) );
  NAND U12222 ( .A(n11628), .B(n11627), .Z(n11772) );
  XOR U12223 ( .A(n11770), .B(n11771), .Z(n11767) );
  XOR U12224 ( .A(n11766), .B(n11767), .Z(n11765) );
  NAND U12225 ( .A(n11630), .B(n11629), .Z(n11633) );
  NAND U12226 ( .A(n11784), .B(n11631), .Z(n11632) );
  NAND U12227 ( .A(n11633), .B(n11632), .Z(n11875) );
  NAND U12228 ( .A(n11635), .B(n11634), .Z(n11638) );
  NAND U12229 ( .A(n11636), .B(n11841), .Z(n11637) );
  NAND U12230 ( .A(n11638), .B(n11637), .Z(n11874) );
  XOR U12231 ( .A(n11875), .B(n11874), .Z(n11873) );
  AND U12232 ( .A(y[113]), .B(x[101]), .Z(n11790) );
  NANDN U12233 ( .A(n11639), .B(n11790), .Z(n11643) );
  NANDN U12234 ( .A(n11641), .B(n11640), .Z(n11642) );
  AND U12235 ( .A(n11643), .B(n11642), .Z(n11861) );
  AND U12236 ( .A(x[85]), .B(y[33]), .Z(n11645) );
  NAND U12237 ( .A(x[84]), .B(y[34]), .Z(n11644) );
  XNOR U12238 ( .A(n11645), .B(n11644), .Z(n11839) );
  AND U12239 ( .A(y[152]), .B(x[110]), .Z(n11838) );
  XOR U12240 ( .A(n11839), .B(n11838), .Z(n11863) );
  AND U12241 ( .A(y[197]), .B(x[113]), .Z(n11960) );
  AND U12242 ( .A(x[116]), .B(y[194]), .Z(n11715) );
  AND U12243 ( .A(n11646), .B(n11715), .Z(n11962) );
  AND U12244 ( .A(y[196]), .B(x[114]), .Z(n11961) );
  XOR U12245 ( .A(n11962), .B(n11961), .Z(n11959) );
  XNOR U12246 ( .A(n11960), .B(n11959), .Z(n11862) );
  XNOR U12247 ( .A(n11861), .B(n11860), .Z(n11872) );
  XOR U12248 ( .A(n11873), .B(n11872), .Z(n11764) );
  XOR U12249 ( .A(n11765), .B(n11764), .Z(n11743) );
  NANDN U12250 ( .A(n11656), .B(n11655), .Z(n11660) );
  NAND U12251 ( .A(n11658), .B(n11657), .Z(n11659) );
  AND U12252 ( .A(n11660), .B(n11659), .Z(n11758) );
  XOR U12253 ( .A(n11759), .B(n11758), .Z(n11757) );
  NAND U12254 ( .A(n11662), .B(n11661), .Z(n11666) );
  NAND U12255 ( .A(n11664), .B(n11663), .Z(n11665) );
  AND U12256 ( .A(n11666), .B(n11665), .Z(n11756) );
  XOR U12257 ( .A(n11757), .B(n11756), .Z(n11740) );
  XOR U12258 ( .A(n11741), .B(n11740), .Z(n12026) );
  XOR U12259 ( .A(n12027), .B(n12026), .Z(n12029) );
  NANDN U12260 ( .A(n11668), .B(n11667), .Z(n11672) );
  NANDN U12261 ( .A(n11670), .B(n11669), .Z(n11671) );
  AND U12262 ( .A(n11672), .B(n11671), .Z(n12005) );
  NANDN U12263 ( .A(n11674), .B(n11673), .Z(n11678) );
  OR U12264 ( .A(n11676), .B(n11675), .Z(n11677) );
  NAND U12265 ( .A(n11678), .B(n11677), .Z(n12007) );
  NAND U12266 ( .A(n11680), .B(n11679), .Z(n11684) );
  NAND U12267 ( .A(n11682), .B(n11681), .Z(n11683) );
  AND U12268 ( .A(n11684), .B(n11683), .Z(n12014) );
  AND U12269 ( .A(y[118]), .B(x[96]), .Z(n11801) );
  AND U12270 ( .A(y[32]), .B(x[86]), .Z(n11800) );
  XOR U12271 ( .A(n11801), .B(n11800), .Z(n11799) );
  AND U12272 ( .A(y[153]), .B(x[109]), .Z(n11798) );
  XOR U12273 ( .A(n11799), .B(n11798), .Z(n11857) );
  AND U12274 ( .A(y[73]), .B(x[93]), .Z(n11822) );
  AND U12275 ( .A(y[76]), .B(x[90]), .Z(n11821) );
  XOR U12276 ( .A(n11822), .B(n11821), .Z(n11820) );
  AND U12277 ( .A(y[77]), .B(x[89]), .Z(n11819) );
  XOR U12278 ( .A(n11820), .B(n11819), .Z(n11968) );
  AND U12279 ( .A(x[92]), .B(y[74]), .Z(n11686) );
  NAND U12280 ( .A(x[91]), .B(y[75]), .Z(n11685) );
  XNOR U12281 ( .A(n11686), .B(n11685), .Z(n11967) );
  XOR U12282 ( .A(n11968), .B(n11967), .Z(n11856) );
  XOR U12283 ( .A(n11857), .B(n11856), .Z(n11855) );
  AND U12284 ( .A(y[198]), .B(x[112]), .Z(n11789) );
  XOR U12285 ( .A(n11790), .B(n11789), .Z(n11788) );
  AND U12286 ( .A(y[112]), .B(x[102]), .Z(n11787) );
  XOR U12287 ( .A(n11788), .B(n11787), .Z(n11854) );
  XOR U12288 ( .A(n11855), .B(n11854), .Z(n11753) );
  NAND U12289 ( .A(n11688), .B(n11687), .Z(n11692) );
  NAND U12290 ( .A(n11690), .B(n11689), .Z(n11691) );
  AND U12291 ( .A(n11692), .B(n11691), .Z(n11776) );
  AND U12292 ( .A(y[154]), .B(x[108]), .Z(n11834) );
  AND U12293 ( .A(x[97]), .B(y[117]), .Z(n11694) );
  AND U12294 ( .A(x[98]), .B(y[116]), .Z(n11693) );
  XOR U12295 ( .A(n11694), .B(n11693), .Z(n11833) );
  XOR U12296 ( .A(n11834), .B(n11833), .Z(n11779) );
  AND U12297 ( .A(y[38]), .B(x[80]), .Z(n11783) );
  AND U12298 ( .A(y[158]), .B(x[104]), .Z(n11696) );
  AND U12299 ( .A(x[105]), .B(y[157]), .Z(n11695) );
  XOR U12300 ( .A(n11696), .B(n11695), .Z(n11782) );
  XNOR U12301 ( .A(n11783), .B(n11782), .Z(n11778) );
  XNOR U12302 ( .A(n11776), .B(n11777), .Z(n11752) );
  NAND U12303 ( .A(n11698), .B(n11697), .Z(n11702) );
  NAND U12304 ( .A(n11700), .B(n11699), .Z(n11701) );
  AND U12305 ( .A(n11702), .B(n11701), .Z(n11750) );
  XOR U12306 ( .A(n11751), .B(n11750), .Z(n12013) );
  XOR U12307 ( .A(n12014), .B(n12013), .Z(n12012) );
  NAND U12308 ( .A(n11703), .B(n11835), .Z(n11707) );
  NAND U12309 ( .A(n11705), .B(n11704), .Z(n11706) );
  NAND U12310 ( .A(n11707), .B(n11706), .Z(n11744) );
  NAND U12311 ( .A(n11709), .B(n11708), .Z(n11713) );
  NAND U12312 ( .A(n11711), .B(n11710), .Z(n11712) );
  AND U12313 ( .A(n11713), .B(n11712), .Z(n11947) );
  AND U12314 ( .A(y[37]), .B(x[81]), .Z(n11956) );
  AND U12315 ( .A(y[72]), .B(x[94]), .Z(n11955) );
  XOR U12316 ( .A(n11956), .B(n11955), .Z(n11954) );
  AND U12317 ( .A(y[78]), .B(x[88]), .Z(n11953) );
  XOR U12318 ( .A(n11954), .B(n11953), .Z(n11950) );
  NAND U12319 ( .A(x[117]), .B(y[193]), .Z(n11714) );
  XNOR U12320 ( .A(n11715), .B(n11714), .Z(n11881) );
  AND U12321 ( .A(y[192]), .B(x[118]), .Z(n11880) );
  XOR U12322 ( .A(n11881), .B(n11880), .Z(n11878) );
  XNOR U12323 ( .A(n11879), .B(n11878), .Z(n11949) );
  XNOR U12324 ( .A(n11947), .B(n11948), .Z(n11747) );
  NANDN U12325 ( .A(n11716), .B(n11960), .Z(n11720) );
  NAND U12326 ( .A(n11718), .B(n11717), .Z(n11719) );
  NAND U12327 ( .A(n11720), .B(n11719), .Z(n11746) );
  XOR U12328 ( .A(n11744), .B(n11745), .Z(n12011) );
  XOR U12329 ( .A(n12012), .B(n12011), .Z(n12008) );
  XNOR U12330 ( .A(n12007), .B(n12008), .Z(n12006) );
  XNOR U12331 ( .A(n12005), .B(n12006), .Z(n12028) );
  XNOR U12332 ( .A(n12029), .B(n12028), .Z(n12021) );
  NANDN U12333 ( .A(n11722), .B(n11721), .Z(n11726) );
  NANDN U12334 ( .A(n11724), .B(n11723), .Z(n11725) );
  NAND U12335 ( .A(n11726), .B(n11725), .Z(n12020) );
  NANDN U12336 ( .A(n11728), .B(n11727), .Z(n11732) );
  NANDN U12337 ( .A(n11730), .B(n11729), .Z(n11731) );
  AND U12338 ( .A(n11732), .B(n11731), .Z(n12019) );
  XOR U12339 ( .A(n12020), .B(n12019), .Z(n11733) );
  XNOR U12340 ( .A(n12021), .B(n11733), .Z(n12023) );
  XNOR U12341 ( .A(n12022), .B(n12023), .Z(n12025) );
  NANDN U12342 ( .A(n11735), .B(n11734), .Z(n11739) );
  NAND U12343 ( .A(n11737), .B(n11736), .Z(n11738) );
  NAND U12344 ( .A(n11739), .B(n11738), .Z(n12024) );
  XOR U12345 ( .A(n12025), .B(n12024), .Z(o[118]) );
  NANDN U12346 ( .A(n11745), .B(n11744), .Z(n11749) );
  NANDN U12347 ( .A(n11747), .B(n11746), .Z(n11748) );
  AND U12348 ( .A(n11749), .B(n11748), .Z(n12004) );
  NAND U12349 ( .A(n11751), .B(n11750), .Z(n11755) );
  NANDN U12350 ( .A(n11753), .B(n11752), .Z(n11754) );
  AND U12351 ( .A(n11755), .B(n11754), .Z(n11763) );
  NAND U12352 ( .A(n11757), .B(n11756), .Z(n11761) );
  NAND U12353 ( .A(n11759), .B(n11758), .Z(n11760) );
  NAND U12354 ( .A(n11761), .B(n11760), .Z(n11762) );
  XNOR U12355 ( .A(n11763), .B(n11762), .Z(n12002) );
  NAND U12356 ( .A(n11765), .B(n11764), .Z(n11769) );
  AND U12357 ( .A(n11767), .B(n11766), .Z(n11768) );
  ANDN U12358 ( .B(n11769), .A(n11768), .Z(n12000) );
  NAND U12359 ( .A(n11771), .B(n11770), .Z(n11775) );
  NANDN U12360 ( .A(n11773), .B(n11772), .Z(n11774) );
  AND U12361 ( .A(n11775), .B(n11774), .Z(n11871) );
  NANDN U12362 ( .A(n11777), .B(n11776), .Z(n11781) );
  NANDN U12363 ( .A(n11779), .B(n11778), .Z(n11780) );
  AND U12364 ( .A(n11781), .B(n11780), .Z(n11853) );
  NAND U12365 ( .A(n11783), .B(n11782), .Z(n11786) );
  AND U12366 ( .A(y[158]), .B(x[105]), .Z(n11934) );
  NAND U12367 ( .A(n11784), .B(n11934), .Z(n11785) );
  AND U12368 ( .A(n11786), .B(n11785), .Z(n11794) );
  NAND U12369 ( .A(n11788), .B(n11787), .Z(n11792) );
  NAND U12370 ( .A(n11790), .B(n11789), .Z(n11791) );
  NAND U12371 ( .A(n11792), .B(n11791), .Z(n11793) );
  XNOR U12372 ( .A(n11794), .B(n11793), .Z(n11851) );
  AND U12373 ( .A(x[96]), .B(y[119]), .Z(n11796) );
  NAND U12374 ( .A(x[107]), .B(y[156]), .Z(n11795) );
  XNOR U12375 ( .A(n11796), .B(n11795), .Z(n11818) );
  AND U12376 ( .A(y[193]), .B(x[116]), .Z(n11797) );
  AND U12377 ( .A(y[194]), .B(x[117]), .Z(n11901) );
  AND U12378 ( .A(n11797), .B(n11901), .Z(n11813) );
  NAND U12379 ( .A(n11799), .B(n11798), .Z(n11803) );
  NAND U12380 ( .A(n11801), .B(n11800), .Z(n11802) );
  AND U12381 ( .A(n11803), .B(n11802), .Z(n11811) );
  AND U12382 ( .A(x[111]), .B(y[152]), .Z(n11805) );
  NAND U12383 ( .A(x[87]), .B(y[32]), .Z(n11804) );
  XNOR U12384 ( .A(n11805), .B(n11804), .Z(n11809) );
  AND U12385 ( .A(x[119]), .B(y[192]), .Z(n11807) );
  NAND U12386 ( .A(x[108]), .B(y[155]), .Z(n11806) );
  XNOR U12387 ( .A(n11807), .B(n11806), .Z(n11808) );
  XNOR U12388 ( .A(n11809), .B(n11808), .Z(n11810) );
  XNOR U12389 ( .A(n11811), .B(n11810), .Z(n11812) );
  XOR U12390 ( .A(n11813), .B(n11812), .Z(n11816) );
  AND U12391 ( .A(y[34]), .B(x[85]), .Z(n11840) );
  XNOR U12392 ( .A(n11840), .B(n11814), .Z(n11815) );
  XNOR U12393 ( .A(n11816), .B(n11815), .Z(n11817) );
  XOR U12394 ( .A(n11818), .B(n11817), .Z(n11849) );
  NAND U12395 ( .A(n11820), .B(n11819), .Z(n11824) );
  NAND U12396 ( .A(n11822), .B(n11821), .Z(n11823) );
  AND U12397 ( .A(n11824), .B(n11823), .Z(n11832) );
  NAND U12398 ( .A(n11826), .B(n11825), .Z(n11830) );
  NAND U12399 ( .A(n11828), .B(n11827), .Z(n11829) );
  NAND U12400 ( .A(n11830), .B(n11829), .Z(n11831) );
  XNOR U12401 ( .A(n11832), .B(n11831), .Z(n11847) );
  NAND U12402 ( .A(n11834), .B(n11833), .Z(n11837) );
  AND U12403 ( .A(y[117]), .B(x[98]), .Z(n11935) );
  NAND U12404 ( .A(n11835), .B(n11935), .Z(n11836) );
  AND U12405 ( .A(n11837), .B(n11836), .Z(n11845) );
  NAND U12406 ( .A(n11839), .B(n11838), .Z(n11843) );
  NAND U12407 ( .A(n11841), .B(n11840), .Z(n11842) );
  NAND U12408 ( .A(n11843), .B(n11842), .Z(n11844) );
  XNOR U12409 ( .A(n11845), .B(n11844), .Z(n11846) );
  XNOR U12410 ( .A(n11847), .B(n11846), .Z(n11848) );
  XNOR U12411 ( .A(n11849), .B(n11848), .Z(n11850) );
  XNOR U12412 ( .A(n11851), .B(n11850), .Z(n11852) );
  XNOR U12413 ( .A(n11853), .B(n11852), .Z(n11869) );
  NAND U12414 ( .A(n11855), .B(n11854), .Z(n11859) );
  NAND U12415 ( .A(n11857), .B(n11856), .Z(n11858) );
  AND U12416 ( .A(n11859), .B(n11858), .Z(n11867) );
  NAND U12417 ( .A(n11861), .B(n11860), .Z(n11865) );
  NANDN U12418 ( .A(n11863), .B(n11862), .Z(n11864) );
  NAND U12419 ( .A(n11865), .B(n11864), .Z(n11866) );
  XNOR U12420 ( .A(n11867), .B(n11866), .Z(n11868) );
  XNOR U12421 ( .A(n11869), .B(n11868), .Z(n11870) );
  XNOR U12422 ( .A(n11871), .B(n11870), .Z(n11998) );
  NAND U12423 ( .A(n11873), .B(n11872), .Z(n11877) );
  NAND U12424 ( .A(n11875), .B(n11874), .Z(n11876) );
  AND U12425 ( .A(n11877), .B(n11876), .Z(n11996) );
  NAND U12426 ( .A(n11879), .B(n11878), .Z(n11883) );
  NAND U12427 ( .A(n11881), .B(n11880), .Z(n11882) );
  AND U12428 ( .A(n11883), .B(n11882), .Z(n11946) );
  AND U12429 ( .A(x[88]), .B(y[79]), .Z(n11885) );
  NAND U12430 ( .A(x[94]), .B(y[73]), .Z(n11884) );
  XNOR U12431 ( .A(n11885), .B(n11884), .Z(n11889) );
  AND U12432 ( .A(x[80]), .B(y[39]), .Z(n11887) );
  NAND U12433 ( .A(x[83]), .B(y[36]), .Z(n11886) );
  XNOR U12434 ( .A(n11887), .B(n11886), .Z(n11888) );
  XOR U12435 ( .A(n11889), .B(n11888), .Z(n11897) );
  AND U12436 ( .A(x[115]), .B(y[196]), .Z(n11891) );
  NAND U12437 ( .A(x[100]), .B(y[115]), .Z(n11890) );
  XNOR U12438 ( .A(n11891), .B(n11890), .Z(n11895) );
  AND U12439 ( .A(x[114]), .B(y[197]), .Z(n11893) );
  NAND U12440 ( .A(x[84]), .B(y[35]), .Z(n11892) );
  XNOR U12441 ( .A(n11893), .B(n11892), .Z(n11894) );
  XNOR U12442 ( .A(n11895), .B(n11894), .Z(n11896) );
  XNOR U12443 ( .A(n11897), .B(n11896), .Z(n11944) );
  AND U12444 ( .A(x[106]), .B(y[157]), .Z(n11903) );
  AND U12445 ( .A(x[104]), .B(y[159]), .Z(n11899) );
  NAND U12446 ( .A(x[89]), .B(y[78]), .Z(n11898) );
  XNOR U12447 ( .A(n11899), .B(n11898), .Z(n11900) );
  XNOR U12448 ( .A(n11901), .B(n11900), .Z(n11902) );
  XNOR U12449 ( .A(n11903), .B(n11902), .Z(n11919) );
  AND U12450 ( .A(x[97]), .B(y[118]), .Z(n11905) );
  NAND U12451 ( .A(x[99]), .B(y[116]), .Z(n11904) );
  XNOR U12452 ( .A(n11905), .B(n11904), .Z(n11909) );
  AND U12453 ( .A(x[81]), .B(y[38]), .Z(n11907) );
  NAND U12454 ( .A(x[101]), .B(y[114]), .Z(n11906) );
  XNOR U12455 ( .A(n11907), .B(n11906), .Z(n11908) );
  XOR U12456 ( .A(n11909), .B(n11908), .Z(n11917) );
  AND U12457 ( .A(x[90]), .B(y[77]), .Z(n11911) );
  NAND U12458 ( .A(x[109]), .B(y[154]), .Z(n11910) );
  XNOR U12459 ( .A(n11911), .B(n11910), .Z(n11915) );
  AND U12460 ( .A(x[93]), .B(y[74]), .Z(n11913) );
  NAND U12461 ( .A(x[95]), .B(y[72]), .Z(n11912) );
  XNOR U12462 ( .A(n11913), .B(n11912), .Z(n11914) );
  XNOR U12463 ( .A(n11915), .B(n11914), .Z(n11916) );
  XNOR U12464 ( .A(n11917), .B(n11916), .Z(n11918) );
  XOR U12465 ( .A(n11919), .B(n11918), .Z(n11942) );
  AND U12466 ( .A(x[113]), .B(y[198]), .Z(n11921) );
  NAND U12467 ( .A(x[86]), .B(y[33]), .Z(n11920) );
  XNOR U12468 ( .A(n11921), .B(n11920), .Z(n11925) );
  AND U12469 ( .A(x[118]), .B(y[193]), .Z(n11923) );
  NAND U12470 ( .A(x[102]), .B(y[113]), .Z(n11922) );
  XNOR U12471 ( .A(n11923), .B(n11922), .Z(n11924) );
  XOR U12472 ( .A(n11925), .B(n11924), .Z(n11933) );
  AND U12473 ( .A(x[112]), .B(y[199]), .Z(n11927) );
  NAND U12474 ( .A(x[103]), .B(y[112]), .Z(n11926) );
  XNOR U12475 ( .A(n11927), .B(n11926), .Z(n11931) );
  AND U12476 ( .A(x[82]), .B(y[37]), .Z(n11929) );
  NAND U12477 ( .A(x[110]), .B(y[153]), .Z(n11928) );
  XNOR U12478 ( .A(n11929), .B(n11928), .Z(n11930) );
  XNOR U12479 ( .A(n11931), .B(n11930), .Z(n11932) );
  XNOR U12480 ( .A(n11933), .B(n11932), .Z(n11940) );
  XOR U12481 ( .A(n11935), .B(n11934), .Z(n11938) );
  AND U12482 ( .A(y[75]), .B(x[92]), .Z(n11969) );
  XNOR U12483 ( .A(n11936), .B(n11969), .Z(n11937) );
  XNOR U12484 ( .A(n11938), .B(n11937), .Z(n11939) );
  XNOR U12485 ( .A(n11940), .B(n11939), .Z(n11941) );
  XNOR U12486 ( .A(n11942), .B(n11941), .Z(n11943) );
  XNOR U12487 ( .A(n11944), .B(n11943), .Z(n11945) );
  XNOR U12488 ( .A(n11946), .B(n11945), .Z(n11994) );
  NANDN U12489 ( .A(n11948), .B(n11947), .Z(n11952) );
  NANDN U12490 ( .A(n11950), .B(n11949), .Z(n11951) );
  AND U12491 ( .A(n11952), .B(n11951), .Z(n11984) );
  NAND U12492 ( .A(n11954), .B(n11953), .Z(n11958) );
  NAND U12493 ( .A(n11956), .B(n11955), .Z(n11957) );
  AND U12494 ( .A(n11958), .B(n11957), .Z(n11966) );
  NAND U12495 ( .A(n11960), .B(n11959), .Z(n11964) );
  NAND U12496 ( .A(n11962), .B(n11961), .Z(n11963) );
  NAND U12497 ( .A(n11964), .B(n11963), .Z(n11965) );
  XNOR U12498 ( .A(n11966), .B(n11965), .Z(n11982) );
  NAND U12499 ( .A(n11968), .B(n11967), .Z(n11972) );
  NAND U12500 ( .A(n11970), .B(n11969), .Z(n11971) );
  AND U12501 ( .A(n11972), .B(n11971), .Z(n11980) );
  NAND U12502 ( .A(n11974), .B(n11973), .Z(n11978) );
  NAND U12503 ( .A(n11976), .B(n11975), .Z(n11977) );
  NAND U12504 ( .A(n11978), .B(n11977), .Z(n11979) );
  XNOR U12505 ( .A(n11980), .B(n11979), .Z(n11981) );
  XNOR U12506 ( .A(n11982), .B(n11981), .Z(n11983) );
  XNOR U12507 ( .A(n11984), .B(n11983), .Z(n11992) );
  NANDN U12508 ( .A(n11986), .B(n11985), .Z(n11990) );
  NANDN U12509 ( .A(n11988), .B(n11987), .Z(n11989) );
  NAND U12510 ( .A(n11990), .B(n11989), .Z(n11991) );
  XNOR U12511 ( .A(n11992), .B(n11991), .Z(n11993) );
  XNOR U12512 ( .A(n11994), .B(n11993), .Z(n11995) );
  XNOR U12513 ( .A(n11996), .B(n11995), .Z(n11997) );
  XNOR U12514 ( .A(n11998), .B(n11997), .Z(n11999) );
  XNOR U12515 ( .A(n12000), .B(n11999), .Z(n12001) );
  XNOR U12516 ( .A(n12002), .B(n12001), .Z(n12003) );
  NANDN U12517 ( .A(n12006), .B(n12005), .Z(n12010) );
  NAND U12518 ( .A(n12008), .B(n12007), .Z(n12009) );
  AND U12519 ( .A(n12010), .B(n12009), .Z(n12018) );
  NAND U12520 ( .A(n12012), .B(n12011), .Z(n12016) );
  NAND U12521 ( .A(n12014), .B(n12013), .Z(n12015) );
  NAND U12522 ( .A(n12016), .B(n12015), .Z(n12017) );
  NAND U12523 ( .A(y[160]), .B(x[152]), .Z(n12144) );
  NAND U12524 ( .A(y[40]), .B(x[128]), .Z(n12032) );
  XOR U12525 ( .A(n12144), .B(n12032), .Z(n12033) );
  AND U12526 ( .A(y[0]), .B(x[120]), .Z(n12040) );
  AND U12527 ( .A(y[80]), .B(x[136]), .Z(n12037) );
  XOR U12528 ( .A(n12040), .B(n12037), .Z(n12036) );
  AND U12529 ( .A(y[120]), .B(x[144]), .Z(n12035) );
  XNOR U12530 ( .A(n12036), .B(n12035), .Z(n12034) );
  XNOR U12531 ( .A(n12033), .B(n12034), .Z(o[120]) );
  AND U12532 ( .A(x[120]), .B(y[1]), .Z(n12031) );
  NAND U12533 ( .A(x[121]), .B(y[0]), .Z(n12030) );
  XNOR U12534 ( .A(n12031), .B(n12030), .Z(n12042) );
  AND U12535 ( .A(y[40]), .B(x[129]), .Z(n12041) );
  XOR U12536 ( .A(n12042), .B(n12041), .Z(n12059) );
  AND U12537 ( .A(y[160]), .B(x[153]), .Z(n12268) );
  NAND U12538 ( .A(y[81]), .B(x[136]), .Z(n12045) );
  XNOR U12539 ( .A(n12268), .B(n12045), .Z(n12047) );
  AND U12540 ( .A(y[161]), .B(x[152]), .Z(n12069) );
  NAND U12541 ( .A(y[80]), .B(x[137]), .Z(n12068) );
  XNOR U12542 ( .A(n12069), .B(n12068), .Z(n12046) );
  XOR U12543 ( .A(n12047), .B(n12046), .Z(n12057) );
  AND U12544 ( .A(y[41]), .B(x[128]), .Z(n12295) );
  AND U12545 ( .A(y[121]), .B(x[144]), .Z(n12062) );
  XOR U12546 ( .A(n12295), .B(n12062), .Z(n12064) );
  AND U12547 ( .A(y[120]), .B(x[145]), .Z(n12063) );
  XNOR U12548 ( .A(n12064), .B(n12063), .Z(n12056) );
  XNOR U12549 ( .A(n12057), .B(n12056), .Z(n12058) );
  XNOR U12550 ( .A(n12059), .B(n12058), .Z(n12053) );
  NAND U12551 ( .A(n12036), .B(n12035), .Z(n12039) );
  AND U12552 ( .A(n12040), .B(n12037), .Z(n12038) );
  ANDN U12553 ( .B(n12039), .A(n12038), .Z(n12050) );
  XNOR U12554 ( .A(n12051), .B(n12050), .Z(n12052) );
  XNOR U12555 ( .A(n12053), .B(n12052), .Z(o[121]) );
  NAND U12556 ( .A(y[1]), .B(x[121]), .Z(n12091) );
  NANDN U12557 ( .A(n12091), .B(n12040), .Z(n12044) );
  NAND U12558 ( .A(n12042), .B(n12041), .Z(n12043) );
  AND U12559 ( .A(n12044), .B(n12043), .Z(n12112) );
  NANDN U12560 ( .A(n12045), .B(n12268), .Z(n12049) );
  NAND U12561 ( .A(n12047), .B(n12046), .Z(n12048) );
  AND U12562 ( .A(n12049), .B(n12048), .Z(n12111) );
  AND U12563 ( .A(y[122]), .B(x[144]), .Z(n12116) );
  NAND U12564 ( .A(y[2]), .B(x[120]), .Z(n12117) );
  XNOR U12565 ( .A(n12116), .B(n12117), .Z(n12118) );
  NAND U12566 ( .A(y[40]), .B(x[130]), .Z(n12119) );
  XNOR U12567 ( .A(n12118), .B(n12119), .Z(n12110) );
  XOR U12568 ( .A(n12111), .B(n12110), .Z(n12113) );
  XOR U12569 ( .A(n12112), .B(n12113), .Z(n12071) );
  NANDN U12570 ( .A(n12051), .B(n12050), .Z(n12055) );
  NAND U12571 ( .A(n12053), .B(n12052), .Z(n12054) );
  NAND U12572 ( .A(n12055), .B(n12054), .Z(n12070) );
  XNOR U12573 ( .A(n12071), .B(n12070), .Z(n12073) );
  NANDN U12574 ( .A(n12057), .B(n12056), .Z(n12061) );
  NANDN U12575 ( .A(n12059), .B(n12058), .Z(n12060) );
  AND U12576 ( .A(n12061), .B(n12060), .Z(n12079) );
  AND U12577 ( .A(y[0]), .B(x[122]), .Z(n12088) );
  NAND U12578 ( .A(y[82]), .B(x[136]), .Z(n12089) );
  XNOR U12579 ( .A(n12088), .B(n12089), .Z(n12090) );
  NAND U12580 ( .A(y[120]), .B(x[146]), .Z(n12125) );
  XNOR U12581 ( .A(n12124), .B(n12125), .Z(n12126) );
  AND U12582 ( .A(y[80]), .B(x[138]), .Z(n12174) );
  AND U12583 ( .A(y[162]), .B(x[152]), .Z(n12101) );
  XOR U12584 ( .A(n12174), .B(n12101), .Z(n12103) );
  NAND U12585 ( .A(y[81]), .B(x[137]), .Z(n12102) );
  XOR U12586 ( .A(n12103), .B(n12102), .Z(n12127) );
  XNOR U12587 ( .A(n12126), .B(n12127), .Z(n12076) );
  NAND U12588 ( .A(n12295), .B(n12062), .Z(n12066) );
  AND U12589 ( .A(n12064), .B(n12063), .Z(n12065) );
  ANDN U12590 ( .B(n12066), .A(n12065), .Z(n12085) );
  AND U12591 ( .A(x[153]), .B(y[161]), .Z(n12149) );
  NAND U12592 ( .A(x[154]), .B(y[160]), .Z(n12067) );
  XNOR U12593 ( .A(n12149), .B(n12067), .Z(n12123) );
  ANDN U12594 ( .B(n12069), .A(n12068), .Z(n12122) );
  XOR U12595 ( .A(n12123), .B(n12122), .Z(n12082) );
  AND U12596 ( .A(y[121]), .B(x[145]), .Z(n12094) );
  NAND U12597 ( .A(y[41]), .B(x[129]), .Z(n12095) );
  XNOR U12598 ( .A(n12094), .B(n12095), .Z(n12096) );
  NAND U12599 ( .A(y[42]), .B(x[128]), .Z(n12097) );
  XOR U12600 ( .A(n12096), .B(n12097), .Z(n12083) );
  XNOR U12601 ( .A(n12082), .B(n12083), .Z(n12084) );
  XOR U12602 ( .A(n12085), .B(n12084), .Z(n12077) );
  XNOR U12603 ( .A(n12076), .B(n12077), .Z(n12078) );
  XNOR U12604 ( .A(n12079), .B(n12078), .Z(n12072) );
  XNOR U12605 ( .A(n12073), .B(n12072), .Z(o[122]) );
  NANDN U12606 ( .A(n12071), .B(n12070), .Z(n12075) );
  NAND U12607 ( .A(n12073), .B(n12072), .Z(n12074) );
  AND U12608 ( .A(n12075), .B(n12074), .Z(n12216) );
  NANDN U12609 ( .A(n12077), .B(n12076), .Z(n12081) );
  NAND U12610 ( .A(n12079), .B(n12078), .Z(n12080) );
  AND U12611 ( .A(n12081), .B(n12080), .Z(n12201) );
  NANDN U12612 ( .A(n12083), .B(n12082), .Z(n12087) );
  NANDN U12613 ( .A(n12085), .B(n12084), .Z(n12086) );
  AND U12614 ( .A(n12087), .B(n12086), .Z(n12199) );
  NANDN U12615 ( .A(n12089), .B(n12088), .Z(n12093) );
  NANDN U12616 ( .A(n12091), .B(n12090), .Z(n12092) );
  AND U12617 ( .A(n12093), .B(n12092), .Z(n12211) );
  NANDN U12618 ( .A(n12095), .B(n12094), .Z(n12099) );
  NANDN U12619 ( .A(n12097), .B(n12096), .Z(n12098) );
  AND U12620 ( .A(n12099), .B(n12098), .Z(n12165) );
  AND U12621 ( .A(y[123]), .B(x[144]), .Z(n12194) );
  AND U12622 ( .A(y[83]), .B(x[136]), .Z(n12193) );
  NAND U12623 ( .A(y[0]), .B(x[123]), .Z(n12192) );
  XOR U12624 ( .A(n12193), .B(n12192), .Z(n12195) );
  XOR U12625 ( .A(n12194), .B(n12195), .Z(n12163) );
  AND U12626 ( .A(y[81]), .B(x[138]), .Z(n12248) );
  NAND U12627 ( .A(x[139]), .B(y[80]), .Z(n12100) );
  XNOR U12628 ( .A(n12248), .B(n12100), .Z(n12176) );
  NAND U12629 ( .A(y[82]), .B(x[137]), .Z(n12177) );
  XNOR U12630 ( .A(n12176), .B(n12177), .Z(n12162) );
  XNOR U12631 ( .A(n12163), .B(n12162), .Z(n12164) );
  XNOR U12632 ( .A(n12165), .B(n12164), .Z(n12210) );
  XNOR U12633 ( .A(n12211), .B(n12210), .Z(n12212) );
  NAND U12634 ( .A(n12174), .B(n12101), .Z(n12105) );
  ANDN U12635 ( .B(n12103), .A(n12102), .Z(n12104) );
  ANDN U12636 ( .B(n12105), .A(n12104), .Z(n12171) );
  AND U12637 ( .A(y[2]), .B(x[121]), .Z(n12140) );
  AND U12638 ( .A(y[1]), .B(x[122]), .Z(n12139) );
  NAND U12639 ( .A(y[122]), .B(x[145]), .Z(n12138) );
  XOR U12640 ( .A(n12139), .B(n12138), .Z(n12141) );
  XOR U12641 ( .A(n12140), .B(n12141), .Z(n12169) );
  AND U12642 ( .A(x[155]), .B(y[160]), .Z(n12107) );
  NAND U12643 ( .A(x[152]), .B(y[163]), .Z(n12106) );
  XNOR U12644 ( .A(n12107), .B(n12106), .Z(n12145) );
  AND U12645 ( .A(x[153]), .B(y[162]), .Z(n12109) );
  NAND U12646 ( .A(x[154]), .B(y[161]), .Z(n12108) );
  XOR U12647 ( .A(n12109), .B(n12108), .Z(n12146) );
  XNOR U12648 ( .A(n12145), .B(n12146), .Z(n12168) );
  XNOR U12649 ( .A(n12169), .B(n12168), .Z(n12170) );
  XOR U12650 ( .A(n12171), .B(n12170), .Z(n12213) );
  XNOR U12651 ( .A(n12212), .B(n12213), .Z(n12198) );
  XNOR U12652 ( .A(n12199), .B(n12198), .Z(n12200) );
  XOR U12653 ( .A(n12201), .B(n12200), .Z(n12217) );
  XNOR U12654 ( .A(n12216), .B(n12217), .Z(n12219) );
  NANDN U12655 ( .A(n12111), .B(n12110), .Z(n12115) );
  OR U12656 ( .A(n12113), .B(n12112), .Z(n12114) );
  AND U12657 ( .A(n12115), .B(n12114), .Z(n12207) );
  NANDN U12658 ( .A(n12117), .B(n12116), .Z(n12121) );
  NANDN U12659 ( .A(n12119), .B(n12118), .Z(n12120) );
  AND U12660 ( .A(n12121), .B(n12120), .Z(n12131) );
  AND U12661 ( .A(y[161]), .B(x[154]), .Z(n12265) );
  XNOR U12662 ( .A(n12131), .B(n12130), .Z(n12133) );
  NAND U12663 ( .A(y[40]), .B(x[131]), .Z(n12185) );
  NAND U12664 ( .A(y[3]), .B(x[120]), .Z(n12183) );
  NAND U12665 ( .A(y[121]), .B(x[146]), .Z(n12182) );
  XOR U12666 ( .A(n12183), .B(n12182), .Z(n12184) );
  XNOR U12667 ( .A(n12185), .B(n12184), .Z(n12159) );
  NAND U12668 ( .A(y[43]), .B(x[128]), .Z(n12153) );
  NAND U12669 ( .A(y[41]), .B(x[130]), .Z(n12151) );
  NAND U12670 ( .A(y[120]), .B(x[147]), .Z(n12150) );
  XOR U12671 ( .A(n12151), .B(n12150), .Z(n12152) );
  XNOR U12672 ( .A(n12153), .B(n12152), .Z(n12157) );
  AND U12673 ( .A(y[42]), .B(x[129]), .Z(n12156) );
  XOR U12674 ( .A(n12157), .B(n12156), .Z(n12158) );
  XOR U12675 ( .A(n12159), .B(n12158), .Z(n12132) );
  XOR U12676 ( .A(n12133), .B(n12132), .Z(n12205) );
  NANDN U12677 ( .A(n12125), .B(n12124), .Z(n12129) );
  NANDN U12678 ( .A(n12127), .B(n12126), .Z(n12128) );
  AND U12679 ( .A(n12129), .B(n12128), .Z(n12204) );
  XNOR U12680 ( .A(n12205), .B(n12204), .Z(n12206) );
  XNOR U12681 ( .A(n12207), .B(n12206), .Z(n12218) );
  XOR U12682 ( .A(n12219), .B(n12218), .Z(o[123]) );
  NANDN U12683 ( .A(n12131), .B(n12130), .Z(n12135) );
  NAND U12684 ( .A(n12133), .B(n12132), .Z(n12134) );
  AND U12685 ( .A(n12135), .B(n12134), .Z(n12233) );
  AND U12686 ( .A(x[131]), .B(y[41]), .Z(n12137) );
  NAND U12687 ( .A(x[128]), .B(y[44]), .Z(n12136) );
  XNOR U12688 ( .A(n12137), .B(n12136), .Z(n12296) );
  NAND U12689 ( .A(y[42]), .B(x[130]), .Z(n12367) );
  NAND U12690 ( .A(y[43]), .B(x[129]), .Z(n12300) );
  AND U12691 ( .A(y[120]), .B(x[148]), .Z(n12254) );
  AND U12692 ( .A(y[3]), .B(x[121]), .Z(n12253) );
  XOR U12693 ( .A(n12254), .B(n12253), .Z(n12256) );
  AND U12694 ( .A(y[4]), .B(x[120]), .Z(n12255) );
  XOR U12695 ( .A(n12256), .B(n12255), .Z(n12301) );
  XOR U12696 ( .A(n12302), .B(n12301), .Z(n12314) );
  NANDN U12697 ( .A(n12139), .B(n12138), .Z(n12143) );
  OR U12698 ( .A(n12141), .B(n12140), .Z(n12142) );
  AND U12699 ( .A(n12143), .B(n12142), .Z(n12312) );
  AND U12700 ( .A(y[163]), .B(x[155]), .Z(n12539) );
  NANDN U12701 ( .A(n12144), .B(n12539), .Z(n12148) );
  NANDN U12702 ( .A(n12146), .B(n12145), .Z(n12147) );
  AND U12703 ( .A(n12148), .B(n12147), .Z(n12311) );
  AND U12704 ( .A(y[0]), .B(x[124]), .Z(n12281) );
  AND U12705 ( .A(y[122]), .B(x[146]), .Z(n12279) );
  NAND U12706 ( .A(y[84]), .B(x[136]), .Z(n12278) );
  AND U12707 ( .A(y[162]), .B(x[154]), .Z(n12191) );
  AND U12708 ( .A(n12149), .B(n12191), .Z(n12275) );
  AND U12709 ( .A(y[80]), .B(x[140]), .Z(n12273) );
  IV U12710 ( .A(n12273), .Z(n12388) );
  NAND U12711 ( .A(y[164]), .B(x[152]), .Z(n12445) );
  XOR U12712 ( .A(n12275), .B(n12274), .Z(n12236) );
  XOR U12713 ( .A(n12237), .B(n12236), .Z(n12239) );
  NAND U12714 ( .A(n12151), .B(n12150), .Z(n12155) );
  NAND U12715 ( .A(n12153), .B(n12152), .Z(n12154) );
  AND U12716 ( .A(n12155), .B(n12154), .Z(n12238) );
  XOR U12717 ( .A(n12239), .B(n12238), .Z(n12326) );
  NAND U12718 ( .A(n12157), .B(n12156), .Z(n12161) );
  NAND U12719 ( .A(n12159), .B(n12158), .Z(n12160) );
  AND U12720 ( .A(n12161), .B(n12160), .Z(n12325) );
  XNOR U12721 ( .A(n12326), .B(n12325), .Z(n12327) );
  XNOR U12722 ( .A(n12328), .B(n12327), .Z(n12232) );
  XNOR U12723 ( .A(n12233), .B(n12232), .Z(n12235) );
  NANDN U12724 ( .A(n12163), .B(n12162), .Z(n12167) );
  NANDN U12725 ( .A(n12165), .B(n12164), .Z(n12166) );
  AND U12726 ( .A(n12167), .B(n12166), .Z(n12318) );
  NANDN U12727 ( .A(n12169), .B(n12168), .Z(n12173) );
  NANDN U12728 ( .A(n12171), .B(n12170), .Z(n12172) );
  NAND U12729 ( .A(n12173), .B(n12172), .Z(n12317) );
  XNOR U12730 ( .A(n12318), .B(n12317), .Z(n12320) );
  AND U12731 ( .A(y[81]), .B(x[139]), .Z(n12175) );
  NAND U12732 ( .A(n12175), .B(n12174), .Z(n12179) );
  NANDN U12733 ( .A(n12177), .B(n12176), .Z(n12178) );
  AND U12734 ( .A(n12179), .B(n12178), .Z(n12322) );
  AND U12735 ( .A(y[40]), .B(x[132]), .Z(n12259) );
  NAND U12736 ( .A(y[124]), .B(x[144]), .Z(n12260) );
  NAND U12737 ( .A(y[123]), .B(x[145]), .Z(n12262) );
  AND U12738 ( .A(x[138]), .B(y[82]), .Z(n12181) );
  NAND U12739 ( .A(x[139]), .B(y[81]), .Z(n12180) );
  XNOR U12740 ( .A(n12181), .B(n12180), .Z(n12250) );
  AND U12741 ( .A(y[83]), .B(x[137]), .Z(n12249) );
  XOR U12742 ( .A(n12250), .B(n12249), .Z(n12305) );
  XOR U12743 ( .A(n12306), .B(n12305), .Z(n12307) );
  NAND U12744 ( .A(n12183), .B(n12182), .Z(n12187) );
  NAND U12745 ( .A(n12185), .B(n12184), .Z(n12186) );
  NAND U12746 ( .A(n12187), .B(n12186), .Z(n12308) );
  XNOR U12747 ( .A(n12322), .B(n12321), .Z(n12324) );
  AND U12748 ( .A(y[2]), .B(x[122]), .Z(n12292) );
  AND U12749 ( .A(y[121]), .B(x[147]), .Z(n12290) );
  NAND U12750 ( .A(y[1]), .B(x[123]), .Z(n12289) );
  AND U12751 ( .A(x[156]), .B(y[160]), .Z(n12189) );
  NAND U12752 ( .A(x[153]), .B(y[163]), .Z(n12188) );
  XNOR U12753 ( .A(n12189), .B(n12188), .Z(n12269) );
  NAND U12754 ( .A(x[155]), .B(y[161]), .Z(n12190) );
  XOR U12755 ( .A(n12191), .B(n12190), .Z(n12270) );
  XOR U12756 ( .A(n12242), .B(n12243), .Z(n12244) );
  NANDN U12757 ( .A(n12193), .B(n12192), .Z(n12197) );
  OR U12758 ( .A(n12195), .B(n12194), .Z(n12196) );
  NAND U12759 ( .A(n12197), .B(n12196), .Z(n12245) );
  XOR U12760 ( .A(n12324), .B(n12323), .Z(n12319) );
  XOR U12761 ( .A(n12320), .B(n12319), .Z(n12234) );
  XOR U12762 ( .A(n12235), .B(n12234), .Z(n12225) );
  NANDN U12763 ( .A(n12199), .B(n12198), .Z(n12203) );
  NANDN U12764 ( .A(n12201), .B(n12200), .Z(n12202) );
  AND U12765 ( .A(n12203), .B(n12202), .Z(n12229) );
  NANDN U12766 ( .A(n12205), .B(n12204), .Z(n12209) );
  NAND U12767 ( .A(n12207), .B(n12206), .Z(n12208) );
  AND U12768 ( .A(n12209), .B(n12208), .Z(n12227) );
  NANDN U12769 ( .A(n12211), .B(n12210), .Z(n12215) );
  NANDN U12770 ( .A(n12213), .B(n12212), .Z(n12214) );
  AND U12771 ( .A(n12215), .B(n12214), .Z(n12226) );
  XNOR U12772 ( .A(n12227), .B(n12226), .Z(n12228) );
  XOR U12773 ( .A(n12229), .B(n12228), .Z(n12224) );
  NANDN U12774 ( .A(n12217), .B(n12216), .Z(n12221) );
  NAND U12775 ( .A(n12219), .B(n12218), .Z(n12220) );
  AND U12776 ( .A(n12221), .B(n12220), .Z(n12223) );
  XNOR U12777 ( .A(n12224), .B(n12223), .Z(n12222) );
  XNOR U12778 ( .A(n12225), .B(n12222), .Z(o[124]) );
  NANDN U12779 ( .A(n12227), .B(n12226), .Z(n12231) );
  NAND U12780 ( .A(n12229), .B(n12228), .Z(n12230) );
  AND U12781 ( .A(n12231), .B(n12230), .Z(n12474) );
  XNOR U12782 ( .A(n12475), .B(n12474), .Z(n12477) );
  NAND U12783 ( .A(n12237), .B(n12236), .Z(n12241) );
  NAND U12784 ( .A(n12239), .B(n12238), .Z(n12240) );
  AND U12785 ( .A(n12241), .B(n12240), .Z(n12332) );
  NAND U12786 ( .A(n12243), .B(n12242), .Z(n12247) );
  NANDN U12787 ( .A(n12245), .B(n12244), .Z(n12246) );
  NAND U12788 ( .A(n12247), .B(n12246), .Z(n12331) );
  AND U12789 ( .A(y[82]), .B(x[139]), .Z(n12390) );
  NAND U12790 ( .A(n12248), .B(n12390), .Z(n12252) );
  NAND U12791 ( .A(n12250), .B(n12249), .Z(n12251) );
  NAND U12792 ( .A(n12252), .B(n12251), .Z(n12398) );
  NAND U12793 ( .A(n12254), .B(n12253), .Z(n12258) );
  NAND U12794 ( .A(n12256), .B(n12255), .Z(n12257) );
  AND U12795 ( .A(n12258), .B(n12257), .Z(n12375) );
  AND U12796 ( .A(y[40]), .B(x[133]), .Z(n12378) );
  NAND U12797 ( .A(y[83]), .B(x[138]), .Z(n12379) );
  NAND U12798 ( .A(y[125]), .B(x[144]), .Z(n12566) );
  AND U12799 ( .A(y[121]), .B(x[148]), .Z(n12383) );
  NAND U12800 ( .A(y[0]), .B(x[125]), .Z(n12384) );
  NAND U12801 ( .A(y[1]), .B(x[124]), .Z(n12591) );
  XOR U12802 ( .A(n12373), .B(n12372), .Z(n12374) );
  XOR U12803 ( .A(n12398), .B(n12399), .Z(n12400) );
  NANDN U12804 ( .A(n12260), .B(n12259), .Z(n12264) );
  NANDN U12805 ( .A(n12262), .B(n12261), .Z(n12263) );
  AND U12806 ( .A(n12264), .B(n12263), .Z(n12425) );
  AND U12807 ( .A(y[162]), .B(x[155]), .Z(n12286) );
  AND U12808 ( .A(n12286), .B(n12265), .Z(n12447) );
  AND U12809 ( .A(x[152]), .B(y[165]), .Z(n12267) );
  AND U12810 ( .A(x[153]), .B(y[164]), .Z(n12266) );
  XOR U12811 ( .A(n12267), .B(n12266), .Z(n12446) );
  XOR U12812 ( .A(n12447), .B(n12446), .Z(n12423) );
  AND U12813 ( .A(y[45]), .B(x[128]), .Z(n12431) );
  AND U12814 ( .A(y[4]), .B(x[121]), .Z(n12430) );
  XOR U12815 ( .A(n12431), .B(n12430), .Z(n12433) );
  AND U12816 ( .A(y[41]), .B(x[132]), .Z(n12432) );
  XOR U12817 ( .A(n12433), .B(n12432), .Z(n12422) );
  XOR U12818 ( .A(n12423), .B(n12422), .Z(n12424) );
  XNOR U12819 ( .A(n12400), .B(n12401), .Z(n12333) );
  XOR U12820 ( .A(n12334), .B(n12333), .Z(n12467) );
  AND U12821 ( .A(y[163]), .B(x[156]), .Z(n12680) );
  NAND U12822 ( .A(n12680), .B(n12268), .Z(n12272) );
  NANDN U12823 ( .A(n12270), .B(n12269), .Z(n12271) );
  NAND U12824 ( .A(n12272), .B(n12271), .Z(n12343) );
  NANDN U12825 ( .A(n12273), .B(n12445), .Z(n12277) );
  NANDN U12826 ( .A(n12275), .B(n12274), .Z(n12276) );
  AND U12827 ( .A(n12277), .B(n12276), .Z(n12344) );
  XOR U12828 ( .A(n12343), .B(n12344), .Z(n12346) );
  NANDN U12829 ( .A(n12279), .B(n12278), .Z(n12283) );
  NANDN U12830 ( .A(n12281), .B(n12280), .Z(n12282) );
  AND U12831 ( .A(n12283), .B(n12282), .Z(n12352) );
  AND U12832 ( .A(x[130]), .B(y[43]), .Z(n12285) );
  NAND U12833 ( .A(x[131]), .B(y[42]), .Z(n12284) );
  XNOR U12834 ( .A(n12285), .B(n12284), .Z(n12369) );
  AND U12835 ( .A(y[44]), .B(x[129]), .Z(n12368) );
  XOR U12836 ( .A(n12369), .B(n12368), .Z(n12350) );
  AND U12837 ( .A(y[163]), .B(x[154]), .Z(n12356) );
  AND U12838 ( .A(y[160]), .B(x[157]), .Z(n12355) );
  XOR U12839 ( .A(n12356), .B(n12355), .Z(n12358) );
  AND U12840 ( .A(y[161]), .B(x[156]), .Z(n12537) );
  XOR U12841 ( .A(n12286), .B(n12537), .Z(n12357) );
  XOR U12842 ( .A(n12358), .B(n12357), .Z(n12349) );
  XOR U12843 ( .A(n12350), .B(n12349), .Z(n12351) );
  XOR U12844 ( .A(n12352), .B(n12351), .Z(n12345) );
  XOR U12845 ( .A(n12346), .B(n12345), .Z(n12413) );
  AND U12846 ( .A(y[81]), .B(x[140]), .Z(n12288) );
  AND U12847 ( .A(x[141]), .B(y[80]), .Z(n12287) );
  XOR U12848 ( .A(n12288), .B(n12287), .Z(n12389) );
  XOR U12849 ( .A(n12390), .B(n12389), .Z(n12417) );
  AND U12850 ( .A(y[120]), .B(x[149]), .Z(n12362) );
  AND U12851 ( .A(y[2]), .B(x[123]), .Z(n12361) );
  XOR U12852 ( .A(n12362), .B(n12361), .Z(n12364) );
  AND U12853 ( .A(y[3]), .B(x[122]), .Z(n12363) );
  XOR U12854 ( .A(n12364), .B(n12363), .Z(n12416) );
  XOR U12855 ( .A(n12417), .B(n12416), .Z(n12419) );
  NANDN U12856 ( .A(n12290), .B(n12289), .Z(n12294) );
  NANDN U12857 ( .A(n12292), .B(n12291), .Z(n12293) );
  AND U12858 ( .A(n12294), .B(n12293), .Z(n12418) );
  XOR U12859 ( .A(n12419), .B(n12418), .Z(n12411) );
  AND U12860 ( .A(y[44]), .B(x[131]), .Z(n12679) );
  NAND U12861 ( .A(n12679), .B(n12295), .Z(n12298) );
  NANDN U12862 ( .A(n12367), .B(n12296), .Z(n12297) );
  NAND U12863 ( .A(n12298), .B(n12297), .Z(n12339) );
  AND U12864 ( .A(y[122]), .B(x[147]), .Z(n12440) );
  NAND U12865 ( .A(y[84]), .B(x[137]), .Z(n12549) );
  NAND U12866 ( .A(y[85]), .B(x[136]), .Z(n12442) );
  AND U12867 ( .A(y[5]), .B(x[120]), .Z(n12450) );
  NAND U12868 ( .A(y[124]), .B(x[145]), .Z(n12451) );
  NAND U12869 ( .A(y[123]), .B(x[146]), .Z(n12453) );
  XOR U12870 ( .A(n12338), .B(n12337), .Z(n12340) );
  XNOR U12871 ( .A(n12339), .B(n12340), .Z(n12410) );
  NANDN U12872 ( .A(n12300), .B(n12299), .Z(n12304) );
  NAND U12873 ( .A(n12302), .B(n12301), .Z(n12303) );
  AND U12874 ( .A(n12304), .B(n12303), .Z(n12405) );
  NAND U12875 ( .A(n12306), .B(n12305), .Z(n12310) );
  NANDN U12876 ( .A(n12308), .B(n12307), .Z(n12309) );
  NAND U12877 ( .A(n12310), .B(n12309), .Z(n12404) );
  NANDN U12878 ( .A(n12312), .B(n12311), .Z(n12316) );
  NANDN U12879 ( .A(n12314), .B(n12313), .Z(n12315) );
  NAND U12880 ( .A(n12316), .B(n12315), .Z(n12407) );
  XOR U12881 ( .A(n12465), .B(n12464), .Z(n12466) );
  XOR U12882 ( .A(n12467), .B(n12466), .Z(n12468) );
  XNOR U12883 ( .A(n12469), .B(n12468), .Z(n12470) );
  NANDN U12884 ( .A(n12326), .B(n12325), .Z(n12330) );
  NAND U12885 ( .A(n12328), .B(n12327), .Z(n12329) );
  AND U12886 ( .A(n12330), .B(n12329), .Z(n12458) );
  XNOR U12887 ( .A(n12459), .B(n12458), .Z(n12460) );
  XOR U12888 ( .A(n12461), .B(n12460), .Z(n12471) );
  XNOR U12889 ( .A(n12470), .B(n12471), .Z(n12476) );
  XOR U12890 ( .A(n12477), .B(n12476), .Z(o[125]) );
  NANDN U12891 ( .A(n12332), .B(n12331), .Z(n12336) );
  NAND U12892 ( .A(n12334), .B(n12333), .Z(n12335) );
  AND U12893 ( .A(n12336), .B(n12335), .Z(n12762) );
  NAND U12894 ( .A(n12338), .B(n12337), .Z(n12342) );
  NAND U12895 ( .A(n12340), .B(n12339), .Z(n12341) );
  AND U12896 ( .A(n12342), .B(n12341), .Z(n12506) );
  NAND U12897 ( .A(n12344), .B(n12343), .Z(n12348) );
  NAND U12898 ( .A(n12346), .B(n12345), .Z(n12347) );
  NAND U12899 ( .A(n12348), .B(n12347), .Z(n12505) );
  NAND U12900 ( .A(n12350), .B(n12349), .Z(n12354) );
  NAND U12901 ( .A(n12352), .B(n12351), .Z(n12353) );
  AND U12902 ( .A(n12354), .B(n12353), .Z(n12507) );
  XOR U12903 ( .A(n12508), .B(n12507), .Z(n12764) );
  IV U12904 ( .A(n12764), .Z(n12397) );
  NAND U12905 ( .A(n12356), .B(n12355), .Z(n12360) );
  NAND U12906 ( .A(n12358), .B(n12357), .Z(n12359) );
  AND U12907 ( .A(n12360), .B(n12359), .Z(n12514) );
  NAND U12908 ( .A(n12362), .B(n12361), .Z(n12366) );
  NAND U12909 ( .A(n12364), .B(n12363), .Z(n12365) );
  AND U12910 ( .A(n12366), .B(n12365), .Z(n12516) );
  AND U12911 ( .A(x[131]), .B(y[43]), .Z(n12429) );
  NANDN U12912 ( .A(n12367), .B(n12429), .Z(n12371) );
  NAND U12913 ( .A(n12369), .B(n12368), .Z(n12370) );
  AND U12914 ( .A(n12371), .B(n12370), .Z(n12726) );
  AND U12915 ( .A(y[123]), .B(x[147]), .Z(n12528) );
  AND U12916 ( .A(y[83]), .B(x[139]), .Z(n12527) );
  XOR U12917 ( .A(n12528), .B(n12527), .Z(n12526) );
  AND U12918 ( .A(y[3]), .B(x[123]), .Z(n12525) );
  XOR U12919 ( .A(n12526), .B(n12525), .Z(n12728) );
  AND U12920 ( .A(y[124]), .B(x[146]), .Z(n12555) );
  AND U12921 ( .A(y[82]), .B(x[140]), .Z(n12554) );
  XOR U12922 ( .A(n12555), .B(n12554), .Z(n12553) );
  AND U12923 ( .A(y[4]), .B(x[122]), .Z(n12552) );
  XNOR U12924 ( .A(n12553), .B(n12552), .Z(n12727) );
  XNOR U12925 ( .A(n12726), .B(n12725), .Z(n12515) );
  NAND U12926 ( .A(n12373), .B(n12372), .Z(n12377) );
  NANDN U12927 ( .A(n12375), .B(n12374), .Z(n12376) );
  AND U12928 ( .A(n12377), .B(n12376), .Z(n12747) );
  NANDN U12929 ( .A(n12379), .B(n12378), .Z(n12382) );
  NANDN U12930 ( .A(n12566), .B(n12380), .Z(n12381) );
  AND U12931 ( .A(n12382), .B(n12381), .Z(n12702) );
  NANDN U12932 ( .A(n12384), .B(n12383), .Z(n12387) );
  NANDN U12933 ( .A(n12591), .B(n12385), .Z(n12386) );
  NAND U12934 ( .A(n12387), .B(n12386), .Z(n12701) );
  AND U12935 ( .A(y[81]), .B(x[141]), .Z(n12572) );
  NANDN U12936 ( .A(n12388), .B(n12572), .Z(n12392) );
  NAND U12937 ( .A(n12390), .B(n12389), .Z(n12391) );
  AND U12938 ( .A(n12392), .B(n12391), .Z(n12714) );
  AND U12939 ( .A(x[125]), .B(y[1]), .Z(n12394) );
  NAND U12940 ( .A(x[124]), .B(y[2]), .Z(n12393) );
  XNOR U12941 ( .A(n12394), .B(n12393), .Z(n12589) );
  NAND U12942 ( .A(y[120]), .B(x[150]), .Z(n12590) );
  IV U12943 ( .A(n12590), .Z(n12395) );
  XOR U12944 ( .A(n12589), .B(n12395), .Z(n12711) );
  AND U12945 ( .A(y[165]), .B(x[153]), .Z(n12615) );
  AND U12946 ( .A(y[161]), .B(x[155]), .Z(n12396) );
  AND U12947 ( .A(x[156]), .B(y[162]), .Z(n12457) );
  AND U12948 ( .A(n12396), .B(n12457), .Z(n12616) );
  NAND U12949 ( .A(y[164]), .B(x[154]), .Z(n12617) );
  XNOR U12950 ( .A(n12615), .B(n12614), .Z(n12712) );
  XOR U12951 ( .A(n12714), .B(n12713), .Z(n12700) );
  XOR U12952 ( .A(n12750), .B(n12749), .Z(n12763) );
  XOR U12953 ( .A(n12397), .B(n12763), .Z(n12761) );
  NAND U12954 ( .A(n12399), .B(n12398), .Z(n12403) );
  NANDN U12955 ( .A(n12401), .B(n12400), .Z(n12402) );
  AND U12956 ( .A(n12403), .B(n12402), .Z(n12487) );
  NANDN U12957 ( .A(n12405), .B(n12404), .Z(n12409) );
  NANDN U12958 ( .A(n12407), .B(n12406), .Z(n12408) );
  AND U12959 ( .A(n12409), .B(n12408), .Z(n12494) );
  NANDN U12960 ( .A(n12411), .B(n12410), .Z(n12415) );
  NANDN U12961 ( .A(n12413), .B(n12412), .Z(n12414) );
  AND U12962 ( .A(n12415), .B(n12414), .Z(n12496) );
  NAND U12963 ( .A(n12417), .B(n12416), .Z(n12421) );
  NAND U12964 ( .A(n12419), .B(n12418), .Z(n12420) );
  AND U12965 ( .A(n12421), .B(n12420), .Z(n12768) );
  NAND U12966 ( .A(n12423), .B(n12422), .Z(n12427) );
  NANDN U12967 ( .A(n12425), .B(n12424), .Z(n12426) );
  AND U12968 ( .A(n12427), .B(n12426), .Z(n12500) );
  AND U12969 ( .A(y[86]), .B(x[136]), .Z(n12586) );
  AND U12970 ( .A(y[0]), .B(x[126]), .Z(n12585) );
  XOR U12971 ( .A(n12586), .B(n12585), .Z(n12584) );
  AND U12972 ( .A(y[121]), .B(x[149]), .Z(n12583) );
  XOR U12973 ( .A(n12584), .B(n12583), .Z(n12522) );
  AND U12974 ( .A(y[41]), .B(x[133]), .Z(n12580) );
  AND U12975 ( .A(y[44]), .B(x[130]), .Z(n12579) );
  XOR U12976 ( .A(n12580), .B(n12579), .Z(n12578) );
  AND U12977 ( .A(y[45]), .B(x[129]), .Z(n12577) );
  XOR U12978 ( .A(n12578), .B(n12577), .Z(n12639) );
  NAND U12979 ( .A(x[132]), .B(y[42]), .Z(n12428) );
  XNOR U12980 ( .A(n12429), .B(n12428), .Z(n12638) );
  XOR U12981 ( .A(n12639), .B(n12638), .Z(n12521) );
  XOR U12982 ( .A(n12522), .B(n12521), .Z(n12520) );
  AND U12983 ( .A(y[166]), .B(x[152]), .Z(n12571) );
  XOR U12984 ( .A(n12572), .B(n12571), .Z(n12570) );
  AND U12985 ( .A(y[80]), .B(x[142]), .Z(n12569) );
  XOR U12986 ( .A(n12570), .B(n12569), .Z(n12519) );
  XOR U12987 ( .A(n12520), .B(n12519), .Z(n12502) );
  NAND U12988 ( .A(n12431), .B(n12430), .Z(n12435) );
  NAND U12989 ( .A(n12433), .B(n12432), .Z(n12434) );
  AND U12990 ( .A(n12435), .B(n12434), .Z(n12719) );
  AND U12991 ( .A(x[137]), .B(y[85]), .Z(n12437) );
  NAND U12992 ( .A(x[138]), .B(y[84]), .Z(n12436) );
  XNOR U12993 ( .A(n12437), .B(n12436), .Z(n12548) );
  AND U12994 ( .A(y[122]), .B(x[148]), .Z(n12547) );
  XOR U12995 ( .A(n12548), .B(n12547), .Z(n12722) );
  AND U12996 ( .A(x[144]), .B(y[126]), .Z(n12439) );
  NAND U12997 ( .A(x[145]), .B(y[125]), .Z(n12438) );
  XNOR U12998 ( .A(n12439), .B(n12438), .Z(n12565) );
  AND U12999 ( .A(y[6]), .B(x[120]), .Z(n12564) );
  XNOR U13000 ( .A(n12565), .B(n12564), .Z(n12721) );
  XNOR U13001 ( .A(n12719), .B(n12720), .Z(n12501) );
  XOR U13002 ( .A(n12500), .B(n12499), .Z(n12767) );
  XOR U13003 ( .A(n12768), .B(n12767), .Z(n12769) );
  NANDN U13004 ( .A(n12549), .B(n12440), .Z(n12444) );
  NANDN U13005 ( .A(n12442), .B(n12441), .Z(n12443) );
  NAND U13006 ( .A(n12444), .B(n12443), .Z(n12741) );
  NANDN U13007 ( .A(n12445), .B(n12615), .Z(n12449) );
  NAND U13008 ( .A(n12447), .B(n12446), .Z(n12448) );
  NAND U13009 ( .A(n12449), .B(n12448), .Z(n12744) );
  NANDN U13010 ( .A(n12451), .B(n12450), .Z(n12455) );
  NANDN U13011 ( .A(n12453), .B(n12452), .Z(n12454) );
  AND U13012 ( .A(n12455), .B(n12454), .Z(n12706) );
  AND U13013 ( .A(y[5]), .B(x[121]), .Z(n12534) );
  AND U13014 ( .A(y[40]), .B(x[134]), .Z(n12533) );
  XOR U13015 ( .A(n12534), .B(n12533), .Z(n12532) );
  AND U13016 ( .A(y[46]), .B(x[128]), .Z(n12531) );
  XOR U13017 ( .A(n12532), .B(n12531), .Z(n12707) );
  NAND U13018 ( .A(x[157]), .B(y[161]), .Z(n12456) );
  XNOR U13019 ( .A(n12457), .B(n12456), .Z(n12542) );
  AND U13020 ( .A(y[160]), .B(x[158]), .Z(n12541) );
  XOR U13021 ( .A(n12542), .B(n12541), .Z(n12538) );
  XNOR U13022 ( .A(n12539), .B(n12538), .Z(n12708) );
  XNOR U13023 ( .A(n12706), .B(n12705), .Z(n12743) );
  XOR U13024 ( .A(n12744), .B(n12743), .Z(n12742) );
  XOR U13025 ( .A(n12741), .B(n12742), .Z(n12770) );
  XOR U13026 ( .A(n12494), .B(n12493), .Z(n12485) );
  XOR U13027 ( .A(n12486), .B(n12485), .Z(n12481) );
  NANDN U13028 ( .A(n12459), .B(n12458), .Z(n12463) );
  NANDN U13029 ( .A(n12461), .B(n12460), .Z(n12462) );
  NAND U13030 ( .A(n12463), .B(n12462), .Z(n12484) );
  XNOR U13031 ( .A(n12484), .B(n12483), .Z(n12482) );
  XNOR U13032 ( .A(n12481), .B(n12482), .Z(n12492) );
  NANDN U13033 ( .A(n12469), .B(n12468), .Z(n12473) );
  NANDN U13034 ( .A(n12471), .B(n12470), .Z(n12472) );
  AND U13035 ( .A(n12473), .B(n12472), .Z(n12491) );
  NANDN U13036 ( .A(n12475), .B(n12474), .Z(n12479) );
  NAND U13037 ( .A(n12477), .B(n12476), .Z(n12478) );
  AND U13038 ( .A(n12479), .B(n12478), .Z(n12489) );
  XOR U13039 ( .A(n12491), .B(n12489), .Z(n12480) );
  XNOR U13040 ( .A(n12492), .B(n12480), .Z(o[126]) );
  IV U13041 ( .A(n12489), .Z(n12490) );
  NAND U13042 ( .A(n12494), .B(n12493), .Z(n12498) );
  NANDN U13043 ( .A(n12496), .B(n12495), .Z(n12497) );
  NAND U13044 ( .A(n12500), .B(n12499), .Z(n12504) );
  NANDN U13045 ( .A(n12502), .B(n12501), .Z(n12503) );
  AND U13046 ( .A(n12504), .B(n12503), .Z(n12512) );
  ANDN U13047 ( .B(n12506), .A(n12505), .Z(n12510) );
  AND U13048 ( .A(n12508), .B(n12507), .Z(n12509) );
  OR U13049 ( .A(n12510), .B(n12509), .Z(n12511) );
  XNOR U13050 ( .A(n12512), .B(n12511), .Z(n12760) );
  NANDN U13051 ( .A(n12514), .B(n12513), .Z(n12518) );
  NANDN U13052 ( .A(n12516), .B(n12515), .Z(n12517) );
  AND U13053 ( .A(n12518), .B(n12517), .Z(n12758) );
  NAND U13054 ( .A(n12520), .B(n12519), .Z(n12524) );
  NAND U13055 ( .A(n12522), .B(n12521), .Z(n12523) );
  AND U13056 ( .A(n12524), .B(n12523), .Z(n12740) );
  NAND U13057 ( .A(n12526), .B(n12525), .Z(n12530) );
  NAND U13058 ( .A(n12528), .B(n12527), .Z(n12529) );
  AND U13059 ( .A(n12530), .B(n12529), .Z(n12698) );
  NAND U13060 ( .A(n12532), .B(n12531), .Z(n12536) );
  NAND U13061 ( .A(n12534), .B(n12533), .Z(n12535) );
  AND U13062 ( .A(n12536), .B(n12535), .Z(n12563) );
  AND U13063 ( .A(y[162]), .B(x[157]), .Z(n12658) );
  NAND U13064 ( .A(n12537), .B(n12658), .Z(n12544) );
  NAND U13065 ( .A(n12539), .B(n12538), .Z(n12540) );
  XNOR U13066 ( .A(n12544), .B(n12540), .Z(n12546) );
  AND U13067 ( .A(n12542), .B(n12541), .Z(n12543) );
  NAND U13068 ( .A(n12544), .B(n12543), .Z(n12545) );
  NAND U13069 ( .A(n12546), .B(n12545), .Z(n12561) );
  NAND U13070 ( .A(n12548), .B(n12547), .Z(n12551) );
  AND U13071 ( .A(y[85]), .B(x[138]), .Z(n12684) );
  NANDN U13072 ( .A(n12549), .B(n12684), .Z(n12550) );
  AND U13073 ( .A(n12551), .B(n12550), .Z(n12559) );
  NAND U13074 ( .A(n12553), .B(n12552), .Z(n12557) );
  NAND U13075 ( .A(n12555), .B(n12554), .Z(n12556) );
  NAND U13076 ( .A(n12557), .B(n12556), .Z(n12558) );
  XNOR U13077 ( .A(n12559), .B(n12558), .Z(n12560) );
  XNOR U13078 ( .A(n12561), .B(n12560), .Z(n12562) );
  XNOR U13079 ( .A(n12563), .B(n12562), .Z(n12696) );
  NAND U13080 ( .A(n12565), .B(n12564), .Z(n12568) );
  AND U13081 ( .A(y[126]), .B(x[145]), .Z(n12657) );
  NANDN U13082 ( .A(n12566), .B(n12657), .Z(n12567) );
  AND U13083 ( .A(n12568), .B(n12567), .Z(n12576) );
  NAND U13084 ( .A(n12570), .B(n12569), .Z(n12574) );
  NAND U13085 ( .A(n12572), .B(n12571), .Z(n12573) );
  NAND U13086 ( .A(n12574), .B(n12573), .Z(n12575) );
  XNOR U13087 ( .A(n12576), .B(n12575), .Z(n12623) );
  NAND U13088 ( .A(n12578), .B(n12577), .Z(n12582) );
  NAND U13089 ( .A(n12580), .B(n12579), .Z(n12581) );
  AND U13090 ( .A(n12582), .B(n12581), .Z(n12613) );
  NAND U13091 ( .A(n12584), .B(n12583), .Z(n12588) );
  NAND U13092 ( .A(n12586), .B(n12585), .Z(n12587) );
  AND U13093 ( .A(n12588), .B(n12587), .Z(n12595) );
  NANDN U13094 ( .A(n12590), .B(n12589), .Z(n12593) );
  AND U13095 ( .A(y[2]), .B(x[125]), .Z(n12678) );
  NANDN U13096 ( .A(n12591), .B(n12678), .Z(n12592) );
  NAND U13097 ( .A(n12593), .B(n12592), .Z(n12594) );
  XNOR U13098 ( .A(n12595), .B(n12594), .Z(n12611) );
  AND U13099 ( .A(x[152]), .B(y[167]), .Z(n12597) );
  NAND U13100 ( .A(x[142]), .B(y[81]), .Z(n12596) );
  XNOR U13101 ( .A(n12597), .B(n12596), .Z(n12601) );
  AND U13102 ( .A(x[153]), .B(y[166]), .Z(n12599) );
  NAND U13103 ( .A(x[126]), .B(y[1]), .Z(n12598) );
  XNOR U13104 ( .A(n12599), .B(n12598), .Z(n12600) );
  XOR U13105 ( .A(n12601), .B(n12600), .Z(n12609) );
  AND U13106 ( .A(x[136]), .B(y[87]), .Z(n12603) );
  NAND U13107 ( .A(x[143]), .B(y[80]), .Z(n12602) );
  XNOR U13108 ( .A(n12603), .B(n12602), .Z(n12607) );
  AND U13109 ( .A(x[128]), .B(y[47]), .Z(n12605) );
  NAND U13110 ( .A(x[147]), .B(y[124]), .Z(n12604) );
  XNOR U13111 ( .A(n12605), .B(n12604), .Z(n12606) );
  XNOR U13112 ( .A(n12607), .B(n12606), .Z(n12608) );
  XNOR U13113 ( .A(n12609), .B(n12608), .Z(n12610) );
  XNOR U13114 ( .A(n12611), .B(n12610), .Z(n12612) );
  XNOR U13115 ( .A(n12613), .B(n12612), .Z(n12621) );
  NAND U13116 ( .A(n12615), .B(n12614), .Z(n12619) );
  NANDN U13117 ( .A(n12617), .B(n12616), .Z(n12618) );
  NAND U13118 ( .A(n12619), .B(n12618), .Z(n12620) );
  XNOR U13119 ( .A(n12621), .B(n12620), .Z(n12622) );
  XOR U13120 ( .A(n12623), .B(n12622), .Z(n12694) );
  AND U13121 ( .A(x[123]), .B(y[4]), .Z(n12625) );
  NAND U13122 ( .A(x[134]), .B(y[41]), .Z(n12624) );
  XNOR U13123 ( .A(n12625), .B(n12624), .Z(n12629) );
  AND U13124 ( .A(x[137]), .B(y[86]), .Z(n12627) );
  NAND U13125 ( .A(x[150]), .B(y[121]), .Z(n12626) );
  XNOR U13126 ( .A(n12627), .B(n12626), .Z(n12628) );
  XOR U13127 ( .A(n12629), .B(n12628), .Z(n12637) );
  AND U13128 ( .A(x[144]), .B(y[127]), .Z(n12631) );
  NAND U13129 ( .A(x[129]), .B(y[46]), .Z(n12630) );
  XNOR U13130 ( .A(n12631), .B(n12630), .Z(n12635) );
  AND U13131 ( .A(x[122]), .B(y[5]), .Z(n12633) );
  NAND U13132 ( .A(x[151]), .B(y[120]), .Z(n12632) );
  XNOR U13133 ( .A(n12633), .B(n12632), .Z(n12634) );
  XNOR U13134 ( .A(n12635), .B(n12634), .Z(n12636) );
  XNOR U13135 ( .A(n12637), .B(n12636), .Z(n12692) );
  NAND U13136 ( .A(n12639), .B(n12638), .Z(n12642) );
  AND U13137 ( .A(y[42]), .B(x[131]), .Z(n12640) );
  AND U13138 ( .A(y[43]), .B(x[132]), .Z(n12677) );
  NAND U13139 ( .A(n12640), .B(n12677), .Z(n12641) );
  AND U13140 ( .A(n12642), .B(n12641), .Z(n12690) );
  AND U13141 ( .A(x[148]), .B(y[123]), .Z(n12644) );
  NAND U13142 ( .A(x[141]), .B(y[82]), .Z(n12643) );
  XNOR U13143 ( .A(n12644), .B(n12643), .Z(n12648) );
  AND U13144 ( .A(x[120]), .B(y[7]), .Z(n12646) );
  NAND U13145 ( .A(x[127]), .B(y[0]), .Z(n12645) );
  XNOR U13146 ( .A(n12646), .B(n12645), .Z(n12647) );
  XOR U13147 ( .A(n12648), .B(n12647), .Z(n12656) );
  AND U13148 ( .A(x[139]), .B(y[84]), .Z(n12650) );
  NAND U13149 ( .A(x[149]), .B(y[122]), .Z(n12649) );
  XNOR U13150 ( .A(n12650), .B(n12649), .Z(n12654) );
  AND U13151 ( .A(x[121]), .B(y[6]), .Z(n12652) );
  NAND U13152 ( .A(x[140]), .B(y[83]), .Z(n12651) );
  XNOR U13153 ( .A(n12652), .B(n12651), .Z(n12653) );
  XNOR U13154 ( .A(n12654), .B(n12653), .Z(n12655) );
  XNOR U13155 ( .A(n12656), .B(n12655), .Z(n12688) );
  AND U13156 ( .A(x[158]), .B(y[161]), .Z(n12660) );
  XNOR U13157 ( .A(n12658), .B(n12657), .Z(n12659) );
  XNOR U13158 ( .A(n12660), .B(n12659), .Z(n12676) );
  AND U13159 ( .A(x[146]), .B(y[125]), .Z(n12662) );
  NAND U13160 ( .A(x[135]), .B(y[40]), .Z(n12661) );
  XNOR U13161 ( .A(n12662), .B(n12661), .Z(n12666) );
  AND U13162 ( .A(x[130]), .B(y[45]), .Z(n12664) );
  NAND U13163 ( .A(x[133]), .B(y[42]), .Z(n12663) );
  XNOR U13164 ( .A(n12664), .B(n12663), .Z(n12665) );
  XOR U13165 ( .A(n12666), .B(n12665), .Z(n12674) );
  AND U13166 ( .A(x[124]), .B(y[3]), .Z(n12668) );
  NAND U13167 ( .A(x[155]), .B(y[164]), .Z(n12667) );
  XNOR U13168 ( .A(n12668), .B(n12667), .Z(n12672) );
  AND U13169 ( .A(x[154]), .B(y[165]), .Z(n12670) );
  NAND U13170 ( .A(x[159]), .B(y[160]), .Z(n12669) );
  XNOR U13171 ( .A(n12670), .B(n12669), .Z(n12671) );
  XNOR U13172 ( .A(n12672), .B(n12671), .Z(n12673) );
  XNOR U13173 ( .A(n12674), .B(n12673), .Z(n12675) );
  XOR U13174 ( .A(n12676), .B(n12675), .Z(n12686) );
  XOR U13175 ( .A(n12678), .B(n12677), .Z(n12682) );
  XNOR U13176 ( .A(n12680), .B(n12679), .Z(n12681) );
  XNOR U13177 ( .A(n12682), .B(n12681), .Z(n12683) );
  XNOR U13178 ( .A(n12684), .B(n12683), .Z(n12685) );
  XNOR U13179 ( .A(n12686), .B(n12685), .Z(n12687) );
  XNOR U13180 ( .A(n12688), .B(n12687), .Z(n12689) );
  XNOR U13181 ( .A(n12690), .B(n12689), .Z(n12691) );
  XNOR U13182 ( .A(n12692), .B(n12691), .Z(n12693) );
  XNOR U13183 ( .A(n12694), .B(n12693), .Z(n12695) );
  XNOR U13184 ( .A(n12696), .B(n12695), .Z(n12697) );
  XNOR U13185 ( .A(n12698), .B(n12697), .Z(n12738) );
  NANDN U13186 ( .A(n12700), .B(n12699), .Z(n12704) );
  NANDN U13187 ( .A(n12702), .B(n12701), .Z(n12703) );
  AND U13188 ( .A(n12704), .B(n12703), .Z(n12736) );
  NAND U13189 ( .A(n12706), .B(n12705), .Z(n12710) );
  ANDN U13190 ( .B(n12708), .A(n12707), .Z(n12709) );
  ANDN U13191 ( .B(n12710), .A(n12709), .Z(n12718) );
  ANDN U13192 ( .B(n12712), .A(n12711), .Z(n12716) );
  AND U13193 ( .A(n12714), .B(n12713), .Z(n12715) );
  OR U13194 ( .A(n12716), .B(n12715), .Z(n12717) );
  XNOR U13195 ( .A(n12718), .B(n12717), .Z(n12734) );
  NANDN U13196 ( .A(n12720), .B(n12719), .Z(n12724) );
  NANDN U13197 ( .A(n12722), .B(n12721), .Z(n12723) );
  AND U13198 ( .A(n12724), .B(n12723), .Z(n12732) );
  NAND U13199 ( .A(n12726), .B(n12725), .Z(n12730) );
  NANDN U13200 ( .A(n12728), .B(n12727), .Z(n12729) );
  NAND U13201 ( .A(n12730), .B(n12729), .Z(n12731) );
  XNOR U13202 ( .A(n12732), .B(n12731), .Z(n12733) );
  XNOR U13203 ( .A(n12734), .B(n12733), .Z(n12735) );
  XNOR U13204 ( .A(n12736), .B(n12735), .Z(n12737) );
  XNOR U13205 ( .A(n12738), .B(n12737), .Z(n12739) );
  XNOR U13206 ( .A(n12740), .B(n12739), .Z(n12756) );
  NAND U13207 ( .A(n12742), .B(n12741), .Z(n12746) );
  AND U13208 ( .A(n12744), .B(n12743), .Z(n12745) );
  ANDN U13209 ( .B(n12746), .A(n12745), .Z(n12754) );
  ANDN U13210 ( .B(n12748), .A(n12747), .Z(n12752) );
  AND U13211 ( .A(n12750), .B(n12749), .Z(n12751) );
  OR U13212 ( .A(n12752), .B(n12751), .Z(n12753) );
  XNOR U13213 ( .A(n12754), .B(n12753), .Z(n12755) );
  XNOR U13214 ( .A(n12756), .B(n12755), .Z(n12757) );
  XNOR U13215 ( .A(n12758), .B(n12757), .Z(n12759) );
  NANDN U13216 ( .A(n12762), .B(n12761), .Z(n12766) );
  NANDN U13217 ( .A(n12764), .B(n12763), .Z(n12765) );
  NAND U13218 ( .A(n12768), .B(n12767), .Z(n12772) );
  NANDN U13219 ( .A(n12770), .B(n12769), .Z(n12771) );
  NAND U13220 ( .A(y[168]), .B(x[152]), .Z(n12907) );
  NAND U13221 ( .A(y[48]), .B(x[128]), .Z(n12775) );
  XOR U13222 ( .A(n12907), .B(n12775), .Z(n12776) );
  AND U13223 ( .A(y[8]), .B(x[120]), .Z(n12783) );
  AND U13224 ( .A(y[88]), .B(x[136]), .Z(n12780) );
  XOR U13225 ( .A(n12783), .B(n12780), .Z(n12779) );
  AND U13226 ( .A(y[128]), .B(x[144]), .Z(n12778) );
  XNOR U13227 ( .A(n12779), .B(n12778), .Z(n12777) );
  XNOR U13228 ( .A(n12776), .B(n12777), .Z(o[128]) );
  AND U13229 ( .A(x[120]), .B(y[9]), .Z(n12774) );
  NAND U13230 ( .A(x[121]), .B(y[8]), .Z(n12773) );
  XNOR U13231 ( .A(n12774), .B(n12773), .Z(n12784) );
  NAND U13232 ( .A(y[48]), .B(x[129]), .Z(n12785) );
  XOR U13233 ( .A(n12784), .B(n12785), .Z(n12801) );
  AND U13234 ( .A(y[168]), .B(x[153]), .Z(n13008) );
  NAND U13235 ( .A(y[89]), .B(x[136]), .Z(n12788) );
  XNOR U13236 ( .A(n13008), .B(n12788), .Z(n12789) );
  AND U13237 ( .A(y[169]), .B(x[152]), .Z(n12812) );
  NAND U13238 ( .A(y[88]), .B(x[137]), .Z(n12811) );
  XOR U13239 ( .A(n12812), .B(n12811), .Z(n12790) );
  XOR U13240 ( .A(n12789), .B(n12790), .Z(n12800) );
  AND U13241 ( .A(y[49]), .B(x[128]), .Z(n13032) );
  AND U13242 ( .A(y[129]), .B(x[144]), .Z(n12805) );
  XOR U13243 ( .A(n13032), .B(n12805), .Z(n12807) );
  AND U13244 ( .A(y[128]), .B(x[145]), .Z(n12806) );
  XNOR U13245 ( .A(n12807), .B(n12806), .Z(n12799) );
  XOR U13246 ( .A(n12800), .B(n12799), .Z(n12802) );
  XOR U13247 ( .A(n12801), .B(n12802), .Z(n12796) );
  NAND U13248 ( .A(n12779), .B(n12778), .Z(n12782) );
  AND U13249 ( .A(n12783), .B(n12780), .Z(n12781) );
  ANDN U13250 ( .B(n12782), .A(n12781), .Z(n12793) );
  XNOR U13251 ( .A(n12794), .B(n12793), .Z(n12795) );
  XNOR U13252 ( .A(n12796), .B(n12795), .Z(o[129]) );
  AND U13253 ( .A(y[9]), .B(x[121]), .Z(n12842) );
  NAND U13254 ( .A(n12842), .B(n12783), .Z(n12787) );
  NANDN U13255 ( .A(n12785), .B(n12784), .Z(n12786) );
  NAND U13256 ( .A(n12787), .B(n12786), .Z(n12854) );
  NANDN U13257 ( .A(n12788), .B(n13008), .Z(n12792) );
  NANDN U13258 ( .A(n12790), .B(n12789), .Z(n12791) );
  NAND U13259 ( .A(n12792), .B(n12791), .Z(n12852) );
  AND U13260 ( .A(y[130]), .B(x[144]), .Z(n12858) );
  NAND U13261 ( .A(y[10]), .B(x[120]), .Z(n12859) );
  XNOR U13262 ( .A(n12858), .B(n12859), .Z(n12861) );
  AND U13263 ( .A(y[48]), .B(x[130]), .Z(n12860) );
  XOR U13264 ( .A(n12861), .B(n12860), .Z(n12853) );
  XOR U13265 ( .A(n12852), .B(n12853), .Z(n12855) );
  XNOR U13266 ( .A(n12854), .B(n12855), .Z(n12814) );
  NANDN U13267 ( .A(n12794), .B(n12793), .Z(n12798) );
  NAND U13268 ( .A(n12796), .B(n12795), .Z(n12797) );
  NAND U13269 ( .A(n12798), .B(n12797), .Z(n12813) );
  XOR U13270 ( .A(n12814), .B(n12813), .Z(n12816) );
  NAND U13271 ( .A(n12800), .B(n12799), .Z(n12804) );
  NAND U13272 ( .A(n12802), .B(n12801), .Z(n12803) );
  AND U13273 ( .A(n12804), .B(n12803), .Z(n12822) );
  AND U13274 ( .A(y[8]), .B(x[122]), .Z(n12840) );
  AND U13275 ( .A(y[90]), .B(x[136]), .Z(n12839) );
  XOR U13276 ( .A(n12840), .B(n12839), .Z(n12841) );
  XOR U13277 ( .A(n12842), .B(n12841), .Z(n12867) );
  AND U13278 ( .A(y[128]), .B(x[146]), .Z(n12866) );
  XOR U13279 ( .A(n12867), .B(n12866), .Z(n12869) );
  AND U13280 ( .A(y[88]), .B(x[138]), .Z(n12946) );
  AND U13281 ( .A(y[170]), .B(x[152]), .Z(n12831) );
  XOR U13282 ( .A(n12946), .B(n12831), .Z(n12833) );
  AND U13283 ( .A(y[89]), .B(x[137]), .Z(n12832) );
  XOR U13284 ( .A(n12833), .B(n12832), .Z(n12868) );
  XOR U13285 ( .A(n12869), .B(n12868), .Z(n12819) );
  AND U13286 ( .A(n13032), .B(n12805), .Z(n12809) );
  NAND U13287 ( .A(n12807), .B(n12806), .Z(n12808) );
  NANDN U13288 ( .A(n12809), .B(n12808), .Z(n12827) );
  AND U13289 ( .A(x[153]), .B(y[169]), .Z(n12912) );
  NAND U13290 ( .A(x[154]), .B(y[168]), .Z(n12810) );
  XNOR U13291 ( .A(n12912), .B(n12810), .Z(n12865) );
  ANDN U13292 ( .B(n12812), .A(n12811), .Z(n12864) );
  XOR U13293 ( .A(n12865), .B(n12864), .Z(n12826) );
  AND U13294 ( .A(y[129]), .B(x[145]), .Z(n12845) );
  NAND U13295 ( .A(y[49]), .B(x[129]), .Z(n12846) );
  XNOR U13296 ( .A(n12845), .B(n12846), .Z(n12847) );
  NAND U13297 ( .A(y[50]), .B(x[128]), .Z(n12848) );
  XNOR U13298 ( .A(n12847), .B(n12848), .Z(n12825) );
  XOR U13299 ( .A(n12826), .B(n12825), .Z(n12828) );
  XOR U13300 ( .A(n12827), .B(n12828), .Z(n12820) );
  XOR U13301 ( .A(n12819), .B(n12820), .Z(n12821) );
  XNOR U13302 ( .A(n12822), .B(n12821), .Z(n12815) );
  XNOR U13303 ( .A(n12816), .B(n12815), .Z(o[130]) );
  NAND U13304 ( .A(n12814), .B(n12813), .Z(n12818) );
  NAND U13305 ( .A(n12816), .B(n12815), .Z(n12817) );
  AND U13306 ( .A(n12818), .B(n12817), .Z(n12873) );
  NAND U13307 ( .A(n12820), .B(n12819), .Z(n12824) );
  NAND U13308 ( .A(n12822), .B(n12821), .Z(n12823) );
  NAND U13309 ( .A(n12824), .B(n12823), .Z(n12878) );
  NAND U13310 ( .A(n12826), .B(n12825), .Z(n12830) );
  NAND U13311 ( .A(n12828), .B(n12827), .Z(n12829) );
  NAND U13312 ( .A(n12830), .B(n12829), .Z(n12876) );
  NAND U13313 ( .A(n12946), .B(n12831), .Z(n12835) );
  AND U13314 ( .A(n12833), .B(n12832), .Z(n12834) );
  ANDN U13315 ( .B(n12835), .A(n12834), .Z(n12934) );
  AND U13316 ( .A(y[10]), .B(x[121]), .Z(n12903) );
  AND U13317 ( .A(y[9]), .B(x[122]), .Z(n12902) );
  NAND U13318 ( .A(y[130]), .B(x[145]), .Z(n12901) );
  XOR U13319 ( .A(n12902), .B(n12901), .Z(n12904) );
  XOR U13320 ( .A(n12903), .B(n12904), .Z(n12932) );
  AND U13321 ( .A(x[155]), .B(y[168]), .Z(n12837) );
  NAND U13322 ( .A(x[152]), .B(y[171]), .Z(n12836) );
  XNOR U13323 ( .A(n12837), .B(n12836), .Z(n12908) );
  AND U13324 ( .A(y[169]), .B(x[154]), .Z(n13005) );
  NAND U13325 ( .A(x[153]), .B(y[170]), .Z(n12838) );
  XOR U13326 ( .A(n13005), .B(n12838), .Z(n12909) );
  XNOR U13327 ( .A(n12908), .B(n12909), .Z(n12931) );
  XNOR U13328 ( .A(n12932), .B(n12931), .Z(n12933) );
  XNOR U13329 ( .A(n12934), .B(n12933), .Z(n12890) );
  NAND U13330 ( .A(n12840), .B(n12839), .Z(n12844) );
  NAND U13331 ( .A(n12842), .B(n12841), .Z(n12843) );
  NAND U13332 ( .A(n12844), .B(n12843), .Z(n12888) );
  NANDN U13333 ( .A(n12846), .B(n12845), .Z(n12850) );
  NANDN U13334 ( .A(n12848), .B(n12847), .Z(n12849) );
  AND U13335 ( .A(n12850), .B(n12849), .Z(n12927) );
  AND U13336 ( .A(y[131]), .B(x[144]), .Z(n12942) );
  AND U13337 ( .A(y[91]), .B(x[136]), .Z(n12941) );
  NAND U13338 ( .A(y[8]), .B(x[123]), .Z(n12940) );
  XOR U13339 ( .A(n12941), .B(n12940), .Z(n12943) );
  XOR U13340 ( .A(n12942), .B(n12943), .Z(n12926) );
  AND U13341 ( .A(y[89]), .B(x[138]), .Z(n12987) );
  NAND U13342 ( .A(x[139]), .B(y[88]), .Z(n12851) );
  XNOR U13343 ( .A(n12987), .B(n12851), .Z(n12947) );
  NAND U13344 ( .A(y[90]), .B(x[137]), .Z(n12948) );
  XNOR U13345 ( .A(n12947), .B(n12948), .Z(n12925) );
  XOR U13346 ( .A(n12926), .B(n12925), .Z(n12928) );
  XOR U13347 ( .A(n12927), .B(n12928), .Z(n12889) );
  XOR U13348 ( .A(n12888), .B(n12889), .Z(n12891) );
  XOR U13349 ( .A(n12890), .B(n12891), .Z(n12877) );
  XOR U13350 ( .A(n12876), .B(n12877), .Z(n12879) );
  XOR U13351 ( .A(n12878), .B(n12879), .Z(n12872) );
  XOR U13352 ( .A(n12873), .B(n12872), .Z(n12875) );
  NAND U13353 ( .A(n12853), .B(n12852), .Z(n12857) );
  NAND U13354 ( .A(n12855), .B(n12854), .Z(n12856) );
  AND U13355 ( .A(n12857), .B(n12856), .Z(n12885) );
  NANDN U13356 ( .A(n12859), .B(n12858), .Z(n12863) );
  NAND U13357 ( .A(n12861), .B(n12860), .Z(n12862) );
  AND U13358 ( .A(n12863), .B(n12862), .Z(n12895) );
  XNOR U13359 ( .A(n12895), .B(n12894), .Z(n12897) );
  NAND U13360 ( .A(y[48]), .B(x[131]), .Z(n12956) );
  NAND U13361 ( .A(y[11]), .B(x[120]), .Z(n12954) );
  NAND U13362 ( .A(y[129]), .B(x[146]), .Z(n12953) );
  XOR U13363 ( .A(n12954), .B(n12953), .Z(n12955) );
  XNOR U13364 ( .A(n12956), .B(n12955), .Z(n12922) );
  NAND U13365 ( .A(y[51]), .B(x[128]), .Z(n12916) );
  NAND U13366 ( .A(y[49]), .B(x[130]), .Z(n12914) );
  NAND U13367 ( .A(y[128]), .B(x[147]), .Z(n12913) );
  XOR U13368 ( .A(n12914), .B(n12913), .Z(n12915) );
  XNOR U13369 ( .A(n12916), .B(n12915), .Z(n12920) );
  AND U13370 ( .A(y[50]), .B(x[129]), .Z(n12919) );
  XOR U13371 ( .A(n12920), .B(n12919), .Z(n12921) );
  XOR U13372 ( .A(n12922), .B(n12921), .Z(n12896) );
  XNOR U13373 ( .A(n12897), .B(n12896), .Z(n12883) );
  NAND U13374 ( .A(n12867), .B(n12866), .Z(n12871) );
  NAND U13375 ( .A(n12869), .B(n12868), .Z(n12870) );
  AND U13376 ( .A(n12871), .B(n12870), .Z(n12882) );
  XOR U13377 ( .A(n12883), .B(n12882), .Z(n12884) );
  XNOR U13378 ( .A(n12885), .B(n12884), .Z(n12874) );
  XOR U13379 ( .A(n12875), .B(n12874), .Z(o[131]) );
  NAND U13380 ( .A(n12877), .B(n12876), .Z(n12881) );
  NAND U13381 ( .A(n12879), .B(n12878), .Z(n12880) );
  AND U13382 ( .A(n12881), .B(n12880), .Z(n12965) );
  NAND U13383 ( .A(n12883), .B(n12882), .Z(n12887) );
  NAND U13384 ( .A(n12885), .B(n12884), .Z(n12886) );
  NAND U13385 ( .A(n12887), .B(n12886), .Z(n12963) );
  NAND U13386 ( .A(n12889), .B(n12888), .Z(n12893) );
  NAND U13387 ( .A(n12891), .B(n12890), .Z(n12892) );
  AND U13388 ( .A(n12893), .B(n12892), .Z(n12964) );
  XOR U13389 ( .A(n12963), .B(n12964), .Z(n12966) );
  XOR U13390 ( .A(n12965), .B(n12966), .Z(n12959) );
  XOR U13391 ( .A(n12960), .B(n12959), .Z(n12962) );
  AND U13392 ( .A(y[50]), .B(x[130]), .Z(n13096) );
  AND U13393 ( .A(x[131]), .B(y[49]), .Z(n12899) );
  NAND U13394 ( .A(x[128]), .B(y[52]), .Z(n12898) );
  XOR U13395 ( .A(n12899), .B(n12898), .Z(n13033) );
  IV U13396 ( .A(n13033), .Z(n12900) );
  XOR U13397 ( .A(n13096), .B(n12900), .Z(n13036) );
  NAND U13398 ( .A(y[51]), .B(x[129]), .Z(n13037) );
  AND U13399 ( .A(y[128]), .B(x[148]), .Z(n12992) );
  NAND U13400 ( .A(y[11]), .B(x[121]), .Z(n12993) );
  NAND U13401 ( .A(y[12]), .B(x[120]), .Z(n12995) );
  XOR U13402 ( .A(n13039), .B(n13038), .Z(n13051) );
  NANDN U13403 ( .A(n12902), .B(n12901), .Z(n12906) );
  OR U13404 ( .A(n12904), .B(n12903), .Z(n12905) );
  AND U13405 ( .A(n12906), .B(n12905), .Z(n13049) );
  AND U13406 ( .A(y[171]), .B(x[155]), .Z(n13265) );
  NANDN U13407 ( .A(n12907), .B(n13265), .Z(n12911) );
  NANDN U13408 ( .A(n12909), .B(n12908), .Z(n12910) );
  AND U13409 ( .A(n12911), .B(n12910), .Z(n13048) );
  NAND U13410 ( .A(y[8]), .B(x[124]), .Z(n13017) );
  NAND U13411 ( .A(y[130]), .B(x[146]), .Z(n13016) );
  NAND U13412 ( .A(y[92]), .B(x[136]), .Z(n13015) );
  XNOR U13413 ( .A(n13016), .B(n13015), .Z(n13018) );
  AND U13414 ( .A(y[170]), .B(x[154]), .Z(n12939) );
  NAND U13415 ( .A(n12939), .B(n12912), .Z(n13013) );
  NAND U13416 ( .A(y[172]), .B(x[152]), .Z(n13162) );
  NAND U13417 ( .A(y[88]), .B(x[140]), .Z(n13107) );
  XNOR U13418 ( .A(n13162), .B(n13107), .Z(n13014) );
  XOR U13419 ( .A(n13013), .B(n13014), .Z(n12975) );
  XOR U13420 ( .A(n12976), .B(n12975), .Z(n12978) );
  NAND U13421 ( .A(n12914), .B(n12913), .Z(n12918) );
  NAND U13422 ( .A(n12916), .B(n12915), .Z(n12917) );
  AND U13423 ( .A(n12918), .B(n12917), .Z(n12977) );
  XOR U13424 ( .A(n12978), .B(n12977), .Z(n13067) );
  NAND U13425 ( .A(n12920), .B(n12919), .Z(n12924) );
  NAND U13426 ( .A(n12922), .B(n12921), .Z(n12923) );
  AND U13427 ( .A(n12924), .B(n12923), .Z(n13066) );
  XNOR U13428 ( .A(n13067), .B(n13066), .Z(n13068) );
  XNOR U13429 ( .A(n13069), .B(n13068), .Z(n12969) );
  XNOR U13430 ( .A(n12970), .B(n12969), .Z(n12972) );
  NANDN U13431 ( .A(n12926), .B(n12925), .Z(n12930) );
  OR U13432 ( .A(n12928), .B(n12927), .Z(n12929) );
  AND U13433 ( .A(n12930), .B(n12929), .Z(n13055) );
  NANDN U13434 ( .A(n12932), .B(n12931), .Z(n12936) );
  NANDN U13435 ( .A(n12934), .B(n12933), .Z(n12935) );
  NAND U13436 ( .A(n12936), .B(n12935), .Z(n13054) );
  XNOR U13437 ( .A(n13055), .B(n13054), .Z(n13056) );
  NAND U13438 ( .A(y[10]), .B(x[122]), .Z(n13028) );
  NAND U13439 ( .A(y[129]), .B(x[147]), .Z(n13027) );
  NAND U13440 ( .A(y[9]), .B(x[123]), .Z(n13026) );
  XNOR U13441 ( .A(n13027), .B(n13026), .Z(n13029) );
  AND U13442 ( .A(x[156]), .B(y[168]), .Z(n12938) );
  NAND U13443 ( .A(x[153]), .B(y[171]), .Z(n12937) );
  XNOR U13444 ( .A(n12938), .B(n12937), .Z(n13010) );
  AND U13445 ( .A(y[169]), .B(x[155]), .Z(n13115) );
  XOR U13446 ( .A(n13115), .B(n12939), .Z(n13009) );
  XOR U13447 ( .A(n13010), .B(n13009), .Z(n12981) );
  NANDN U13448 ( .A(n12941), .B(n12940), .Z(n12945) );
  OR U13449 ( .A(n12943), .B(n12942), .Z(n12944) );
  NAND U13450 ( .A(n12945), .B(n12944), .Z(n12982) );
  XOR U13451 ( .A(n12983), .B(n12984), .Z(n13062) );
  AND U13452 ( .A(x[139]), .B(y[89]), .Z(n12952) );
  NAND U13453 ( .A(n12952), .B(n12946), .Z(n12950) );
  NANDN U13454 ( .A(n12948), .B(n12947), .Z(n12949) );
  AND U13455 ( .A(n12950), .B(n12949), .Z(n13061) );
  AND U13456 ( .A(y[48]), .B(x[132]), .Z(n12998) );
  NAND U13457 ( .A(y[132]), .B(x[144]), .Z(n12999) );
  NAND U13458 ( .A(y[131]), .B(x[145]), .Z(n13001) );
  NAND U13459 ( .A(x[138]), .B(y[90]), .Z(n12951) );
  XNOR U13460 ( .A(n12952), .B(n12951), .Z(n12988) );
  NAND U13461 ( .A(y[91]), .B(x[137]), .Z(n12989) );
  XOR U13462 ( .A(n13043), .B(n13042), .Z(n13044) );
  NAND U13463 ( .A(n12954), .B(n12953), .Z(n12958) );
  NAND U13464 ( .A(n12956), .B(n12955), .Z(n12957) );
  NAND U13465 ( .A(n12958), .B(n12957), .Z(n13045) );
  XOR U13466 ( .A(n13061), .B(n13060), .Z(n13063) );
  XOR U13467 ( .A(n13062), .B(n13063), .Z(n13057) );
  XNOR U13468 ( .A(n13056), .B(n13057), .Z(n12971) );
  XNOR U13469 ( .A(n12972), .B(n12971), .Z(n12961) );
  XNOR U13470 ( .A(n12962), .B(n12961), .Z(o[132]) );
  NAND U13471 ( .A(n12964), .B(n12963), .Z(n12968) );
  NAND U13472 ( .A(n12966), .B(n12965), .Z(n12967) );
  NAND U13473 ( .A(n12968), .B(n12967), .Z(n13216) );
  XNOR U13474 ( .A(n13215), .B(n13216), .Z(n13218) );
  NANDN U13475 ( .A(n12970), .B(n12969), .Z(n12974) );
  NAND U13476 ( .A(n12972), .B(n12971), .Z(n12973) );
  AND U13477 ( .A(n12974), .B(n12973), .Z(n13073) );
  NAND U13478 ( .A(n12976), .B(n12975), .Z(n12980) );
  NAND U13479 ( .A(n12978), .B(n12977), .Z(n12979) );
  AND U13480 ( .A(n12980), .B(n12979), .Z(n13127) );
  NANDN U13481 ( .A(n12982), .B(n12981), .Z(n12986) );
  NAND U13482 ( .A(n12984), .B(n12983), .Z(n12985) );
  NAND U13483 ( .A(n12986), .B(n12985), .Z(n13126) );
  AND U13484 ( .A(y[90]), .B(x[139]), .Z(n13108) );
  NAND U13485 ( .A(n13108), .B(n12987), .Z(n12991) );
  NANDN U13486 ( .A(n12989), .B(n12988), .Z(n12990) );
  AND U13487 ( .A(n12991), .B(n12990), .Z(n13079) );
  NANDN U13488 ( .A(n12993), .B(n12992), .Z(n12997) );
  NANDN U13489 ( .A(n12995), .B(n12994), .Z(n12996) );
  NAND U13490 ( .A(n12997), .B(n12996), .Z(n13086) );
  AND U13491 ( .A(y[133]), .B(x[144]), .Z(n13404) );
  AND U13492 ( .A(y[48]), .B(x[133]), .Z(n13122) );
  AND U13493 ( .A(y[91]), .B(x[138]), .Z(n13121) );
  XOR U13494 ( .A(n13122), .B(n13121), .Z(n13123) );
  XOR U13495 ( .A(n13404), .B(n13123), .Z(n13085) );
  AND U13496 ( .A(y[129]), .B(x[148]), .Z(n13117) );
  AND U13497 ( .A(y[8]), .B(x[125]), .Z(n13116) );
  XOR U13498 ( .A(n13117), .B(n13116), .Z(n13118) );
  AND U13499 ( .A(y[9]), .B(x[124]), .Z(n13392) );
  XOR U13500 ( .A(n13118), .B(n13392), .Z(n13084) );
  XOR U13501 ( .A(n13085), .B(n13084), .Z(n13087) );
  XOR U13502 ( .A(n13086), .B(n13087), .Z(n13078) );
  NANDN U13503 ( .A(n12999), .B(n12998), .Z(n13003) );
  NANDN U13504 ( .A(n13001), .B(n13000), .Z(n13002) );
  NAND U13505 ( .A(n13003), .B(n13002), .Z(n13200) );
  AND U13506 ( .A(y[170]), .B(x[155]), .Z(n13004) );
  AND U13507 ( .A(n13005), .B(n13004), .Z(n13164) );
  AND U13508 ( .A(x[152]), .B(y[173]), .Z(n13007) );
  AND U13509 ( .A(x[153]), .B(y[172]), .Z(n13006) );
  XOR U13510 ( .A(n13007), .B(n13006), .Z(n13163) );
  XOR U13511 ( .A(n13164), .B(n13163), .Z(n13199) );
  AND U13512 ( .A(y[53]), .B(x[128]), .Z(n13189) );
  AND U13513 ( .A(y[12]), .B(x[121]), .Z(n13188) );
  XOR U13514 ( .A(n13189), .B(n13188), .Z(n13191) );
  AND U13515 ( .A(y[49]), .B(x[132]), .Z(n13190) );
  XOR U13516 ( .A(n13191), .B(n13190), .Z(n13198) );
  XOR U13517 ( .A(n13199), .B(n13198), .Z(n13201) );
  XOR U13518 ( .A(n13200), .B(n13201), .Z(n13080) );
  XOR U13519 ( .A(n13081), .B(n13080), .Z(n13128) );
  XOR U13520 ( .A(n13129), .B(n13128), .Z(n13213) );
  AND U13521 ( .A(y[171]), .B(x[156]), .Z(n13418) );
  NAND U13522 ( .A(n13418), .B(n13008), .Z(n13012) );
  NAND U13523 ( .A(n13010), .B(n13009), .Z(n13011) );
  AND U13524 ( .A(n13012), .B(n13011), .Z(n13145) );
  NAND U13525 ( .A(n13016), .B(n13015), .Z(n13020) );
  NANDN U13526 ( .A(n13018), .B(n13017), .Z(n13019) );
  AND U13527 ( .A(n13020), .B(n13019), .Z(n13135) );
  AND U13528 ( .A(x[130]), .B(y[51]), .Z(n13022) );
  NAND U13529 ( .A(x[131]), .B(y[50]), .Z(n13021) );
  XNOR U13530 ( .A(n13022), .B(n13021), .Z(n13097) );
  NAND U13531 ( .A(y[52]), .B(x[129]), .Z(n13098) );
  AND U13532 ( .A(y[171]), .B(x[154]), .Z(n13090) );
  NAND U13533 ( .A(y[168]), .B(x[157]), .Z(n13091) );
  AND U13534 ( .A(y[169]), .B(x[156]), .Z(n13400) );
  NAND U13535 ( .A(x[155]), .B(y[170]), .Z(n13023) );
  XOR U13536 ( .A(n13400), .B(n13023), .Z(n13093) );
  XOR U13537 ( .A(n13133), .B(n13132), .Z(n13134) );
  XOR U13538 ( .A(n13135), .B(n13134), .Z(n13146) );
  XOR U13539 ( .A(n13147), .B(n13146), .Z(n13159) );
  AND U13540 ( .A(x[140]), .B(y[89]), .Z(n13025) );
  NAND U13541 ( .A(x[141]), .B(y[88]), .Z(n13024) );
  XOR U13542 ( .A(n13025), .B(n13024), .Z(n13109) );
  AND U13543 ( .A(y[128]), .B(x[149]), .Z(n13101) );
  NAND U13544 ( .A(y[10]), .B(x[123]), .Z(n13102) );
  AND U13545 ( .A(y[11]), .B(x[122]), .Z(n13103) );
  XOR U13546 ( .A(n13104), .B(n13103), .Z(n13180) );
  XOR U13547 ( .A(n13181), .B(n13180), .Z(n13183) );
  NAND U13548 ( .A(n13027), .B(n13026), .Z(n13031) );
  NANDN U13549 ( .A(n13029), .B(n13028), .Z(n13030) );
  AND U13550 ( .A(n13031), .B(n13030), .Z(n13182) );
  XOR U13551 ( .A(n13183), .B(n13182), .Z(n13157) );
  AND U13552 ( .A(y[52]), .B(x[131]), .Z(n13417) );
  NAND U13553 ( .A(n13417), .B(n13032), .Z(n13035) );
  NANDN U13554 ( .A(n13033), .B(n13096), .Z(n13034) );
  AND U13555 ( .A(n13035), .B(n13034), .Z(n13141) );
  AND U13556 ( .A(y[92]), .B(x[137]), .Z(n13338) );
  AND U13557 ( .A(y[130]), .B(x[147]), .Z(n13175) );
  XOR U13558 ( .A(n13338), .B(n13175), .Z(n13177) );
  AND U13559 ( .A(y[93]), .B(x[136]), .Z(n13176) );
  XOR U13560 ( .A(n13177), .B(n13176), .Z(n13139) );
  AND U13561 ( .A(y[13]), .B(x[120]), .Z(n13168) );
  AND U13562 ( .A(y[132]), .B(x[145]), .Z(n13167) );
  XOR U13563 ( .A(n13168), .B(n13167), .Z(n13170) );
  AND U13564 ( .A(y[131]), .B(x[146]), .Z(n13169) );
  XOR U13565 ( .A(n13170), .B(n13169), .Z(n13138) );
  XOR U13566 ( .A(n13139), .B(n13138), .Z(n13140) );
  XOR U13567 ( .A(n13141), .B(n13140), .Z(n13156) );
  NANDN U13568 ( .A(n13037), .B(n13036), .Z(n13041) );
  NAND U13569 ( .A(n13039), .B(n13038), .Z(n13040) );
  AND U13570 ( .A(n13041), .B(n13040), .Z(n13151) );
  NAND U13571 ( .A(n13043), .B(n13042), .Z(n13047) );
  NANDN U13572 ( .A(n13045), .B(n13044), .Z(n13046) );
  NAND U13573 ( .A(n13047), .B(n13046), .Z(n13150) );
  NANDN U13574 ( .A(n13049), .B(n13048), .Z(n13053) );
  NANDN U13575 ( .A(n13051), .B(n13050), .Z(n13052) );
  NAND U13576 ( .A(n13053), .B(n13052), .Z(n13153) );
  XOR U13577 ( .A(n13211), .B(n13210), .Z(n13212) );
  XOR U13578 ( .A(n13213), .B(n13212), .Z(n13072) );
  XNOR U13579 ( .A(n13073), .B(n13072), .Z(n13074) );
  NANDN U13580 ( .A(n13055), .B(n13054), .Z(n13059) );
  NANDN U13581 ( .A(n13057), .B(n13056), .Z(n13058) );
  AND U13582 ( .A(n13059), .B(n13058), .Z(n13207) );
  NANDN U13583 ( .A(n13061), .B(n13060), .Z(n13065) );
  NANDN U13584 ( .A(n13063), .B(n13062), .Z(n13064) );
  AND U13585 ( .A(n13065), .B(n13064), .Z(n13205) );
  NANDN U13586 ( .A(n13067), .B(n13066), .Z(n13071) );
  NAND U13587 ( .A(n13069), .B(n13068), .Z(n13070) );
  AND U13588 ( .A(n13071), .B(n13070), .Z(n13204) );
  XNOR U13589 ( .A(n13205), .B(n13204), .Z(n13206) );
  XOR U13590 ( .A(n13207), .B(n13206), .Z(n13075) );
  XNOR U13591 ( .A(n13074), .B(n13075), .Z(n13217) );
  XOR U13592 ( .A(n13218), .B(n13217), .Z(o[133]) );
  NANDN U13593 ( .A(n13073), .B(n13072), .Z(n13077) );
  NANDN U13594 ( .A(n13075), .B(n13074), .Z(n13076) );
  AND U13595 ( .A(n13077), .B(n13076), .Z(n13502) );
  NANDN U13596 ( .A(n13079), .B(n13078), .Z(n13083) );
  NAND U13597 ( .A(n13081), .B(n13080), .Z(n13082) );
  AND U13598 ( .A(n13083), .B(n13082), .Z(n13507) );
  NAND U13599 ( .A(n13085), .B(n13084), .Z(n13089) );
  NAND U13600 ( .A(n13087), .B(n13086), .Z(n13088) );
  NAND U13601 ( .A(n13089), .B(n13088), .Z(n13230) );
  NANDN U13602 ( .A(n13091), .B(n13090), .Z(n13095) );
  NANDN U13603 ( .A(n13093), .B(n13092), .Z(n13094) );
  NAND U13604 ( .A(n13095), .B(n13094), .Z(n13371) );
  AND U13605 ( .A(x[131]), .B(y[51]), .Z(n13187) );
  NAND U13606 ( .A(n13096), .B(n13187), .Z(n13100) );
  NANDN U13607 ( .A(n13098), .B(n13097), .Z(n13099) );
  AND U13608 ( .A(n13100), .B(n13099), .Z(n13465) );
  AND U13609 ( .A(y[131]), .B(x[147]), .Z(n13432) );
  AND U13610 ( .A(y[91]), .B(x[139]), .Z(n13431) );
  XOR U13611 ( .A(n13432), .B(n13431), .Z(n13430) );
  AND U13612 ( .A(y[11]), .B(x[123]), .Z(n13429) );
  XOR U13613 ( .A(n13430), .B(n13429), .Z(n13468) );
  AND U13614 ( .A(y[132]), .B(x[146]), .Z(n13426) );
  AND U13615 ( .A(y[90]), .B(x[140]), .Z(n13425) );
  XOR U13616 ( .A(n13426), .B(n13425), .Z(n13424) );
  AND U13617 ( .A(y[12]), .B(x[122]), .Z(n13423) );
  XNOR U13618 ( .A(n13424), .B(n13423), .Z(n13467) );
  XNOR U13619 ( .A(n13465), .B(n13466), .Z(n13374) );
  NANDN U13620 ( .A(n13102), .B(n13101), .Z(n13106) );
  NAND U13621 ( .A(n13104), .B(n13103), .Z(n13105) );
  NAND U13622 ( .A(n13106), .B(n13105), .Z(n13373) );
  XOR U13623 ( .A(n13371), .B(n13372), .Z(n13231) );
  XOR U13624 ( .A(n13230), .B(n13231), .Z(n13228) );
  AND U13625 ( .A(y[89]), .B(x[141]), .Z(n13352) );
  NANDN U13626 ( .A(n13107), .B(n13352), .Z(n13111) );
  NANDN U13627 ( .A(n13109), .B(n13108), .Z(n13110) );
  AND U13628 ( .A(n13111), .B(n13110), .Z(n13377) );
  AND U13629 ( .A(x[125]), .B(y[9]), .Z(n13113) );
  NAND U13630 ( .A(x[124]), .B(y[10]), .Z(n13112) );
  XNOR U13631 ( .A(n13113), .B(n13112), .Z(n13390) );
  AND U13632 ( .A(y[128]), .B(x[150]), .Z(n13389) );
  XOR U13633 ( .A(n13390), .B(n13389), .Z(n13380) );
  AND U13634 ( .A(y[173]), .B(x[153]), .Z(n13356) );
  AND U13635 ( .A(y[170]), .B(x[156]), .Z(n13114) );
  AND U13636 ( .A(n13115), .B(n13114), .Z(n13358) );
  AND U13637 ( .A(y[172]), .B(x[154]), .Z(n13357) );
  XOR U13638 ( .A(n13358), .B(n13357), .Z(n13355) );
  XNOR U13639 ( .A(n13356), .B(n13355), .Z(n13379) );
  XOR U13640 ( .A(n13377), .B(n13378), .Z(n13252) );
  NAND U13641 ( .A(n13117), .B(n13116), .Z(n13120) );
  NAND U13642 ( .A(n13118), .B(n13392), .Z(n13119) );
  NAND U13643 ( .A(n13120), .B(n13119), .Z(n13255) );
  NAND U13644 ( .A(n13122), .B(n13121), .Z(n13125) );
  NAND U13645 ( .A(n13404), .B(n13123), .Z(n13124) );
  NAND U13646 ( .A(n13125), .B(n13124), .Z(n13254) );
  XNOR U13647 ( .A(n13255), .B(n13254), .Z(n13253) );
  XNOR U13648 ( .A(n13228), .B(n13229), .Z(n13227) );
  NANDN U13649 ( .A(n13127), .B(n13126), .Z(n13131) );
  NAND U13650 ( .A(n13129), .B(n13128), .Z(n13130) );
  AND U13651 ( .A(n13131), .B(n13130), .Z(n13226) );
  NAND U13652 ( .A(n13133), .B(n13132), .Z(n13137) );
  NAND U13653 ( .A(n13135), .B(n13134), .Z(n13136) );
  AND U13654 ( .A(n13137), .B(n13136), .Z(n13233) );
  NAND U13655 ( .A(n13139), .B(n13138), .Z(n13143) );
  NANDN U13656 ( .A(n13141), .B(n13140), .Z(n13142) );
  AND U13657 ( .A(n13143), .B(n13142), .Z(n13235) );
  NANDN U13658 ( .A(n13145), .B(n13144), .Z(n13149) );
  NAND U13659 ( .A(n13147), .B(n13146), .Z(n13148) );
  AND U13660 ( .A(n13149), .B(n13148), .Z(n13234) );
  XOR U13661 ( .A(n13235), .B(n13234), .Z(n13232) );
  XOR U13662 ( .A(n13233), .B(n13232), .Z(n13224) );
  XOR U13663 ( .A(n13225), .B(n13224), .Z(n13506) );
  XOR U13664 ( .A(n13507), .B(n13506), .Z(n13509) );
  NANDN U13665 ( .A(n13151), .B(n13150), .Z(n13155) );
  NANDN U13666 ( .A(n13153), .B(n13152), .Z(n13154) );
  AND U13667 ( .A(n13155), .B(n13154), .Z(n13486) );
  NANDN U13668 ( .A(n13157), .B(n13156), .Z(n13161) );
  NANDN U13669 ( .A(n13159), .B(n13158), .Z(n13160) );
  NAND U13670 ( .A(n13161), .B(n13160), .Z(n13487) );
  NANDN U13671 ( .A(n13162), .B(n13356), .Z(n13166) );
  NAND U13672 ( .A(n13164), .B(n13163), .Z(n13165) );
  NAND U13673 ( .A(n13166), .B(n13165), .Z(n13247) );
  NAND U13674 ( .A(n13168), .B(n13167), .Z(n13172) );
  NAND U13675 ( .A(n13170), .B(n13169), .Z(n13171) );
  AND U13676 ( .A(n13172), .B(n13171), .Z(n13460) );
  AND U13677 ( .A(y[13]), .B(x[121]), .Z(n13446) );
  AND U13678 ( .A(y[48]), .B(x[134]), .Z(n13445) );
  XOR U13679 ( .A(n13446), .B(n13445), .Z(n13444) );
  AND U13680 ( .A(y[54]), .B(x[128]), .Z(n13443) );
  XOR U13681 ( .A(n13444), .B(n13443), .Z(n13462) );
  AND U13682 ( .A(x[157]), .B(y[169]), .Z(n13174) );
  NAND U13683 ( .A(x[156]), .B(y[170]), .Z(n13173) );
  XNOR U13684 ( .A(n13174), .B(n13173), .Z(n13267) );
  AND U13685 ( .A(y[168]), .B(x[158]), .Z(n13266) );
  XOR U13686 ( .A(n13267), .B(n13266), .Z(n13264) );
  XNOR U13687 ( .A(n13265), .B(n13264), .Z(n13461) );
  XNOR U13688 ( .A(n13460), .B(n13459), .Z(n13246) );
  XOR U13689 ( .A(n13247), .B(n13246), .Z(n13245) );
  AND U13690 ( .A(n13338), .B(n13175), .Z(n13179) );
  NAND U13691 ( .A(n13177), .B(n13176), .Z(n13178) );
  NANDN U13692 ( .A(n13179), .B(n13178), .Z(n13244) );
  XOR U13693 ( .A(n13245), .B(n13244), .Z(n13493) );
  NAND U13694 ( .A(n13181), .B(n13180), .Z(n13185) );
  NAND U13695 ( .A(n13183), .B(n13182), .Z(n13184) );
  AND U13696 ( .A(n13185), .B(n13184), .Z(n13492) );
  AND U13697 ( .A(y[94]), .B(x[136]), .Z(n13386) );
  AND U13698 ( .A(y[8]), .B(x[126]), .Z(n13385) );
  XOR U13699 ( .A(n13386), .B(n13385), .Z(n13384) );
  AND U13700 ( .A(y[129]), .B(x[149]), .Z(n13383) );
  XOR U13701 ( .A(n13384), .B(n13383), .Z(n13261) );
  AND U13702 ( .A(y[49]), .B(x[133]), .Z(n13440) );
  AND U13703 ( .A(y[52]), .B(x[130]), .Z(n13439) );
  XOR U13704 ( .A(n13440), .B(n13439), .Z(n13438) );
  AND U13705 ( .A(y[53]), .B(x[129]), .Z(n13437) );
  XOR U13706 ( .A(n13438), .B(n13437), .Z(n13342) );
  NAND U13707 ( .A(x[132]), .B(y[50]), .Z(n13186) );
  XNOR U13708 ( .A(n13187), .B(n13186), .Z(n13341) );
  XOR U13709 ( .A(n13342), .B(n13341), .Z(n13260) );
  XOR U13710 ( .A(n13261), .B(n13260), .Z(n13259) );
  AND U13711 ( .A(y[174]), .B(x[152]), .Z(n13351) );
  XOR U13712 ( .A(n13352), .B(n13351), .Z(n13350) );
  AND U13713 ( .A(y[88]), .B(x[142]), .Z(n13349) );
  XOR U13714 ( .A(n13350), .B(n13349), .Z(n13258) );
  XOR U13715 ( .A(n13259), .B(n13258), .Z(n13241) );
  NAND U13716 ( .A(n13189), .B(n13188), .Z(n13193) );
  NAND U13717 ( .A(n13191), .B(n13190), .Z(n13192) );
  AND U13718 ( .A(n13193), .B(n13192), .Z(n13329) );
  AND U13719 ( .A(y[130]), .B(x[148]), .Z(n13336) );
  AND U13720 ( .A(x[137]), .B(y[93]), .Z(n13195) );
  AND U13721 ( .A(x[138]), .B(y[92]), .Z(n13194) );
  XOR U13722 ( .A(n13195), .B(n13194), .Z(n13335) );
  XOR U13723 ( .A(n13336), .B(n13335), .Z(n13332) );
  AND U13724 ( .A(y[14]), .B(x[120]), .Z(n13402) );
  AND U13725 ( .A(y[134]), .B(x[144]), .Z(n13197) );
  AND U13726 ( .A(x[145]), .B(y[133]), .Z(n13196) );
  XOR U13727 ( .A(n13197), .B(n13196), .Z(n13401) );
  XNOR U13728 ( .A(n13402), .B(n13401), .Z(n13331) );
  XNOR U13729 ( .A(n13329), .B(n13330), .Z(n13240) );
  NAND U13730 ( .A(n13199), .B(n13198), .Z(n13203) );
  NAND U13731 ( .A(n13201), .B(n13200), .Z(n13202) );
  AND U13732 ( .A(n13203), .B(n13202), .Z(n13238) );
  XOR U13733 ( .A(n13239), .B(n13238), .Z(n13491) );
  XOR U13734 ( .A(n13492), .B(n13491), .Z(n13494) );
  XOR U13735 ( .A(n13487), .B(n13488), .Z(n13485) );
  XOR U13736 ( .A(n13486), .B(n13485), .Z(n13508) );
  XOR U13737 ( .A(n13509), .B(n13508), .Z(n13223) );
  NANDN U13738 ( .A(n13205), .B(n13204), .Z(n13209) );
  NANDN U13739 ( .A(n13207), .B(n13206), .Z(n13208) );
  AND U13740 ( .A(n13209), .B(n13208), .Z(n13222) );
  XOR U13741 ( .A(n13222), .B(n13221), .Z(n13214) );
  XOR U13742 ( .A(n13223), .B(n13214), .Z(n13503) );
  NANDN U13743 ( .A(n13216), .B(n13215), .Z(n13220) );
  NAND U13744 ( .A(n13218), .B(n13217), .Z(n13219) );
  NAND U13745 ( .A(n13220), .B(n13219), .Z(n13500) );
  XOR U13746 ( .A(n13501), .B(n13500), .Z(o[134]) );
  NAND U13747 ( .A(n13233), .B(n13232), .Z(n13237) );
  NAND U13748 ( .A(n13235), .B(n13234), .Z(n13236) );
  AND U13749 ( .A(n13237), .B(n13236), .Z(n13484) );
  NAND U13750 ( .A(n13239), .B(n13238), .Z(n13243) );
  NANDN U13751 ( .A(n13241), .B(n13240), .Z(n13242) );
  AND U13752 ( .A(n13243), .B(n13242), .Z(n13251) );
  NAND U13753 ( .A(n13245), .B(n13244), .Z(n13249) );
  NAND U13754 ( .A(n13247), .B(n13246), .Z(n13248) );
  NAND U13755 ( .A(n13249), .B(n13248), .Z(n13250) );
  XNOR U13756 ( .A(n13251), .B(n13250), .Z(n13482) );
  NANDN U13757 ( .A(n13253), .B(n13252), .Z(n13257) );
  NAND U13758 ( .A(n13255), .B(n13254), .Z(n13256) );
  AND U13759 ( .A(n13257), .B(n13256), .Z(n13480) );
  NAND U13760 ( .A(n13259), .B(n13258), .Z(n13263) );
  NAND U13761 ( .A(n13261), .B(n13260), .Z(n13262) );
  AND U13762 ( .A(n13263), .B(n13262), .Z(n13370) );
  NAND U13763 ( .A(n13265), .B(n13264), .Z(n13269) );
  NAND U13764 ( .A(n13267), .B(n13266), .Z(n13268) );
  AND U13765 ( .A(n13269), .B(n13268), .Z(n13328) );
  AND U13766 ( .A(x[148]), .B(y[131]), .Z(n13271) );
  NAND U13767 ( .A(x[126]), .B(y[9]), .Z(n13270) );
  XNOR U13768 ( .A(n13271), .B(n13270), .Z(n13275) );
  AND U13769 ( .A(x[127]), .B(y[8]), .Z(n13273) );
  NAND U13770 ( .A(x[159]), .B(y[168]), .Z(n13272) );
  XNOR U13771 ( .A(n13273), .B(n13272), .Z(n13274) );
  XOR U13772 ( .A(n13275), .B(n13274), .Z(n13283) );
  AND U13773 ( .A(x[137]), .B(y[94]), .Z(n13277) );
  NAND U13774 ( .A(x[135]), .B(y[48]), .Z(n13276) );
  XNOR U13775 ( .A(n13277), .B(n13276), .Z(n13281) );
  AND U13776 ( .A(x[136]), .B(y[95]), .Z(n13279) );
  NAND U13777 ( .A(x[147]), .B(y[132]), .Z(n13278) );
  XNOR U13778 ( .A(n13279), .B(n13278), .Z(n13280) );
  XNOR U13779 ( .A(n13281), .B(n13280), .Z(n13282) );
  XNOR U13780 ( .A(n13283), .B(n13282), .Z(n13326) );
  AND U13781 ( .A(x[155]), .B(y[172]), .Z(n13288) );
  AND U13782 ( .A(y[10]), .B(x[125]), .Z(n13391) );
  AND U13783 ( .A(x[154]), .B(y[173]), .Z(n13285) );
  NAND U13784 ( .A(x[133]), .B(y[50]), .Z(n13284) );
  XNOR U13785 ( .A(n13285), .B(n13284), .Z(n13286) );
  XNOR U13786 ( .A(n13391), .B(n13286), .Z(n13287) );
  XNOR U13787 ( .A(n13288), .B(n13287), .Z(n13304) );
  AND U13788 ( .A(x[140]), .B(y[91]), .Z(n13290) );
  NAND U13789 ( .A(x[139]), .B(y[92]), .Z(n13289) );
  XNOR U13790 ( .A(n13290), .B(n13289), .Z(n13294) );
  AND U13791 ( .A(x[144]), .B(y[135]), .Z(n13292) );
  NAND U13792 ( .A(x[129]), .B(y[54]), .Z(n13291) );
  XNOR U13793 ( .A(n13292), .B(n13291), .Z(n13293) );
  XOR U13794 ( .A(n13294), .B(n13293), .Z(n13302) );
  AND U13795 ( .A(x[121]), .B(y[14]), .Z(n13296) );
  NAND U13796 ( .A(x[141]), .B(y[90]), .Z(n13295) );
  XNOR U13797 ( .A(n13296), .B(n13295), .Z(n13300) );
  AND U13798 ( .A(x[124]), .B(y[11]), .Z(n13298) );
  NAND U13799 ( .A(x[149]), .B(y[130]), .Z(n13297) );
  XNOR U13800 ( .A(n13298), .B(n13297), .Z(n13299) );
  XNOR U13801 ( .A(n13300), .B(n13299), .Z(n13301) );
  XNOR U13802 ( .A(n13302), .B(n13301), .Z(n13303) );
  XOR U13803 ( .A(n13304), .B(n13303), .Z(n13324) );
  AND U13804 ( .A(x[120]), .B(y[15]), .Z(n13306) );
  NAND U13805 ( .A(x[153]), .B(y[174]), .Z(n13305) );
  XNOR U13806 ( .A(n13306), .B(n13305), .Z(n13310) );
  AND U13807 ( .A(x[122]), .B(y[13]), .Z(n13308) );
  NAND U13808 ( .A(x[150]), .B(y[129]), .Z(n13307) );
  XNOR U13809 ( .A(n13308), .B(n13307), .Z(n13309) );
  XOR U13810 ( .A(n13310), .B(n13309), .Z(n13318) );
  AND U13811 ( .A(x[123]), .B(y[12]), .Z(n13312) );
  NAND U13812 ( .A(x[134]), .B(y[49]), .Z(n13311) );
  XNOR U13813 ( .A(n13312), .B(n13311), .Z(n13316) );
  AND U13814 ( .A(x[152]), .B(y[175]), .Z(n13314) );
  NAND U13815 ( .A(x[143]), .B(y[88]), .Z(n13313) );
  XNOR U13816 ( .A(n13314), .B(n13313), .Z(n13315) );
  XNOR U13817 ( .A(n13316), .B(n13315), .Z(n13317) );
  XNOR U13818 ( .A(n13318), .B(n13317), .Z(n13322) );
  AND U13819 ( .A(y[93]), .B(x[138]), .Z(n13337) );
  AND U13820 ( .A(y[134]), .B(x[145]), .Z(n13403) );
  XOR U13821 ( .A(n13337), .B(n13403), .Z(n13320) );
  AND U13822 ( .A(y[170]), .B(x[157]), .Z(n13399) );
  AND U13823 ( .A(y[51]), .B(x[132]), .Z(n13343) );
  XNOR U13824 ( .A(n13399), .B(n13343), .Z(n13319) );
  XNOR U13825 ( .A(n13320), .B(n13319), .Z(n13321) );
  XNOR U13826 ( .A(n13322), .B(n13321), .Z(n13323) );
  XNOR U13827 ( .A(n13324), .B(n13323), .Z(n13325) );
  XNOR U13828 ( .A(n13326), .B(n13325), .Z(n13327) );
  XNOR U13829 ( .A(n13328), .B(n13327), .Z(n13368) );
  NANDN U13830 ( .A(n13330), .B(n13329), .Z(n13334) );
  NANDN U13831 ( .A(n13332), .B(n13331), .Z(n13333) );
  AND U13832 ( .A(n13334), .B(n13333), .Z(n13366) );
  NAND U13833 ( .A(n13336), .B(n13335), .Z(n13340) );
  NAND U13834 ( .A(n13338), .B(n13337), .Z(n13339) );
  AND U13835 ( .A(n13340), .B(n13339), .Z(n13348) );
  NAND U13836 ( .A(n13342), .B(n13341), .Z(n13346) );
  AND U13837 ( .A(y[50]), .B(x[131]), .Z(n13344) );
  NAND U13838 ( .A(n13344), .B(n13343), .Z(n13345) );
  NAND U13839 ( .A(n13346), .B(n13345), .Z(n13347) );
  XNOR U13840 ( .A(n13348), .B(n13347), .Z(n13364) );
  NAND U13841 ( .A(n13350), .B(n13349), .Z(n13354) );
  NAND U13842 ( .A(n13352), .B(n13351), .Z(n13353) );
  AND U13843 ( .A(n13354), .B(n13353), .Z(n13362) );
  NAND U13844 ( .A(n13356), .B(n13355), .Z(n13360) );
  NAND U13845 ( .A(n13358), .B(n13357), .Z(n13359) );
  NAND U13846 ( .A(n13360), .B(n13359), .Z(n13361) );
  XNOR U13847 ( .A(n13362), .B(n13361), .Z(n13363) );
  XNOR U13848 ( .A(n13364), .B(n13363), .Z(n13365) );
  XNOR U13849 ( .A(n13366), .B(n13365), .Z(n13367) );
  XNOR U13850 ( .A(n13368), .B(n13367), .Z(n13369) );
  XNOR U13851 ( .A(n13370), .B(n13369), .Z(n13478) );
  NAND U13852 ( .A(n13372), .B(n13371), .Z(n13376) );
  NANDN U13853 ( .A(n13374), .B(n13373), .Z(n13375) );
  AND U13854 ( .A(n13376), .B(n13375), .Z(n13476) );
  NANDN U13855 ( .A(n13378), .B(n13377), .Z(n13382) );
  NANDN U13856 ( .A(n13380), .B(n13379), .Z(n13381) );
  AND U13857 ( .A(n13382), .B(n13381), .Z(n13458) );
  NAND U13858 ( .A(n13384), .B(n13383), .Z(n13388) );
  NAND U13859 ( .A(n13386), .B(n13385), .Z(n13387) );
  AND U13860 ( .A(n13388), .B(n13387), .Z(n13396) );
  NAND U13861 ( .A(n13390), .B(n13389), .Z(n13394) );
  NAND U13862 ( .A(n13392), .B(n13391), .Z(n13393) );
  NAND U13863 ( .A(n13394), .B(n13393), .Z(n13395) );
  XNOR U13864 ( .A(n13396), .B(n13395), .Z(n13456) );
  AND U13865 ( .A(x[130]), .B(y[53]), .Z(n13398) );
  NAND U13866 ( .A(x[146]), .B(y[133]), .Z(n13397) );
  XNOR U13867 ( .A(n13398), .B(n13397), .Z(n13422) );
  AND U13868 ( .A(n13400), .B(n13399), .Z(n13416) );
  NAND U13869 ( .A(n13402), .B(n13401), .Z(n13406) );
  NAND U13870 ( .A(n13404), .B(n13403), .Z(n13405) );
  AND U13871 ( .A(n13406), .B(n13405), .Z(n13414) );
  AND U13872 ( .A(x[128]), .B(y[55]), .Z(n13408) );
  NAND U13873 ( .A(x[158]), .B(y[169]), .Z(n13407) );
  XNOR U13874 ( .A(n13408), .B(n13407), .Z(n13412) );
  AND U13875 ( .A(x[151]), .B(y[128]), .Z(n13410) );
  NAND U13876 ( .A(x[142]), .B(y[89]), .Z(n13409) );
  XNOR U13877 ( .A(n13410), .B(n13409), .Z(n13411) );
  XNOR U13878 ( .A(n13412), .B(n13411), .Z(n13413) );
  XNOR U13879 ( .A(n13414), .B(n13413), .Z(n13415) );
  XOR U13880 ( .A(n13416), .B(n13415), .Z(n13420) );
  XNOR U13881 ( .A(n13418), .B(n13417), .Z(n13419) );
  XNOR U13882 ( .A(n13420), .B(n13419), .Z(n13421) );
  XOR U13883 ( .A(n13422), .B(n13421), .Z(n13454) );
  NAND U13884 ( .A(n13424), .B(n13423), .Z(n13428) );
  NAND U13885 ( .A(n13426), .B(n13425), .Z(n13427) );
  AND U13886 ( .A(n13428), .B(n13427), .Z(n13436) );
  NAND U13887 ( .A(n13430), .B(n13429), .Z(n13434) );
  NAND U13888 ( .A(n13432), .B(n13431), .Z(n13433) );
  NAND U13889 ( .A(n13434), .B(n13433), .Z(n13435) );
  XNOR U13890 ( .A(n13436), .B(n13435), .Z(n13452) );
  NAND U13891 ( .A(n13438), .B(n13437), .Z(n13442) );
  NAND U13892 ( .A(n13440), .B(n13439), .Z(n13441) );
  AND U13893 ( .A(n13442), .B(n13441), .Z(n13450) );
  NAND U13894 ( .A(n13444), .B(n13443), .Z(n13448) );
  NAND U13895 ( .A(n13446), .B(n13445), .Z(n13447) );
  NAND U13896 ( .A(n13448), .B(n13447), .Z(n13449) );
  XNOR U13897 ( .A(n13450), .B(n13449), .Z(n13451) );
  XNOR U13898 ( .A(n13452), .B(n13451), .Z(n13453) );
  XNOR U13899 ( .A(n13454), .B(n13453), .Z(n13455) );
  XNOR U13900 ( .A(n13456), .B(n13455), .Z(n13457) );
  XNOR U13901 ( .A(n13458), .B(n13457), .Z(n13474) );
  NAND U13902 ( .A(n13460), .B(n13459), .Z(n13464) );
  NANDN U13903 ( .A(n13462), .B(n13461), .Z(n13463) );
  AND U13904 ( .A(n13464), .B(n13463), .Z(n13472) );
  NANDN U13905 ( .A(n13466), .B(n13465), .Z(n13470) );
  NANDN U13906 ( .A(n13468), .B(n13467), .Z(n13469) );
  NAND U13907 ( .A(n13470), .B(n13469), .Z(n13471) );
  XNOR U13908 ( .A(n13472), .B(n13471), .Z(n13473) );
  XNOR U13909 ( .A(n13474), .B(n13473), .Z(n13475) );
  XNOR U13910 ( .A(n13476), .B(n13475), .Z(n13477) );
  XNOR U13911 ( .A(n13478), .B(n13477), .Z(n13479) );
  XNOR U13912 ( .A(n13480), .B(n13479), .Z(n13481) );
  XNOR U13913 ( .A(n13482), .B(n13481), .Z(n13483) );
  NAND U13914 ( .A(n13486), .B(n13485), .Z(n13490) );
  AND U13915 ( .A(n13488), .B(n13487), .Z(n13489) );
  ANDN U13916 ( .B(n13490), .A(n13489), .Z(n13498) );
  AND U13917 ( .A(n13492), .B(n13491), .Z(n13496) );
  ANDN U13918 ( .B(n13494), .A(n13493), .Z(n13495) );
  OR U13919 ( .A(n13496), .B(n13495), .Z(n13497) );
  XNOR U13920 ( .A(n13498), .B(n13497), .Z(n13499) );
  NAND U13921 ( .A(n13501), .B(n13500), .Z(n13505) );
  ANDN U13922 ( .B(n13503), .A(n13502), .Z(n13504) );
  AND U13923 ( .A(n13507), .B(n13506), .Z(n13511) );
  AND U13924 ( .A(n13509), .B(n13508), .Z(n13510) );
  AND U13925 ( .A(y[176]), .B(x[152]), .Z(n13515) );
  IV U13926 ( .A(n13515), .Z(n13628) );
  NAND U13927 ( .A(y[56]), .B(x[128]), .Z(n13514) );
  XOR U13928 ( .A(n13628), .B(n13514), .Z(n13516) );
  AND U13929 ( .A(y[16]), .B(x[120]), .Z(n13525) );
  AND U13930 ( .A(y[96]), .B(x[136]), .Z(n13522) );
  XOR U13931 ( .A(n13525), .B(n13522), .Z(n13521) );
  AND U13932 ( .A(y[136]), .B(x[144]), .Z(n13520) );
  XNOR U13933 ( .A(n13521), .B(n13520), .Z(n13517) );
  XNOR U13934 ( .A(n13516), .B(n13517), .Z(o[136]) );
  AND U13935 ( .A(x[121]), .B(y[16]), .Z(n13513) );
  NAND U13936 ( .A(x[120]), .B(y[17]), .Z(n13512) );
  XNOR U13937 ( .A(n13513), .B(n13512), .Z(n13527) );
  AND U13938 ( .A(y[56]), .B(x[129]), .Z(n13526) );
  XNOR U13939 ( .A(n13527), .B(n13526), .Z(n13542) );
  AND U13940 ( .A(y[176]), .B(x[153]), .Z(n13738) );
  AND U13941 ( .A(y[97]), .B(x[136]), .Z(n13530) );
  XOR U13942 ( .A(n13738), .B(n13530), .Z(n13532) );
  AND U13943 ( .A(y[177]), .B(x[152]), .Z(n13551) );
  AND U13944 ( .A(y[96]), .B(x[137]), .Z(n13550) );
  XOR U13945 ( .A(n13551), .B(n13550), .Z(n13531) );
  XNOR U13946 ( .A(n13532), .B(n13531), .Z(n13540) );
  AND U13947 ( .A(y[57]), .B(x[128]), .Z(n13762) );
  AND U13948 ( .A(y[137]), .B(x[144]), .Z(n13547) );
  XOR U13949 ( .A(n13762), .B(n13547), .Z(n13546) );
  AND U13950 ( .A(y[136]), .B(x[145]), .Z(n13545) );
  XNOR U13951 ( .A(n13546), .B(n13545), .Z(n13539) );
  XOR U13952 ( .A(n13540), .B(n13539), .Z(n13541) );
  XOR U13953 ( .A(n13542), .B(n13541), .Z(n13536) );
  NANDN U13954 ( .A(n13515), .B(n13514), .Z(n13519) );
  NAND U13955 ( .A(n13517), .B(n13516), .Z(n13518) );
  AND U13956 ( .A(n13519), .B(n13518), .Z(n13534) );
  NAND U13957 ( .A(n13521), .B(n13520), .Z(n13524) );
  AND U13958 ( .A(n13525), .B(n13522), .Z(n13523) );
  ANDN U13959 ( .B(n13524), .A(n13523), .Z(n13533) );
  XNOR U13960 ( .A(n13534), .B(n13533), .Z(n13535) );
  XNOR U13961 ( .A(n13536), .B(n13535), .Z(o[137]) );
  AND U13962 ( .A(y[17]), .B(x[121]), .Z(n13568) );
  NAND U13963 ( .A(n13568), .B(n13525), .Z(n13529) );
  NAND U13964 ( .A(n13527), .B(n13526), .Z(n13528) );
  NAND U13965 ( .A(n13529), .B(n13528), .Z(n13596) );
  AND U13966 ( .A(y[138]), .B(x[144]), .Z(n13599) );
  AND U13967 ( .A(y[18]), .B(x[120]), .Z(n13600) );
  XOR U13968 ( .A(n13599), .B(n13600), .Z(n13601) );
  AND U13969 ( .A(y[56]), .B(x[130]), .Z(n13602) );
  XOR U13970 ( .A(n13601), .B(n13602), .Z(n13593) );
  XOR U13971 ( .A(n13594), .B(n13593), .Z(n13595) );
  XNOR U13972 ( .A(n13596), .B(n13595), .Z(n13588) );
  NANDN U13973 ( .A(n13534), .B(n13533), .Z(n13538) );
  NAND U13974 ( .A(n13536), .B(n13535), .Z(n13537) );
  NAND U13975 ( .A(n13538), .B(n13537), .Z(n13587) );
  XOR U13976 ( .A(n13588), .B(n13587), .Z(n13590) );
  NAND U13977 ( .A(n13540), .B(n13539), .Z(n13544) );
  NAND U13978 ( .A(n13542), .B(n13541), .Z(n13543) );
  AND U13979 ( .A(n13544), .B(n13543), .Z(n13556) );
  AND U13980 ( .A(y[16]), .B(x[122]), .Z(n13565) );
  AND U13981 ( .A(y[98]), .B(x[136]), .Z(n13566) );
  XOR U13982 ( .A(n13565), .B(n13566), .Z(n13567) );
  XOR U13983 ( .A(n13568), .B(n13567), .Z(n13610) );
  AND U13984 ( .A(y[136]), .B(x[146]), .Z(n13609) );
  XOR U13985 ( .A(n13610), .B(n13609), .Z(n13612) );
  AND U13986 ( .A(y[96]), .B(x[138]), .Z(n13654) );
  AND U13987 ( .A(y[178]), .B(x[152]), .Z(n13579) );
  XOR U13988 ( .A(n13654), .B(n13579), .Z(n13581) );
  AND U13989 ( .A(y[97]), .B(x[137]), .Z(n13580) );
  XOR U13990 ( .A(n13581), .B(n13580), .Z(n13611) );
  XOR U13991 ( .A(n13612), .B(n13611), .Z(n13554) );
  AND U13992 ( .A(n13546), .B(n13545), .Z(n13549) );
  NAND U13993 ( .A(n13762), .B(n13547), .Z(n13548) );
  NANDN U13994 ( .A(n13549), .B(n13548), .Z(n13562) );
  AND U13995 ( .A(n13551), .B(n13550), .Z(n13606) );
  AND U13996 ( .A(x[154]), .B(y[176]), .Z(n13552) );
  AND U13997 ( .A(x[153]), .B(y[177]), .Z(n13633) );
  XOR U13998 ( .A(n13552), .B(n13633), .Z(n13605) );
  XOR U13999 ( .A(n13606), .B(n13605), .Z(n13559) );
  AND U14000 ( .A(y[137]), .B(x[145]), .Z(n13571) );
  NAND U14001 ( .A(y[57]), .B(x[129]), .Z(n13572) );
  XNOR U14002 ( .A(n13571), .B(n13572), .Z(n13573) );
  NAND U14003 ( .A(y[58]), .B(x[128]), .Z(n13574) );
  XNOR U14004 ( .A(n13573), .B(n13574), .Z(n13560) );
  XOR U14005 ( .A(n13559), .B(n13560), .Z(n13561) );
  XOR U14006 ( .A(n13562), .B(n13561), .Z(n13553) );
  XOR U14007 ( .A(n13554), .B(n13553), .Z(n13555) );
  XNOR U14008 ( .A(n13556), .B(n13555), .Z(n13589) );
  XNOR U14009 ( .A(n13590), .B(n13589), .Z(o[138]) );
  NAND U14010 ( .A(n13554), .B(n13553), .Z(n13558) );
  NAND U14011 ( .A(n13556), .B(n13555), .Z(n13557) );
  NAND U14012 ( .A(n13558), .B(n13557), .Z(n13676) );
  NAND U14013 ( .A(n13560), .B(n13559), .Z(n13564) );
  NAND U14014 ( .A(n13562), .B(n13561), .Z(n13563) );
  NAND U14015 ( .A(n13564), .B(n13563), .Z(n13674) );
  NAND U14016 ( .A(n13566), .B(n13565), .Z(n13570) );
  NAND U14017 ( .A(n13568), .B(n13567), .Z(n13569) );
  NAND U14018 ( .A(n13570), .B(n13569), .Z(n13685) );
  NANDN U14019 ( .A(n13572), .B(n13571), .Z(n13576) );
  NANDN U14020 ( .A(n13574), .B(n13573), .Z(n13575) );
  NAND U14021 ( .A(n13576), .B(n13575), .Z(n13646) );
  NAND U14022 ( .A(y[139]), .B(x[144]), .Z(n13668) );
  NAND U14023 ( .A(y[99]), .B(x[136]), .Z(n13666) );
  NAND U14024 ( .A(y[16]), .B(x[123]), .Z(n13667) );
  XOR U14025 ( .A(n13666), .B(n13667), .Z(n13669) );
  XOR U14026 ( .A(n13668), .B(n13669), .Z(n13645) );
  AND U14027 ( .A(x[139]), .B(y[96]), .Z(n13578) );
  NAND U14028 ( .A(x[138]), .B(y[97]), .Z(n13577) );
  XNOR U14029 ( .A(n13578), .B(n13577), .Z(n13656) );
  AND U14030 ( .A(y[98]), .B(x[137]), .Z(n13655) );
  XOR U14031 ( .A(n13656), .B(n13655), .Z(n13644) );
  XNOR U14032 ( .A(n13645), .B(n13644), .Z(n13647) );
  XOR U14033 ( .A(n13646), .B(n13647), .Z(n13686) );
  XOR U14034 ( .A(n13685), .B(n13686), .Z(n13687) );
  AND U14035 ( .A(n13654), .B(n13579), .Z(n13583) );
  NAND U14036 ( .A(n13581), .B(n13580), .Z(n13582) );
  NANDN U14037 ( .A(n13583), .B(n13582), .Z(n13650) );
  NAND U14038 ( .A(y[18]), .B(x[121]), .Z(n13626) );
  NAND U14039 ( .A(y[17]), .B(x[122]), .Z(n13624) );
  NAND U14040 ( .A(y[138]), .B(x[145]), .Z(n13625) );
  XOR U14041 ( .A(n13624), .B(n13625), .Z(n13627) );
  XOR U14042 ( .A(n13626), .B(n13627), .Z(n13649) );
  AND U14043 ( .A(x[155]), .B(y[176]), .Z(n13585) );
  NAND U14044 ( .A(x[152]), .B(y[179]), .Z(n13584) );
  XNOR U14045 ( .A(n13585), .B(n13584), .Z(n13630) );
  AND U14046 ( .A(x[154]), .B(y[177]), .Z(n13734) );
  NAND U14047 ( .A(x[153]), .B(y[178]), .Z(n13586) );
  XNOR U14048 ( .A(n13734), .B(n13586), .Z(n13629) );
  XOR U14049 ( .A(n13630), .B(n13629), .Z(n13648) );
  XOR U14050 ( .A(n13649), .B(n13648), .Z(n13651) );
  XNOR U14051 ( .A(n13650), .B(n13651), .Z(n13688) );
  XOR U14052 ( .A(n13687), .B(n13688), .Z(n13673) );
  XOR U14053 ( .A(n13674), .B(n13673), .Z(n13675) );
  XNOR U14054 ( .A(n13676), .B(n13675), .Z(n13671) );
  NAND U14055 ( .A(n13588), .B(n13587), .Z(n13592) );
  NAND U14056 ( .A(n13590), .B(n13589), .Z(n13591) );
  AND U14057 ( .A(n13592), .B(n13591), .Z(n13670) );
  NAND U14058 ( .A(n13594), .B(n13593), .Z(n13598) );
  NAND U14059 ( .A(n13596), .B(n13595), .Z(n13597) );
  AND U14060 ( .A(n13598), .B(n13597), .Z(n13682) );
  NAND U14061 ( .A(n13600), .B(n13599), .Z(n13604) );
  NAND U14062 ( .A(n13602), .B(n13601), .Z(n13603) );
  NAND U14063 ( .A(n13604), .B(n13603), .Z(n13617) );
  AND U14064 ( .A(n13606), .B(n13605), .Z(n13608) );
  NAND U14065 ( .A(n13734), .B(n13738), .Z(n13607) );
  NANDN U14066 ( .A(n13608), .B(n13607), .Z(n13616) );
  XOR U14067 ( .A(n13617), .B(n13616), .Z(n13619) );
  NAND U14068 ( .A(y[56]), .B(x[131]), .Z(n13661) );
  NAND U14069 ( .A(y[19]), .B(x[120]), .Z(n13659) );
  NAND U14070 ( .A(y[137]), .B(x[146]), .Z(n13660) );
  XOR U14071 ( .A(n13659), .B(n13660), .Z(n13662) );
  XOR U14072 ( .A(n13661), .B(n13662), .Z(n13641) );
  NAND U14073 ( .A(y[59]), .B(x[128]), .Z(n13636) );
  NAND U14074 ( .A(y[57]), .B(x[130]), .Z(n13634) );
  NAND U14075 ( .A(y[136]), .B(x[147]), .Z(n13635) );
  XOR U14076 ( .A(n13634), .B(n13635), .Z(n13637) );
  XOR U14077 ( .A(n13636), .B(n13637), .Z(n13639) );
  AND U14078 ( .A(y[58]), .B(x[129]), .Z(n13638) );
  XNOR U14079 ( .A(n13639), .B(n13638), .Z(n13640) );
  XNOR U14080 ( .A(n13641), .B(n13640), .Z(n13618) );
  XNOR U14081 ( .A(n13619), .B(n13618), .Z(n13680) );
  NAND U14082 ( .A(n13610), .B(n13609), .Z(n13614) );
  NAND U14083 ( .A(n13612), .B(n13611), .Z(n13613) );
  AND U14084 ( .A(n13614), .B(n13613), .Z(n13679) );
  XOR U14085 ( .A(n13680), .B(n13679), .Z(n13681) );
  XOR U14086 ( .A(n13682), .B(n13681), .Z(n13672) );
  XNOR U14087 ( .A(n13670), .B(n13672), .Z(n13615) );
  XNOR U14088 ( .A(n13671), .B(n13615), .Z(o[139]) );
  NAND U14089 ( .A(n13617), .B(n13616), .Z(n13621) );
  NAND U14090 ( .A(n13619), .B(n13618), .Z(n13620) );
  NAND U14091 ( .A(n13621), .B(n13620), .Z(n13706) );
  AND U14092 ( .A(y[58]), .B(x[130]), .Z(n13804) );
  AND U14093 ( .A(y[60]), .B(x[128]), .Z(n13623) );
  AND U14094 ( .A(x[131]), .B(y[57]), .Z(n13622) );
  XOR U14095 ( .A(n13623), .B(n13622), .Z(n13763) );
  XOR U14096 ( .A(n13804), .B(n13763), .Z(n13769) );
  AND U14097 ( .A(y[59]), .B(x[129]), .Z(n13768) );
  XOR U14098 ( .A(n13769), .B(n13768), .Z(n13771) );
  AND U14099 ( .A(y[136]), .B(x[148]), .Z(n13727) );
  AND U14100 ( .A(y[19]), .B(x[121]), .Z(n13726) );
  XOR U14101 ( .A(n13727), .B(n13726), .Z(n13729) );
  AND U14102 ( .A(y[20]), .B(x[120]), .Z(n13728) );
  XOR U14103 ( .A(n13729), .B(n13728), .Z(n13770) );
  XOR U14104 ( .A(n13771), .B(n13770), .Z(n13767) );
  AND U14105 ( .A(y[179]), .B(x[155]), .Z(n14008) );
  NANDN U14106 ( .A(n13628), .B(n14008), .Z(n13632) );
  NAND U14107 ( .A(n13630), .B(n13629), .Z(n13631) );
  AND U14108 ( .A(n13632), .B(n13631), .Z(n13765) );
  XOR U14109 ( .A(n13764), .B(n13765), .Z(n13766) );
  XNOR U14110 ( .A(n13767), .B(n13766), .Z(n13787) );
  NAND U14111 ( .A(y[16]), .B(x[124]), .Z(n13747) );
  NAND U14112 ( .A(y[138]), .B(x[146]), .Z(n13746) );
  NAND U14113 ( .A(y[100]), .B(x[136]), .Z(n13745) );
  XOR U14114 ( .A(n13746), .B(n13745), .Z(n13748) );
  XOR U14115 ( .A(n13747), .B(n13748), .Z(n13712) );
  AND U14116 ( .A(x[154]), .B(y[178]), .Z(n13665) );
  NAND U14117 ( .A(n13665), .B(n13633), .Z(n13743) );
  NAND U14118 ( .A(y[180]), .B(x[152]), .Z(n13881) );
  NAND U14119 ( .A(y[96]), .B(x[140]), .Z(n13821) );
  XNOR U14120 ( .A(n13881), .B(n13821), .Z(n13744) );
  XOR U14121 ( .A(n13743), .B(n13744), .Z(n13711) );
  XNOR U14122 ( .A(n13712), .B(n13711), .Z(n13714) );
  XOR U14123 ( .A(n13714), .B(n13713), .Z(n13785) );
  NANDN U14124 ( .A(n13639), .B(n13638), .Z(n13643) );
  NANDN U14125 ( .A(n13641), .B(n13640), .Z(n13642) );
  AND U14126 ( .A(n13643), .B(n13642), .Z(n13784) );
  XNOR U14127 ( .A(n13785), .B(n13784), .Z(n13786) );
  XNOR U14128 ( .A(n13787), .B(n13786), .Z(n13705) );
  XOR U14129 ( .A(n13706), .B(n13705), .Z(n13708) );
  NANDN U14130 ( .A(n13649), .B(n13648), .Z(n13653) );
  NANDN U14131 ( .A(n13651), .B(n13650), .Z(n13652) );
  NAND U14132 ( .A(n13653), .B(n13652), .Z(n13777) );
  XOR U14133 ( .A(n13776), .B(n13777), .Z(n13779) );
  AND U14134 ( .A(y[97]), .B(x[139]), .Z(n13658) );
  AND U14135 ( .A(y[56]), .B(x[132]), .Z(n13731) );
  AND U14136 ( .A(y[140]), .B(x[144]), .Z(n13730) );
  XOR U14137 ( .A(n13731), .B(n13730), .Z(n13733) );
  AND U14138 ( .A(y[139]), .B(x[145]), .Z(n13732) );
  XOR U14139 ( .A(n13733), .B(n13732), .Z(n13773) );
  NAND U14140 ( .A(x[138]), .B(y[98]), .Z(n13657) );
  XNOR U14141 ( .A(n13658), .B(n13657), .Z(n13723) );
  AND U14142 ( .A(y[99]), .B(x[137]), .Z(n13722) );
  XOR U14143 ( .A(n13723), .B(n13722), .Z(n13772) );
  XOR U14144 ( .A(n13773), .B(n13772), .Z(n13775) );
  XOR U14145 ( .A(n13775), .B(n13774), .Z(n13781) );
  XOR U14146 ( .A(n13780), .B(n13781), .Z(n13783) );
  NAND U14147 ( .A(y[18]), .B(x[122]), .Z(n13758) );
  NAND U14148 ( .A(y[137]), .B(x[147]), .Z(n13757) );
  NAND U14149 ( .A(y[17]), .B(x[123]), .Z(n13756) );
  XOR U14150 ( .A(n13757), .B(n13756), .Z(n13759) );
  XOR U14151 ( .A(n13758), .B(n13759), .Z(n13716) );
  AND U14152 ( .A(x[156]), .B(y[176]), .Z(n13664) );
  NAND U14153 ( .A(x[153]), .B(y[179]), .Z(n13663) );
  XNOR U14154 ( .A(n13664), .B(n13663), .Z(n13740) );
  AND U14155 ( .A(x[155]), .B(y[177]), .Z(n13826) );
  XOR U14156 ( .A(n13826), .B(n13665), .Z(n13739) );
  XOR U14157 ( .A(n13740), .B(n13739), .Z(n13715) );
  XNOR U14158 ( .A(n13716), .B(n13715), .Z(n13718) );
  XOR U14159 ( .A(n13718), .B(n13717), .Z(n13782) );
  XOR U14160 ( .A(n13783), .B(n13782), .Z(n13778) );
  XOR U14161 ( .A(n13779), .B(n13778), .Z(n13707) );
  XOR U14162 ( .A(n13708), .B(n13707), .Z(n13695) );
  NAND U14163 ( .A(n13674), .B(n13673), .Z(n13678) );
  NAND U14164 ( .A(n13676), .B(n13675), .Z(n13677) );
  AND U14165 ( .A(n13678), .B(n13677), .Z(n13702) );
  NAND U14166 ( .A(n13680), .B(n13679), .Z(n13684) );
  NAND U14167 ( .A(n13682), .B(n13681), .Z(n13683) );
  NAND U14168 ( .A(n13684), .B(n13683), .Z(n13699) );
  NAND U14169 ( .A(n13686), .B(n13685), .Z(n13690) );
  NAND U14170 ( .A(n13688), .B(n13687), .Z(n13689) );
  AND U14171 ( .A(n13690), .B(n13689), .Z(n13700) );
  XOR U14172 ( .A(n13699), .B(n13700), .Z(n13701) );
  XOR U14173 ( .A(n13702), .B(n13701), .Z(n13694) );
  IV U14174 ( .A(n13694), .Z(n13692) );
  XOR U14175 ( .A(n13693), .B(n13692), .Z(n13691) );
  XNOR U14176 ( .A(n13695), .B(n13691), .Z(o[140]) );
  NANDN U14177 ( .A(n13692), .B(n13693), .Z(n13698) );
  NOR U14178 ( .A(n13694), .B(n13693), .Z(n13696) );
  OR U14179 ( .A(n13696), .B(n13695), .Z(n13697) );
  AND U14180 ( .A(n13698), .B(n13697), .Z(n13907) );
  NAND U14181 ( .A(n13700), .B(n13699), .Z(n13704) );
  NAND U14182 ( .A(n13702), .B(n13701), .Z(n13703) );
  NAND U14183 ( .A(n13704), .B(n13703), .Z(n13908) );
  XNOR U14184 ( .A(n13907), .B(n13908), .Z(n13910) );
  NAND U14185 ( .A(n13706), .B(n13705), .Z(n13710) );
  NAND U14186 ( .A(n13708), .B(n13707), .Z(n13709) );
  NAND U14187 ( .A(n13710), .B(n13709), .Z(n13913) );
  NANDN U14188 ( .A(n13716), .B(n13715), .Z(n13720) );
  NAND U14189 ( .A(n13718), .B(n13717), .Z(n13719) );
  NAND U14190 ( .A(n13720), .B(n13719), .Z(n13828) );
  XOR U14191 ( .A(n13827), .B(n13828), .Z(n13830) );
  AND U14192 ( .A(y[98]), .B(x[139]), .Z(n13823) );
  AND U14193 ( .A(y[97]), .B(x[138]), .Z(n13721) );
  NAND U14194 ( .A(n13823), .B(n13721), .Z(n13725) );
  NAND U14195 ( .A(n13723), .B(n13722), .Z(n13724) );
  NAND U14196 ( .A(n13725), .B(n13724), .Z(n13790) );
  AND U14197 ( .A(y[141]), .B(x[144]), .Z(n13973) );
  AND U14198 ( .A(y[56]), .B(x[133]), .Z(n13812) );
  AND U14199 ( .A(y[99]), .B(x[138]), .Z(n13811) );
  XOR U14200 ( .A(n13812), .B(n13811), .Z(n13813) );
  XOR U14201 ( .A(n13973), .B(n13813), .Z(n13808) );
  AND U14202 ( .A(y[17]), .B(x[124]), .Z(n13951) );
  AND U14203 ( .A(y[137]), .B(x[148]), .Z(n13817) );
  AND U14204 ( .A(y[16]), .B(x[125]), .Z(n13816) );
  XOR U14205 ( .A(n13817), .B(n13816), .Z(n13818) );
  XOR U14206 ( .A(n13951), .B(n13818), .Z(n13807) );
  XOR U14207 ( .A(n13808), .B(n13807), .Z(n13810) );
  XOR U14208 ( .A(n13810), .B(n13809), .Z(n13791) );
  XOR U14209 ( .A(n13790), .B(n13791), .Z(n13793) );
  AND U14210 ( .A(y[178]), .B(x[155]), .Z(n13735) );
  AND U14211 ( .A(n13735), .B(n13734), .Z(n13883) );
  AND U14212 ( .A(x[152]), .B(y[181]), .Z(n13737) );
  AND U14213 ( .A(x[153]), .B(y[180]), .Z(n13736) );
  XOR U14214 ( .A(n13737), .B(n13736), .Z(n13882) );
  XOR U14215 ( .A(n13883), .B(n13882), .Z(n13864) );
  AND U14216 ( .A(y[61]), .B(x[128]), .Z(n13872) );
  AND U14217 ( .A(y[20]), .B(x[121]), .Z(n13871) );
  XOR U14218 ( .A(n13872), .B(n13871), .Z(n13874) );
  AND U14219 ( .A(y[57]), .B(x[132]), .Z(n13873) );
  XOR U14220 ( .A(n13874), .B(n13873), .Z(n13863) );
  XOR U14221 ( .A(n13864), .B(n13863), .Z(n13866) );
  XOR U14222 ( .A(n13865), .B(n13866), .Z(n13792) );
  XOR U14223 ( .A(n13793), .B(n13792), .Z(n13829) );
  XOR U14224 ( .A(n13830), .B(n13829), .Z(n13905) );
  AND U14225 ( .A(y[179]), .B(x[156]), .Z(n14075) );
  NAND U14226 ( .A(n14075), .B(n13738), .Z(n13742) );
  NAND U14227 ( .A(n13740), .B(n13739), .Z(n13741) );
  NAND U14228 ( .A(n13742), .B(n13741), .Z(n13837) );
  XOR U14229 ( .A(n13837), .B(n13838), .Z(n13840) );
  NAND U14230 ( .A(n13746), .B(n13745), .Z(n13750) );
  NAND U14231 ( .A(n13748), .B(n13747), .Z(n13749) );
  AND U14232 ( .A(n13750), .B(n13749), .Z(n13844) );
  AND U14233 ( .A(y[58]), .B(x[131]), .Z(n14004) );
  NAND U14234 ( .A(x[130]), .B(y[59]), .Z(n13751) );
  XNOR U14235 ( .A(n14004), .B(n13751), .Z(n13806) );
  AND U14236 ( .A(y[60]), .B(x[129]), .Z(n13805) );
  XOR U14237 ( .A(n13806), .B(n13805), .Z(n13842) );
  AND U14238 ( .A(y[179]), .B(x[154]), .Z(n13797) );
  AND U14239 ( .A(y[176]), .B(x[157]), .Z(n13796) );
  XOR U14240 ( .A(n13797), .B(n13796), .Z(n13799) );
  AND U14241 ( .A(x[156]), .B(y[177]), .Z(n13753) );
  NAND U14242 ( .A(x[155]), .B(y[178]), .Z(n13752) );
  XNOR U14243 ( .A(n13753), .B(n13752), .Z(n13798) );
  XOR U14244 ( .A(n13799), .B(n13798), .Z(n13841) );
  XOR U14245 ( .A(n13842), .B(n13841), .Z(n13843) );
  XOR U14246 ( .A(n13844), .B(n13843), .Z(n13839) );
  XOR U14247 ( .A(n13840), .B(n13839), .Z(n13854) );
  AND U14248 ( .A(x[141]), .B(y[96]), .Z(n13755) );
  AND U14249 ( .A(x[140]), .B(y[97]), .Z(n13754) );
  XOR U14250 ( .A(n13755), .B(n13754), .Z(n13822) );
  XOR U14251 ( .A(n13823), .B(n13822), .Z(n13858) );
  AND U14252 ( .A(y[136]), .B(x[149]), .Z(n13801) );
  AND U14253 ( .A(y[18]), .B(x[123]), .Z(n13800) );
  XOR U14254 ( .A(n13801), .B(n13800), .Z(n13803) );
  AND U14255 ( .A(y[19]), .B(x[122]), .Z(n13802) );
  XOR U14256 ( .A(n13803), .B(n13802), .Z(n13857) );
  XOR U14257 ( .A(n13858), .B(n13857), .Z(n13860) );
  NAND U14258 ( .A(n13757), .B(n13756), .Z(n13761) );
  NAND U14259 ( .A(n13759), .B(n13758), .Z(n13760) );
  AND U14260 ( .A(n13761), .B(n13760), .Z(n13859) );
  XOR U14261 ( .A(n13860), .B(n13859), .Z(n13852) );
  AND U14262 ( .A(y[60]), .B(x[131]), .Z(n14074) );
  AND U14263 ( .A(y[138]), .B(x[147]), .Z(n13894) );
  AND U14264 ( .A(y[100]), .B(x[137]), .Z(n13958) );
  XOR U14265 ( .A(n13894), .B(n13958), .Z(n13896) );
  AND U14266 ( .A(y[101]), .B(x[136]), .Z(n13895) );
  XOR U14267 ( .A(n13896), .B(n13895), .Z(n13832) );
  AND U14268 ( .A(y[21]), .B(x[120]), .Z(n13887) );
  AND U14269 ( .A(y[140]), .B(x[145]), .Z(n13886) );
  XOR U14270 ( .A(n13887), .B(n13886), .Z(n13889) );
  AND U14271 ( .A(y[139]), .B(x[146]), .Z(n13888) );
  XOR U14272 ( .A(n13889), .B(n13888), .Z(n13831) );
  XNOR U14273 ( .A(n13832), .B(n13831), .Z(n13834) );
  XOR U14274 ( .A(n13833), .B(n13834), .Z(n13851) );
  XNOR U14275 ( .A(n13852), .B(n13851), .Z(n13853) );
  XOR U14276 ( .A(n13854), .B(n13853), .Z(n13904) );
  XOR U14277 ( .A(n13847), .B(n13848), .Z(n13849) );
  XOR U14278 ( .A(n13850), .B(n13849), .Z(n13903) );
  XNOR U14279 ( .A(n13904), .B(n13903), .Z(n13906) );
  XNOR U14280 ( .A(n13905), .B(n13906), .Z(n13914) );
  XOR U14281 ( .A(n13913), .B(n13914), .Z(n13915) );
  NANDN U14282 ( .A(n13785), .B(n13784), .Z(n13789) );
  NAND U14283 ( .A(n13787), .B(n13786), .Z(n13788) );
  AND U14284 ( .A(n13789), .B(n13788), .Z(n13899) );
  XNOR U14285 ( .A(n13900), .B(n13899), .Z(n13902) );
  XOR U14286 ( .A(n13901), .B(n13902), .Z(n13916) );
  XOR U14287 ( .A(n13910), .B(n13909), .Z(o[141]) );
  NAND U14288 ( .A(n13791), .B(n13790), .Z(n13795) );
  NAND U14289 ( .A(n13793), .B(n13792), .Z(n13794) );
  AND U14290 ( .A(n13795), .B(n13794), .Z(n14198) );
  AND U14291 ( .A(y[139]), .B(x[147]), .Z(n14024) );
  AND U14292 ( .A(y[99]), .B(x[139]), .Z(n14023) );
  XOR U14293 ( .A(n14024), .B(n14023), .Z(n14022) );
  AND U14294 ( .A(y[19]), .B(x[123]), .Z(n14021) );
  XOR U14295 ( .A(n14022), .B(n14021), .Z(n13999) );
  AND U14296 ( .A(y[140]), .B(x[146]), .Z(n13979) );
  AND U14297 ( .A(y[98]), .B(x[140]), .Z(n13978) );
  XOR U14298 ( .A(n13979), .B(n13978), .Z(n13977) );
  AND U14299 ( .A(y[20]), .B(x[122]), .Z(n13976) );
  XNOR U14300 ( .A(n13977), .B(n13976), .Z(n13998) );
  XNOR U14301 ( .A(n13997), .B(n13996), .Z(n14157) );
  XOR U14302 ( .A(n14158), .B(n14157), .Z(n14156) );
  XOR U14303 ( .A(n14155), .B(n14156), .Z(n13928) );
  XOR U14304 ( .A(n13928), .B(n13927), .Z(n13926) );
  NAND U14305 ( .A(n13812), .B(n13811), .Z(n13815) );
  NAND U14306 ( .A(n13973), .B(n13813), .Z(n13814) );
  NAND U14307 ( .A(n13815), .B(n13814), .Z(n14118) );
  NAND U14308 ( .A(n13817), .B(n13816), .Z(n13820) );
  NAND U14309 ( .A(n13951), .B(n13818), .Z(n13819) );
  NAND U14310 ( .A(n13820), .B(n13819), .Z(n14117) );
  XOR U14311 ( .A(n14118), .B(n14117), .Z(n14120) );
  AND U14312 ( .A(y[97]), .B(x[141]), .Z(n13964) );
  AND U14313 ( .A(x[124]), .B(y[18]), .Z(n13825) );
  NAND U14314 ( .A(x[125]), .B(y[17]), .Z(n13824) );
  XNOR U14315 ( .A(n13825), .B(n13824), .Z(n13950) );
  AND U14316 ( .A(y[136]), .B(x[150]), .Z(n13949) );
  XOR U14317 ( .A(n13950), .B(n13949), .Z(n14144) );
  AND U14318 ( .A(y[181]), .B(x[153]), .Z(n14016) );
  AND U14319 ( .A(y[178]), .B(x[156]), .Z(n13893) );
  AND U14320 ( .A(n13893), .B(n13826), .Z(n14014) );
  AND U14321 ( .A(y[180]), .B(x[154]), .Z(n14013) );
  XOR U14322 ( .A(n14014), .B(n14013), .Z(n14015) );
  XNOR U14323 ( .A(n14016), .B(n14015), .Z(n14143) );
  XNOR U14324 ( .A(n14142), .B(n14141), .Z(n14119) );
  XOR U14325 ( .A(n14120), .B(n14119), .Z(n13925) );
  XOR U14326 ( .A(n13926), .B(n13925), .Z(n13922) );
  NAND U14327 ( .A(n13832), .B(n13831), .Z(n13836) );
  NANDN U14328 ( .A(n13834), .B(n13833), .Z(n13835) );
  AND U14329 ( .A(n13836), .B(n13835), .Z(n14152) );
  XOR U14330 ( .A(n14152), .B(n14151), .Z(n14150) );
  NAND U14331 ( .A(n13842), .B(n13841), .Z(n13846) );
  NAND U14332 ( .A(n13844), .B(n13843), .Z(n13845) );
  AND U14333 ( .A(n13846), .B(n13845), .Z(n14149) );
  XOR U14334 ( .A(n14150), .B(n14149), .Z(n13919) );
  XOR U14335 ( .A(n13920), .B(n13919), .Z(n14197) );
  XOR U14336 ( .A(n14198), .B(n14197), .Z(n14196) );
  NANDN U14337 ( .A(n13852), .B(n13851), .Z(n13856) );
  NANDN U14338 ( .A(n13854), .B(n13853), .Z(n13855) );
  NAND U14339 ( .A(n13856), .B(n13855), .Z(n14173) );
  NAND U14340 ( .A(n13858), .B(n13857), .Z(n13862) );
  NAND U14341 ( .A(n13860), .B(n13859), .Z(n13861) );
  AND U14342 ( .A(n13862), .B(n13861), .Z(n14178) );
  NAND U14343 ( .A(n13864), .B(n13863), .Z(n13868) );
  NAND U14344 ( .A(n13866), .B(n13865), .Z(n13867) );
  AND U14345 ( .A(n13868), .B(n13867), .Z(n13932) );
  AND U14346 ( .A(y[102]), .B(x[136]), .Z(n13991) );
  AND U14347 ( .A(y[16]), .B(x[126]), .Z(n13990) );
  XOR U14348 ( .A(n13991), .B(n13990), .Z(n13989) );
  AND U14349 ( .A(y[137]), .B(x[149]), .Z(n13988) );
  XOR U14350 ( .A(n13989), .B(n13988), .Z(n14132) );
  AND U14351 ( .A(y[57]), .B(x[133]), .Z(n13946) );
  AND U14352 ( .A(y[60]), .B(x[130]), .Z(n13945) );
  XOR U14353 ( .A(n13946), .B(n13945), .Z(n13944) );
  AND U14354 ( .A(y[61]), .B(x[129]), .Z(n13943) );
  XOR U14355 ( .A(n13944), .B(n13943), .Z(n14003) );
  AND U14356 ( .A(x[132]), .B(y[58]), .Z(n13870) );
  NAND U14357 ( .A(x[131]), .B(y[59]), .Z(n13869) );
  XNOR U14358 ( .A(n13870), .B(n13869), .Z(n14002) );
  XOR U14359 ( .A(n14003), .B(n14002), .Z(n14131) );
  XOR U14360 ( .A(n14132), .B(n14131), .Z(n14130) );
  AND U14361 ( .A(y[182]), .B(x[152]), .Z(n13963) );
  XOR U14362 ( .A(n13964), .B(n13963), .Z(n13962) );
  AND U14363 ( .A(y[96]), .B(x[142]), .Z(n13961) );
  XOR U14364 ( .A(n13962), .B(n13961), .Z(n14129) );
  XOR U14365 ( .A(n14130), .B(n14129), .Z(n13934) );
  NAND U14366 ( .A(n13872), .B(n13871), .Z(n13876) );
  NAND U14367 ( .A(n13874), .B(n13873), .Z(n13875) );
  AND U14368 ( .A(n13876), .B(n13875), .Z(n13937) );
  AND U14369 ( .A(y[138]), .B(x[148]), .Z(n13957) );
  AND U14370 ( .A(x[137]), .B(y[101]), .Z(n13878) );
  AND U14371 ( .A(x[138]), .B(y[100]), .Z(n13877) );
  XOR U14372 ( .A(n13878), .B(n13877), .Z(n13956) );
  XOR U14373 ( .A(n13957), .B(n13956), .Z(n13940) );
  AND U14374 ( .A(y[22]), .B(x[120]), .Z(n13972) );
  AND U14375 ( .A(y[142]), .B(x[144]), .Z(n13880) );
  AND U14376 ( .A(x[145]), .B(y[141]), .Z(n13879) );
  XOR U14377 ( .A(n13880), .B(n13879), .Z(n13971) );
  XNOR U14378 ( .A(n13972), .B(n13971), .Z(n13939) );
  XNOR U14379 ( .A(n13937), .B(n13938), .Z(n13933) );
  XOR U14380 ( .A(n13932), .B(n13931), .Z(n14177) );
  XOR U14381 ( .A(n14178), .B(n14177), .Z(n14180) );
  NANDN U14382 ( .A(n13881), .B(n14016), .Z(n13885) );
  NAND U14383 ( .A(n13883), .B(n13882), .Z(n13884) );
  NAND U14384 ( .A(n13885), .B(n13884), .Z(n14116) );
  NAND U14385 ( .A(n13887), .B(n13886), .Z(n13891) );
  NAND U14386 ( .A(n13889), .B(n13888), .Z(n13890) );
  AND U14387 ( .A(n13891), .B(n13890), .Z(n14136) );
  AND U14388 ( .A(y[21]), .B(x[121]), .Z(n13987) );
  AND U14389 ( .A(y[56]), .B(x[134]), .Z(n13986) );
  XOR U14390 ( .A(n13987), .B(n13986), .Z(n13985) );
  AND U14391 ( .A(y[62]), .B(x[128]), .Z(n13984) );
  XOR U14392 ( .A(n13985), .B(n13984), .Z(n14138) );
  NAND U14393 ( .A(x[157]), .B(y[177]), .Z(n13892) );
  XNOR U14394 ( .A(n13893), .B(n13892), .Z(n14010) );
  AND U14395 ( .A(y[176]), .B(x[158]), .Z(n14009) );
  XOR U14396 ( .A(n14010), .B(n14009), .Z(n14007) );
  XNOR U14397 ( .A(n14008), .B(n14007), .Z(n14137) );
  XNOR U14398 ( .A(n14136), .B(n14135), .Z(n14115) );
  XOR U14399 ( .A(n14116), .B(n14115), .Z(n14114) );
  NAND U14400 ( .A(n13894), .B(n13958), .Z(n13898) );
  NAND U14401 ( .A(n13896), .B(n13895), .Z(n13897) );
  NAND U14402 ( .A(n13898), .B(n13897), .Z(n14113) );
  XOR U14403 ( .A(n14114), .B(n14113), .Z(n14179) );
  XOR U14404 ( .A(n14173), .B(n14174), .Z(n14171) );
  XOR U14405 ( .A(n14172), .B(n14171), .Z(n14195) );
  XOR U14406 ( .A(n14196), .B(n14195), .Z(n14189) );
  XNOR U14407 ( .A(n14192), .B(n14191), .Z(n14190) );
  XOR U14408 ( .A(n14189), .B(n14190), .Z(n14210) );
  NANDN U14409 ( .A(n13908), .B(n13907), .Z(n13912) );
  NAND U14410 ( .A(n13910), .B(n13909), .Z(n13911) );
  AND U14411 ( .A(n13912), .B(n13911), .Z(n14209) );
  NAND U14412 ( .A(n13914), .B(n13913), .Z(n13918) );
  NANDN U14413 ( .A(n13916), .B(n13915), .Z(n13917) );
  AND U14414 ( .A(n13918), .B(n13917), .Z(n14207) );
  XNOR U14415 ( .A(n14208), .B(n14207), .Z(o[142]) );
  NAND U14416 ( .A(n13920), .B(n13919), .Z(n13924) );
  NANDN U14417 ( .A(n13922), .B(n13921), .Z(n13923) );
  AND U14418 ( .A(n13924), .B(n13923), .Z(n14206) );
  NAND U14419 ( .A(n13926), .B(n13925), .Z(n13930) );
  NAND U14420 ( .A(n13928), .B(n13927), .Z(n13929) );
  AND U14421 ( .A(n13930), .B(n13929), .Z(n14188) );
  NAND U14422 ( .A(n13932), .B(n13931), .Z(n13936) );
  NANDN U14423 ( .A(n13934), .B(n13933), .Z(n13935) );
  AND U14424 ( .A(n13936), .B(n13935), .Z(n14170) );
  NANDN U14425 ( .A(n13938), .B(n13937), .Z(n13942) );
  NANDN U14426 ( .A(n13940), .B(n13939), .Z(n13941) );
  AND U14427 ( .A(n13942), .B(n13941), .Z(n14128) );
  NAND U14428 ( .A(n13944), .B(n13943), .Z(n13948) );
  NAND U14429 ( .A(n13946), .B(n13945), .Z(n13947) );
  AND U14430 ( .A(n13948), .B(n13947), .Z(n13955) );
  NAND U14431 ( .A(n13950), .B(n13949), .Z(n13953) );
  AND U14432 ( .A(y[18]), .B(x[125]), .Z(n14076) );
  NAND U14433 ( .A(n13951), .B(n14076), .Z(n13952) );
  NAND U14434 ( .A(n13953), .B(n13952), .Z(n13954) );
  XNOR U14435 ( .A(n13955), .B(n13954), .Z(n13970) );
  NAND U14436 ( .A(n13957), .B(n13956), .Z(n13960) );
  AND U14437 ( .A(y[101]), .B(x[138]), .Z(n14080) );
  NAND U14438 ( .A(n13958), .B(n14080), .Z(n13959) );
  AND U14439 ( .A(n13960), .B(n13959), .Z(n13968) );
  NAND U14440 ( .A(n13962), .B(n13961), .Z(n13966) );
  NAND U14441 ( .A(n13964), .B(n13963), .Z(n13965) );
  NAND U14442 ( .A(n13966), .B(n13965), .Z(n13967) );
  XNOR U14443 ( .A(n13968), .B(n13967), .Z(n13969) );
  XOR U14444 ( .A(n13970), .B(n13969), .Z(n13995) );
  NAND U14445 ( .A(n13972), .B(n13971), .Z(n13975) );
  AND U14446 ( .A(y[142]), .B(x[145]), .Z(n14079) );
  NAND U14447 ( .A(n13973), .B(n14079), .Z(n13974) );
  AND U14448 ( .A(n13975), .B(n13974), .Z(n13983) );
  NAND U14449 ( .A(n13977), .B(n13976), .Z(n13981) );
  NAND U14450 ( .A(n13979), .B(n13978), .Z(n13980) );
  NAND U14451 ( .A(n13981), .B(n13980), .Z(n13982) );
  XNOR U14452 ( .A(n13983), .B(n13982), .Z(n13993) );
  XNOR U14453 ( .A(n13993), .B(n13992), .Z(n13994) );
  XNOR U14454 ( .A(n13995), .B(n13994), .Z(n14126) );
  NAND U14455 ( .A(n13997), .B(n13996), .Z(n14001) );
  NANDN U14456 ( .A(n13999), .B(n13998), .Z(n14000) );
  AND U14457 ( .A(n14001), .B(n14000), .Z(n14124) );
  NAND U14458 ( .A(n14003), .B(n14002), .Z(n14006) );
  AND U14459 ( .A(y[59]), .B(x[132]), .Z(n14073) );
  NAND U14460 ( .A(n14004), .B(n14073), .Z(n14005) );
  AND U14461 ( .A(n14006), .B(n14005), .Z(n14112) );
  NAND U14462 ( .A(n14008), .B(n14007), .Z(n14012) );
  AND U14463 ( .A(n14010), .B(n14009), .Z(n14011) );
  ANDN U14464 ( .B(n14012), .A(n14011), .Z(n14020) );
  AND U14465 ( .A(n14014), .B(n14013), .Z(n14018) );
  AND U14466 ( .A(n14016), .B(n14015), .Z(n14017) );
  OR U14467 ( .A(n14018), .B(n14017), .Z(n14019) );
  XNOR U14468 ( .A(n14020), .B(n14019), .Z(n14110) );
  NAND U14469 ( .A(n14022), .B(n14021), .Z(n14026) );
  NAND U14470 ( .A(n14024), .B(n14023), .Z(n14025) );
  AND U14471 ( .A(n14026), .B(n14025), .Z(n14108) );
  AND U14472 ( .A(x[129]), .B(y[62]), .Z(n14028) );
  NAND U14473 ( .A(x[130]), .B(y[61]), .Z(n14027) );
  XNOR U14474 ( .A(n14028), .B(n14027), .Z(n14034) );
  AND U14475 ( .A(x[144]), .B(y[143]), .Z(n14032) );
  NAND U14476 ( .A(y[177]), .B(x[156]), .Z(n14029) );
  AND U14477 ( .A(x[157]), .B(n14029), .Z(n14030) );
  NAND U14478 ( .A(n14030), .B(y[178]), .Z(n14031) );
  XNOR U14479 ( .A(n14032), .B(n14031), .Z(n14033) );
  XOR U14480 ( .A(n14034), .B(n14033), .Z(n14042) );
  AND U14481 ( .A(x[134]), .B(y[57]), .Z(n14036) );
  NAND U14482 ( .A(x[146]), .B(y[141]), .Z(n14035) );
  XNOR U14483 ( .A(n14036), .B(n14035), .Z(n14040) );
  AND U14484 ( .A(x[133]), .B(y[58]), .Z(n14038) );
  NAND U14485 ( .A(x[135]), .B(y[56]), .Z(n14037) );
  XNOR U14486 ( .A(n14038), .B(n14037), .Z(n14039) );
  XNOR U14487 ( .A(n14040), .B(n14039), .Z(n14041) );
  XNOR U14488 ( .A(n14042), .B(n14041), .Z(n14106) );
  AND U14489 ( .A(x[139]), .B(y[100]), .Z(n14044) );
  NAND U14490 ( .A(x[123]), .B(y[20]), .Z(n14043) );
  XNOR U14491 ( .A(n14044), .B(n14043), .Z(n14048) );
  AND U14492 ( .A(x[150]), .B(y[137]), .Z(n14046) );
  NAND U14493 ( .A(x[140]), .B(y[99]), .Z(n14045) );
  XNOR U14494 ( .A(n14046), .B(n14045), .Z(n14047) );
  XOR U14495 ( .A(n14048), .B(n14047), .Z(n14056) );
  AND U14496 ( .A(x[122]), .B(y[21]), .Z(n14050) );
  NAND U14497 ( .A(x[154]), .B(y[181]), .Z(n14049) );
  XNOR U14498 ( .A(n14050), .B(n14049), .Z(n14054) );
  AND U14499 ( .A(x[155]), .B(y[180]), .Z(n14052) );
  NAND U14500 ( .A(x[124]), .B(y[19]), .Z(n14051) );
  XNOR U14501 ( .A(n14052), .B(n14051), .Z(n14053) );
  XNOR U14502 ( .A(n14054), .B(n14053), .Z(n14055) );
  XNOR U14503 ( .A(n14056), .B(n14055), .Z(n14072) );
  AND U14504 ( .A(x[152]), .B(y[183]), .Z(n14058) );
  NAND U14505 ( .A(x[128]), .B(y[63]), .Z(n14057) );
  XNOR U14506 ( .A(n14058), .B(n14057), .Z(n14062) );
  AND U14507 ( .A(x[148]), .B(y[139]), .Z(n14060) );
  NAND U14508 ( .A(x[127]), .B(y[16]), .Z(n14059) );
  XNOR U14509 ( .A(n14060), .B(n14059), .Z(n14061) );
  XOR U14510 ( .A(n14062), .B(n14061), .Z(n14070) );
  AND U14511 ( .A(x[143]), .B(y[96]), .Z(n14064) );
  NAND U14512 ( .A(x[151]), .B(y[136]), .Z(n14063) );
  XNOR U14513 ( .A(n14064), .B(n14063), .Z(n14068) );
  AND U14514 ( .A(x[121]), .B(y[22]), .Z(n14066) );
  NAND U14515 ( .A(x[141]), .B(y[98]), .Z(n14065) );
  XNOR U14516 ( .A(n14066), .B(n14065), .Z(n14067) );
  XNOR U14517 ( .A(n14068), .B(n14067), .Z(n14069) );
  XNOR U14518 ( .A(n14070), .B(n14069), .Z(n14071) );
  XOR U14519 ( .A(n14072), .B(n14071), .Z(n14104) );
  XOR U14520 ( .A(n14074), .B(n14073), .Z(n14078) );
  XNOR U14521 ( .A(n14076), .B(n14075), .Z(n14077) );
  XNOR U14522 ( .A(n14078), .B(n14077), .Z(n14102) );
  AND U14523 ( .A(x[147]), .B(y[140]), .Z(n14100) );
  AND U14524 ( .A(x[136]), .B(y[103]), .Z(n14082) );
  XNOR U14525 ( .A(n14080), .B(n14079), .Z(n14081) );
  XNOR U14526 ( .A(n14082), .B(n14081), .Z(n14098) );
  AND U14527 ( .A(x[137]), .B(y[102]), .Z(n14084) );
  NAND U14528 ( .A(x[158]), .B(y[177]), .Z(n14083) );
  XNOR U14529 ( .A(n14084), .B(n14083), .Z(n14088) );
  AND U14530 ( .A(x[159]), .B(y[176]), .Z(n14086) );
  NAND U14531 ( .A(x[142]), .B(y[97]), .Z(n14085) );
  XNOR U14532 ( .A(n14086), .B(n14085), .Z(n14087) );
  XOR U14533 ( .A(n14088), .B(n14087), .Z(n14096) );
  AND U14534 ( .A(x[153]), .B(y[182]), .Z(n14090) );
  NAND U14535 ( .A(x[126]), .B(y[17]), .Z(n14089) );
  XNOR U14536 ( .A(n14090), .B(n14089), .Z(n14094) );
  AND U14537 ( .A(x[120]), .B(y[23]), .Z(n14092) );
  NAND U14538 ( .A(x[149]), .B(y[138]), .Z(n14091) );
  XNOR U14539 ( .A(n14092), .B(n14091), .Z(n14093) );
  XNOR U14540 ( .A(n14094), .B(n14093), .Z(n14095) );
  XNOR U14541 ( .A(n14096), .B(n14095), .Z(n14097) );
  XNOR U14542 ( .A(n14098), .B(n14097), .Z(n14099) );
  XNOR U14543 ( .A(n14100), .B(n14099), .Z(n14101) );
  XNOR U14544 ( .A(n14102), .B(n14101), .Z(n14103) );
  XNOR U14545 ( .A(n14104), .B(n14103), .Z(n14105) );
  XNOR U14546 ( .A(n14106), .B(n14105), .Z(n14107) );
  XNOR U14547 ( .A(n14108), .B(n14107), .Z(n14109) );
  XNOR U14548 ( .A(n14110), .B(n14109), .Z(n14111) );
  XNOR U14549 ( .A(n14112), .B(n14111), .Z(n14122) );
  XNOR U14550 ( .A(n14122), .B(n14121), .Z(n14123) );
  XNOR U14551 ( .A(n14124), .B(n14123), .Z(n14125) );
  XNOR U14552 ( .A(n14126), .B(n14125), .Z(n14127) );
  XNOR U14553 ( .A(n14128), .B(n14127), .Z(n14168) );
  NAND U14554 ( .A(n14130), .B(n14129), .Z(n14134) );
  NAND U14555 ( .A(n14132), .B(n14131), .Z(n14133) );
  AND U14556 ( .A(n14134), .B(n14133), .Z(n14166) );
  NAND U14557 ( .A(n14136), .B(n14135), .Z(n14140) );
  NANDN U14558 ( .A(n14138), .B(n14137), .Z(n14139) );
  AND U14559 ( .A(n14140), .B(n14139), .Z(n14148) );
  NAND U14560 ( .A(n14142), .B(n14141), .Z(n14146) );
  NANDN U14561 ( .A(n14144), .B(n14143), .Z(n14145) );
  NAND U14562 ( .A(n14146), .B(n14145), .Z(n14147) );
  XNOR U14563 ( .A(n14148), .B(n14147), .Z(n14164) );
  NAND U14564 ( .A(n14150), .B(n14149), .Z(n14154) );
  NAND U14565 ( .A(n14152), .B(n14151), .Z(n14153) );
  AND U14566 ( .A(n14154), .B(n14153), .Z(n14162) );
  NAND U14567 ( .A(n14156), .B(n14155), .Z(n14160) );
  NAND U14568 ( .A(n14158), .B(n14157), .Z(n14159) );
  NAND U14569 ( .A(n14160), .B(n14159), .Z(n14161) );
  XNOR U14570 ( .A(n14162), .B(n14161), .Z(n14163) );
  XNOR U14571 ( .A(n14164), .B(n14163), .Z(n14165) );
  XNOR U14572 ( .A(n14166), .B(n14165), .Z(n14167) );
  XNOR U14573 ( .A(n14168), .B(n14167), .Z(n14169) );
  XNOR U14574 ( .A(n14170), .B(n14169), .Z(n14186) );
  NAND U14575 ( .A(n14172), .B(n14171), .Z(n14176) );
  AND U14576 ( .A(n14174), .B(n14173), .Z(n14175) );
  ANDN U14577 ( .B(n14176), .A(n14175), .Z(n14184) );
  AND U14578 ( .A(n14178), .B(n14177), .Z(n14182) );
  ANDN U14579 ( .B(n14180), .A(n14179), .Z(n14181) );
  OR U14580 ( .A(n14182), .B(n14181), .Z(n14183) );
  XNOR U14581 ( .A(n14184), .B(n14183), .Z(n14185) );
  XNOR U14582 ( .A(n14186), .B(n14185), .Z(n14187) );
  XNOR U14583 ( .A(n14188), .B(n14187), .Z(n14204) );
  OR U14584 ( .A(n14190), .B(n14189), .Z(n14194) );
  NAND U14585 ( .A(n14192), .B(n14191), .Z(n14193) );
  AND U14586 ( .A(n14194), .B(n14193), .Z(n14202) );
  NAND U14587 ( .A(n14196), .B(n14195), .Z(n14200) );
  NAND U14588 ( .A(n14198), .B(n14197), .Z(n14199) );
  NAND U14589 ( .A(n14200), .B(n14199), .Z(n14201) );
  XNOR U14590 ( .A(n14202), .B(n14201), .Z(n14203) );
  XNOR U14591 ( .A(n14204), .B(n14203), .Z(n14205) );
  XNOR U14592 ( .A(n14206), .B(n14205), .Z(n14214) );
  NAND U14593 ( .A(n14208), .B(n14207), .Z(n14212) );
  NANDN U14594 ( .A(n14210), .B(n14209), .Z(n14211) );
  NAND U14595 ( .A(n14212), .B(n14211), .Z(n14213) );
  XNOR U14596 ( .A(n14214), .B(n14213), .Z(o[143]) );
  NAND U14597 ( .A(y[184]), .B(x[152]), .Z(n14328) );
  NAND U14598 ( .A(y[64]), .B(x[128]), .Z(n14217) );
  XOR U14599 ( .A(n14328), .B(n14217), .Z(n14218) );
  AND U14600 ( .A(y[24]), .B(x[120]), .Z(n14225) );
  AND U14601 ( .A(y[104]), .B(x[136]), .Z(n14222) );
  XOR U14602 ( .A(n14225), .B(n14222), .Z(n14221) );
  AND U14603 ( .A(y[144]), .B(x[144]), .Z(n14220) );
  XNOR U14604 ( .A(n14221), .B(n14220), .Z(n14219) );
  XNOR U14605 ( .A(n14218), .B(n14219), .Z(o[144]) );
  AND U14606 ( .A(x[121]), .B(y[24]), .Z(n14216) );
  NAND U14607 ( .A(x[120]), .B(y[25]), .Z(n14215) );
  XNOR U14608 ( .A(n14216), .B(n14215), .Z(n14227) );
  AND U14609 ( .A(y[64]), .B(x[129]), .Z(n14226) );
  XOR U14610 ( .A(n14227), .B(n14226), .Z(n14244) );
  AND U14611 ( .A(y[184]), .B(x[153]), .Z(n14451) );
  AND U14612 ( .A(y[105]), .B(x[136]), .Z(n14230) );
  XOR U14613 ( .A(n14451), .B(n14230), .Z(n14232) );
  AND U14614 ( .A(y[185]), .B(x[152]), .Z(n14254) );
  NAND U14615 ( .A(y[104]), .B(x[137]), .Z(n14253) );
  XNOR U14616 ( .A(n14254), .B(n14253), .Z(n14231) );
  XOR U14617 ( .A(n14232), .B(n14231), .Z(n14242) );
  AND U14618 ( .A(y[65]), .B(x[128]), .Z(n14474) );
  AND U14619 ( .A(y[145]), .B(x[144]), .Z(n14247) );
  XOR U14620 ( .A(n14474), .B(n14247), .Z(n14249) );
  AND U14621 ( .A(y[144]), .B(x[145]), .Z(n14248) );
  XNOR U14622 ( .A(n14249), .B(n14248), .Z(n14241) );
  XNOR U14623 ( .A(n14242), .B(n14241), .Z(n14243) );
  XNOR U14624 ( .A(n14244), .B(n14243), .Z(n14238) );
  NAND U14625 ( .A(n14221), .B(n14220), .Z(n14224) );
  AND U14626 ( .A(n14225), .B(n14222), .Z(n14223) );
  ANDN U14627 ( .B(n14224), .A(n14223), .Z(n14235) );
  XNOR U14628 ( .A(n14236), .B(n14235), .Z(n14237) );
  XNOR U14629 ( .A(n14238), .B(n14237), .Z(o[145]) );
  NAND U14630 ( .A(y[25]), .B(x[121]), .Z(n14276) );
  NANDN U14631 ( .A(n14276), .B(n14225), .Z(n14229) );
  NAND U14632 ( .A(n14227), .B(n14226), .Z(n14228) );
  AND U14633 ( .A(n14229), .B(n14228), .Z(n14296) );
  NAND U14634 ( .A(n14451), .B(n14230), .Z(n14234) );
  NAND U14635 ( .A(n14232), .B(n14231), .Z(n14233) );
  AND U14636 ( .A(n14234), .B(n14233), .Z(n14295) );
  AND U14637 ( .A(y[146]), .B(x[144]), .Z(n14300) );
  NAND U14638 ( .A(y[26]), .B(x[120]), .Z(n14301) );
  XNOR U14639 ( .A(n14300), .B(n14301), .Z(n14302) );
  NAND U14640 ( .A(y[64]), .B(x[130]), .Z(n14303) );
  XNOR U14641 ( .A(n14302), .B(n14303), .Z(n14294) );
  XOR U14642 ( .A(n14295), .B(n14294), .Z(n14297) );
  XOR U14643 ( .A(n14296), .B(n14297), .Z(n14256) );
  NANDN U14644 ( .A(n14236), .B(n14235), .Z(n14240) );
  NAND U14645 ( .A(n14238), .B(n14237), .Z(n14239) );
  NAND U14646 ( .A(n14240), .B(n14239), .Z(n14255) );
  XNOR U14647 ( .A(n14256), .B(n14255), .Z(n14258) );
  NANDN U14648 ( .A(n14242), .B(n14241), .Z(n14246) );
  NANDN U14649 ( .A(n14244), .B(n14243), .Z(n14245) );
  AND U14650 ( .A(n14246), .B(n14245), .Z(n14264) );
  AND U14651 ( .A(y[24]), .B(x[122]), .Z(n14273) );
  NAND U14652 ( .A(y[106]), .B(x[136]), .Z(n14274) );
  XNOR U14653 ( .A(n14273), .B(n14274), .Z(n14275) );
  AND U14654 ( .A(y[144]), .B(x[146]), .Z(n14308) );
  XOR U14655 ( .A(n14309), .B(n14308), .Z(n14311) );
  AND U14656 ( .A(y[104]), .B(x[138]), .Z(n14368) );
  AND U14657 ( .A(y[186]), .B(x[152]), .Z(n14286) );
  XOR U14658 ( .A(n14368), .B(n14286), .Z(n14288) );
  AND U14659 ( .A(y[105]), .B(x[137]), .Z(n14287) );
  XOR U14660 ( .A(n14288), .B(n14287), .Z(n14310) );
  XOR U14661 ( .A(n14311), .B(n14310), .Z(n14261) );
  NAND U14662 ( .A(n14474), .B(n14247), .Z(n14251) );
  AND U14663 ( .A(n14249), .B(n14248), .Z(n14250) );
  ANDN U14664 ( .B(n14251), .A(n14250), .Z(n14270) );
  AND U14665 ( .A(x[153]), .B(y[185]), .Z(n14333) );
  NAND U14666 ( .A(x[154]), .B(y[184]), .Z(n14252) );
  XNOR U14667 ( .A(n14333), .B(n14252), .Z(n14307) );
  ANDN U14668 ( .B(n14254), .A(n14253), .Z(n14306) );
  XOR U14669 ( .A(n14307), .B(n14306), .Z(n14267) );
  AND U14670 ( .A(y[145]), .B(x[145]), .Z(n14279) );
  NAND U14671 ( .A(y[65]), .B(x[129]), .Z(n14280) );
  XNOR U14672 ( .A(n14279), .B(n14280), .Z(n14281) );
  NAND U14673 ( .A(y[66]), .B(x[128]), .Z(n14282) );
  XOR U14674 ( .A(n14281), .B(n14282), .Z(n14268) );
  XNOR U14675 ( .A(n14267), .B(n14268), .Z(n14269) );
  XOR U14676 ( .A(n14270), .B(n14269), .Z(n14262) );
  XNOR U14677 ( .A(n14261), .B(n14262), .Z(n14263) );
  XNOR U14678 ( .A(n14264), .B(n14263), .Z(n14257) );
  XNOR U14679 ( .A(n14258), .B(n14257), .Z(o[146]) );
  NANDN U14680 ( .A(n14256), .B(n14255), .Z(n14260) );
  NAND U14681 ( .A(n14258), .B(n14257), .Z(n14259) );
  AND U14682 ( .A(n14260), .B(n14259), .Z(n14399) );
  NANDN U14683 ( .A(n14262), .B(n14261), .Z(n14266) );
  NAND U14684 ( .A(n14264), .B(n14263), .Z(n14265) );
  AND U14685 ( .A(n14266), .B(n14265), .Z(n14384) );
  NANDN U14686 ( .A(n14268), .B(n14267), .Z(n14272) );
  NANDN U14687 ( .A(n14270), .B(n14269), .Z(n14271) );
  AND U14688 ( .A(n14272), .B(n14271), .Z(n14382) );
  NANDN U14689 ( .A(n14274), .B(n14273), .Z(n14278) );
  NANDN U14690 ( .A(n14276), .B(n14275), .Z(n14277) );
  NAND U14691 ( .A(n14278), .B(n14277), .Z(n14393) );
  NANDN U14692 ( .A(n14280), .B(n14279), .Z(n14284) );
  NANDN U14693 ( .A(n14282), .B(n14281), .Z(n14283) );
  AND U14694 ( .A(n14284), .B(n14283), .Z(n14349) );
  AND U14695 ( .A(y[147]), .B(x[144]), .Z(n14363) );
  AND U14696 ( .A(y[107]), .B(x[136]), .Z(n14362) );
  NAND U14697 ( .A(y[24]), .B(x[123]), .Z(n14361) );
  XOR U14698 ( .A(n14362), .B(n14361), .Z(n14364) );
  XOR U14699 ( .A(n14363), .B(n14364), .Z(n14347) );
  AND U14700 ( .A(x[138]), .B(y[105]), .Z(n14421) );
  NAND U14701 ( .A(x[139]), .B(y[104]), .Z(n14285) );
  XNOR U14702 ( .A(n14421), .B(n14285), .Z(n14369) );
  NAND U14703 ( .A(y[106]), .B(x[137]), .Z(n14370) );
  XNOR U14704 ( .A(n14369), .B(n14370), .Z(n14346) );
  XNOR U14705 ( .A(n14347), .B(n14346), .Z(n14348) );
  XNOR U14706 ( .A(n14349), .B(n14348), .Z(n14394) );
  XOR U14707 ( .A(n14393), .B(n14394), .Z(n14396) );
  NAND U14708 ( .A(n14368), .B(n14286), .Z(n14290) );
  AND U14709 ( .A(n14288), .B(n14287), .Z(n14289) );
  ANDN U14710 ( .B(n14290), .A(n14289), .Z(n14354) );
  AND U14711 ( .A(y[26]), .B(x[121]), .Z(n14324) );
  AND U14712 ( .A(y[25]), .B(x[122]), .Z(n14323) );
  NAND U14713 ( .A(y[146]), .B(x[145]), .Z(n14322) );
  XOR U14714 ( .A(n14323), .B(n14322), .Z(n14325) );
  XOR U14715 ( .A(n14324), .B(n14325), .Z(n14353) );
  AND U14716 ( .A(x[155]), .B(y[184]), .Z(n14292) );
  NAND U14717 ( .A(x[152]), .B(y[187]), .Z(n14291) );
  XNOR U14718 ( .A(n14292), .B(n14291), .Z(n14329) );
  AND U14719 ( .A(x[154]), .B(y[185]), .Z(n14438) );
  NAND U14720 ( .A(x[153]), .B(y[186]), .Z(n14293) );
  XOR U14721 ( .A(n14438), .B(n14293), .Z(n14330) );
  XNOR U14722 ( .A(n14329), .B(n14330), .Z(n14352) );
  XOR U14723 ( .A(n14353), .B(n14352), .Z(n14355) );
  XOR U14724 ( .A(n14354), .B(n14355), .Z(n14395) );
  XOR U14725 ( .A(n14396), .B(n14395), .Z(n14381) );
  XNOR U14726 ( .A(n14382), .B(n14381), .Z(n14383) );
  XOR U14727 ( .A(n14384), .B(n14383), .Z(n14400) );
  XNOR U14728 ( .A(n14399), .B(n14400), .Z(n14402) );
  NANDN U14729 ( .A(n14295), .B(n14294), .Z(n14299) );
  OR U14730 ( .A(n14297), .B(n14296), .Z(n14298) );
  AND U14731 ( .A(n14299), .B(n14298), .Z(n14390) );
  NANDN U14732 ( .A(n14301), .B(n14300), .Z(n14305) );
  NANDN U14733 ( .A(n14303), .B(n14302), .Z(n14304) );
  AND U14734 ( .A(n14305), .B(n14304), .Z(n14315) );
  XNOR U14735 ( .A(n14315), .B(n14314), .Z(n14317) );
  AND U14736 ( .A(y[64]), .B(x[131]), .Z(n14377) );
  AND U14737 ( .A(y[27]), .B(x[120]), .Z(n14376) );
  NAND U14738 ( .A(y[145]), .B(x[146]), .Z(n14375) );
  XOR U14739 ( .A(n14376), .B(n14375), .Z(n14378) );
  XOR U14740 ( .A(n14377), .B(n14378), .Z(n14343) );
  AND U14741 ( .A(y[67]), .B(x[128]), .Z(n14336) );
  AND U14742 ( .A(y[65]), .B(x[130]), .Z(n14335) );
  NAND U14743 ( .A(y[144]), .B(x[147]), .Z(n14334) );
  XOR U14744 ( .A(n14335), .B(n14334), .Z(n14337) );
  XOR U14745 ( .A(n14336), .B(n14337), .Z(n14341) );
  AND U14746 ( .A(y[66]), .B(x[129]), .Z(n14340) );
  XNOR U14747 ( .A(n14341), .B(n14340), .Z(n14342) );
  XNOR U14748 ( .A(n14343), .B(n14342), .Z(n14316) );
  XOR U14749 ( .A(n14317), .B(n14316), .Z(n14388) );
  NAND U14750 ( .A(n14309), .B(n14308), .Z(n14313) );
  NAND U14751 ( .A(n14311), .B(n14310), .Z(n14312) );
  AND U14752 ( .A(n14313), .B(n14312), .Z(n14387) );
  XNOR U14753 ( .A(n14388), .B(n14387), .Z(n14389) );
  XNOR U14754 ( .A(n14390), .B(n14389), .Z(n14401) );
  XOR U14755 ( .A(n14402), .B(n14401), .Z(o[147]) );
  NANDN U14756 ( .A(n14315), .B(n14314), .Z(n14319) );
  NAND U14757 ( .A(n14317), .B(n14316), .Z(n14318) );
  AND U14758 ( .A(n14319), .B(n14318), .Z(n14416) );
  AND U14759 ( .A(x[128]), .B(y[68]), .Z(n14321) );
  NAND U14760 ( .A(x[131]), .B(y[65]), .Z(n14320) );
  XNOR U14761 ( .A(n14321), .B(n14320), .Z(n14475) );
  NAND U14762 ( .A(y[66]), .B(x[130]), .Z(n14549) );
  XNOR U14763 ( .A(n14475), .B(n14549), .Z(n14484) );
  NAND U14764 ( .A(y[67]), .B(x[129]), .Z(n14485) );
  XNOR U14765 ( .A(n14484), .B(n14485), .Z(n14487) );
  AND U14766 ( .A(y[144]), .B(x[148]), .Z(n14426) );
  NAND U14767 ( .A(y[27]), .B(x[121]), .Z(n14427) );
  XNOR U14768 ( .A(n14426), .B(n14427), .Z(n14428) );
  NAND U14769 ( .A(y[28]), .B(x[120]), .Z(n14429) );
  XNOR U14770 ( .A(n14428), .B(n14429), .Z(n14486) );
  XOR U14771 ( .A(n14487), .B(n14486), .Z(n14481) );
  NANDN U14772 ( .A(n14323), .B(n14322), .Z(n14327) );
  OR U14773 ( .A(n14325), .B(n14324), .Z(n14326) );
  AND U14774 ( .A(n14327), .B(n14326), .Z(n14479) );
  AND U14775 ( .A(y[187]), .B(x[155]), .Z(n14695) );
  NANDN U14776 ( .A(n14328), .B(n14695), .Z(n14332) );
  NANDN U14777 ( .A(n14330), .B(n14329), .Z(n14331) );
  AND U14778 ( .A(n14332), .B(n14331), .Z(n14478) );
  XNOR U14779 ( .A(n14479), .B(n14478), .Z(n14480) );
  XNOR U14780 ( .A(n14481), .B(n14480), .Z(n14511) );
  NAND U14781 ( .A(y[24]), .B(x[124]), .Z(n14460) );
  AND U14782 ( .A(y[146]), .B(x[146]), .Z(n14459) );
  NAND U14783 ( .A(y[108]), .B(x[136]), .Z(n14458) );
  XOR U14784 ( .A(n14459), .B(n14458), .Z(n14461) );
  XOR U14785 ( .A(n14460), .B(n14461), .Z(n14441) );
  AND U14786 ( .A(x[154]), .B(y[186]), .Z(n14360) );
  NAND U14787 ( .A(n14360), .B(n14333), .Z(n14456) );
  NAND U14788 ( .A(y[104]), .B(x[140]), .Z(n14570) );
  NAND U14789 ( .A(y[188]), .B(x[152]), .Z(n14626) );
  XNOR U14790 ( .A(n14570), .B(n14626), .Z(n14457) );
  XOR U14791 ( .A(n14456), .B(n14457), .Z(n14442) );
  XOR U14792 ( .A(n14441), .B(n14442), .Z(n14444) );
  NANDN U14793 ( .A(n14335), .B(n14334), .Z(n14339) );
  OR U14794 ( .A(n14337), .B(n14336), .Z(n14338) );
  AND U14795 ( .A(n14339), .B(n14338), .Z(n14443) );
  XOR U14796 ( .A(n14444), .B(n14443), .Z(n14509) );
  NANDN U14797 ( .A(n14341), .B(n14340), .Z(n14345) );
  NANDN U14798 ( .A(n14343), .B(n14342), .Z(n14344) );
  AND U14799 ( .A(n14345), .B(n14344), .Z(n14508) );
  XNOR U14800 ( .A(n14509), .B(n14508), .Z(n14510) );
  XNOR U14801 ( .A(n14511), .B(n14510), .Z(n14415) );
  XNOR U14802 ( .A(n14416), .B(n14415), .Z(n14418) );
  NANDN U14803 ( .A(n14347), .B(n14346), .Z(n14351) );
  NANDN U14804 ( .A(n14349), .B(n14348), .Z(n14350) );
  AND U14805 ( .A(n14351), .B(n14350), .Z(n14497) );
  NANDN U14806 ( .A(n14353), .B(n14352), .Z(n14357) );
  OR U14807 ( .A(n14355), .B(n14354), .Z(n14356) );
  NAND U14808 ( .A(n14357), .B(n14356), .Z(n14496) );
  XNOR U14809 ( .A(n14497), .B(n14496), .Z(n14498) );
  NAND U14810 ( .A(y[26]), .B(x[122]), .Z(n14470) );
  NAND U14811 ( .A(y[145]), .B(x[147]), .Z(n14469) );
  NAND U14812 ( .A(y[25]), .B(x[123]), .Z(n14468) );
  XNOR U14813 ( .A(n14469), .B(n14468), .Z(n14471) );
  AND U14814 ( .A(x[156]), .B(y[184]), .Z(n14359) );
  NAND U14815 ( .A(x[153]), .B(y[187]), .Z(n14358) );
  XNOR U14816 ( .A(n14359), .B(n14358), .Z(n14452) );
  AND U14817 ( .A(y[185]), .B(x[155]), .Z(n14578) );
  XNOR U14818 ( .A(n14578), .B(n14360), .Z(n14453) );
  XNOR U14819 ( .A(n14452), .B(n14453), .Z(n14445) );
  XOR U14820 ( .A(n14446), .B(n14445), .Z(n14447) );
  NANDN U14821 ( .A(n14362), .B(n14361), .Z(n14366) );
  OR U14822 ( .A(n14364), .B(n14363), .Z(n14365) );
  NAND U14823 ( .A(n14366), .B(n14365), .Z(n14448) );
  XNOR U14824 ( .A(n14447), .B(n14448), .Z(n14504) );
  AND U14825 ( .A(y[105]), .B(x[139]), .Z(n14367) );
  NAND U14826 ( .A(n14368), .B(n14367), .Z(n14372) );
  NANDN U14827 ( .A(n14370), .B(n14369), .Z(n14371) );
  AND U14828 ( .A(n14372), .B(n14371), .Z(n14503) );
  AND U14829 ( .A(y[64]), .B(x[132]), .Z(n14432) );
  NAND U14830 ( .A(y[148]), .B(x[144]), .Z(n14433) );
  XNOR U14831 ( .A(n14432), .B(n14433), .Z(n14434) );
  NAND U14832 ( .A(y[147]), .B(x[145]), .Z(n14435) );
  XNOR U14833 ( .A(n14434), .B(n14435), .Z(n14490) );
  AND U14834 ( .A(x[138]), .B(y[106]), .Z(n14374) );
  NAND U14835 ( .A(x[139]), .B(y[105]), .Z(n14373) );
  XNOR U14836 ( .A(n14374), .B(n14373), .Z(n14422) );
  NAND U14837 ( .A(y[107]), .B(x[137]), .Z(n14423) );
  XOR U14838 ( .A(n14422), .B(n14423), .Z(n14491) );
  XNOR U14839 ( .A(n14490), .B(n14491), .Z(n14492) );
  NANDN U14840 ( .A(n14376), .B(n14375), .Z(n14380) );
  OR U14841 ( .A(n14378), .B(n14377), .Z(n14379) );
  NAND U14842 ( .A(n14380), .B(n14379), .Z(n14493) );
  XNOR U14843 ( .A(n14492), .B(n14493), .Z(n14502) );
  XOR U14844 ( .A(n14503), .B(n14502), .Z(n14505) );
  XOR U14845 ( .A(n14504), .B(n14505), .Z(n14499) );
  XNOR U14846 ( .A(n14498), .B(n14499), .Z(n14417) );
  XNOR U14847 ( .A(n14418), .B(n14417), .Z(n14408) );
  NANDN U14848 ( .A(n14382), .B(n14381), .Z(n14386) );
  NANDN U14849 ( .A(n14384), .B(n14383), .Z(n14385) );
  AND U14850 ( .A(n14386), .B(n14385), .Z(n14411) );
  NANDN U14851 ( .A(n14388), .B(n14387), .Z(n14392) );
  NAND U14852 ( .A(n14390), .B(n14389), .Z(n14391) );
  NAND U14853 ( .A(n14392), .B(n14391), .Z(n14409) );
  NAND U14854 ( .A(n14394), .B(n14393), .Z(n14398) );
  NAND U14855 ( .A(n14396), .B(n14395), .Z(n14397) );
  AND U14856 ( .A(n14398), .B(n14397), .Z(n14410) );
  XNOR U14857 ( .A(n14409), .B(n14410), .Z(n14412) );
  NANDN U14858 ( .A(n14400), .B(n14399), .Z(n14404) );
  NAND U14859 ( .A(n14402), .B(n14401), .Z(n14403) );
  NAND U14860 ( .A(n14404), .B(n14403), .Z(n14406) );
  XNOR U14861 ( .A(n14407), .B(n14406), .Z(n14405) );
  XNOR U14862 ( .A(n14408), .B(n14405), .Z(o[148]) );
  NAND U14863 ( .A(n14410), .B(n14409), .Z(n14414) );
  NANDN U14864 ( .A(n14412), .B(n14411), .Z(n14413) );
  AND U14865 ( .A(n14414), .B(n14413), .Z(n14657) );
  XNOR U14866 ( .A(n14658), .B(n14657), .Z(n14660) );
  NANDN U14867 ( .A(n14416), .B(n14415), .Z(n14420) );
  NAND U14868 ( .A(n14418), .B(n14417), .Z(n14419) );
  AND U14869 ( .A(n14420), .B(n14419), .Z(n14652) );
  AND U14870 ( .A(y[106]), .B(x[139]), .Z(n14571) );
  NAND U14871 ( .A(n14421), .B(n14571), .Z(n14425) );
  NANDN U14872 ( .A(n14423), .B(n14422), .Z(n14424) );
  NAND U14873 ( .A(n14425), .B(n14424), .Z(n14579) );
  NANDN U14874 ( .A(n14427), .B(n14426), .Z(n14431) );
  NANDN U14875 ( .A(n14429), .B(n14428), .Z(n14430) );
  AND U14876 ( .A(n14431), .B(n14430), .Z(n14557) );
  AND U14877 ( .A(y[64]), .B(x[133]), .Z(n14561) );
  AND U14878 ( .A(y[107]), .B(x[138]), .Z(n14560) );
  XOR U14879 ( .A(n14561), .B(n14560), .Z(n14562) );
  AND U14880 ( .A(y[149]), .B(x[144]), .Z(n14834) );
  XOR U14881 ( .A(n14562), .B(n14834), .Z(n14554) );
  AND U14882 ( .A(y[145]), .B(x[148]), .Z(n14566) );
  AND U14883 ( .A(y[24]), .B(x[125]), .Z(n14565) );
  XOR U14884 ( .A(n14566), .B(n14565), .Z(n14567) );
  AND U14885 ( .A(y[25]), .B(x[124]), .Z(n14822) );
  XNOR U14886 ( .A(n14567), .B(n14822), .Z(n14555) );
  XNOR U14887 ( .A(n14554), .B(n14555), .Z(n14556) );
  XNOR U14888 ( .A(n14557), .B(n14556), .Z(n14580) );
  XOR U14889 ( .A(n14579), .B(n14580), .Z(n14581) );
  NANDN U14890 ( .A(n14433), .B(n14432), .Z(n14437) );
  NANDN U14891 ( .A(n14435), .B(n14434), .Z(n14436) );
  NAND U14892 ( .A(n14437), .B(n14436), .Z(n14617) );
  AND U14893 ( .A(x[155]), .B(y[186]), .Z(n14465) );
  AND U14894 ( .A(n14465), .B(n14438), .Z(n14628) );
  AND U14895 ( .A(x[152]), .B(y[189]), .Z(n14440) );
  AND U14896 ( .A(x[153]), .B(y[188]), .Z(n14439) );
  XOR U14897 ( .A(n14440), .B(n14439), .Z(n14627) );
  XOR U14898 ( .A(n14628), .B(n14627), .Z(n14616) );
  AND U14899 ( .A(y[65]), .B(x[132]), .Z(n14608) );
  AND U14900 ( .A(y[69]), .B(x[128]), .Z(n14606) );
  AND U14901 ( .A(y[28]), .B(x[121]), .Z(n14605) );
  XOR U14902 ( .A(n14606), .B(n14605), .Z(n14607) );
  XOR U14903 ( .A(n14608), .B(n14607), .Z(n14615) );
  XOR U14904 ( .A(n14616), .B(n14615), .Z(n14618) );
  XNOR U14905 ( .A(n14617), .B(n14618), .Z(n14582) );
  NAND U14906 ( .A(n14446), .B(n14445), .Z(n14450) );
  NANDN U14907 ( .A(n14448), .B(n14447), .Z(n14449) );
  NAND U14908 ( .A(n14450), .B(n14449), .Z(n14514) );
  XOR U14909 ( .A(n14515), .B(n14514), .Z(n14517) );
  XNOR U14910 ( .A(n14516), .B(n14517), .Z(n14647) );
  AND U14911 ( .A(y[187]), .B(x[156]), .Z(n14848) );
  NAND U14912 ( .A(n14848), .B(n14451), .Z(n14455) );
  NANDN U14913 ( .A(n14453), .B(n14452), .Z(n14454) );
  AND U14914 ( .A(n14455), .B(n14454), .Z(n14525) );
  XNOR U14915 ( .A(n14525), .B(n14524), .Z(n14527) );
  NANDN U14916 ( .A(n14459), .B(n14458), .Z(n14463) );
  NANDN U14917 ( .A(n14461), .B(n14460), .Z(n14462) );
  AND U14918 ( .A(n14463), .B(n14462), .Z(n14533) );
  AND U14919 ( .A(y[66]), .B(x[131]), .Z(n14768) );
  NAND U14920 ( .A(x[130]), .B(y[67]), .Z(n14464) );
  XNOR U14921 ( .A(n14768), .B(n14464), .Z(n14551) );
  AND U14922 ( .A(y[68]), .B(x[129]), .Z(n14550) );
  XOR U14923 ( .A(n14551), .B(n14550), .Z(n14531) );
  AND U14924 ( .A(y[187]), .B(x[154]), .Z(n14537) );
  AND U14925 ( .A(y[184]), .B(x[157]), .Z(n14536) );
  XOR U14926 ( .A(n14537), .B(n14536), .Z(n14539) );
  AND U14927 ( .A(y[185]), .B(x[156]), .Z(n14830) );
  XOR U14928 ( .A(n14830), .B(n14465), .Z(n14538) );
  XOR U14929 ( .A(n14539), .B(n14538), .Z(n14530) );
  XOR U14930 ( .A(n14531), .B(n14530), .Z(n14532) );
  XOR U14931 ( .A(n14533), .B(n14532), .Z(n14526) );
  XOR U14932 ( .A(n14527), .B(n14526), .Z(n14593) );
  AND U14933 ( .A(x[140]), .B(y[105]), .Z(n14467) );
  NAND U14934 ( .A(x[141]), .B(y[104]), .Z(n14466) );
  XOR U14935 ( .A(n14467), .B(n14466), .Z(n14572) );
  XNOR U14936 ( .A(n14571), .B(n14572), .Z(n14598) );
  AND U14937 ( .A(y[144]), .B(x[149]), .Z(n14542) );
  NAND U14938 ( .A(y[26]), .B(x[123]), .Z(n14543) );
  XNOR U14939 ( .A(n14542), .B(n14543), .Z(n14545) );
  AND U14940 ( .A(y[27]), .B(x[122]), .Z(n14544) );
  XOR U14941 ( .A(n14545), .B(n14544), .Z(n14597) );
  XOR U14942 ( .A(n14598), .B(n14597), .Z(n14600) );
  NAND U14943 ( .A(n14469), .B(n14468), .Z(n14473) );
  NANDN U14944 ( .A(n14471), .B(n14470), .Z(n14472) );
  AND U14945 ( .A(n14473), .B(n14472), .Z(n14599) );
  XOR U14946 ( .A(n14600), .B(n14599), .Z(n14592) );
  AND U14947 ( .A(y[68]), .B(x[131]), .Z(n14847) );
  NAND U14948 ( .A(n14847), .B(n14474), .Z(n14477) );
  NANDN U14949 ( .A(n14549), .B(n14475), .Z(n14476) );
  AND U14950 ( .A(n14477), .B(n14476), .Z(n14523) );
  AND U14951 ( .A(y[146]), .B(x[147]), .Z(n14621) );
  AND U14952 ( .A(y[108]), .B(x[137]), .Z(n14862) );
  XOR U14953 ( .A(n14621), .B(n14862), .Z(n14623) );
  AND U14954 ( .A(y[109]), .B(x[136]), .Z(n14622) );
  XOR U14955 ( .A(n14623), .B(n14622), .Z(n14521) );
  AND U14956 ( .A(y[29]), .B(x[120]), .Z(n14632) );
  AND U14957 ( .A(y[148]), .B(x[145]), .Z(n14631) );
  XOR U14958 ( .A(n14632), .B(n14631), .Z(n14634) );
  AND U14959 ( .A(y[147]), .B(x[146]), .Z(n14633) );
  XOR U14960 ( .A(n14634), .B(n14633), .Z(n14520) );
  XOR U14961 ( .A(n14521), .B(n14520), .Z(n14522) );
  XOR U14962 ( .A(n14523), .B(n14522), .Z(n14591) );
  XOR U14963 ( .A(n14592), .B(n14591), .Z(n14594) );
  XOR U14964 ( .A(n14593), .B(n14594), .Z(n14646) );
  NANDN U14965 ( .A(n14479), .B(n14478), .Z(n14483) );
  NANDN U14966 ( .A(n14481), .B(n14480), .Z(n14482) );
  AND U14967 ( .A(n14483), .B(n14482), .Z(n14587) );
  NANDN U14968 ( .A(n14485), .B(n14484), .Z(n14489) );
  NAND U14969 ( .A(n14487), .B(n14486), .Z(n14488) );
  AND U14970 ( .A(n14489), .B(n14488), .Z(n14586) );
  NANDN U14971 ( .A(n14491), .B(n14490), .Z(n14495) );
  NANDN U14972 ( .A(n14493), .B(n14492), .Z(n14494) );
  NAND U14973 ( .A(n14495), .B(n14494), .Z(n14585) );
  XOR U14974 ( .A(n14586), .B(n14585), .Z(n14588) );
  XNOR U14975 ( .A(n14587), .B(n14588), .Z(n14645) );
  XOR U14976 ( .A(n14646), .B(n14645), .Z(n14648) );
  XNOR U14977 ( .A(n14647), .B(n14648), .Z(n14651) );
  XNOR U14978 ( .A(n14652), .B(n14651), .Z(n14653) );
  NANDN U14979 ( .A(n14497), .B(n14496), .Z(n14501) );
  NANDN U14980 ( .A(n14499), .B(n14498), .Z(n14500) );
  AND U14981 ( .A(n14501), .B(n14500), .Z(n14642) );
  NANDN U14982 ( .A(n14503), .B(n14502), .Z(n14507) );
  NANDN U14983 ( .A(n14505), .B(n14504), .Z(n14506) );
  AND U14984 ( .A(n14507), .B(n14506), .Z(n14640) );
  NANDN U14985 ( .A(n14509), .B(n14508), .Z(n14513) );
  NAND U14986 ( .A(n14511), .B(n14510), .Z(n14512) );
  AND U14987 ( .A(n14513), .B(n14512), .Z(n14639) );
  XNOR U14988 ( .A(n14640), .B(n14639), .Z(n14641) );
  XOR U14989 ( .A(n14642), .B(n14641), .Z(n14654) );
  XNOR U14990 ( .A(n14653), .B(n14654), .Z(n14659) );
  XOR U14991 ( .A(n14660), .B(n14659), .Z(o[149]) );
  NANDN U14992 ( .A(n14515), .B(n14514), .Z(n14519) );
  NANDN U14993 ( .A(n14517), .B(n14516), .Z(n14518) );
  NAND U14994 ( .A(n14519), .B(n14518), .Z(n14664) );
  NANDN U14995 ( .A(n14525), .B(n14524), .Z(n14529) );
  NAND U14996 ( .A(n14527), .B(n14526), .Z(n14528) );
  AND U14997 ( .A(n14529), .B(n14528), .Z(n14670) );
  XOR U14998 ( .A(n14671), .B(n14670), .Z(n14669) );
  NAND U14999 ( .A(n14531), .B(n14530), .Z(n14535) );
  NAND U15000 ( .A(n14533), .B(n14532), .Z(n14534) );
  AND U15001 ( .A(n14535), .B(n14534), .Z(n14668) );
  XOR U15002 ( .A(n14669), .B(n14668), .Z(n14667) );
  NAND U15003 ( .A(n14537), .B(n14536), .Z(n14541) );
  NAND U15004 ( .A(n14539), .B(n14538), .Z(n14540) );
  NAND U15005 ( .A(n14541), .B(n14540), .Z(n14801) );
  NANDN U15006 ( .A(n14543), .B(n14542), .Z(n14547) );
  NAND U15007 ( .A(n14545), .B(n14544), .Z(n14546) );
  NAND U15008 ( .A(n14547), .B(n14546), .Z(n14804) );
  AND U15009 ( .A(y[67]), .B(x[131]), .Z(n14548) );
  NANDN U15010 ( .A(n14549), .B(n14548), .Z(n14553) );
  NAND U15011 ( .A(n14551), .B(n14550), .Z(n14552) );
  AND U15012 ( .A(n14553), .B(n14552), .Z(n14808) );
  AND U15013 ( .A(y[147]), .B(x[147]), .Z(n14774) );
  AND U15014 ( .A(y[107]), .B(x[139]), .Z(n14773) );
  XOR U15015 ( .A(n14774), .B(n14773), .Z(n14772) );
  AND U15016 ( .A(y[27]), .B(x[123]), .Z(n14771) );
  XOR U15017 ( .A(n14772), .B(n14771), .Z(n14810) );
  AND U15018 ( .A(y[148]), .B(x[146]), .Z(n14876) );
  AND U15019 ( .A(y[106]), .B(x[140]), .Z(n14875) );
  XOR U15020 ( .A(n14876), .B(n14875), .Z(n14874) );
  AND U15021 ( .A(y[28]), .B(x[122]), .Z(n14873) );
  XNOR U15022 ( .A(n14874), .B(n14873), .Z(n14809) );
  XNOR U15023 ( .A(n14808), .B(n14807), .Z(n14803) );
  XOR U15024 ( .A(n14804), .B(n14803), .Z(n14802) );
  XOR U15025 ( .A(n14801), .B(n14802), .Z(n14675) );
  NANDN U15026 ( .A(n14555), .B(n14554), .Z(n14559) );
  NANDN U15027 ( .A(n14557), .B(n14556), .Z(n14558) );
  NAND U15028 ( .A(n14559), .B(n14558), .Z(n14674) );
  XOR U15029 ( .A(n14675), .B(n14674), .Z(n14673) );
  NAND U15030 ( .A(n14561), .B(n14560), .Z(n14564) );
  NAND U15031 ( .A(n14562), .B(n14834), .Z(n14563) );
  NAND U15032 ( .A(n14564), .B(n14563), .Z(n14687) );
  NAND U15033 ( .A(n14566), .B(n14565), .Z(n14569) );
  NAND U15034 ( .A(n14567), .B(n14822), .Z(n14568) );
  NAND U15035 ( .A(n14569), .B(n14568), .Z(n14686) );
  XOR U15036 ( .A(n14687), .B(n14686), .Z(n14685) );
  AND U15037 ( .A(y[105]), .B(x[141]), .Z(n14816) );
  NANDN U15038 ( .A(n14570), .B(n14816), .Z(n14574) );
  NANDN U15039 ( .A(n14572), .B(n14571), .Z(n14573) );
  AND U15040 ( .A(n14574), .B(n14573), .Z(n14898) );
  AND U15041 ( .A(x[125]), .B(y[25]), .Z(n14576) );
  NAND U15042 ( .A(x[124]), .B(y[26]), .Z(n14575) );
  XNOR U15043 ( .A(n14576), .B(n14575), .Z(n14820) );
  AND U15044 ( .A(y[144]), .B(x[150]), .Z(n14819) );
  XOR U15045 ( .A(n14820), .B(n14819), .Z(n14895) );
  AND U15046 ( .A(y[189]), .B(x[153]), .Z(n14786) );
  AND U15047 ( .A(y[186]), .B(x[156]), .Z(n14577) );
  AND U15048 ( .A(n14578), .B(n14577), .Z(n14788) );
  AND U15049 ( .A(y[188]), .B(x[154]), .Z(n14787) );
  XOR U15050 ( .A(n14788), .B(n14787), .Z(n14785) );
  XNOR U15051 ( .A(n14786), .B(n14785), .Z(n14896) );
  XNOR U15052 ( .A(n14898), .B(n14897), .Z(n14684) );
  XOR U15053 ( .A(n14685), .B(n14684), .Z(n14672) );
  XOR U15054 ( .A(n14673), .B(n14672), .Z(n14666) );
  XOR U15055 ( .A(n14664), .B(n14665), .Z(n14926) );
  NAND U15056 ( .A(n14580), .B(n14579), .Z(n14584) );
  NANDN U15057 ( .A(n14582), .B(n14581), .Z(n14583) );
  AND U15058 ( .A(n14584), .B(n14583), .Z(n14925) );
  NANDN U15059 ( .A(n14586), .B(n14585), .Z(n14590) );
  NANDN U15060 ( .A(n14588), .B(n14587), .Z(n14589) );
  AND U15061 ( .A(n14590), .B(n14589), .Z(n14908) );
  NANDN U15062 ( .A(n14592), .B(n14591), .Z(n14596) );
  OR U15063 ( .A(n14594), .B(n14593), .Z(n14595) );
  NAND U15064 ( .A(n14596), .B(n14595), .Z(n14909) );
  NAND U15065 ( .A(n14598), .B(n14597), .Z(n14602) );
  NAND U15066 ( .A(n14600), .B(n14599), .Z(n14601) );
  AND U15067 ( .A(n14602), .B(n14601), .Z(n14914) );
  AND U15068 ( .A(y[110]), .B(x[136]), .Z(n14782) );
  AND U15069 ( .A(y[24]), .B(x[126]), .Z(n14781) );
  XOR U15070 ( .A(n14782), .B(n14781), .Z(n14780) );
  AND U15071 ( .A(y[145]), .B(x[149]), .Z(n14779) );
  XOR U15072 ( .A(n14780), .B(n14779), .Z(n14691) );
  AND U15073 ( .A(y[65]), .B(x[133]), .Z(n14870) );
  AND U15074 ( .A(y[68]), .B(x[130]), .Z(n14869) );
  XOR U15075 ( .A(n14870), .B(n14869), .Z(n14868) );
  AND U15076 ( .A(y[69]), .B(x[129]), .Z(n14867) );
  XOR U15077 ( .A(n14868), .B(n14867), .Z(n14766) );
  AND U15078 ( .A(x[132]), .B(y[66]), .Z(n14604) );
  NAND U15079 ( .A(x[131]), .B(y[67]), .Z(n14603) );
  XNOR U15080 ( .A(n14604), .B(n14603), .Z(n14765) );
  XOR U15081 ( .A(n14766), .B(n14765), .Z(n14690) );
  XOR U15082 ( .A(n14691), .B(n14690), .Z(n14689) );
  AND U15083 ( .A(y[190]), .B(x[152]), .Z(n14815) );
  XOR U15084 ( .A(n14816), .B(n14815), .Z(n14814) );
  AND U15085 ( .A(y[104]), .B(x[142]), .Z(n14813) );
  XOR U15086 ( .A(n14814), .B(n14813), .Z(n14688) );
  XOR U15087 ( .A(n14689), .B(n14688), .Z(n14680) );
  NAND U15088 ( .A(n14606), .B(n14605), .Z(n14610) );
  NAND U15089 ( .A(n14608), .B(n14607), .Z(n14609) );
  AND U15090 ( .A(n14610), .B(n14609), .Z(n14759) );
  AND U15091 ( .A(y[146]), .B(x[148]), .Z(n14860) );
  AND U15092 ( .A(x[137]), .B(y[109]), .Z(n14612) );
  AND U15093 ( .A(x[138]), .B(y[108]), .Z(n14611) );
  XOR U15094 ( .A(n14612), .B(n14611), .Z(n14859) );
  XOR U15095 ( .A(n14860), .B(n14859), .Z(n14762) );
  AND U15096 ( .A(y[30]), .B(x[120]), .Z(n14832) );
  AND U15097 ( .A(y[150]), .B(x[144]), .Z(n14614) );
  AND U15098 ( .A(x[145]), .B(y[149]), .Z(n14613) );
  XOR U15099 ( .A(n14614), .B(n14613), .Z(n14831) );
  XNOR U15100 ( .A(n14832), .B(n14831), .Z(n14761) );
  XNOR U15101 ( .A(n14759), .B(n14760), .Z(n14681) );
  XNOR U15102 ( .A(n14680), .B(n14681), .Z(n14683) );
  NAND U15103 ( .A(n14616), .B(n14615), .Z(n14620) );
  NAND U15104 ( .A(n14618), .B(n14617), .Z(n14619) );
  AND U15105 ( .A(n14620), .B(n14619), .Z(n14682) );
  XOR U15106 ( .A(n14683), .B(n14682), .Z(n14913) );
  XOR U15107 ( .A(n14914), .B(n14913), .Z(n14916) );
  NAND U15108 ( .A(n14621), .B(n14862), .Z(n14625) );
  NAND U15109 ( .A(n14623), .B(n14622), .Z(n14624) );
  NAND U15110 ( .A(n14625), .B(n14624), .Z(n14676) );
  NANDN U15111 ( .A(n14626), .B(n14786), .Z(n14630) );
  NAND U15112 ( .A(n14628), .B(n14627), .Z(n14629) );
  NAND U15113 ( .A(n14630), .B(n14629), .Z(n14679) );
  NAND U15114 ( .A(n14632), .B(n14631), .Z(n14636) );
  NAND U15115 ( .A(n14634), .B(n14633), .Z(n14635) );
  AND U15116 ( .A(n14636), .B(n14635), .Z(n14890) );
  AND U15117 ( .A(y[29]), .B(x[121]), .Z(n14856) );
  AND U15118 ( .A(y[64]), .B(x[134]), .Z(n14855) );
  XOR U15119 ( .A(n14856), .B(n14855), .Z(n14854) );
  AND U15120 ( .A(y[70]), .B(x[128]), .Z(n14853) );
  XOR U15121 ( .A(n14854), .B(n14853), .Z(n14891) );
  AND U15122 ( .A(x[157]), .B(y[185]), .Z(n14638) );
  NAND U15123 ( .A(x[156]), .B(y[186]), .Z(n14637) );
  XNOR U15124 ( .A(n14638), .B(n14637), .Z(n14697) );
  AND U15125 ( .A(y[184]), .B(x[158]), .Z(n14696) );
  XOR U15126 ( .A(n14697), .B(n14696), .Z(n14694) );
  XNOR U15127 ( .A(n14695), .B(n14694), .Z(n14892) );
  XNOR U15128 ( .A(n14890), .B(n14889), .Z(n14678) );
  XOR U15129 ( .A(n14679), .B(n14678), .Z(n14677) );
  XOR U15130 ( .A(n14676), .B(n14677), .Z(n14915) );
  XOR U15131 ( .A(n14909), .B(n14910), .Z(n14907) );
  XOR U15132 ( .A(n14908), .B(n14907), .Z(n14923) );
  XOR U15133 ( .A(n14924), .B(n14923), .Z(n14929) );
  NANDN U15134 ( .A(n14640), .B(n14639), .Z(n14644) );
  NANDN U15135 ( .A(n14642), .B(n14641), .Z(n14643) );
  NAND U15136 ( .A(n14644), .B(n14643), .Z(n14932) );
  NANDN U15137 ( .A(n14646), .B(n14645), .Z(n14650) );
  NANDN U15138 ( .A(n14648), .B(n14647), .Z(n14649) );
  NAND U15139 ( .A(n14650), .B(n14649), .Z(n14931) );
  XNOR U15140 ( .A(n14932), .B(n14931), .Z(n14930) );
  XNOR U15141 ( .A(n14929), .B(n14930), .Z(n14937) );
  NANDN U15142 ( .A(n14652), .B(n14651), .Z(n14656) );
  NANDN U15143 ( .A(n14654), .B(n14653), .Z(n14655) );
  AND U15144 ( .A(n14656), .B(n14655), .Z(n14936) );
  NANDN U15145 ( .A(n14658), .B(n14657), .Z(n14662) );
  NAND U15146 ( .A(n14660), .B(n14659), .Z(n14661) );
  AND U15147 ( .A(n14662), .B(n14661), .Z(n14935) );
  XOR U15148 ( .A(n14936), .B(n14935), .Z(n14663) );
  XNOR U15149 ( .A(n14937), .B(n14663), .Z(o[150]) );
  NAND U15150 ( .A(n14689), .B(n14688), .Z(n14693) );
  NAND U15151 ( .A(n14691), .B(n14690), .Z(n14692) );
  AND U15152 ( .A(n14693), .B(n14692), .Z(n14800) );
  NAND U15153 ( .A(n14695), .B(n14694), .Z(n14699) );
  NAND U15154 ( .A(n14697), .B(n14696), .Z(n14698) );
  AND U15155 ( .A(n14699), .B(n14698), .Z(n14758) );
  AND U15156 ( .A(x[120]), .B(y[31]), .Z(n14701) );
  NAND U15157 ( .A(x[153]), .B(y[190]), .Z(n14700) );
  XNOR U15158 ( .A(n14701), .B(n14700), .Z(n14705) );
  AND U15159 ( .A(x[152]), .B(y[191]), .Z(n14703) );
  NAND U15160 ( .A(x[143]), .B(y[104]), .Z(n14702) );
  XNOR U15161 ( .A(n14703), .B(n14702), .Z(n14704) );
  XOR U15162 ( .A(n14705), .B(n14704), .Z(n14713) );
  AND U15163 ( .A(x[126]), .B(y[25]), .Z(n14707) );
  NAND U15164 ( .A(x[142]), .B(y[105]), .Z(n14706) );
  XNOR U15165 ( .A(n14707), .B(n14706), .Z(n14711) );
  AND U15166 ( .A(x[127]), .B(y[24]), .Z(n14709) );
  NAND U15167 ( .A(x[148]), .B(y[147]), .Z(n14708) );
  XNOR U15168 ( .A(n14709), .B(n14708), .Z(n14710) );
  XNOR U15169 ( .A(n14711), .B(n14710), .Z(n14712) );
  XNOR U15170 ( .A(n14713), .B(n14712), .Z(n14756) );
  AND U15171 ( .A(x[140]), .B(y[107]), .Z(n14718) );
  AND U15172 ( .A(y[186]), .B(x[157]), .Z(n14829) );
  AND U15173 ( .A(x[136]), .B(y[111]), .Z(n14715) );
  NAND U15174 ( .A(x[151]), .B(y[144]), .Z(n14714) );
  XNOR U15175 ( .A(n14715), .B(n14714), .Z(n14716) );
  XNOR U15176 ( .A(n14829), .B(n14716), .Z(n14717) );
  XNOR U15177 ( .A(n14718), .B(n14717), .Z(n14734) );
  AND U15178 ( .A(x[122]), .B(y[29]), .Z(n14720) );
  NAND U15179 ( .A(x[150]), .B(y[145]), .Z(n14719) );
  XNOR U15180 ( .A(n14720), .B(n14719), .Z(n14724) );
  AND U15181 ( .A(x[123]), .B(y[28]), .Z(n14722) );
  NAND U15182 ( .A(x[134]), .B(y[65]), .Z(n14721) );
  XNOR U15183 ( .A(n14722), .B(n14721), .Z(n14723) );
  XOR U15184 ( .A(n14724), .B(n14723), .Z(n14732) );
  AND U15185 ( .A(x[139]), .B(y[108]), .Z(n14726) );
  NAND U15186 ( .A(x[147]), .B(y[148]), .Z(n14725) );
  XNOR U15187 ( .A(n14726), .B(n14725), .Z(n14730) );
  AND U15188 ( .A(x[128]), .B(y[71]), .Z(n14728) );
  NAND U15189 ( .A(x[137]), .B(y[110]), .Z(n14727) );
  XNOR U15190 ( .A(n14728), .B(n14727), .Z(n14729) );
  XNOR U15191 ( .A(n14730), .B(n14729), .Z(n14731) );
  XNOR U15192 ( .A(n14732), .B(n14731), .Z(n14733) );
  XOR U15193 ( .A(n14734), .B(n14733), .Z(n14754) );
  AND U15194 ( .A(x[155]), .B(y[188]), .Z(n14736) );
  NAND U15195 ( .A(x[124]), .B(y[27]), .Z(n14735) );
  XNOR U15196 ( .A(n14736), .B(n14735), .Z(n14740) );
  AND U15197 ( .A(x[158]), .B(y[185]), .Z(n14738) );
  NAND U15198 ( .A(x[159]), .B(y[184]), .Z(n14737) );
  XNOR U15199 ( .A(n14738), .B(n14737), .Z(n14739) );
  XOR U15200 ( .A(n14740), .B(n14739), .Z(n14748) );
  AND U15201 ( .A(x[121]), .B(y[30]), .Z(n14742) );
  NAND U15202 ( .A(x[141]), .B(y[106]), .Z(n14741) );
  XNOR U15203 ( .A(n14742), .B(n14741), .Z(n14746) );
  AND U15204 ( .A(x[154]), .B(y[189]), .Z(n14744) );
  NAND U15205 ( .A(x[149]), .B(y[146]), .Z(n14743) );
  XNOR U15206 ( .A(n14744), .B(n14743), .Z(n14745) );
  XNOR U15207 ( .A(n14746), .B(n14745), .Z(n14747) );
  XNOR U15208 ( .A(n14748), .B(n14747), .Z(n14752) );
  AND U15209 ( .A(y[109]), .B(x[138]), .Z(n14861) );
  AND U15210 ( .A(y[150]), .B(x[145]), .Z(n14833) );
  XOR U15211 ( .A(n14861), .B(n14833), .Z(n14750) );
  AND U15212 ( .A(y[26]), .B(x[125]), .Z(n14821) );
  AND U15213 ( .A(y[67]), .B(x[132]), .Z(n14767) );
  XNOR U15214 ( .A(n14821), .B(n14767), .Z(n14749) );
  XNOR U15215 ( .A(n14750), .B(n14749), .Z(n14751) );
  XNOR U15216 ( .A(n14752), .B(n14751), .Z(n14753) );
  XNOR U15217 ( .A(n14754), .B(n14753), .Z(n14755) );
  XNOR U15218 ( .A(n14756), .B(n14755), .Z(n14757) );
  XNOR U15219 ( .A(n14758), .B(n14757), .Z(n14798) );
  NANDN U15220 ( .A(n14760), .B(n14759), .Z(n14764) );
  NANDN U15221 ( .A(n14762), .B(n14761), .Z(n14763) );
  AND U15222 ( .A(n14764), .B(n14763), .Z(n14796) );
  NAND U15223 ( .A(n14766), .B(n14765), .Z(n14770) );
  NAND U15224 ( .A(n14768), .B(n14767), .Z(n14769) );
  AND U15225 ( .A(n14770), .B(n14769), .Z(n14778) );
  NAND U15226 ( .A(n14772), .B(n14771), .Z(n14776) );
  NAND U15227 ( .A(n14774), .B(n14773), .Z(n14775) );
  NAND U15228 ( .A(n14776), .B(n14775), .Z(n14777) );
  XNOR U15229 ( .A(n14778), .B(n14777), .Z(n14794) );
  NAND U15230 ( .A(n14780), .B(n14779), .Z(n14784) );
  NAND U15231 ( .A(n14782), .B(n14781), .Z(n14783) );
  AND U15232 ( .A(n14784), .B(n14783), .Z(n14792) );
  NAND U15233 ( .A(n14786), .B(n14785), .Z(n14790) );
  NAND U15234 ( .A(n14788), .B(n14787), .Z(n14789) );
  NAND U15235 ( .A(n14790), .B(n14789), .Z(n14791) );
  XNOR U15236 ( .A(n14792), .B(n14791), .Z(n14793) );
  XNOR U15237 ( .A(n14794), .B(n14793), .Z(n14795) );
  XNOR U15238 ( .A(n14796), .B(n14795), .Z(n14797) );
  XNOR U15239 ( .A(n14798), .B(n14797), .Z(n14799) );
  NAND U15240 ( .A(n14802), .B(n14801), .Z(n14806) );
  NAND U15241 ( .A(n14804), .B(n14803), .Z(n14805) );
  AND U15242 ( .A(n14806), .B(n14805), .Z(n14906) );
  NAND U15243 ( .A(n14808), .B(n14807), .Z(n14812) );
  NANDN U15244 ( .A(n14810), .B(n14809), .Z(n14811) );
  AND U15245 ( .A(n14812), .B(n14811), .Z(n14888) );
  NAND U15246 ( .A(n14814), .B(n14813), .Z(n14818) );
  NAND U15247 ( .A(n14816), .B(n14815), .Z(n14817) );
  AND U15248 ( .A(n14818), .B(n14817), .Z(n14826) );
  NAND U15249 ( .A(n14820), .B(n14819), .Z(n14824) );
  NAND U15250 ( .A(n14822), .B(n14821), .Z(n14823) );
  NAND U15251 ( .A(n14824), .B(n14823), .Z(n14825) );
  XNOR U15252 ( .A(n14826), .B(n14825), .Z(n14886) );
  AND U15253 ( .A(x[146]), .B(y[149]), .Z(n14828) );
  NAND U15254 ( .A(x[135]), .B(y[64]), .Z(n14827) );
  XNOR U15255 ( .A(n14828), .B(n14827), .Z(n14852) );
  AND U15256 ( .A(n14830), .B(n14829), .Z(n14846) );
  NAND U15257 ( .A(n14832), .B(n14831), .Z(n14836) );
  NAND U15258 ( .A(n14834), .B(n14833), .Z(n14835) );
  AND U15259 ( .A(n14836), .B(n14835), .Z(n14844) );
  AND U15260 ( .A(x[130]), .B(y[69]), .Z(n14838) );
  NAND U15261 ( .A(x[133]), .B(y[66]), .Z(n14837) );
  XNOR U15262 ( .A(n14838), .B(n14837), .Z(n14842) );
  AND U15263 ( .A(x[144]), .B(y[151]), .Z(n14840) );
  NAND U15264 ( .A(x[129]), .B(y[70]), .Z(n14839) );
  XNOR U15265 ( .A(n14840), .B(n14839), .Z(n14841) );
  XNOR U15266 ( .A(n14842), .B(n14841), .Z(n14843) );
  XNOR U15267 ( .A(n14844), .B(n14843), .Z(n14845) );
  XOR U15268 ( .A(n14846), .B(n14845), .Z(n14850) );
  XNOR U15269 ( .A(n14848), .B(n14847), .Z(n14849) );
  XNOR U15270 ( .A(n14850), .B(n14849), .Z(n14851) );
  XOR U15271 ( .A(n14852), .B(n14851), .Z(n14884) );
  NAND U15272 ( .A(n14854), .B(n14853), .Z(n14858) );
  NAND U15273 ( .A(n14856), .B(n14855), .Z(n14857) );
  AND U15274 ( .A(n14858), .B(n14857), .Z(n14866) );
  NAND U15275 ( .A(n14860), .B(n14859), .Z(n14864) );
  NAND U15276 ( .A(n14862), .B(n14861), .Z(n14863) );
  NAND U15277 ( .A(n14864), .B(n14863), .Z(n14865) );
  XNOR U15278 ( .A(n14866), .B(n14865), .Z(n14882) );
  NAND U15279 ( .A(n14868), .B(n14867), .Z(n14872) );
  NAND U15280 ( .A(n14870), .B(n14869), .Z(n14871) );
  AND U15281 ( .A(n14872), .B(n14871), .Z(n14880) );
  NAND U15282 ( .A(n14874), .B(n14873), .Z(n14878) );
  NAND U15283 ( .A(n14876), .B(n14875), .Z(n14877) );
  NAND U15284 ( .A(n14878), .B(n14877), .Z(n14879) );
  XNOR U15285 ( .A(n14880), .B(n14879), .Z(n14881) );
  XNOR U15286 ( .A(n14882), .B(n14881), .Z(n14883) );
  XNOR U15287 ( .A(n14884), .B(n14883), .Z(n14885) );
  XNOR U15288 ( .A(n14886), .B(n14885), .Z(n14887) );
  XNOR U15289 ( .A(n14888), .B(n14887), .Z(n14904) );
  NAND U15290 ( .A(n14890), .B(n14889), .Z(n14894) );
  ANDN U15291 ( .B(n14892), .A(n14891), .Z(n14893) );
  ANDN U15292 ( .B(n14894), .A(n14893), .Z(n14902) );
  ANDN U15293 ( .B(n14896), .A(n14895), .Z(n14900) );
  AND U15294 ( .A(n14898), .B(n14897), .Z(n14899) );
  OR U15295 ( .A(n14900), .B(n14899), .Z(n14901) );
  XNOR U15296 ( .A(n14902), .B(n14901), .Z(n14903) );
  XNOR U15297 ( .A(n14904), .B(n14903), .Z(n14905) );
  NAND U15298 ( .A(n14908), .B(n14907), .Z(n14912) );
  AND U15299 ( .A(n14910), .B(n14909), .Z(n14911) );
  ANDN U15300 ( .B(n14912), .A(n14911), .Z(n14920) );
  AND U15301 ( .A(n14914), .B(n14913), .Z(n14918) );
  ANDN U15302 ( .B(n14916), .A(n14915), .Z(n14917) );
  OR U15303 ( .A(n14918), .B(n14917), .Z(n14919) );
  XNOR U15304 ( .A(n14920), .B(n14919), .Z(n14921) );
  NANDN U15305 ( .A(n14926), .B(n14925), .Z(n14927) );
  OR U15306 ( .A(n14930), .B(n14929), .Z(n14934) );
  NAND U15307 ( .A(n14932), .B(n14931), .Z(n14933) );
  NAND U15308 ( .A(y[192]), .B(x[152]), .Z(n15054) );
  NAND U15309 ( .A(y[72]), .B(x[128]), .Z(n14940) );
  XOR U15310 ( .A(n15054), .B(n14940), .Z(n14941) );
  AND U15311 ( .A(y[32]), .B(x[120]), .Z(n14948) );
  AND U15312 ( .A(y[112]), .B(x[136]), .Z(n14945) );
  XOR U15313 ( .A(n14948), .B(n14945), .Z(n14944) );
  AND U15314 ( .A(y[152]), .B(x[144]), .Z(n14943) );
  XNOR U15315 ( .A(n14944), .B(n14943), .Z(n14942) );
  XNOR U15316 ( .A(n14941), .B(n14942), .Z(o[152]) );
  AND U15317 ( .A(x[121]), .B(y[32]), .Z(n14939) );
  NAND U15318 ( .A(x[120]), .B(y[33]), .Z(n14938) );
  XNOR U15319 ( .A(n14939), .B(n14938), .Z(n14949) );
  NAND U15320 ( .A(y[72]), .B(x[129]), .Z(n14950) );
  XOR U15321 ( .A(n14949), .B(n14950), .Z(n14966) );
  AND U15322 ( .A(y[192]), .B(x[153]), .Z(n15172) );
  NAND U15323 ( .A(y[113]), .B(x[136]), .Z(n14953) );
  XNOR U15324 ( .A(n15172), .B(n14953), .Z(n14954) );
  AND U15325 ( .A(y[193]), .B(x[152]), .Z(n14976) );
  AND U15326 ( .A(y[112]), .B(x[137]), .Z(n14975) );
  XNOR U15327 ( .A(n14976), .B(n14975), .Z(n14955) );
  XOR U15328 ( .A(n14954), .B(n14955), .Z(n14965) );
  AND U15329 ( .A(y[73]), .B(x[128]), .Z(n15196) );
  AND U15330 ( .A(y[153]), .B(x[144]), .Z(n14970) );
  XOR U15331 ( .A(n15196), .B(n14970), .Z(n14972) );
  AND U15332 ( .A(y[152]), .B(x[145]), .Z(n14971) );
  XNOR U15333 ( .A(n14972), .B(n14971), .Z(n14964) );
  XOR U15334 ( .A(n14965), .B(n14964), .Z(n14967) );
  XOR U15335 ( .A(n14966), .B(n14967), .Z(n14961) );
  NAND U15336 ( .A(n14944), .B(n14943), .Z(n14947) );
  AND U15337 ( .A(n14948), .B(n14945), .Z(n14946) );
  ANDN U15338 ( .B(n14947), .A(n14946), .Z(n14958) );
  XNOR U15339 ( .A(n14959), .B(n14958), .Z(n14960) );
  XNOR U15340 ( .A(n14961), .B(n14960), .Z(o[153]) );
  AND U15341 ( .A(y[33]), .B(x[121]), .Z(n14999) );
  NAND U15342 ( .A(n14999), .B(n14948), .Z(n14952) );
  NANDN U15343 ( .A(n14950), .B(n14949), .Z(n14951) );
  NAND U15344 ( .A(n14952), .B(n14951), .Z(n15036) );
  NANDN U15345 ( .A(n14953), .B(n15172), .Z(n14957) );
  NANDN U15346 ( .A(n14955), .B(n14954), .Z(n14956) );
  NAND U15347 ( .A(n14957), .B(n14956), .Z(n15034) );
  AND U15348 ( .A(y[154]), .B(x[144]), .Z(n15018) );
  NAND U15349 ( .A(y[34]), .B(x[120]), .Z(n15019) );
  AND U15350 ( .A(y[72]), .B(x[130]), .Z(n15020) );
  XOR U15351 ( .A(n15021), .B(n15020), .Z(n15035) );
  XNOR U15352 ( .A(n15034), .B(n15035), .Z(n15037) );
  NANDN U15353 ( .A(n14959), .B(n14958), .Z(n14963) );
  NAND U15354 ( .A(n14961), .B(n14960), .Z(n14962) );
  NAND U15355 ( .A(n14963), .B(n14962), .Z(n14978) );
  XOR U15356 ( .A(n14979), .B(n14978), .Z(n14981) );
  NAND U15357 ( .A(n14965), .B(n14964), .Z(n14969) );
  NAND U15358 ( .A(n14967), .B(n14966), .Z(n14968) );
  AND U15359 ( .A(n14969), .B(n14968), .Z(n14987) );
  AND U15360 ( .A(y[32]), .B(x[122]), .Z(n14997) );
  AND U15361 ( .A(y[114]), .B(x[136]), .Z(n14996) );
  XOR U15362 ( .A(n14997), .B(n14996), .Z(n14998) );
  XOR U15363 ( .A(n14999), .B(n14998), .Z(n15029) );
  AND U15364 ( .A(y[152]), .B(x[146]), .Z(n15028) );
  XOR U15365 ( .A(n15029), .B(n15028), .Z(n15031) );
  AND U15366 ( .A(y[112]), .B(x[138]), .Z(n15082) );
  AND U15367 ( .A(y[194]), .B(x[152]), .Z(n15009) );
  XOR U15368 ( .A(n15082), .B(n15009), .Z(n15011) );
  AND U15369 ( .A(y[113]), .B(x[137]), .Z(n15010) );
  XOR U15370 ( .A(n15011), .B(n15010), .Z(n15030) );
  XOR U15371 ( .A(n15031), .B(n15030), .Z(n14984) );
  AND U15372 ( .A(n15196), .B(n14970), .Z(n14974) );
  NAND U15373 ( .A(n14972), .B(n14971), .Z(n14973) );
  NANDN U15374 ( .A(n14974), .B(n14973), .Z(n14992) );
  AND U15375 ( .A(n14976), .B(n14975), .Z(n15025) );
  AND U15376 ( .A(x[153]), .B(y[193]), .Z(n15059) );
  NAND U15377 ( .A(x[154]), .B(y[192]), .Z(n14977) );
  XOR U15378 ( .A(n15059), .B(n14977), .Z(n15024) );
  AND U15379 ( .A(y[153]), .B(x[145]), .Z(n15002) );
  NAND U15380 ( .A(y[73]), .B(x[129]), .Z(n15003) );
  XNOR U15381 ( .A(n15002), .B(n15003), .Z(n15004) );
  NAND U15382 ( .A(y[74]), .B(x[128]), .Z(n15005) );
  XNOR U15383 ( .A(n15004), .B(n15005), .Z(n14990) );
  XOR U15384 ( .A(n14991), .B(n14990), .Z(n14993) );
  XOR U15385 ( .A(n14992), .B(n14993), .Z(n14985) );
  XOR U15386 ( .A(n14984), .B(n14985), .Z(n14986) );
  XNOR U15387 ( .A(n14987), .B(n14986), .Z(n14980) );
  XNOR U15388 ( .A(n14981), .B(n14980), .Z(o[154]) );
  NAND U15389 ( .A(n14979), .B(n14978), .Z(n14983) );
  NAND U15390 ( .A(n14981), .B(n14980), .Z(n14982) );
  AND U15391 ( .A(n14983), .B(n14982), .Z(n15103) );
  NAND U15392 ( .A(n14985), .B(n14984), .Z(n14989) );
  NAND U15393 ( .A(n14987), .B(n14986), .Z(n14988) );
  NAND U15394 ( .A(n14989), .B(n14988), .Z(n15108) );
  NAND U15395 ( .A(n14991), .B(n14990), .Z(n14995) );
  NAND U15396 ( .A(n14993), .B(n14992), .Z(n14994) );
  NAND U15397 ( .A(n14995), .B(n14994), .Z(n15106) );
  NAND U15398 ( .A(n14997), .B(n14996), .Z(n15001) );
  NAND U15399 ( .A(n14999), .B(n14998), .Z(n15000) );
  NAND U15400 ( .A(n15001), .B(n15000), .Z(n15118) );
  NANDN U15401 ( .A(n15003), .B(n15002), .Z(n15007) );
  NANDN U15402 ( .A(n15005), .B(n15004), .Z(n15006) );
  AND U15403 ( .A(n15007), .B(n15006), .Z(n15073) );
  AND U15404 ( .A(y[155]), .B(x[144]), .Z(n15098) );
  AND U15405 ( .A(y[115]), .B(x[136]), .Z(n15097) );
  NAND U15406 ( .A(y[32]), .B(x[123]), .Z(n15096) );
  XOR U15407 ( .A(n15097), .B(n15096), .Z(n15099) );
  XOR U15408 ( .A(n15098), .B(n15099), .Z(n15071) );
  AND U15409 ( .A(x[138]), .B(y[113]), .Z(n15152) );
  NAND U15410 ( .A(x[139]), .B(y[112]), .Z(n15008) );
  XNOR U15411 ( .A(n15152), .B(n15008), .Z(n15084) );
  AND U15412 ( .A(y[114]), .B(x[137]), .Z(n15083) );
  XOR U15413 ( .A(n15084), .B(n15083), .Z(n15070) );
  XNOR U15414 ( .A(n15071), .B(n15070), .Z(n15072) );
  XNOR U15415 ( .A(n15073), .B(n15072), .Z(n15119) );
  XOR U15416 ( .A(n15118), .B(n15119), .Z(n15121) );
  NAND U15417 ( .A(n15082), .B(n15009), .Z(n15013) );
  AND U15418 ( .A(n15011), .B(n15010), .Z(n15012) );
  ANDN U15419 ( .B(n15013), .A(n15012), .Z(n15078) );
  AND U15420 ( .A(y[34]), .B(x[121]), .Z(n15050) );
  AND U15421 ( .A(y[33]), .B(x[122]), .Z(n15049) );
  NAND U15422 ( .A(y[154]), .B(x[145]), .Z(n15048) );
  XOR U15423 ( .A(n15049), .B(n15048), .Z(n15051) );
  XOR U15424 ( .A(n15050), .B(n15051), .Z(n15077) );
  AND U15425 ( .A(x[155]), .B(y[192]), .Z(n15015) );
  NAND U15426 ( .A(x[152]), .B(y[195]), .Z(n15014) );
  XNOR U15427 ( .A(n15015), .B(n15014), .Z(n15055) );
  AND U15428 ( .A(x[153]), .B(y[194]), .Z(n15017) );
  NAND U15429 ( .A(x[154]), .B(y[193]), .Z(n15016) );
  XOR U15430 ( .A(n15017), .B(n15016), .Z(n15056) );
  XNOR U15431 ( .A(n15055), .B(n15056), .Z(n15076) );
  XOR U15432 ( .A(n15077), .B(n15076), .Z(n15079) );
  XOR U15433 ( .A(n15078), .B(n15079), .Z(n15120) );
  XOR U15434 ( .A(n15121), .B(n15120), .Z(n15107) );
  XOR U15435 ( .A(n15106), .B(n15107), .Z(n15109) );
  XOR U15436 ( .A(n15108), .B(n15109), .Z(n15102) );
  XOR U15437 ( .A(n15103), .B(n15102), .Z(n15105) );
  NANDN U15438 ( .A(n15019), .B(n15018), .Z(n15023) );
  NAND U15439 ( .A(n15021), .B(n15020), .Z(n15022) );
  AND U15440 ( .A(n15023), .B(n15022), .Z(n15041) );
  ANDN U15441 ( .B(n15025), .A(n15024), .Z(n15027) );
  AND U15442 ( .A(y[193]), .B(x[154]), .Z(n15169) );
  NAND U15443 ( .A(n15169), .B(n15172), .Z(n15026) );
  NANDN U15444 ( .A(n15027), .B(n15026), .Z(n15040) );
  AND U15445 ( .A(y[72]), .B(x[131]), .Z(n15090) );
  AND U15446 ( .A(y[35]), .B(x[120]), .Z(n15088) );
  NAND U15447 ( .A(y[153]), .B(x[146]), .Z(n15087) );
  XNOR U15448 ( .A(n15088), .B(n15087), .Z(n15089) );
  XOR U15449 ( .A(n15090), .B(n15089), .Z(n15068) );
  AND U15450 ( .A(y[75]), .B(x[128]), .Z(n15063) );
  AND U15451 ( .A(y[73]), .B(x[130]), .Z(n15061) );
  NAND U15452 ( .A(y[152]), .B(x[147]), .Z(n15060) );
  XNOR U15453 ( .A(n15061), .B(n15060), .Z(n15062) );
  XOR U15454 ( .A(n15063), .B(n15062), .Z(n15066) );
  AND U15455 ( .A(y[74]), .B(x[129]), .Z(n15067) );
  XOR U15456 ( .A(n15066), .B(n15067), .Z(n15069) );
  XOR U15457 ( .A(n15068), .B(n15069), .Z(n15042) );
  XOR U15458 ( .A(n15043), .B(n15042), .Z(n15113) );
  NAND U15459 ( .A(n15029), .B(n15028), .Z(n15033) );
  NAND U15460 ( .A(n15031), .B(n15030), .Z(n15032) );
  AND U15461 ( .A(n15033), .B(n15032), .Z(n15112) );
  NAND U15462 ( .A(n15035), .B(n15034), .Z(n15039) );
  NANDN U15463 ( .A(n15037), .B(n15036), .Z(n15038) );
  AND U15464 ( .A(n15039), .B(n15038), .Z(n15114) );
  XNOR U15465 ( .A(n15115), .B(n15114), .Z(n15104) );
  XOR U15466 ( .A(n15105), .B(n15104), .Z(o[155]) );
  NANDN U15467 ( .A(n15041), .B(n15040), .Z(n15045) );
  NAND U15468 ( .A(n15043), .B(n15042), .Z(n15044) );
  AND U15469 ( .A(n15045), .B(n15044), .Z(n15135) );
  AND U15470 ( .A(y[74]), .B(x[130]), .Z(n15263) );
  AND U15471 ( .A(x[128]), .B(y[76]), .Z(n15047) );
  NAND U15472 ( .A(x[131]), .B(y[73]), .Z(n15046) );
  XOR U15473 ( .A(n15047), .B(n15046), .Z(n15197) );
  XNOR U15474 ( .A(n15263), .B(n15197), .Z(n15200) );
  NAND U15475 ( .A(y[75]), .B(x[129]), .Z(n15201) );
  XNOR U15476 ( .A(n15200), .B(n15201), .Z(n15203) );
  AND U15477 ( .A(y[152]), .B(x[148]), .Z(n15157) );
  NAND U15478 ( .A(y[35]), .B(x[121]), .Z(n15158) );
  XNOR U15479 ( .A(n15157), .B(n15158), .Z(n15159) );
  NAND U15480 ( .A(y[36]), .B(x[120]), .Z(n15160) );
  XNOR U15481 ( .A(n15159), .B(n15160), .Z(n15202) );
  XOR U15482 ( .A(n15203), .B(n15202), .Z(n15215) );
  NANDN U15483 ( .A(n15049), .B(n15048), .Z(n15053) );
  OR U15484 ( .A(n15051), .B(n15050), .Z(n15052) );
  AND U15485 ( .A(n15053), .B(n15052), .Z(n15213) );
  AND U15486 ( .A(y[195]), .B(x[155]), .Z(n15484) );
  NANDN U15487 ( .A(n15054), .B(n15484), .Z(n15058) );
  NANDN U15488 ( .A(n15056), .B(n15055), .Z(n15057) );
  AND U15489 ( .A(n15058), .B(n15057), .Z(n15212) );
  XNOR U15490 ( .A(n15213), .B(n15212), .Z(n15214) );
  XNOR U15491 ( .A(n15215), .B(n15214), .Z(n15229) );
  NAND U15492 ( .A(y[32]), .B(x[124]), .Z(n15184) );
  NAND U15493 ( .A(y[154]), .B(x[146]), .Z(n15183) );
  NAND U15494 ( .A(y[116]), .B(x[136]), .Z(n15182) );
  XOR U15495 ( .A(n15183), .B(n15182), .Z(n15185) );
  XNOR U15496 ( .A(n15184), .B(n15185), .Z(n15141) );
  AND U15497 ( .A(y[194]), .B(x[154]), .Z(n15095) );
  NAND U15498 ( .A(n15095), .B(n15059), .Z(n15177) );
  NAND U15499 ( .A(y[196]), .B(x[152]), .Z(n15318) );
  NAND U15500 ( .A(y[112]), .B(x[140]), .Z(n15278) );
  XNOR U15501 ( .A(n15318), .B(n15278), .Z(n15178) );
  XOR U15502 ( .A(n15177), .B(n15178), .Z(n15140) );
  XOR U15503 ( .A(n15141), .B(n15140), .Z(n15142) );
  NANDN U15504 ( .A(n15061), .B(n15060), .Z(n15065) );
  NANDN U15505 ( .A(n15063), .B(n15062), .Z(n15064) );
  NAND U15506 ( .A(n15065), .B(n15064), .Z(n15143) );
  XOR U15507 ( .A(n15142), .B(n15143), .Z(n15226) );
  XOR U15508 ( .A(n15226), .B(n15227), .Z(n15228) );
  XNOR U15509 ( .A(n15229), .B(n15228), .Z(n15134) );
  NANDN U15510 ( .A(n15071), .B(n15070), .Z(n15075) );
  NANDN U15511 ( .A(n15073), .B(n15072), .Z(n15074) );
  NAND U15512 ( .A(n15075), .B(n15074), .Z(n15218) );
  NANDN U15513 ( .A(n15077), .B(n15076), .Z(n15081) );
  OR U15514 ( .A(n15079), .B(n15078), .Z(n15080) );
  NAND U15515 ( .A(n15081), .B(n15080), .Z(n15219) );
  XOR U15516 ( .A(n15218), .B(n15219), .Z(n15221) );
  AND U15517 ( .A(y[72]), .B(x[132]), .Z(n15163) );
  NAND U15518 ( .A(y[156]), .B(x[144]), .Z(n15164) );
  XNOR U15519 ( .A(n15163), .B(n15164), .Z(n15165) );
  NAND U15520 ( .A(y[155]), .B(x[145]), .Z(n15166) );
  XNOR U15521 ( .A(n15165), .B(n15166), .Z(n15206) );
  AND U15522 ( .A(x[138]), .B(y[114]), .Z(n15086) );
  NAND U15523 ( .A(x[139]), .B(y[113]), .Z(n15085) );
  XNOR U15524 ( .A(n15086), .B(n15085), .Z(n15153) );
  NAND U15525 ( .A(y[115]), .B(x[137]), .Z(n15154) );
  XOR U15526 ( .A(n15153), .B(n15154), .Z(n15207) );
  XNOR U15527 ( .A(n15206), .B(n15207), .Z(n15208) );
  NANDN U15528 ( .A(n15088), .B(n15087), .Z(n15092) );
  NANDN U15529 ( .A(n15090), .B(n15089), .Z(n15091) );
  NAND U15530 ( .A(n15092), .B(n15091), .Z(n15209) );
  XNOR U15531 ( .A(n15208), .B(n15209), .Z(n15223) );
  XOR U15532 ( .A(n15222), .B(n15223), .Z(n15225) );
  NAND U15533 ( .A(y[34]), .B(x[122]), .Z(n15192) );
  NAND U15534 ( .A(y[153]), .B(x[147]), .Z(n15191) );
  NAND U15535 ( .A(y[33]), .B(x[123]), .Z(n15190) );
  XNOR U15536 ( .A(n15191), .B(n15190), .Z(n15193) );
  AND U15537 ( .A(x[156]), .B(y[192]), .Z(n15094) );
  NAND U15538 ( .A(x[153]), .B(y[195]), .Z(n15093) );
  XNOR U15539 ( .A(n15094), .B(n15093), .Z(n15174) );
  AND U15540 ( .A(y[193]), .B(x[155]), .Z(n15285) );
  XOR U15541 ( .A(n15095), .B(n15285), .Z(n15173) );
  XOR U15542 ( .A(n15174), .B(n15173), .Z(n15146) );
  XOR U15543 ( .A(n15147), .B(n15146), .Z(n15148) );
  NANDN U15544 ( .A(n15097), .B(n15096), .Z(n15101) );
  OR U15545 ( .A(n15099), .B(n15098), .Z(n15100) );
  NAND U15546 ( .A(n15101), .B(n15100), .Z(n15149) );
  XNOR U15547 ( .A(n15148), .B(n15149), .Z(n15224) );
  XOR U15548 ( .A(n15225), .B(n15224), .Z(n15220) );
  XOR U15549 ( .A(n15221), .B(n15220), .Z(n15136) );
  XNOR U15550 ( .A(n15137), .B(n15136), .Z(n15127) );
  NAND U15551 ( .A(n15107), .B(n15106), .Z(n15111) );
  NAND U15552 ( .A(n15109), .B(n15108), .Z(n15110) );
  AND U15553 ( .A(n15111), .B(n15110), .Z(n15130) );
  NANDN U15554 ( .A(n15113), .B(n15112), .Z(n15117) );
  NAND U15555 ( .A(n15115), .B(n15114), .Z(n15116) );
  NAND U15556 ( .A(n15117), .B(n15116), .Z(n15128) );
  NAND U15557 ( .A(n15119), .B(n15118), .Z(n15123) );
  NAND U15558 ( .A(n15121), .B(n15120), .Z(n15122) );
  AND U15559 ( .A(n15123), .B(n15122), .Z(n15129) );
  XOR U15560 ( .A(n15128), .B(n15129), .Z(n15131) );
  XNOR U15561 ( .A(n15130), .B(n15131), .Z(n15126) );
  XOR U15562 ( .A(n15125), .B(n15126), .Z(n15124) );
  XNOR U15563 ( .A(n15127), .B(n15124), .Z(o[156]) );
  NAND U15564 ( .A(n15129), .B(n15128), .Z(n15133) );
  NAND U15565 ( .A(n15131), .B(n15130), .Z(n15132) );
  AND U15566 ( .A(n15133), .B(n15132), .Z(n15365) );
  XNOR U15567 ( .A(n15366), .B(n15365), .Z(n15368) );
  NANDN U15568 ( .A(n15135), .B(n15134), .Z(n15139) );
  NAND U15569 ( .A(n15137), .B(n15136), .Z(n15138) );
  AND U15570 ( .A(n15139), .B(n15138), .Z(n15231) );
  NAND U15571 ( .A(n15141), .B(n15140), .Z(n15145) );
  NANDN U15572 ( .A(n15143), .B(n15142), .Z(n15144) );
  AND U15573 ( .A(n15145), .B(n15144), .Z(n15287) );
  NAND U15574 ( .A(n15147), .B(n15146), .Z(n15151) );
  NANDN U15575 ( .A(n15149), .B(n15148), .Z(n15150) );
  NAND U15576 ( .A(n15151), .B(n15150), .Z(n15286) );
  XNOR U15577 ( .A(n15287), .B(n15286), .Z(n15289) );
  AND U15578 ( .A(y[114]), .B(x[139]), .Z(n15279) );
  NAND U15579 ( .A(n15152), .B(n15279), .Z(n15156) );
  NANDN U15580 ( .A(n15154), .B(n15153), .Z(n15155) );
  AND U15581 ( .A(n15156), .B(n15155), .Z(n15241) );
  NANDN U15582 ( .A(n15158), .B(n15157), .Z(n15162) );
  NANDN U15583 ( .A(n15160), .B(n15159), .Z(n15161) );
  NAND U15584 ( .A(n15162), .B(n15161), .Z(n15248) );
  AND U15585 ( .A(y[72]), .B(x[133]), .Z(n15269) );
  AND U15586 ( .A(y[115]), .B(x[138]), .Z(n15268) );
  XOR U15587 ( .A(n15269), .B(n15268), .Z(n15270) );
  AND U15588 ( .A(y[157]), .B(x[144]), .Z(n15541) );
  XOR U15589 ( .A(n15270), .B(n15541), .Z(n15247) );
  AND U15590 ( .A(y[153]), .B(x[148]), .Z(n15274) );
  AND U15591 ( .A(y[32]), .B(x[125]), .Z(n15273) );
  XOR U15592 ( .A(n15274), .B(n15273), .Z(n15275) );
  AND U15593 ( .A(y[33]), .B(x[124]), .Z(n15505) );
  XOR U15594 ( .A(n15275), .B(n15505), .Z(n15246) );
  XOR U15595 ( .A(n15247), .B(n15246), .Z(n15249) );
  XOR U15596 ( .A(n15248), .B(n15249), .Z(n15240) );
  NANDN U15597 ( .A(n15164), .B(n15163), .Z(n15168) );
  NANDN U15598 ( .A(n15166), .B(n15165), .Z(n15167) );
  NAND U15599 ( .A(n15168), .B(n15167), .Z(n15356) );
  AND U15600 ( .A(y[194]), .B(x[155]), .Z(n15180) );
  AND U15601 ( .A(n15180), .B(n15169), .Z(n15320) );
  AND U15602 ( .A(x[152]), .B(y[197]), .Z(n15171) );
  AND U15603 ( .A(x[153]), .B(y[196]), .Z(n15170) );
  XOR U15604 ( .A(n15171), .B(n15170), .Z(n15319) );
  XOR U15605 ( .A(n15320), .B(n15319), .Z(n15355) );
  AND U15606 ( .A(y[73]), .B(x[132]), .Z(n15347) );
  AND U15607 ( .A(y[77]), .B(x[128]), .Z(n15345) );
  AND U15608 ( .A(y[36]), .B(x[121]), .Z(n15344) );
  XOR U15609 ( .A(n15345), .B(n15344), .Z(n15346) );
  XOR U15610 ( .A(n15347), .B(n15346), .Z(n15354) );
  XOR U15611 ( .A(n15355), .B(n15354), .Z(n15357) );
  XOR U15612 ( .A(n15356), .B(n15357), .Z(n15242) );
  XOR U15613 ( .A(n15243), .B(n15242), .Z(n15288) );
  XOR U15614 ( .A(n15289), .B(n15288), .Z(n15238) );
  AND U15615 ( .A(y[195]), .B(x[156]), .Z(n15572) );
  NAND U15616 ( .A(n15572), .B(n15172), .Z(n15176) );
  NAND U15617 ( .A(n15174), .B(n15173), .Z(n15175) );
  AND U15618 ( .A(n15176), .B(n15175), .Z(n15301) );
  XNOR U15619 ( .A(n15301), .B(n15300), .Z(n15303) );
  AND U15620 ( .A(y[195]), .B(x[154]), .Z(n15250) );
  NAND U15621 ( .A(y[192]), .B(x[157]), .Z(n15251) );
  XNOR U15622 ( .A(n15250), .B(n15251), .Z(n15252) );
  NAND U15623 ( .A(x[156]), .B(y[193]), .Z(n15179) );
  XOR U15624 ( .A(n15180), .B(n15179), .Z(n15253) );
  XNOR U15625 ( .A(n15252), .B(n15253), .Z(n15290) );
  AND U15626 ( .A(y[74]), .B(x[131]), .Z(n15413) );
  NAND U15627 ( .A(x[130]), .B(y[75]), .Z(n15181) );
  XNOR U15628 ( .A(n15413), .B(n15181), .Z(n15264) );
  NAND U15629 ( .A(y[76]), .B(x[129]), .Z(n15265) );
  XOR U15630 ( .A(n15264), .B(n15265), .Z(n15291) );
  XNOR U15631 ( .A(n15290), .B(n15291), .Z(n15292) );
  NAND U15632 ( .A(n15183), .B(n15182), .Z(n15187) );
  NAND U15633 ( .A(n15185), .B(n15184), .Z(n15186) );
  NAND U15634 ( .A(n15187), .B(n15186), .Z(n15293) );
  XNOR U15635 ( .A(n15292), .B(n15293), .Z(n15302) );
  XOR U15636 ( .A(n15303), .B(n15302), .Z(n15315) );
  AND U15637 ( .A(x[140]), .B(y[113]), .Z(n15189) );
  NAND U15638 ( .A(x[141]), .B(y[112]), .Z(n15188) );
  XOR U15639 ( .A(n15189), .B(n15188), .Z(n15280) );
  XNOR U15640 ( .A(n15279), .B(n15280), .Z(n15337) );
  AND U15641 ( .A(y[152]), .B(x[149]), .Z(n15256) );
  NAND U15642 ( .A(y[34]), .B(x[123]), .Z(n15257) );
  XNOR U15643 ( .A(n15256), .B(n15257), .Z(n15259) );
  AND U15644 ( .A(y[35]), .B(x[122]), .Z(n15258) );
  XOR U15645 ( .A(n15259), .B(n15258), .Z(n15336) );
  XOR U15646 ( .A(n15337), .B(n15336), .Z(n15339) );
  NAND U15647 ( .A(n15191), .B(n15190), .Z(n15195) );
  NANDN U15648 ( .A(n15193), .B(n15192), .Z(n15194) );
  AND U15649 ( .A(n15195), .B(n15194), .Z(n15338) );
  XOR U15650 ( .A(n15339), .B(n15338), .Z(n15313) );
  AND U15651 ( .A(y[76]), .B(x[131]), .Z(n15466) );
  NAND U15652 ( .A(n15466), .B(n15196), .Z(n15199) );
  NANDN U15653 ( .A(n15197), .B(n15263), .Z(n15198) );
  AND U15654 ( .A(n15199), .B(n15198), .Z(n15299) );
  AND U15655 ( .A(y[154]), .B(x[147]), .Z(n15331) );
  AND U15656 ( .A(y[116]), .B(x[137]), .Z(n15559) );
  XOR U15657 ( .A(n15331), .B(n15559), .Z(n15333) );
  AND U15658 ( .A(y[117]), .B(x[136]), .Z(n15332) );
  XOR U15659 ( .A(n15333), .B(n15332), .Z(n15297) );
  AND U15660 ( .A(y[37]), .B(x[120]), .Z(n15324) );
  AND U15661 ( .A(y[156]), .B(x[145]), .Z(n15323) );
  XOR U15662 ( .A(n15324), .B(n15323), .Z(n15326) );
  AND U15663 ( .A(y[155]), .B(x[146]), .Z(n15325) );
  XOR U15664 ( .A(n15326), .B(n15325), .Z(n15296) );
  XOR U15665 ( .A(n15297), .B(n15296), .Z(n15298) );
  XOR U15666 ( .A(n15299), .B(n15298), .Z(n15312) );
  XNOR U15667 ( .A(n15313), .B(n15312), .Z(n15314) );
  XOR U15668 ( .A(n15315), .B(n15314), .Z(n15237) );
  NANDN U15669 ( .A(n15201), .B(n15200), .Z(n15205) );
  NAND U15670 ( .A(n15203), .B(n15202), .Z(n15204) );
  AND U15671 ( .A(n15205), .B(n15204), .Z(n15307) );
  NANDN U15672 ( .A(n15207), .B(n15206), .Z(n15211) );
  NANDN U15673 ( .A(n15209), .B(n15208), .Z(n15210) );
  NAND U15674 ( .A(n15211), .B(n15210), .Z(n15306) );
  XNOR U15675 ( .A(n15307), .B(n15306), .Z(n15309) );
  NANDN U15676 ( .A(n15213), .B(n15212), .Z(n15217) );
  NANDN U15677 ( .A(n15215), .B(n15214), .Z(n15216) );
  AND U15678 ( .A(n15217), .B(n15216), .Z(n15308) );
  XOR U15679 ( .A(n15309), .B(n15308), .Z(n15236) );
  XNOR U15680 ( .A(n15237), .B(n15236), .Z(n15239) );
  XNOR U15681 ( .A(n15238), .B(n15239), .Z(n15230) );
  XOR U15682 ( .A(n15360), .B(n15361), .Z(n15363) );
  XOR U15683 ( .A(n15362), .B(n15363), .Z(n15232) );
  XOR U15684 ( .A(n15233), .B(n15232), .Z(n15367) );
  XOR U15685 ( .A(n15368), .B(n15367), .Z(o[157]) );
  NANDN U15686 ( .A(n15231), .B(n15230), .Z(n15235) );
  NAND U15687 ( .A(n15233), .B(n15232), .Z(n15234) );
  NAND U15688 ( .A(n15235), .B(n15234), .Z(n15661) );
  NANDN U15689 ( .A(n15241), .B(n15240), .Z(n15245) );
  NAND U15690 ( .A(n15243), .B(n15242), .Z(n15244) );
  AND U15691 ( .A(n15245), .B(n15244), .Z(n15665) );
  NANDN U15692 ( .A(n15251), .B(n15250), .Z(n15255) );
  NANDN U15693 ( .A(n15253), .B(n15252), .Z(n15254) );
  NAND U15694 ( .A(n15255), .B(n15254), .Z(n15526) );
  NANDN U15695 ( .A(n15257), .B(n15256), .Z(n15261) );
  NAND U15696 ( .A(n15259), .B(n15258), .Z(n15260) );
  NAND U15697 ( .A(n15261), .B(n15260), .Z(n15529) );
  AND U15698 ( .A(y[75]), .B(x[131]), .Z(n15262) );
  NAND U15699 ( .A(n15263), .B(n15262), .Z(n15267) );
  NANDN U15700 ( .A(n15265), .B(n15264), .Z(n15266) );
  AND U15701 ( .A(n15267), .B(n15266), .Z(n15621) );
  AND U15702 ( .A(y[155]), .B(x[147]), .Z(n15547) );
  AND U15703 ( .A(y[115]), .B(x[139]), .Z(n15546) );
  XOR U15704 ( .A(n15547), .B(n15546), .Z(n15545) );
  AND U15705 ( .A(y[35]), .B(x[123]), .Z(n15544) );
  XOR U15706 ( .A(n15545), .B(n15544), .Z(n15623) );
  AND U15707 ( .A(y[156]), .B(x[146]), .Z(n15601) );
  AND U15708 ( .A(y[114]), .B(x[140]), .Z(n15600) );
  XOR U15709 ( .A(n15601), .B(n15600), .Z(n15599) );
  AND U15710 ( .A(y[36]), .B(x[122]), .Z(n15598) );
  XNOR U15711 ( .A(n15599), .B(n15598), .Z(n15622) );
  XNOR U15712 ( .A(n15621), .B(n15620), .Z(n15528) );
  XOR U15713 ( .A(n15529), .B(n15528), .Z(n15527) );
  XOR U15714 ( .A(n15526), .B(n15527), .Z(n15402) );
  XOR U15715 ( .A(n15401), .B(n15402), .Z(n15400) );
  NAND U15716 ( .A(n15269), .B(n15268), .Z(n15272) );
  NAND U15717 ( .A(n15270), .B(n15541), .Z(n15271) );
  NAND U15718 ( .A(n15272), .B(n15271), .Z(n15408) );
  NAND U15719 ( .A(n15274), .B(n15273), .Z(n15277) );
  NAND U15720 ( .A(n15275), .B(n15505), .Z(n15276) );
  NAND U15721 ( .A(n15277), .B(n15276), .Z(n15407) );
  XOR U15722 ( .A(n15408), .B(n15407), .Z(n15406) );
  AND U15723 ( .A(y[113]), .B(x[141]), .Z(n15595) );
  NANDN U15724 ( .A(n15278), .B(n15595), .Z(n15282) );
  NANDN U15725 ( .A(n15280), .B(n15279), .Z(n15281) );
  AND U15726 ( .A(n15282), .B(n15281), .Z(n15615) );
  AND U15727 ( .A(x[125]), .B(y[33]), .Z(n15284) );
  NAND U15728 ( .A(x[124]), .B(y[34]), .Z(n15283) );
  XNOR U15729 ( .A(n15284), .B(n15283), .Z(n15504) );
  AND U15730 ( .A(y[152]), .B(x[150]), .Z(n15503) );
  XOR U15731 ( .A(n15504), .B(n15503), .Z(n15617) );
  AND U15732 ( .A(y[197]), .B(x[153]), .Z(n15492) );
  AND U15733 ( .A(x[156]), .B(y[194]), .Z(n15330) );
  AND U15734 ( .A(n15330), .B(n15285), .Z(n15490) );
  AND U15735 ( .A(y[196]), .B(x[154]), .Z(n15489) );
  XOR U15736 ( .A(n15490), .B(n15489), .Z(n15491) );
  XNOR U15737 ( .A(n15492), .B(n15491), .Z(n15616) );
  XNOR U15738 ( .A(n15615), .B(n15614), .Z(n15405) );
  XOR U15739 ( .A(n15406), .B(n15405), .Z(n15399) );
  XOR U15740 ( .A(n15400), .B(n15399), .Z(n15376) );
  NANDN U15741 ( .A(n15291), .B(n15290), .Z(n15295) );
  NANDN U15742 ( .A(n15293), .B(n15292), .Z(n15294) );
  AND U15743 ( .A(n15295), .B(n15294), .Z(n15392) );
  NANDN U15744 ( .A(n15301), .B(n15300), .Z(n15305) );
  NAND U15745 ( .A(n15303), .B(n15302), .Z(n15304) );
  AND U15746 ( .A(n15305), .B(n15304), .Z(n15393) );
  XOR U15747 ( .A(n15394), .B(n15393), .Z(n15391) );
  XOR U15748 ( .A(n15392), .B(n15391), .Z(n15372) );
  XOR U15749 ( .A(n15373), .B(n15372), .Z(n15664) );
  XOR U15750 ( .A(n15665), .B(n15664), .Z(n15662) );
  NANDN U15751 ( .A(n15307), .B(n15306), .Z(n15311) );
  NAND U15752 ( .A(n15309), .B(n15308), .Z(n15310) );
  AND U15753 ( .A(n15311), .B(n15310), .Z(n15640) );
  NANDN U15754 ( .A(n15313), .B(n15312), .Z(n15317) );
  NANDN U15755 ( .A(n15315), .B(n15314), .Z(n15316) );
  NAND U15756 ( .A(n15317), .B(n15316), .Z(n15643) );
  NANDN U15757 ( .A(n15318), .B(n15492), .Z(n15322) );
  NAND U15758 ( .A(n15320), .B(n15319), .Z(n15321) );
  NAND U15759 ( .A(n15322), .B(n15321), .Z(n15388) );
  NAND U15760 ( .A(n15324), .B(n15323), .Z(n15328) );
  NAND U15761 ( .A(n15326), .B(n15325), .Z(n15327) );
  AND U15762 ( .A(n15328), .B(n15327), .Z(n15478) );
  AND U15763 ( .A(y[37]), .B(x[121]), .Z(n15587) );
  AND U15764 ( .A(y[72]), .B(x[134]), .Z(n15586) );
  XOR U15765 ( .A(n15587), .B(n15586), .Z(n15585) );
  AND U15766 ( .A(y[78]), .B(x[128]), .Z(n15584) );
  XOR U15767 ( .A(n15585), .B(n15584), .Z(n15479) );
  NAND U15768 ( .A(x[157]), .B(y[193]), .Z(n15329) );
  XNOR U15769 ( .A(n15330), .B(n15329), .Z(n15486) );
  AND U15770 ( .A(y[192]), .B(x[158]), .Z(n15485) );
  XOR U15771 ( .A(n15486), .B(n15485), .Z(n15483) );
  XNOR U15772 ( .A(n15484), .B(n15483), .Z(n15480) );
  XNOR U15773 ( .A(n15478), .B(n15477), .Z(n15387) );
  XOR U15774 ( .A(n15388), .B(n15387), .Z(n15385) );
  NAND U15775 ( .A(n15331), .B(n15559), .Z(n15335) );
  NAND U15776 ( .A(n15333), .B(n15332), .Z(n15334) );
  NAND U15777 ( .A(n15335), .B(n15334), .Z(n15384) );
  XOR U15778 ( .A(n15385), .B(n15384), .Z(n15648) );
  NAND U15779 ( .A(n15337), .B(n15336), .Z(n15341) );
  NAND U15780 ( .A(n15339), .B(n15338), .Z(n15340) );
  AND U15781 ( .A(n15341), .B(n15340), .Z(n15647) );
  AND U15782 ( .A(y[118]), .B(x[136]), .Z(n15500) );
  AND U15783 ( .A(y[32]), .B(x[126]), .Z(n15499) );
  XOR U15784 ( .A(n15500), .B(n15499), .Z(n15498) );
  AND U15785 ( .A(y[153]), .B(x[149]), .Z(n15497) );
  XOR U15786 ( .A(n15498), .B(n15497), .Z(n15535) );
  AND U15787 ( .A(y[73]), .B(x[133]), .Z(n15581) );
  AND U15788 ( .A(y[76]), .B(x[130]), .Z(n15580) );
  XOR U15789 ( .A(n15581), .B(n15580), .Z(n15579) );
  AND U15790 ( .A(y[77]), .B(x[129]), .Z(n15578) );
  XOR U15791 ( .A(n15579), .B(n15578), .Z(n15412) );
  AND U15792 ( .A(x[132]), .B(y[74]), .Z(n15343) );
  NAND U15793 ( .A(x[131]), .B(y[75]), .Z(n15342) );
  XNOR U15794 ( .A(n15343), .B(n15342), .Z(n15411) );
  XOR U15795 ( .A(n15412), .B(n15411), .Z(n15534) );
  XOR U15796 ( .A(n15535), .B(n15534), .Z(n15533) );
  AND U15797 ( .A(y[198]), .B(x[152]), .Z(n15594) );
  XOR U15798 ( .A(n15595), .B(n15594), .Z(n15593) );
  AND U15799 ( .A(y[112]), .B(x[142]), .Z(n15592) );
  XOR U15800 ( .A(n15593), .B(n15592), .Z(n15532) );
  XOR U15801 ( .A(n15533), .B(n15532), .Z(n15381) );
  NAND U15802 ( .A(n15345), .B(n15344), .Z(n15349) );
  NAND U15803 ( .A(n15347), .B(n15346), .Z(n15348) );
  AND U15804 ( .A(n15349), .B(n15348), .Z(n15514) );
  AND U15805 ( .A(y[154]), .B(x[148]), .Z(n15557) );
  AND U15806 ( .A(x[137]), .B(y[117]), .Z(n15351) );
  AND U15807 ( .A(x[138]), .B(y[116]), .Z(n15350) );
  XOR U15808 ( .A(n15351), .B(n15350), .Z(n15556) );
  XOR U15809 ( .A(n15557), .B(n15556), .Z(n15517) );
  AND U15810 ( .A(y[38]), .B(x[120]), .Z(n15539) );
  AND U15811 ( .A(y[158]), .B(x[144]), .Z(n15353) );
  AND U15812 ( .A(x[145]), .B(y[157]), .Z(n15352) );
  XOR U15813 ( .A(n15353), .B(n15352), .Z(n15538) );
  XNOR U15814 ( .A(n15539), .B(n15538), .Z(n15516) );
  XNOR U15815 ( .A(n15514), .B(n15515), .Z(n15380) );
  NAND U15816 ( .A(n15355), .B(n15354), .Z(n15359) );
  NAND U15817 ( .A(n15357), .B(n15356), .Z(n15358) );
  AND U15818 ( .A(n15359), .B(n15358), .Z(n15377) );
  XOR U15819 ( .A(n15378), .B(n15377), .Z(n15646) );
  XOR U15820 ( .A(n15647), .B(n15646), .Z(n15649) );
  XOR U15821 ( .A(n15643), .B(n15642), .Z(n15641) );
  XOR U15822 ( .A(n15640), .B(n15641), .Z(n15663) );
  XOR U15823 ( .A(n15658), .B(n15654), .Z(n15364) );
  XNOR U15824 ( .A(n15655), .B(n15364), .Z(n15660) );
  NANDN U15825 ( .A(n15366), .B(n15365), .Z(n15370) );
  NAND U15826 ( .A(n15368), .B(n15367), .Z(n15369) );
  AND U15827 ( .A(n15370), .B(n15369), .Z(n15659) );
  XOR U15828 ( .A(n15660), .B(n15659), .Z(n15371) );
  XNOR U15829 ( .A(n15661), .B(n15371), .Z(o[158]) );
  IV U15830 ( .A(n15372), .Z(n15374) );
  IV U15831 ( .A(n15377), .Z(n15379) );
  NANDN U15832 ( .A(n15379), .B(n15378), .Z(n15383) );
  NANDN U15833 ( .A(n15381), .B(n15380), .Z(n15382) );
  AND U15834 ( .A(n15383), .B(n15382), .Z(n15639) );
  IV U15835 ( .A(n15384), .Z(n15386) );
  NANDN U15836 ( .A(n15386), .B(n15385), .Z(n15390) );
  NAND U15837 ( .A(n15388), .B(n15387), .Z(n15389) );
  AND U15838 ( .A(n15390), .B(n15389), .Z(n15398) );
  NAND U15839 ( .A(n15392), .B(n15391), .Z(n15396) );
  NAND U15840 ( .A(n15394), .B(n15393), .Z(n15395) );
  NAND U15841 ( .A(n15396), .B(n15395), .Z(n15397) );
  XNOR U15842 ( .A(n15398), .B(n15397), .Z(n15637) );
  NAND U15843 ( .A(n15400), .B(n15399), .Z(n15404) );
  AND U15844 ( .A(n15402), .B(n15401), .Z(n15403) );
  ANDN U15845 ( .B(n15404), .A(n15403), .Z(n15635) );
  NAND U15846 ( .A(n15406), .B(n15405), .Z(n15410) );
  AND U15847 ( .A(n15408), .B(n15407), .Z(n15409) );
  ANDN U15848 ( .B(n15410), .A(n15409), .Z(n15525) );
  NAND U15849 ( .A(n15412), .B(n15411), .Z(n15415) );
  AND U15850 ( .A(y[75]), .B(x[132]), .Z(n15465) );
  NAND U15851 ( .A(n15413), .B(n15465), .Z(n15414) );
  AND U15852 ( .A(n15415), .B(n15414), .Z(n15476) );
  AND U15853 ( .A(x[120]), .B(y[39]), .Z(n15417) );
  NAND U15854 ( .A(x[141]), .B(y[114]), .Z(n15416) );
  XNOR U15855 ( .A(n15417), .B(n15416), .Z(n15421) );
  AND U15856 ( .A(x[153]), .B(y[198]), .Z(n15419) );
  NAND U15857 ( .A(x[148]), .B(y[155]), .Z(n15418) );
  XNOR U15858 ( .A(n15419), .B(n15418), .Z(n15420) );
  XOR U15859 ( .A(n15421), .B(n15420), .Z(n15429) );
  AND U15860 ( .A(x[149]), .B(y[154]), .Z(n15423) );
  NAND U15861 ( .A(x[142]), .B(y[113]), .Z(n15422) );
  XNOR U15862 ( .A(n15423), .B(n15422), .Z(n15427) );
  AND U15863 ( .A(x[128]), .B(y[79]), .Z(n15425) );
  NAND U15864 ( .A(x[151]), .B(y[152]), .Z(n15424) );
  XNOR U15865 ( .A(n15425), .B(n15424), .Z(n15426) );
  XNOR U15866 ( .A(n15427), .B(n15426), .Z(n15428) );
  XNOR U15867 ( .A(n15429), .B(n15428), .Z(n15474) );
  AND U15868 ( .A(x[134]), .B(y[73]), .Z(n15434) );
  AND U15869 ( .A(y[158]), .B(x[145]), .Z(n15540) );
  AND U15870 ( .A(x[122]), .B(y[37]), .Z(n15431) );
  NAND U15871 ( .A(x[123]), .B(y[36]), .Z(n15430) );
  XNOR U15872 ( .A(n15431), .B(n15430), .Z(n15432) );
  XNOR U15873 ( .A(n15540), .B(n15432), .Z(n15433) );
  XNOR U15874 ( .A(n15434), .B(n15433), .Z(n15450) );
  AND U15875 ( .A(x[126]), .B(y[33]), .Z(n15436) );
  NAND U15876 ( .A(x[143]), .B(y[112]), .Z(n15435) );
  XNOR U15877 ( .A(n15436), .B(n15435), .Z(n15440) );
  AND U15878 ( .A(x[152]), .B(y[199]), .Z(n15438) );
  NAND U15879 ( .A(x[140]), .B(y[115]), .Z(n15437) );
  XNOR U15880 ( .A(n15438), .B(n15437), .Z(n15439) );
  XOR U15881 ( .A(n15440), .B(n15439), .Z(n15448) );
  AND U15882 ( .A(x[139]), .B(y[116]), .Z(n15442) );
  NAND U15883 ( .A(x[159]), .B(y[192]), .Z(n15441) );
  XNOR U15884 ( .A(n15442), .B(n15441), .Z(n15446) );
  AND U15885 ( .A(x[158]), .B(y[193]), .Z(n15444) );
  NAND U15886 ( .A(x[150]), .B(y[153]), .Z(n15443) );
  XNOR U15887 ( .A(n15444), .B(n15443), .Z(n15445) );
  XNOR U15888 ( .A(n15446), .B(n15445), .Z(n15447) );
  XNOR U15889 ( .A(n15448), .B(n15447), .Z(n15449) );
  XOR U15890 ( .A(n15450), .B(n15449), .Z(n15472) );
  AND U15891 ( .A(x[121]), .B(y[38]), .Z(n15452) );
  NAND U15892 ( .A(x[155]), .B(y[196]), .Z(n15451) );
  XNOR U15893 ( .A(n15452), .B(n15451), .Z(n15456) );
  AND U15894 ( .A(x[137]), .B(y[118]), .Z(n15454) );
  NAND U15895 ( .A(x[124]), .B(y[35]), .Z(n15453) );
  XNOR U15896 ( .A(n15454), .B(n15453), .Z(n15455) );
  XOR U15897 ( .A(n15456), .B(n15455), .Z(n15464) );
  AND U15898 ( .A(x[127]), .B(y[32]), .Z(n15458) );
  NAND U15899 ( .A(x[147]), .B(y[156]), .Z(n15457) );
  XNOR U15900 ( .A(n15458), .B(n15457), .Z(n15462) );
  AND U15901 ( .A(x[136]), .B(y[119]), .Z(n15460) );
  NAND U15902 ( .A(x[154]), .B(y[197]), .Z(n15459) );
  XNOR U15903 ( .A(n15460), .B(n15459), .Z(n15461) );
  XNOR U15904 ( .A(n15462), .B(n15461), .Z(n15463) );
  XNOR U15905 ( .A(n15464), .B(n15463), .Z(n15470) );
  AND U15906 ( .A(y[117]), .B(x[138]), .Z(n15558) );
  XOR U15907 ( .A(n15465), .B(n15558), .Z(n15468) );
  AND U15908 ( .A(y[194]), .B(x[157]), .Z(n15554) );
  XNOR U15909 ( .A(n15466), .B(n15554), .Z(n15467) );
  XNOR U15910 ( .A(n15468), .B(n15467), .Z(n15469) );
  XNOR U15911 ( .A(n15470), .B(n15469), .Z(n15471) );
  XNOR U15912 ( .A(n15472), .B(n15471), .Z(n15473) );
  XNOR U15913 ( .A(n15474), .B(n15473), .Z(n15475) );
  XNOR U15914 ( .A(n15476), .B(n15475), .Z(n15523) );
  NAND U15915 ( .A(n15478), .B(n15477), .Z(n15482) );
  ANDN U15916 ( .B(n15480), .A(n15479), .Z(n15481) );
  ANDN U15917 ( .B(n15482), .A(n15481), .Z(n15513) );
  NAND U15918 ( .A(n15484), .B(n15483), .Z(n15488) );
  AND U15919 ( .A(n15486), .B(n15485), .Z(n15487) );
  ANDN U15920 ( .B(n15488), .A(n15487), .Z(n15496) );
  AND U15921 ( .A(n15490), .B(n15489), .Z(n15494) );
  AND U15922 ( .A(n15492), .B(n15491), .Z(n15493) );
  OR U15923 ( .A(n15494), .B(n15493), .Z(n15495) );
  XNOR U15924 ( .A(n15496), .B(n15495), .Z(n15511) );
  NAND U15925 ( .A(n15498), .B(n15497), .Z(n15502) );
  NAND U15926 ( .A(n15500), .B(n15499), .Z(n15501) );
  AND U15927 ( .A(n15502), .B(n15501), .Z(n15509) );
  NAND U15928 ( .A(n15504), .B(n15503), .Z(n15507) );
  AND U15929 ( .A(y[34]), .B(x[125]), .Z(n15573) );
  NAND U15930 ( .A(n15505), .B(n15573), .Z(n15506) );
  NAND U15931 ( .A(n15507), .B(n15506), .Z(n15508) );
  XNOR U15932 ( .A(n15509), .B(n15508), .Z(n15510) );
  XNOR U15933 ( .A(n15511), .B(n15510), .Z(n15512) );
  XNOR U15934 ( .A(n15513), .B(n15512), .Z(n15521) );
  NANDN U15935 ( .A(n15515), .B(n15514), .Z(n15519) );
  NANDN U15936 ( .A(n15517), .B(n15516), .Z(n15518) );
  NAND U15937 ( .A(n15519), .B(n15518), .Z(n15520) );
  XNOR U15938 ( .A(n15521), .B(n15520), .Z(n15522) );
  XNOR U15939 ( .A(n15523), .B(n15522), .Z(n15524) );
  XNOR U15940 ( .A(n15525), .B(n15524), .Z(n15633) );
  NAND U15941 ( .A(n15527), .B(n15526), .Z(n15531) );
  NAND U15942 ( .A(n15529), .B(n15528), .Z(n15530) );
  AND U15943 ( .A(n15531), .B(n15530), .Z(n15631) );
  NAND U15944 ( .A(n15533), .B(n15532), .Z(n15537) );
  AND U15945 ( .A(n15535), .B(n15534), .Z(n15536) );
  ANDN U15946 ( .B(n15537), .A(n15536), .Z(n15613) );
  NAND U15947 ( .A(n15539), .B(n15538), .Z(n15543) );
  NAND U15948 ( .A(n15541), .B(n15540), .Z(n15542) );
  AND U15949 ( .A(n15543), .B(n15542), .Z(n15551) );
  NAND U15950 ( .A(n15545), .B(n15544), .Z(n15549) );
  NAND U15951 ( .A(n15547), .B(n15546), .Z(n15548) );
  NAND U15952 ( .A(n15549), .B(n15548), .Z(n15550) );
  XNOR U15953 ( .A(n15551), .B(n15550), .Z(n15611) );
  AND U15954 ( .A(x[144]), .B(y[159]), .Z(n15553) );
  NAND U15955 ( .A(x[129]), .B(y[78]), .Z(n15552) );
  XNOR U15956 ( .A(n15553), .B(n15552), .Z(n15577) );
  AND U15957 ( .A(y[193]), .B(x[156]), .Z(n15555) );
  AND U15958 ( .A(n15555), .B(n15554), .Z(n15571) );
  NAND U15959 ( .A(n15557), .B(n15556), .Z(n15561) );
  NAND U15960 ( .A(n15559), .B(n15558), .Z(n15560) );
  AND U15961 ( .A(n15561), .B(n15560), .Z(n15569) );
  AND U15962 ( .A(x[130]), .B(y[77]), .Z(n15563) );
  NAND U15963 ( .A(x[133]), .B(y[74]), .Z(n15562) );
  XNOR U15964 ( .A(n15563), .B(n15562), .Z(n15567) );
  AND U15965 ( .A(x[146]), .B(y[157]), .Z(n15565) );
  NAND U15966 ( .A(x[135]), .B(y[72]), .Z(n15564) );
  XNOR U15967 ( .A(n15565), .B(n15564), .Z(n15566) );
  XNOR U15968 ( .A(n15567), .B(n15566), .Z(n15568) );
  XNOR U15969 ( .A(n15569), .B(n15568), .Z(n15570) );
  XOR U15970 ( .A(n15571), .B(n15570), .Z(n15575) );
  XNOR U15971 ( .A(n15573), .B(n15572), .Z(n15574) );
  XNOR U15972 ( .A(n15575), .B(n15574), .Z(n15576) );
  XOR U15973 ( .A(n15577), .B(n15576), .Z(n15609) );
  NAND U15974 ( .A(n15579), .B(n15578), .Z(n15583) );
  NAND U15975 ( .A(n15581), .B(n15580), .Z(n15582) );
  AND U15976 ( .A(n15583), .B(n15582), .Z(n15591) );
  NAND U15977 ( .A(n15585), .B(n15584), .Z(n15589) );
  NAND U15978 ( .A(n15587), .B(n15586), .Z(n15588) );
  NAND U15979 ( .A(n15589), .B(n15588), .Z(n15590) );
  XNOR U15980 ( .A(n15591), .B(n15590), .Z(n15607) );
  NAND U15981 ( .A(n15593), .B(n15592), .Z(n15597) );
  NAND U15982 ( .A(n15595), .B(n15594), .Z(n15596) );
  AND U15983 ( .A(n15597), .B(n15596), .Z(n15605) );
  NAND U15984 ( .A(n15599), .B(n15598), .Z(n15603) );
  NAND U15985 ( .A(n15601), .B(n15600), .Z(n15602) );
  NAND U15986 ( .A(n15603), .B(n15602), .Z(n15604) );
  XNOR U15987 ( .A(n15605), .B(n15604), .Z(n15606) );
  XNOR U15988 ( .A(n15607), .B(n15606), .Z(n15608) );
  XNOR U15989 ( .A(n15609), .B(n15608), .Z(n15610) );
  XNOR U15990 ( .A(n15611), .B(n15610), .Z(n15612) );
  XNOR U15991 ( .A(n15613), .B(n15612), .Z(n15629) );
  NAND U15992 ( .A(n15615), .B(n15614), .Z(n15619) );
  NANDN U15993 ( .A(n15617), .B(n15616), .Z(n15618) );
  AND U15994 ( .A(n15619), .B(n15618), .Z(n15627) );
  NAND U15995 ( .A(n15621), .B(n15620), .Z(n15625) );
  NANDN U15996 ( .A(n15623), .B(n15622), .Z(n15624) );
  NAND U15997 ( .A(n15625), .B(n15624), .Z(n15626) );
  XNOR U15998 ( .A(n15627), .B(n15626), .Z(n15628) );
  XNOR U15999 ( .A(n15629), .B(n15628), .Z(n15630) );
  XNOR U16000 ( .A(n15631), .B(n15630), .Z(n15632) );
  XNOR U16001 ( .A(n15633), .B(n15632), .Z(n15634) );
  XNOR U16002 ( .A(n15635), .B(n15634), .Z(n15636) );
  XNOR U16003 ( .A(n15637), .B(n15636), .Z(n15638) );
  NANDN U16004 ( .A(n15641), .B(n15640), .Z(n15645) );
  ANDN U16005 ( .B(n15643), .A(n15642), .Z(n15644) );
  ANDN U16006 ( .B(n15645), .A(n15644), .Z(n15653) );
  AND U16007 ( .A(n15647), .B(n15646), .Z(n15651) );
  ANDN U16008 ( .B(n15649), .A(n15648), .Z(n15650) );
  OR U16009 ( .A(n15651), .B(n15650), .Z(n15652) );
  IV U16010 ( .A(n15654), .Z(n15656) );
  ANDN U16011 ( .B(n15656), .A(n15655), .Z(n15657) );
  NAND U16012 ( .A(y[160]), .B(x[192]), .Z(n15814) );
  NAND U16013 ( .A(y[40]), .B(x[168]), .Z(n15668) );
  XOR U16014 ( .A(n15814), .B(n15668), .Z(n15669) );
  AND U16015 ( .A(y[0]), .B(x[160]), .Z(n15676) );
  AND U16016 ( .A(y[80]), .B(x[176]), .Z(n15673) );
  XOR U16017 ( .A(n15676), .B(n15673), .Z(n15672) );
  AND U16018 ( .A(y[120]), .B(x[184]), .Z(n15671) );
  XNOR U16019 ( .A(n15672), .B(n15671), .Z(n15670) );
  XNOR U16020 ( .A(n15669), .B(n15670), .Z(o[160]) );
  AND U16021 ( .A(x[160]), .B(y[1]), .Z(n15667) );
  NAND U16022 ( .A(x[161]), .B(y[0]), .Z(n15666) );
  XNOR U16023 ( .A(n15667), .B(n15666), .Z(n15677) );
  NAND U16024 ( .A(y[40]), .B(x[169]), .Z(n15678) );
  XOR U16025 ( .A(n15677), .B(n15678), .Z(n15694) );
  AND U16026 ( .A(y[160]), .B(x[193]), .Z(n15902) );
  NAND U16027 ( .A(y[81]), .B(x[176]), .Z(n15681) );
  XNOR U16028 ( .A(n15902), .B(n15681), .Z(n15682) );
  AND U16029 ( .A(y[161]), .B(x[192]), .Z(n15705) );
  NAND U16030 ( .A(y[80]), .B(x[177]), .Z(n15704) );
  XOR U16031 ( .A(n15705), .B(n15704), .Z(n15683) );
  XOR U16032 ( .A(n15682), .B(n15683), .Z(n15693) );
  AND U16033 ( .A(y[41]), .B(x[168]), .Z(n15927) );
  AND U16034 ( .A(y[121]), .B(x[184]), .Z(n15698) );
  XOR U16035 ( .A(n15927), .B(n15698), .Z(n15700) );
  AND U16036 ( .A(y[120]), .B(x[185]), .Z(n15699) );
  XNOR U16037 ( .A(n15700), .B(n15699), .Z(n15692) );
  XOR U16038 ( .A(n15693), .B(n15692), .Z(n15695) );
  XOR U16039 ( .A(n15694), .B(n15695), .Z(n15689) );
  NAND U16040 ( .A(n15672), .B(n15671), .Z(n15675) );
  AND U16041 ( .A(n15676), .B(n15673), .Z(n15674) );
  ANDN U16042 ( .B(n15675), .A(n15674), .Z(n15686) );
  XNOR U16043 ( .A(n15687), .B(n15686), .Z(n15688) );
  XNOR U16044 ( .A(n15689), .B(n15688), .Z(o[161]) );
  AND U16045 ( .A(y[1]), .B(x[161]), .Z(n15736) );
  NAND U16046 ( .A(n15736), .B(n15676), .Z(n15680) );
  NANDN U16047 ( .A(n15678), .B(n15677), .Z(n15679) );
  NAND U16048 ( .A(n15680), .B(n15679), .Z(n15748) );
  NANDN U16049 ( .A(n15681), .B(n15902), .Z(n15685) );
  NANDN U16050 ( .A(n15683), .B(n15682), .Z(n15684) );
  NAND U16051 ( .A(n15685), .B(n15684), .Z(n15746) );
  AND U16052 ( .A(y[122]), .B(x[184]), .Z(n15752) );
  NAND U16053 ( .A(y[2]), .B(x[160]), .Z(n15753) );
  XNOR U16054 ( .A(n15752), .B(n15753), .Z(n15755) );
  AND U16055 ( .A(y[40]), .B(x[170]), .Z(n15754) );
  XOR U16056 ( .A(n15755), .B(n15754), .Z(n15747) );
  XOR U16057 ( .A(n15746), .B(n15747), .Z(n15749) );
  XNOR U16058 ( .A(n15748), .B(n15749), .Z(n15707) );
  NANDN U16059 ( .A(n15687), .B(n15686), .Z(n15691) );
  NAND U16060 ( .A(n15689), .B(n15688), .Z(n15690) );
  NAND U16061 ( .A(n15691), .B(n15690), .Z(n15706) );
  XOR U16062 ( .A(n15707), .B(n15706), .Z(n15709) );
  NAND U16063 ( .A(n15693), .B(n15692), .Z(n15697) );
  NAND U16064 ( .A(n15695), .B(n15694), .Z(n15696) );
  AND U16065 ( .A(n15697), .B(n15696), .Z(n15715) );
  AND U16066 ( .A(y[0]), .B(x[162]), .Z(n15734) );
  AND U16067 ( .A(y[82]), .B(x[176]), .Z(n15733) );
  XOR U16068 ( .A(n15734), .B(n15733), .Z(n15735) );
  XOR U16069 ( .A(n15736), .B(n15735), .Z(n15761) );
  AND U16070 ( .A(y[120]), .B(x[186]), .Z(n15760) );
  XOR U16071 ( .A(n15761), .B(n15760), .Z(n15763) );
  AND U16072 ( .A(y[80]), .B(x[178]), .Z(n15831) );
  AND U16073 ( .A(y[162]), .B(x[192]), .Z(n15724) );
  XOR U16074 ( .A(n15831), .B(n15724), .Z(n15726) );
  AND U16075 ( .A(y[81]), .B(x[177]), .Z(n15725) );
  XOR U16076 ( .A(n15726), .B(n15725), .Z(n15762) );
  XOR U16077 ( .A(n15763), .B(n15762), .Z(n15712) );
  AND U16078 ( .A(n15927), .B(n15698), .Z(n15702) );
  NAND U16079 ( .A(n15700), .B(n15699), .Z(n15701) );
  NANDN U16080 ( .A(n15702), .B(n15701), .Z(n15720) );
  AND U16081 ( .A(x[193]), .B(y[161]), .Z(n15792) );
  NAND U16082 ( .A(x[194]), .B(y[160]), .Z(n15703) );
  XNOR U16083 ( .A(n15792), .B(n15703), .Z(n15759) );
  ANDN U16084 ( .B(n15705), .A(n15704), .Z(n15758) );
  XOR U16085 ( .A(n15759), .B(n15758), .Z(n15719) );
  AND U16086 ( .A(y[121]), .B(x[185]), .Z(n15739) );
  NAND U16087 ( .A(y[41]), .B(x[169]), .Z(n15740) );
  XNOR U16088 ( .A(n15739), .B(n15740), .Z(n15741) );
  NAND U16089 ( .A(y[42]), .B(x[168]), .Z(n15742) );
  XNOR U16090 ( .A(n15741), .B(n15742), .Z(n15718) );
  XOR U16091 ( .A(n15719), .B(n15718), .Z(n15721) );
  XOR U16092 ( .A(n15720), .B(n15721), .Z(n15713) );
  XOR U16093 ( .A(n15712), .B(n15713), .Z(n15714) );
  XNOR U16094 ( .A(n15715), .B(n15714), .Z(n15708) );
  XNOR U16095 ( .A(n15709), .B(n15708), .Z(o[162]) );
  NAND U16096 ( .A(n15707), .B(n15706), .Z(n15711) );
  NAND U16097 ( .A(n15709), .B(n15708), .Z(n15710) );
  AND U16098 ( .A(n15711), .B(n15710), .Z(n15767) );
  NAND U16099 ( .A(n15713), .B(n15712), .Z(n15717) );
  NAND U16100 ( .A(n15715), .B(n15714), .Z(n15716) );
  NAND U16101 ( .A(n15717), .B(n15716), .Z(n15772) );
  NAND U16102 ( .A(n15719), .B(n15718), .Z(n15723) );
  NAND U16103 ( .A(n15721), .B(n15720), .Z(n15722) );
  NAND U16104 ( .A(n15723), .B(n15722), .Z(n15770) );
  NAND U16105 ( .A(n15831), .B(n15724), .Z(n15728) );
  AND U16106 ( .A(n15726), .B(n15725), .Z(n15727) );
  ANDN U16107 ( .B(n15728), .A(n15727), .Z(n15828) );
  AND U16108 ( .A(y[2]), .B(x[161]), .Z(n15810) );
  AND U16109 ( .A(y[1]), .B(x[162]), .Z(n15809) );
  NAND U16110 ( .A(y[122]), .B(x[185]), .Z(n15808) );
  XOR U16111 ( .A(n15809), .B(n15808), .Z(n15811) );
  XOR U16112 ( .A(n15810), .B(n15811), .Z(n15826) );
  AND U16113 ( .A(x[195]), .B(y[160]), .Z(n15730) );
  NAND U16114 ( .A(x[192]), .B(y[163]), .Z(n15729) );
  XNOR U16115 ( .A(n15730), .B(n15729), .Z(n15815) );
  AND U16116 ( .A(x[193]), .B(y[162]), .Z(n15732) );
  NAND U16117 ( .A(x[194]), .B(y[161]), .Z(n15731) );
  XOR U16118 ( .A(n15732), .B(n15731), .Z(n15816) );
  XNOR U16119 ( .A(n15815), .B(n15816), .Z(n15825) );
  XNOR U16120 ( .A(n15826), .B(n15825), .Z(n15827) );
  XNOR U16121 ( .A(n15828), .B(n15827), .Z(n15784) );
  NAND U16122 ( .A(n15734), .B(n15733), .Z(n15738) );
  NAND U16123 ( .A(n15736), .B(n15735), .Z(n15737) );
  NAND U16124 ( .A(n15738), .B(n15737), .Z(n15782) );
  NANDN U16125 ( .A(n15740), .B(n15739), .Z(n15744) );
  NANDN U16126 ( .A(n15742), .B(n15741), .Z(n15743) );
  AND U16127 ( .A(n15744), .B(n15743), .Z(n15821) );
  AND U16128 ( .A(y[123]), .B(x[184]), .Z(n15850) );
  AND U16129 ( .A(y[83]), .B(x[176]), .Z(n15849) );
  NAND U16130 ( .A(y[0]), .B(x[163]), .Z(n15848) );
  XOR U16131 ( .A(n15849), .B(n15848), .Z(n15851) );
  XOR U16132 ( .A(n15850), .B(n15851), .Z(n15820) );
  AND U16133 ( .A(y[81]), .B(x[178]), .Z(n15882) );
  NAND U16134 ( .A(x[179]), .B(y[80]), .Z(n15745) );
  XNOR U16135 ( .A(n15882), .B(n15745), .Z(n15833) );
  NAND U16136 ( .A(y[82]), .B(x[177]), .Z(n15834) );
  XNOR U16137 ( .A(n15833), .B(n15834), .Z(n15819) );
  XOR U16138 ( .A(n15820), .B(n15819), .Z(n15822) );
  XOR U16139 ( .A(n15821), .B(n15822), .Z(n15783) );
  XOR U16140 ( .A(n15782), .B(n15783), .Z(n15785) );
  XOR U16141 ( .A(n15784), .B(n15785), .Z(n15771) );
  XOR U16142 ( .A(n15770), .B(n15771), .Z(n15773) );
  XOR U16143 ( .A(n15772), .B(n15773), .Z(n15766) );
  XOR U16144 ( .A(n15767), .B(n15766), .Z(n15769) );
  NAND U16145 ( .A(n15747), .B(n15746), .Z(n15751) );
  NAND U16146 ( .A(n15749), .B(n15748), .Z(n15750) );
  AND U16147 ( .A(n15751), .B(n15750), .Z(n15779) );
  NANDN U16148 ( .A(n15753), .B(n15752), .Z(n15757) );
  NAND U16149 ( .A(n15755), .B(n15754), .Z(n15756) );
  AND U16150 ( .A(n15757), .B(n15756), .Z(n15789) );
  AND U16151 ( .A(y[161]), .B(x[194]), .Z(n15901) );
  XNOR U16152 ( .A(n15789), .B(n15788), .Z(n15791) );
  NAND U16153 ( .A(y[40]), .B(x[171]), .Z(n15842) );
  NAND U16154 ( .A(y[3]), .B(x[160]), .Z(n15840) );
  NAND U16155 ( .A(y[121]), .B(x[186]), .Z(n15839) );
  XOR U16156 ( .A(n15840), .B(n15839), .Z(n15841) );
  XNOR U16157 ( .A(n15842), .B(n15841), .Z(n15802) );
  NAND U16158 ( .A(y[43]), .B(x[168]), .Z(n15796) );
  NAND U16159 ( .A(y[41]), .B(x[170]), .Z(n15794) );
  NAND U16160 ( .A(y[120]), .B(x[187]), .Z(n15793) );
  XOR U16161 ( .A(n15794), .B(n15793), .Z(n15795) );
  XNOR U16162 ( .A(n15796), .B(n15795), .Z(n15800) );
  AND U16163 ( .A(y[42]), .B(x[169]), .Z(n15799) );
  XOR U16164 ( .A(n15800), .B(n15799), .Z(n15801) );
  XOR U16165 ( .A(n15802), .B(n15801), .Z(n15790) );
  XNOR U16166 ( .A(n15791), .B(n15790), .Z(n15777) );
  NAND U16167 ( .A(n15761), .B(n15760), .Z(n15765) );
  NAND U16168 ( .A(n15763), .B(n15762), .Z(n15764) );
  AND U16169 ( .A(n15765), .B(n15764), .Z(n15776) );
  XOR U16170 ( .A(n15777), .B(n15776), .Z(n15778) );
  XNOR U16171 ( .A(n15779), .B(n15778), .Z(n15768) );
  XOR U16172 ( .A(n15769), .B(n15768), .Z(o[163]) );
  NAND U16173 ( .A(n15771), .B(n15770), .Z(n15775) );
  NAND U16174 ( .A(n15773), .B(n15772), .Z(n15774) );
  AND U16175 ( .A(n15775), .B(n15774), .Z(n15860) );
  NAND U16176 ( .A(n15777), .B(n15776), .Z(n15781) );
  NAND U16177 ( .A(n15779), .B(n15778), .Z(n15780) );
  NAND U16178 ( .A(n15781), .B(n15780), .Z(n15858) );
  NAND U16179 ( .A(n15783), .B(n15782), .Z(n15787) );
  NAND U16180 ( .A(n15785), .B(n15784), .Z(n15786) );
  AND U16181 ( .A(n15787), .B(n15786), .Z(n15859) );
  XOR U16182 ( .A(n15858), .B(n15859), .Z(n15861) );
  XOR U16183 ( .A(n15860), .B(n15861), .Z(n15854) );
  XOR U16184 ( .A(n15855), .B(n15854), .Z(n15857) );
  NAND U16185 ( .A(y[0]), .B(x[164]), .Z(n15911) );
  NAND U16186 ( .A(y[122]), .B(x[186]), .Z(n15910) );
  NAND U16187 ( .A(y[84]), .B(x[176]), .Z(n15909) );
  XNOR U16188 ( .A(n15910), .B(n15909), .Z(n15912) );
  AND U16189 ( .A(y[162]), .B(x[194]), .Z(n15847) );
  NAND U16190 ( .A(n15847), .B(n15792), .Z(n15907) );
  NAND U16191 ( .A(y[164]), .B(x[192]), .Z(n16057) );
  NAND U16192 ( .A(y[80]), .B(x[180]), .Z(n16008) );
  XNOR U16193 ( .A(n16057), .B(n16008), .Z(n15908) );
  XOR U16194 ( .A(n15907), .B(n15908), .Z(n15870) );
  XOR U16195 ( .A(n15871), .B(n15870), .Z(n15873) );
  NAND U16196 ( .A(n15794), .B(n15793), .Z(n15798) );
  NAND U16197 ( .A(n15796), .B(n15795), .Z(n15797) );
  AND U16198 ( .A(n15798), .B(n15797), .Z(n15872) );
  XOR U16199 ( .A(n15873), .B(n15872), .Z(n15958) );
  NAND U16200 ( .A(n15800), .B(n15799), .Z(n15804) );
  NAND U16201 ( .A(n15802), .B(n15801), .Z(n15803) );
  AND U16202 ( .A(n15804), .B(n15803), .Z(n15957) );
  XNOR U16203 ( .A(n15958), .B(n15957), .Z(n15960) );
  AND U16204 ( .A(y[42]), .B(x[170]), .Z(n15993) );
  AND U16205 ( .A(x[171]), .B(y[41]), .Z(n15806) );
  NAND U16206 ( .A(x[168]), .B(y[44]), .Z(n15805) );
  XOR U16207 ( .A(n15806), .B(n15805), .Z(n15928) );
  IV U16208 ( .A(n15928), .Z(n15807) );
  XOR U16209 ( .A(n15993), .B(n15807), .Z(n15931) );
  NAND U16210 ( .A(y[43]), .B(x[169]), .Z(n15932) );
  AND U16211 ( .A(y[120]), .B(x[188]), .Z(n15887) );
  NAND U16212 ( .A(y[3]), .B(x[161]), .Z(n15888) );
  NAND U16213 ( .A(y[4]), .B(x[160]), .Z(n15890) );
  XOR U16214 ( .A(n15934), .B(n15933), .Z(n15946) );
  NANDN U16215 ( .A(n15809), .B(n15808), .Z(n15813) );
  OR U16216 ( .A(n15811), .B(n15810), .Z(n15812) );
  AND U16217 ( .A(n15813), .B(n15812), .Z(n15944) );
  AND U16218 ( .A(y[163]), .B(x[195]), .Z(n16155) );
  NANDN U16219 ( .A(n15814), .B(n16155), .Z(n15818) );
  NANDN U16220 ( .A(n15816), .B(n15815), .Z(n15817) );
  AND U16221 ( .A(n15818), .B(n15817), .Z(n15943) );
  XNOR U16222 ( .A(n15960), .B(n15959), .Z(n15864) );
  XNOR U16223 ( .A(n15865), .B(n15864), .Z(n15867) );
  NANDN U16224 ( .A(n15820), .B(n15819), .Z(n15824) );
  OR U16225 ( .A(n15822), .B(n15821), .Z(n15823) );
  AND U16226 ( .A(n15824), .B(n15823), .Z(n15950) );
  NANDN U16227 ( .A(n15826), .B(n15825), .Z(n15830) );
  NANDN U16228 ( .A(n15828), .B(n15827), .Z(n15829) );
  NAND U16229 ( .A(n15830), .B(n15829), .Z(n15949) );
  XNOR U16230 ( .A(n15950), .B(n15949), .Z(n15952) );
  AND U16231 ( .A(y[81]), .B(x[179]), .Z(n15832) );
  NAND U16232 ( .A(n15832), .B(n15831), .Z(n15836) );
  NANDN U16233 ( .A(n15834), .B(n15833), .Z(n15835) );
  AND U16234 ( .A(n15836), .B(n15835), .Z(n15954) );
  AND U16235 ( .A(y[40]), .B(x[172]), .Z(n15893) );
  NAND U16236 ( .A(y[124]), .B(x[184]), .Z(n15894) );
  NAND U16237 ( .A(y[123]), .B(x[185]), .Z(n15896) );
  AND U16238 ( .A(x[178]), .B(y[82]), .Z(n15838) );
  NAND U16239 ( .A(x[179]), .B(y[81]), .Z(n15837) );
  XNOR U16240 ( .A(n15838), .B(n15837), .Z(n15883) );
  NAND U16241 ( .A(y[83]), .B(x[177]), .Z(n15884) );
  XOR U16242 ( .A(n15938), .B(n15937), .Z(n15939) );
  NAND U16243 ( .A(n15840), .B(n15839), .Z(n15844) );
  NAND U16244 ( .A(n15842), .B(n15841), .Z(n15843) );
  NAND U16245 ( .A(n15844), .B(n15843), .Z(n15940) );
  XNOR U16246 ( .A(n15954), .B(n15953), .Z(n15956) );
  NAND U16247 ( .A(y[2]), .B(x[162]), .Z(n15923) );
  NAND U16248 ( .A(y[121]), .B(x[187]), .Z(n15922) );
  NAND U16249 ( .A(y[1]), .B(x[163]), .Z(n15921) );
  XNOR U16250 ( .A(n15922), .B(n15921), .Z(n15924) );
  AND U16251 ( .A(x[196]), .B(y[160]), .Z(n15846) );
  NAND U16252 ( .A(x[193]), .B(y[163]), .Z(n15845) );
  XNOR U16253 ( .A(n15846), .B(n15845), .Z(n15904) );
  AND U16254 ( .A(y[161]), .B(x[195]), .Z(n16015) );
  XOR U16255 ( .A(n15847), .B(n16015), .Z(n15903) );
  XOR U16256 ( .A(n15904), .B(n15903), .Z(n15877) );
  XOR U16257 ( .A(n15876), .B(n15877), .Z(n15878) );
  NANDN U16258 ( .A(n15849), .B(n15848), .Z(n15853) );
  OR U16259 ( .A(n15851), .B(n15850), .Z(n15852) );
  NAND U16260 ( .A(n15853), .B(n15852), .Z(n15879) );
  XOR U16261 ( .A(n15956), .B(n15955), .Z(n15951) );
  XOR U16262 ( .A(n15952), .B(n15951), .Z(n15866) );
  XNOR U16263 ( .A(n15867), .B(n15866), .Z(n15856) );
  XNOR U16264 ( .A(n15857), .B(n15856), .Z(o[164]) );
  NAND U16265 ( .A(n15859), .B(n15858), .Z(n15863) );
  NAND U16266 ( .A(n15861), .B(n15860), .Z(n15862) );
  NAND U16267 ( .A(n15863), .B(n15862), .Z(n16106) );
  XNOR U16268 ( .A(n16105), .B(n16106), .Z(n16108) );
  NANDN U16269 ( .A(n15865), .B(n15864), .Z(n15869) );
  NAND U16270 ( .A(n15867), .B(n15866), .Z(n15868) );
  AND U16271 ( .A(n15869), .B(n15868), .Z(n15964) );
  NAND U16272 ( .A(n15871), .B(n15870), .Z(n15875) );
  NAND U16273 ( .A(n15873), .B(n15872), .Z(n15874) );
  AND U16274 ( .A(n15875), .B(n15874), .Z(n16017) );
  NAND U16275 ( .A(n15877), .B(n15876), .Z(n15881) );
  NANDN U16276 ( .A(n15879), .B(n15878), .Z(n15880) );
  NAND U16277 ( .A(n15881), .B(n15880), .Z(n16016) );
  AND U16278 ( .A(y[82]), .B(x[179]), .Z(n16009) );
  NAND U16279 ( .A(n16009), .B(n15882), .Z(n15886) );
  NANDN U16280 ( .A(n15884), .B(n15883), .Z(n15885) );
  AND U16281 ( .A(n15886), .B(n15885), .Z(n15970) );
  NANDN U16282 ( .A(n15888), .B(n15887), .Z(n15892) );
  NANDN U16283 ( .A(n15890), .B(n15889), .Z(n15891) );
  NAND U16284 ( .A(n15892), .B(n15891), .Z(n15977) );
  AND U16285 ( .A(y[125]), .B(x[184]), .Z(n16277) );
  AND U16286 ( .A(y[40]), .B(x[173]), .Z(n15999) );
  AND U16287 ( .A(y[83]), .B(x[178]), .Z(n15998) );
  XOR U16288 ( .A(n15999), .B(n15998), .Z(n16000) );
  XOR U16289 ( .A(n16277), .B(n16000), .Z(n15976) );
  AND U16290 ( .A(y[121]), .B(x[188]), .Z(n16004) );
  AND U16291 ( .A(y[0]), .B(x[165]), .Z(n16003) );
  XOR U16292 ( .A(n16004), .B(n16003), .Z(n16005) );
  AND U16293 ( .A(y[1]), .B(x[164]), .Z(n16336) );
  XOR U16294 ( .A(n16005), .B(n16336), .Z(n15975) );
  XOR U16295 ( .A(n15976), .B(n15975), .Z(n15978) );
  XOR U16296 ( .A(n15977), .B(n15978), .Z(n15969) );
  NANDN U16297 ( .A(n15894), .B(n15893), .Z(n15898) );
  NANDN U16298 ( .A(n15896), .B(n15895), .Z(n15897) );
  NAND U16299 ( .A(n15898), .B(n15897), .Z(n16090) );
  AND U16300 ( .A(x[192]), .B(y[165]), .Z(n15900) );
  NAND U16301 ( .A(x[193]), .B(y[164]), .Z(n15899) );
  XNOR U16302 ( .A(n15900), .B(n15899), .Z(n16059) );
  AND U16303 ( .A(y[162]), .B(x[195]), .Z(n15918) );
  AND U16304 ( .A(n15901), .B(n15918), .Z(n16058) );
  XOR U16305 ( .A(n16059), .B(n16058), .Z(n16089) );
  AND U16306 ( .A(y[45]), .B(x[168]), .Z(n16079) );
  AND U16307 ( .A(y[4]), .B(x[161]), .Z(n16078) );
  XOR U16308 ( .A(n16079), .B(n16078), .Z(n16081) );
  AND U16309 ( .A(y[41]), .B(x[172]), .Z(n16080) );
  XOR U16310 ( .A(n16081), .B(n16080), .Z(n16088) );
  XOR U16311 ( .A(n16089), .B(n16088), .Z(n16091) );
  XOR U16312 ( .A(n16090), .B(n16091), .Z(n15971) );
  XOR U16313 ( .A(n15972), .B(n15971), .Z(n16018) );
  XOR U16314 ( .A(n16019), .B(n16018), .Z(n16103) );
  AND U16315 ( .A(y[163]), .B(x[196]), .Z(n16210) );
  NAND U16316 ( .A(n16210), .B(n15902), .Z(n15906) );
  NAND U16317 ( .A(n15904), .B(n15903), .Z(n15905) );
  AND U16318 ( .A(n15906), .B(n15905), .Z(n16035) );
  NAND U16319 ( .A(n15910), .B(n15909), .Z(n15914) );
  NANDN U16320 ( .A(n15912), .B(n15911), .Z(n15913) );
  AND U16321 ( .A(n15914), .B(n15913), .Z(n16025) );
  AND U16322 ( .A(y[44]), .B(x[169]), .Z(n15994) );
  AND U16323 ( .A(x[170]), .B(y[43]), .Z(n15916) );
  NAND U16324 ( .A(x[171]), .B(y[42]), .Z(n15915) );
  XOR U16325 ( .A(n15916), .B(n15915), .Z(n15995) );
  NAND U16326 ( .A(x[196]), .B(y[161]), .Z(n15917) );
  XNOR U16327 ( .A(n15918), .B(n15917), .Z(n15984) );
  AND U16328 ( .A(y[160]), .B(x[197]), .Z(n15981) );
  NAND U16329 ( .A(y[163]), .B(x[194]), .Z(n15982) );
  XOR U16330 ( .A(n15984), .B(n15983), .Z(n16022) );
  XOR U16331 ( .A(n16023), .B(n16022), .Z(n16024) );
  XOR U16332 ( .A(n16025), .B(n16024), .Z(n16036) );
  XOR U16333 ( .A(n16037), .B(n16036), .Z(n16049) );
  AND U16334 ( .A(x[180]), .B(y[81]), .Z(n15920) );
  NAND U16335 ( .A(x[181]), .B(y[80]), .Z(n15919) );
  XOR U16336 ( .A(n15920), .B(n15919), .Z(n16010) );
  AND U16337 ( .A(y[120]), .B(x[189]), .Z(n15987) );
  NAND U16338 ( .A(y[2]), .B(x[163]), .Z(n15988) );
  AND U16339 ( .A(y[3]), .B(x[162]), .Z(n15989) );
  XOR U16340 ( .A(n15990), .B(n15989), .Z(n16070) );
  XOR U16341 ( .A(n16071), .B(n16070), .Z(n16073) );
  NAND U16342 ( .A(n15922), .B(n15921), .Z(n15926) );
  NANDN U16343 ( .A(n15924), .B(n15923), .Z(n15925) );
  AND U16344 ( .A(n15926), .B(n15925), .Z(n16072) );
  XOR U16345 ( .A(n16073), .B(n16072), .Z(n16047) );
  AND U16346 ( .A(y[44]), .B(x[171]), .Z(n16209) );
  NAND U16347 ( .A(n16209), .B(n15927), .Z(n15930) );
  NANDN U16348 ( .A(n15928), .B(n15993), .Z(n15929) );
  AND U16349 ( .A(n15930), .B(n15929), .Z(n16031) );
  AND U16350 ( .A(y[84]), .B(x[177]), .Z(n16292) );
  AND U16351 ( .A(y[122]), .B(x[187]), .Z(n16052) );
  XOR U16352 ( .A(n16292), .B(n16052), .Z(n16054) );
  AND U16353 ( .A(y[85]), .B(x[176]), .Z(n16053) );
  XOR U16354 ( .A(n16054), .B(n16053), .Z(n16029) );
  AND U16355 ( .A(y[5]), .B(x[160]), .Z(n16063) );
  AND U16356 ( .A(y[124]), .B(x[185]), .Z(n16062) );
  XOR U16357 ( .A(n16063), .B(n16062), .Z(n16065) );
  AND U16358 ( .A(y[123]), .B(x[186]), .Z(n16064) );
  XOR U16359 ( .A(n16065), .B(n16064), .Z(n16028) );
  XOR U16360 ( .A(n16029), .B(n16028), .Z(n16030) );
  XOR U16361 ( .A(n16031), .B(n16030), .Z(n16046) );
  NANDN U16362 ( .A(n15932), .B(n15931), .Z(n15936) );
  NAND U16363 ( .A(n15934), .B(n15933), .Z(n15935) );
  AND U16364 ( .A(n15936), .B(n15935), .Z(n16041) );
  NAND U16365 ( .A(n15938), .B(n15937), .Z(n15942) );
  NANDN U16366 ( .A(n15940), .B(n15939), .Z(n15941) );
  NAND U16367 ( .A(n15942), .B(n15941), .Z(n16040) );
  NANDN U16368 ( .A(n15944), .B(n15943), .Z(n15948) );
  NANDN U16369 ( .A(n15946), .B(n15945), .Z(n15947) );
  NAND U16370 ( .A(n15948), .B(n15947), .Z(n16043) );
  XOR U16371 ( .A(n16101), .B(n16100), .Z(n16102) );
  XOR U16372 ( .A(n16103), .B(n16102), .Z(n15963) );
  XNOR U16373 ( .A(n15964), .B(n15963), .Z(n15965) );
  NANDN U16374 ( .A(n15958), .B(n15957), .Z(n15962) );
  NAND U16375 ( .A(n15960), .B(n15959), .Z(n15961) );
  AND U16376 ( .A(n15962), .B(n15961), .Z(n16094) );
  XNOR U16377 ( .A(n16095), .B(n16094), .Z(n16096) );
  XOR U16378 ( .A(n16097), .B(n16096), .Z(n15966) );
  XNOR U16379 ( .A(n15965), .B(n15966), .Z(n16107) );
  XOR U16380 ( .A(n16108), .B(n16107), .Z(o[165]) );
  NANDN U16381 ( .A(n15964), .B(n15963), .Z(n15968) );
  NANDN U16382 ( .A(n15966), .B(n15965), .Z(n15967) );
  AND U16383 ( .A(n15968), .B(n15967), .Z(n16392) );
  NANDN U16384 ( .A(n15970), .B(n15969), .Z(n15974) );
  NAND U16385 ( .A(n15972), .B(n15971), .Z(n15973) );
  AND U16386 ( .A(n15974), .B(n15973), .Z(n16397) );
  NAND U16387 ( .A(n15976), .B(n15975), .Z(n15980) );
  NAND U16388 ( .A(n15978), .B(n15977), .Z(n15979) );
  NAND U16389 ( .A(n15980), .B(n15979), .Z(n16120) );
  NANDN U16390 ( .A(n15982), .B(n15981), .Z(n15986) );
  NAND U16391 ( .A(n15984), .B(n15983), .Z(n15985) );
  NAND U16392 ( .A(n15986), .B(n15985), .Z(n16262) );
  NANDN U16393 ( .A(n15988), .B(n15987), .Z(n15992) );
  NAND U16394 ( .A(n15990), .B(n15989), .Z(n15991) );
  NAND U16395 ( .A(n15992), .B(n15991), .Z(n16265) );
  AND U16396 ( .A(x[171]), .B(y[43]), .Z(n16077) );
  NAND U16397 ( .A(n16077), .B(n15993), .Z(n15997) );
  NANDN U16398 ( .A(n15995), .B(n15994), .Z(n15996) );
  AND U16399 ( .A(n15997), .B(n15996), .Z(n16356) );
  AND U16400 ( .A(y[123]), .B(x[187]), .Z(n16283) );
  AND U16401 ( .A(y[83]), .B(x[179]), .Z(n16282) );
  XOR U16402 ( .A(n16283), .B(n16282), .Z(n16281) );
  AND U16403 ( .A(y[3]), .B(x[163]), .Z(n16280) );
  XOR U16404 ( .A(n16281), .B(n16280), .Z(n16358) );
  AND U16405 ( .A(y[124]), .B(x[186]), .Z(n16249) );
  AND U16406 ( .A(y[82]), .B(x[180]), .Z(n16248) );
  XOR U16407 ( .A(n16249), .B(n16248), .Z(n16247) );
  AND U16408 ( .A(y[4]), .B(x[162]), .Z(n16246) );
  XNOR U16409 ( .A(n16247), .B(n16246), .Z(n16357) );
  XNOR U16410 ( .A(n16356), .B(n16355), .Z(n16264) );
  XOR U16411 ( .A(n16265), .B(n16264), .Z(n16263) );
  XOR U16412 ( .A(n16262), .B(n16263), .Z(n16121) );
  XOR U16413 ( .A(n16120), .B(n16121), .Z(n16119) );
  NAND U16414 ( .A(n15999), .B(n15998), .Z(n16002) );
  NAND U16415 ( .A(n16277), .B(n16000), .Z(n16001) );
  NAND U16416 ( .A(n16002), .B(n16001), .Z(n16145) );
  NAND U16417 ( .A(n16004), .B(n16003), .Z(n16007) );
  NAND U16418 ( .A(n16005), .B(n16336), .Z(n16006) );
  NAND U16419 ( .A(n16007), .B(n16006), .Z(n16144) );
  XOR U16420 ( .A(n16145), .B(n16144), .Z(n16143) );
  AND U16421 ( .A(y[81]), .B(x[181]), .Z(n16330) );
  NANDN U16422 ( .A(n16008), .B(n16330), .Z(n16012) );
  NANDN U16423 ( .A(n16010), .B(n16009), .Z(n16011) );
  AND U16424 ( .A(n16012), .B(n16011), .Z(n16269) );
  AND U16425 ( .A(x[165]), .B(y[1]), .Z(n16014) );
  NAND U16426 ( .A(x[164]), .B(y[2]), .Z(n16013) );
  XNOR U16427 ( .A(n16014), .B(n16013), .Z(n16334) );
  AND U16428 ( .A(y[120]), .B(x[190]), .Z(n16333) );
  XOR U16429 ( .A(n16334), .B(n16333), .Z(n16271) );
  AND U16430 ( .A(y[165]), .B(x[193]), .Z(n16233) );
  AND U16431 ( .A(x[196]), .B(y[162]), .Z(n16069) );
  AND U16432 ( .A(n16069), .B(n16015), .Z(n16235) );
  AND U16433 ( .A(y[164]), .B(x[194]), .Z(n16234) );
  XOR U16434 ( .A(n16235), .B(n16234), .Z(n16232) );
  XNOR U16435 ( .A(n16233), .B(n16232), .Z(n16270) );
  XNOR U16436 ( .A(n16269), .B(n16268), .Z(n16142) );
  XOR U16437 ( .A(n16143), .B(n16142), .Z(n16118) );
  XOR U16438 ( .A(n16119), .B(n16118), .Z(n16117) );
  NANDN U16439 ( .A(n16017), .B(n16016), .Z(n16021) );
  NAND U16440 ( .A(n16019), .B(n16018), .Z(n16020) );
  AND U16441 ( .A(n16021), .B(n16020), .Z(n16116) );
  NAND U16442 ( .A(n16023), .B(n16022), .Z(n16027) );
  NAND U16443 ( .A(n16025), .B(n16024), .Z(n16026) );
  AND U16444 ( .A(n16027), .B(n16026), .Z(n16123) );
  NAND U16445 ( .A(n16029), .B(n16028), .Z(n16033) );
  NANDN U16446 ( .A(n16031), .B(n16030), .Z(n16032) );
  AND U16447 ( .A(n16033), .B(n16032), .Z(n16125) );
  NANDN U16448 ( .A(n16035), .B(n16034), .Z(n16039) );
  NAND U16449 ( .A(n16037), .B(n16036), .Z(n16038) );
  AND U16450 ( .A(n16039), .B(n16038), .Z(n16124) );
  XOR U16451 ( .A(n16125), .B(n16124), .Z(n16122) );
  XOR U16452 ( .A(n16123), .B(n16122), .Z(n16114) );
  XOR U16453 ( .A(n16115), .B(n16114), .Z(n16396) );
  XOR U16454 ( .A(n16397), .B(n16396), .Z(n16399) );
  NANDN U16455 ( .A(n16041), .B(n16040), .Z(n16045) );
  NANDN U16456 ( .A(n16043), .B(n16042), .Z(n16044) );
  AND U16457 ( .A(n16045), .B(n16044), .Z(n16376) );
  NANDN U16458 ( .A(n16047), .B(n16046), .Z(n16051) );
  NANDN U16459 ( .A(n16049), .B(n16048), .Z(n16050) );
  NAND U16460 ( .A(n16051), .B(n16050), .Z(n16377) );
  AND U16461 ( .A(n16292), .B(n16052), .Z(n16056) );
  NAND U16462 ( .A(n16054), .B(n16053), .Z(n16055) );
  NANDN U16463 ( .A(n16056), .B(n16055), .Z(n16134) );
  NANDN U16464 ( .A(n16057), .B(n16233), .Z(n16061) );
  NAND U16465 ( .A(n16059), .B(n16058), .Z(n16060) );
  NAND U16466 ( .A(n16061), .B(n16060), .Z(n16137) );
  NAND U16467 ( .A(n16063), .B(n16062), .Z(n16067) );
  NAND U16468 ( .A(n16065), .B(n16064), .Z(n16066) );
  AND U16469 ( .A(n16067), .B(n16066), .Z(n16350) );
  AND U16470 ( .A(y[5]), .B(x[161]), .Z(n16243) );
  AND U16471 ( .A(y[40]), .B(x[174]), .Z(n16242) );
  XOR U16472 ( .A(n16243), .B(n16242), .Z(n16241) );
  AND U16473 ( .A(y[46]), .B(x[168]), .Z(n16240) );
  XOR U16474 ( .A(n16241), .B(n16240), .Z(n16352) );
  NAND U16475 ( .A(x[197]), .B(y[161]), .Z(n16068) );
  XNOR U16476 ( .A(n16069), .B(n16068), .Z(n16157) );
  AND U16477 ( .A(y[160]), .B(x[198]), .Z(n16156) );
  XOR U16478 ( .A(n16157), .B(n16156), .Z(n16154) );
  XNOR U16479 ( .A(n16155), .B(n16154), .Z(n16351) );
  XNOR U16480 ( .A(n16350), .B(n16349), .Z(n16136) );
  XOR U16481 ( .A(n16137), .B(n16136), .Z(n16135) );
  XOR U16482 ( .A(n16134), .B(n16135), .Z(n16383) );
  NAND U16483 ( .A(n16071), .B(n16070), .Z(n16075) );
  NAND U16484 ( .A(n16073), .B(n16072), .Z(n16074) );
  AND U16485 ( .A(n16075), .B(n16074), .Z(n16382) );
  AND U16486 ( .A(y[86]), .B(x[176]), .Z(n16322) );
  AND U16487 ( .A(y[0]), .B(x[166]), .Z(n16321) );
  XOR U16488 ( .A(n16322), .B(n16321), .Z(n16320) );
  AND U16489 ( .A(y[121]), .B(x[189]), .Z(n16319) );
  XOR U16490 ( .A(n16320), .B(n16319), .Z(n16151) );
  AND U16491 ( .A(y[41]), .B(x[173]), .Z(n16316) );
  AND U16492 ( .A(y[44]), .B(x[170]), .Z(n16315) );
  XOR U16493 ( .A(n16316), .B(n16315), .Z(n16314) );
  AND U16494 ( .A(y[45]), .B(x[169]), .Z(n16313) );
  XOR U16495 ( .A(n16314), .B(n16313), .Z(n16228) );
  NAND U16496 ( .A(x[172]), .B(y[42]), .Z(n16076) );
  XNOR U16497 ( .A(n16077), .B(n16076), .Z(n16227) );
  XOR U16498 ( .A(n16228), .B(n16227), .Z(n16150) );
  XOR U16499 ( .A(n16151), .B(n16150), .Z(n16149) );
  AND U16500 ( .A(y[166]), .B(x[192]), .Z(n16329) );
  XOR U16501 ( .A(n16330), .B(n16329), .Z(n16328) );
  AND U16502 ( .A(y[80]), .B(x[182]), .Z(n16327) );
  XOR U16503 ( .A(n16328), .B(n16327), .Z(n16148) );
  XOR U16504 ( .A(n16149), .B(n16148), .Z(n16131) );
  NAND U16505 ( .A(n16079), .B(n16078), .Z(n16083) );
  NAND U16506 ( .A(n16081), .B(n16080), .Z(n16082) );
  AND U16507 ( .A(n16083), .B(n16082), .Z(n16221) );
  AND U16508 ( .A(y[122]), .B(x[188]), .Z(n16291) );
  AND U16509 ( .A(x[177]), .B(y[85]), .Z(n16085) );
  AND U16510 ( .A(x[178]), .B(y[84]), .Z(n16084) );
  XOR U16511 ( .A(n16085), .B(n16084), .Z(n16290) );
  XOR U16512 ( .A(n16291), .B(n16290), .Z(n16224) );
  AND U16513 ( .A(y[6]), .B(x[160]), .Z(n16275) );
  AND U16514 ( .A(y[126]), .B(x[184]), .Z(n16087) );
  AND U16515 ( .A(x[185]), .B(y[125]), .Z(n16086) );
  XOR U16516 ( .A(n16087), .B(n16086), .Z(n16274) );
  XNOR U16517 ( .A(n16275), .B(n16274), .Z(n16223) );
  XNOR U16518 ( .A(n16221), .B(n16222), .Z(n16130) );
  NAND U16519 ( .A(n16089), .B(n16088), .Z(n16093) );
  NAND U16520 ( .A(n16091), .B(n16090), .Z(n16092) );
  AND U16521 ( .A(n16093), .B(n16092), .Z(n16128) );
  XOR U16522 ( .A(n16129), .B(n16128), .Z(n16381) );
  XOR U16523 ( .A(n16382), .B(n16381), .Z(n16384) );
  XOR U16524 ( .A(n16377), .B(n16378), .Z(n16375) );
  XOR U16525 ( .A(n16376), .B(n16375), .Z(n16398) );
  XOR U16526 ( .A(n16399), .B(n16398), .Z(n16113) );
  NANDN U16527 ( .A(n16095), .B(n16094), .Z(n16099) );
  NANDN U16528 ( .A(n16097), .B(n16096), .Z(n16098) );
  AND U16529 ( .A(n16099), .B(n16098), .Z(n16112) );
  XOR U16530 ( .A(n16112), .B(n16111), .Z(n16104) );
  XOR U16531 ( .A(n16113), .B(n16104), .Z(n16393) );
  NANDN U16532 ( .A(n16106), .B(n16105), .Z(n16110) );
  NAND U16533 ( .A(n16108), .B(n16107), .Z(n16109) );
  NAND U16534 ( .A(n16110), .B(n16109), .Z(n16390) );
  XOR U16535 ( .A(n16391), .B(n16390), .Z(o[166]) );
  NAND U16536 ( .A(n16123), .B(n16122), .Z(n16127) );
  NAND U16537 ( .A(n16125), .B(n16124), .Z(n16126) );
  AND U16538 ( .A(n16127), .B(n16126), .Z(n16374) );
  NAND U16539 ( .A(n16129), .B(n16128), .Z(n16133) );
  NANDN U16540 ( .A(n16131), .B(n16130), .Z(n16132) );
  AND U16541 ( .A(n16133), .B(n16132), .Z(n16141) );
  NAND U16542 ( .A(n16135), .B(n16134), .Z(n16139) );
  NAND U16543 ( .A(n16137), .B(n16136), .Z(n16138) );
  NAND U16544 ( .A(n16139), .B(n16138), .Z(n16140) );
  XNOR U16545 ( .A(n16141), .B(n16140), .Z(n16372) );
  NAND U16546 ( .A(n16143), .B(n16142), .Z(n16147) );
  NAND U16547 ( .A(n16145), .B(n16144), .Z(n16146) );
  AND U16548 ( .A(n16147), .B(n16146), .Z(n16370) );
  NAND U16549 ( .A(n16149), .B(n16148), .Z(n16153) );
  NAND U16550 ( .A(n16151), .B(n16150), .Z(n16152) );
  AND U16551 ( .A(n16153), .B(n16152), .Z(n16261) );
  NAND U16552 ( .A(n16155), .B(n16154), .Z(n16159) );
  NAND U16553 ( .A(n16157), .B(n16156), .Z(n16158) );
  AND U16554 ( .A(n16159), .B(n16158), .Z(n16220) );
  AND U16555 ( .A(x[175]), .B(y[40]), .Z(n16161) );
  NAND U16556 ( .A(x[173]), .B(y[42]), .Z(n16160) );
  XNOR U16557 ( .A(n16161), .B(n16160), .Z(n16165) );
  AND U16558 ( .A(x[192]), .B(y[167]), .Z(n16163) );
  NAND U16559 ( .A(x[170]), .B(y[45]), .Z(n16162) );
  XNOR U16560 ( .A(n16163), .B(n16162), .Z(n16164) );
  XOR U16561 ( .A(n16165), .B(n16164), .Z(n16173) );
  AND U16562 ( .A(x[169]), .B(y[46]), .Z(n16167) );
  NAND U16563 ( .A(x[179]), .B(y[84]), .Z(n16166) );
  XNOR U16564 ( .A(n16167), .B(n16166), .Z(n16171) );
  AND U16565 ( .A(x[184]), .B(y[127]), .Z(n16169) );
  NAND U16566 ( .A(x[186]), .B(y[125]), .Z(n16168) );
  XNOR U16567 ( .A(n16169), .B(n16168), .Z(n16170) );
  XNOR U16568 ( .A(n16171), .B(n16170), .Z(n16172) );
  XNOR U16569 ( .A(n16173), .B(n16172), .Z(n16218) );
  AND U16570 ( .A(x[198]), .B(y[161]), .Z(n16178) );
  AND U16571 ( .A(y[2]), .B(x[165]), .Z(n16335) );
  AND U16572 ( .A(x[168]), .B(y[47]), .Z(n16175) );
  NAND U16573 ( .A(x[191]), .B(y[120]), .Z(n16174) );
  XNOR U16574 ( .A(n16175), .B(n16174), .Z(n16176) );
  XNOR U16575 ( .A(n16335), .B(n16176), .Z(n16177) );
  XNOR U16576 ( .A(n16178), .B(n16177), .Z(n16194) );
  AND U16577 ( .A(x[176]), .B(y[87]), .Z(n16180) );
  NAND U16578 ( .A(x[180]), .B(y[83]), .Z(n16179) );
  XNOR U16579 ( .A(n16180), .B(n16179), .Z(n16184) );
  AND U16580 ( .A(x[187]), .B(y[124]), .Z(n16182) );
  NAND U16581 ( .A(x[190]), .B(y[121]), .Z(n16181) );
  XNOR U16582 ( .A(n16182), .B(n16181), .Z(n16183) );
  XOR U16583 ( .A(n16184), .B(n16183), .Z(n16192) );
  AND U16584 ( .A(x[162]), .B(y[5]), .Z(n16186) );
  NAND U16585 ( .A(x[174]), .B(y[41]), .Z(n16185) );
  XNOR U16586 ( .A(n16186), .B(n16185), .Z(n16190) );
  AND U16587 ( .A(x[163]), .B(y[4]), .Z(n16188) );
  NAND U16588 ( .A(x[199]), .B(y[160]), .Z(n16187) );
  XNOR U16589 ( .A(n16188), .B(n16187), .Z(n16189) );
  XNOR U16590 ( .A(n16190), .B(n16189), .Z(n16191) );
  XNOR U16591 ( .A(n16192), .B(n16191), .Z(n16193) );
  XOR U16592 ( .A(n16194), .B(n16193), .Z(n16216) );
  AND U16593 ( .A(x[194]), .B(y[165]), .Z(n16196) );
  NAND U16594 ( .A(x[166]), .B(y[1]), .Z(n16195) );
  XNOR U16595 ( .A(n16196), .B(n16195), .Z(n16200) );
  AND U16596 ( .A(x[164]), .B(y[3]), .Z(n16198) );
  NAND U16597 ( .A(x[167]), .B(y[0]), .Z(n16197) );
  XNOR U16598 ( .A(n16198), .B(n16197), .Z(n16199) );
  XOR U16599 ( .A(n16200), .B(n16199), .Z(n16208) );
  AND U16600 ( .A(x[189]), .B(y[122]), .Z(n16202) );
  NAND U16601 ( .A(x[195]), .B(y[164]), .Z(n16201) );
  XNOR U16602 ( .A(n16202), .B(n16201), .Z(n16206) );
  AND U16603 ( .A(x[161]), .B(y[6]), .Z(n16204) );
  NAND U16604 ( .A(x[181]), .B(y[82]), .Z(n16203) );
  XNOR U16605 ( .A(n16204), .B(n16203), .Z(n16205) );
  XNOR U16606 ( .A(n16206), .B(n16205), .Z(n16207) );
  XNOR U16607 ( .A(n16208), .B(n16207), .Z(n16214) );
  AND U16608 ( .A(y[162]), .B(x[197]), .Z(n16305) );
  AND U16609 ( .A(y[126]), .B(x[185]), .Z(n16276) );
  XOR U16610 ( .A(n16305), .B(n16276), .Z(n16212) );
  XNOR U16611 ( .A(n16210), .B(n16209), .Z(n16211) );
  XNOR U16612 ( .A(n16212), .B(n16211), .Z(n16213) );
  XNOR U16613 ( .A(n16214), .B(n16213), .Z(n16215) );
  XNOR U16614 ( .A(n16216), .B(n16215), .Z(n16217) );
  XNOR U16615 ( .A(n16218), .B(n16217), .Z(n16219) );
  XNOR U16616 ( .A(n16220), .B(n16219), .Z(n16259) );
  NANDN U16617 ( .A(n16222), .B(n16221), .Z(n16226) );
  NANDN U16618 ( .A(n16224), .B(n16223), .Z(n16225) );
  AND U16619 ( .A(n16226), .B(n16225), .Z(n16257) );
  NAND U16620 ( .A(n16228), .B(n16227), .Z(n16231) );
  AND U16621 ( .A(y[42]), .B(x[171]), .Z(n16229) );
  AND U16622 ( .A(y[43]), .B(x[172]), .Z(n16307) );
  NAND U16623 ( .A(n16229), .B(n16307), .Z(n16230) );
  AND U16624 ( .A(n16231), .B(n16230), .Z(n16239) );
  NAND U16625 ( .A(n16233), .B(n16232), .Z(n16237) );
  NAND U16626 ( .A(n16235), .B(n16234), .Z(n16236) );
  NAND U16627 ( .A(n16237), .B(n16236), .Z(n16238) );
  XNOR U16628 ( .A(n16239), .B(n16238), .Z(n16255) );
  NAND U16629 ( .A(n16241), .B(n16240), .Z(n16245) );
  NAND U16630 ( .A(n16243), .B(n16242), .Z(n16244) );
  AND U16631 ( .A(n16245), .B(n16244), .Z(n16253) );
  NAND U16632 ( .A(n16247), .B(n16246), .Z(n16251) );
  NAND U16633 ( .A(n16249), .B(n16248), .Z(n16250) );
  NAND U16634 ( .A(n16251), .B(n16250), .Z(n16252) );
  XNOR U16635 ( .A(n16253), .B(n16252), .Z(n16254) );
  XNOR U16636 ( .A(n16255), .B(n16254), .Z(n16256) );
  XNOR U16637 ( .A(n16257), .B(n16256), .Z(n16258) );
  XNOR U16638 ( .A(n16259), .B(n16258), .Z(n16260) );
  XNOR U16639 ( .A(n16261), .B(n16260), .Z(n16368) );
  NAND U16640 ( .A(n16263), .B(n16262), .Z(n16267) );
  NAND U16641 ( .A(n16265), .B(n16264), .Z(n16266) );
  AND U16642 ( .A(n16267), .B(n16266), .Z(n16366) );
  NAND U16643 ( .A(n16269), .B(n16268), .Z(n16273) );
  NANDN U16644 ( .A(n16271), .B(n16270), .Z(n16272) );
  AND U16645 ( .A(n16273), .B(n16272), .Z(n16348) );
  NAND U16646 ( .A(n16275), .B(n16274), .Z(n16279) );
  NAND U16647 ( .A(n16277), .B(n16276), .Z(n16278) );
  AND U16648 ( .A(n16279), .B(n16278), .Z(n16287) );
  NAND U16649 ( .A(n16281), .B(n16280), .Z(n16285) );
  NAND U16650 ( .A(n16283), .B(n16282), .Z(n16284) );
  NAND U16651 ( .A(n16285), .B(n16284), .Z(n16286) );
  XNOR U16652 ( .A(n16287), .B(n16286), .Z(n16346) );
  AND U16653 ( .A(x[188]), .B(y[123]), .Z(n16289) );
  NAND U16654 ( .A(x[182]), .B(y[81]), .Z(n16288) );
  XNOR U16655 ( .A(n16289), .B(n16288), .Z(n16312) );
  AND U16656 ( .A(y[85]), .B(x[178]), .Z(n16304) );
  NAND U16657 ( .A(n16291), .B(n16290), .Z(n16294) );
  NAND U16658 ( .A(n16292), .B(n16304), .Z(n16293) );
  AND U16659 ( .A(n16294), .B(n16293), .Z(n16302) );
  AND U16660 ( .A(x[177]), .B(y[86]), .Z(n16296) );
  NAND U16661 ( .A(x[183]), .B(y[80]), .Z(n16295) );
  XNOR U16662 ( .A(n16296), .B(n16295), .Z(n16300) );
  AND U16663 ( .A(x[160]), .B(y[7]), .Z(n16298) );
  NAND U16664 ( .A(x[193]), .B(y[166]), .Z(n16297) );
  XNOR U16665 ( .A(n16298), .B(n16297), .Z(n16299) );
  XNOR U16666 ( .A(n16300), .B(n16299), .Z(n16301) );
  XNOR U16667 ( .A(n16302), .B(n16301), .Z(n16303) );
  XOR U16668 ( .A(n16304), .B(n16303), .Z(n16310) );
  AND U16669 ( .A(y[161]), .B(x[196]), .Z(n16306) );
  AND U16670 ( .A(n16306), .B(n16305), .Z(n16308) );
  XNOR U16671 ( .A(n16308), .B(n16307), .Z(n16309) );
  XNOR U16672 ( .A(n16310), .B(n16309), .Z(n16311) );
  XOR U16673 ( .A(n16312), .B(n16311), .Z(n16344) );
  NAND U16674 ( .A(n16314), .B(n16313), .Z(n16318) );
  NAND U16675 ( .A(n16316), .B(n16315), .Z(n16317) );
  AND U16676 ( .A(n16318), .B(n16317), .Z(n16326) );
  NAND U16677 ( .A(n16320), .B(n16319), .Z(n16324) );
  NAND U16678 ( .A(n16322), .B(n16321), .Z(n16323) );
  NAND U16679 ( .A(n16324), .B(n16323), .Z(n16325) );
  XNOR U16680 ( .A(n16326), .B(n16325), .Z(n16342) );
  NAND U16681 ( .A(n16328), .B(n16327), .Z(n16332) );
  NAND U16682 ( .A(n16330), .B(n16329), .Z(n16331) );
  AND U16683 ( .A(n16332), .B(n16331), .Z(n16340) );
  NAND U16684 ( .A(n16334), .B(n16333), .Z(n16338) );
  NAND U16685 ( .A(n16336), .B(n16335), .Z(n16337) );
  NAND U16686 ( .A(n16338), .B(n16337), .Z(n16339) );
  XNOR U16687 ( .A(n16340), .B(n16339), .Z(n16341) );
  XNOR U16688 ( .A(n16342), .B(n16341), .Z(n16343) );
  XNOR U16689 ( .A(n16344), .B(n16343), .Z(n16345) );
  XNOR U16690 ( .A(n16346), .B(n16345), .Z(n16347) );
  XNOR U16691 ( .A(n16348), .B(n16347), .Z(n16364) );
  NAND U16692 ( .A(n16350), .B(n16349), .Z(n16354) );
  NANDN U16693 ( .A(n16352), .B(n16351), .Z(n16353) );
  AND U16694 ( .A(n16354), .B(n16353), .Z(n16362) );
  NAND U16695 ( .A(n16356), .B(n16355), .Z(n16360) );
  NANDN U16696 ( .A(n16358), .B(n16357), .Z(n16359) );
  NAND U16697 ( .A(n16360), .B(n16359), .Z(n16361) );
  XNOR U16698 ( .A(n16362), .B(n16361), .Z(n16363) );
  XNOR U16699 ( .A(n16364), .B(n16363), .Z(n16365) );
  XNOR U16700 ( .A(n16366), .B(n16365), .Z(n16367) );
  XNOR U16701 ( .A(n16368), .B(n16367), .Z(n16369) );
  XNOR U16702 ( .A(n16370), .B(n16369), .Z(n16371) );
  XNOR U16703 ( .A(n16372), .B(n16371), .Z(n16373) );
  NAND U16704 ( .A(n16376), .B(n16375), .Z(n16380) );
  AND U16705 ( .A(n16378), .B(n16377), .Z(n16379) );
  ANDN U16706 ( .B(n16380), .A(n16379), .Z(n16388) );
  AND U16707 ( .A(n16382), .B(n16381), .Z(n16386) );
  ANDN U16708 ( .B(n16384), .A(n16383), .Z(n16385) );
  OR U16709 ( .A(n16386), .B(n16385), .Z(n16387) );
  XNOR U16710 ( .A(n16388), .B(n16387), .Z(n16389) );
  NAND U16711 ( .A(n16391), .B(n16390), .Z(n16395) );
  ANDN U16712 ( .B(n16393), .A(n16392), .Z(n16394) );
  AND U16713 ( .A(n16397), .B(n16396), .Z(n16401) );
  AND U16714 ( .A(n16399), .B(n16398), .Z(n16400) );
  NAND U16715 ( .A(y[168]), .B(x[192]), .Z(n16539) );
  NAND U16716 ( .A(y[48]), .B(x[168]), .Z(n16404) );
  XOR U16717 ( .A(n16539), .B(n16404), .Z(n16405) );
  AND U16718 ( .A(y[8]), .B(x[160]), .Z(n16412) );
  AND U16719 ( .A(y[88]), .B(x[176]), .Z(n16409) );
  XOR U16720 ( .A(n16412), .B(n16409), .Z(n16408) );
  AND U16721 ( .A(y[128]), .B(x[184]), .Z(n16407) );
  XNOR U16722 ( .A(n16408), .B(n16407), .Z(n16406) );
  XNOR U16723 ( .A(n16405), .B(n16406), .Z(o[168]) );
  AND U16724 ( .A(x[160]), .B(y[9]), .Z(n16403) );
  NAND U16725 ( .A(x[161]), .B(y[8]), .Z(n16402) );
  XNOR U16726 ( .A(n16403), .B(n16402), .Z(n16414) );
  AND U16727 ( .A(y[48]), .B(x[169]), .Z(n16413) );
  XOR U16728 ( .A(n16414), .B(n16413), .Z(n16431) );
  AND U16729 ( .A(y[168]), .B(x[193]), .Z(n16632) );
  AND U16730 ( .A(y[89]), .B(x[176]), .Z(n16417) );
  XOR U16731 ( .A(n16632), .B(n16417), .Z(n16419) );
  AND U16732 ( .A(y[169]), .B(x[192]), .Z(n16441) );
  NAND U16733 ( .A(y[88]), .B(x[177]), .Z(n16440) );
  XNOR U16734 ( .A(n16441), .B(n16440), .Z(n16418) );
  XOR U16735 ( .A(n16419), .B(n16418), .Z(n16429) );
  AND U16736 ( .A(y[49]), .B(x[168]), .Z(n16657) );
  AND U16737 ( .A(y[129]), .B(x[184]), .Z(n16434) );
  XOR U16738 ( .A(n16657), .B(n16434), .Z(n16436) );
  AND U16739 ( .A(y[128]), .B(x[185]), .Z(n16435) );
  XNOR U16740 ( .A(n16436), .B(n16435), .Z(n16428) );
  XNOR U16741 ( .A(n16429), .B(n16428), .Z(n16430) );
  XNOR U16742 ( .A(n16431), .B(n16430), .Z(n16425) );
  NAND U16743 ( .A(n16408), .B(n16407), .Z(n16411) );
  AND U16744 ( .A(n16412), .B(n16409), .Z(n16410) );
  ANDN U16745 ( .B(n16411), .A(n16410), .Z(n16422) );
  XNOR U16746 ( .A(n16423), .B(n16422), .Z(n16424) );
  XNOR U16747 ( .A(n16425), .B(n16424), .Z(o[169]) );
  NAND U16748 ( .A(y[9]), .B(x[161]), .Z(n16463) );
  NANDN U16749 ( .A(n16463), .B(n16412), .Z(n16416) );
  NAND U16750 ( .A(n16414), .B(n16413), .Z(n16415) );
  AND U16751 ( .A(n16416), .B(n16415), .Z(n16497) );
  NAND U16752 ( .A(n16632), .B(n16417), .Z(n16421) );
  NAND U16753 ( .A(n16419), .B(n16418), .Z(n16420) );
  AND U16754 ( .A(n16421), .B(n16420), .Z(n16496) );
  AND U16755 ( .A(y[130]), .B(x[184]), .Z(n16481) );
  NAND U16756 ( .A(y[10]), .B(x[160]), .Z(n16482) );
  XNOR U16757 ( .A(n16481), .B(n16482), .Z(n16483) );
  NAND U16758 ( .A(y[48]), .B(x[170]), .Z(n16484) );
  XNOR U16759 ( .A(n16483), .B(n16484), .Z(n16495) );
  XOR U16760 ( .A(n16496), .B(n16495), .Z(n16498) );
  XOR U16761 ( .A(n16497), .B(n16498), .Z(n16443) );
  NANDN U16762 ( .A(n16423), .B(n16422), .Z(n16427) );
  NAND U16763 ( .A(n16425), .B(n16424), .Z(n16426) );
  NAND U16764 ( .A(n16427), .B(n16426), .Z(n16442) );
  XNOR U16765 ( .A(n16443), .B(n16442), .Z(n16445) );
  NANDN U16766 ( .A(n16429), .B(n16428), .Z(n16433) );
  NANDN U16767 ( .A(n16431), .B(n16430), .Z(n16432) );
  AND U16768 ( .A(n16433), .B(n16432), .Z(n16451) );
  AND U16769 ( .A(y[8]), .B(x[162]), .Z(n16460) );
  NAND U16770 ( .A(y[90]), .B(x[176]), .Z(n16461) );
  XNOR U16771 ( .A(n16460), .B(n16461), .Z(n16462) );
  AND U16772 ( .A(y[128]), .B(x[186]), .Z(n16489) );
  XOR U16773 ( .A(n16490), .B(n16489), .Z(n16492) );
  AND U16774 ( .A(y[88]), .B(x[178]), .Z(n16576) );
  AND U16775 ( .A(y[170]), .B(x[192]), .Z(n16473) );
  XOR U16776 ( .A(n16576), .B(n16473), .Z(n16475) );
  AND U16777 ( .A(y[89]), .B(x[177]), .Z(n16474) );
  XOR U16778 ( .A(n16475), .B(n16474), .Z(n16491) );
  XOR U16779 ( .A(n16492), .B(n16491), .Z(n16448) );
  NAND U16780 ( .A(n16657), .B(n16434), .Z(n16438) );
  AND U16781 ( .A(n16436), .B(n16435), .Z(n16437) );
  ANDN U16782 ( .B(n16438), .A(n16437), .Z(n16457) );
  AND U16783 ( .A(x[193]), .B(y[169]), .Z(n16544) );
  NAND U16784 ( .A(x[194]), .B(y[168]), .Z(n16439) );
  XNOR U16785 ( .A(n16544), .B(n16439), .Z(n16488) );
  ANDN U16786 ( .B(n16441), .A(n16440), .Z(n16487) );
  XOR U16787 ( .A(n16488), .B(n16487), .Z(n16454) );
  AND U16788 ( .A(y[129]), .B(x[185]), .Z(n16466) );
  NAND U16789 ( .A(y[49]), .B(x[169]), .Z(n16467) );
  XNOR U16790 ( .A(n16466), .B(n16467), .Z(n16468) );
  NAND U16791 ( .A(y[50]), .B(x[168]), .Z(n16469) );
  XOR U16792 ( .A(n16468), .B(n16469), .Z(n16455) );
  XNOR U16793 ( .A(n16454), .B(n16455), .Z(n16456) );
  XOR U16794 ( .A(n16457), .B(n16456), .Z(n16449) );
  XNOR U16795 ( .A(n16448), .B(n16449), .Z(n16450) );
  XNOR U16796 ( .A(n16451), .B(n16450), .Z(n16444) );
  XNOR U16797 ( .A(n16445), .B(n16444), .Z(o[170]) );
  NANDN U16798 ( .A(n16443), .B(n16442), .Z(n16447) );
  NAND U16799 ( .A(n16445), .B(n16444), .Z(n16446) );
  AND U16800 ( .A(n16447), .B(n16446), .Z(n16519) );
  NANDN U16801 ( .A(n16449), .B(n16448), .Z(n16453) );
  NAND U16802 ( .A(n16451), .B(n16450), .Z(n16452) );
  AND U16803 ( .A(n16453), .B(n16452), .Z(n16504) );
  NANDN U16804 ( .A(n16455), .B(n16454), .Z(n16459) );
  NANDN U16805 ( .A(n16457), .B(n16456), .Z(n16458) );
  AND U16806 ( .A(n16459), .B(n16458), .Z(n16502) );
  NANDN U16807 ( .A(n16461), .B(n16460), .Z(n16465) );
  NANDN U16808 ( .A(n16463), .B(n16462), .Z(n16464) );
  NAND U16809 ( .A(n16465), .B(n16464), .Z(n16513) );
  NANDN U16810 ( .A(n16467), .B(n16466), .Z(n16471) );
  NANDN U16811 ( .A(n16469), .B(n16468), .Z(n16470) );
  AND U16812 ( .A(n16471), .B(n16470), .Z(n16558) );
  AND U16813 ( .A(y[131]), .B(x[184]), .Z(n16572) );
  AND U16814 ( .A(y[91]), .B(x[176]), .Z(n16571) );
  NAND U16815 ( .A(y[8]), .B(x[163]), .Z(n16570) );
  XOR U16816 ( .A(n16571), .B(n16570), .Z(n16573) );
  XOR U16817 ( .A(n16572), .B(n16573), .Z(n16556) );
  AND U16818 ( .A(x[178]), .B(y[89]), .Z(n16615) );
  NAND U16819 ( .A(x[179]), .B(y[88]), .Z(n16472) );
  XNOR U16820 ( .A(n16615), .B(n16472), .Z(n16577) );
  NAND U16821 ( .A(y[90]), .B(x[177]), .Z(n16578) );
  XNOR U16822 ( .A(n16556), .B(n16555), .Z(n16557) );
  XNOR U16823 ( .A(n16558), .B(n16557), .Z(n16514) );
  XOR U16824 ( .A(n16513), .B(n16514), .Z(n16516) );
  NAND U16825 ( .A(n16576), .B(n16473), .Z(n16477) );
  AND U16826 ( .A(n16475), .B(n16474), .Z(n16476) );
  ANDN U16827 ( .B(n16477), .A(n16476), .Z(n16563) );
  AND U16828 ( .A(y[10]), .B(x[161]), .Z(n16535) );
  AND U16829 ( .A(y[9]), .B(x[162]), .Z(n16534) );
  NAND U16830 ( .A(y[130]), .B(x[185]), .Z(n16533) );
  XOR U16831 ( .A(n16534), .B(n16533), .Z(n16536) );
  XOR U16832 ( .A(n16535), .B(n16536), .Z(n16562) );
  AND U16833 ( .A(x[195]), .B(y[168]), .Z(n16479) );
  NAND U16834 ( .A(x[192]), .B(y[171]), .Z(n16478) );
  XNOR U16835 ( .A(n16479), .B(n16478), .Z(n16540) );
  AND U16836 ( .A(x[194]), .B(y[169]), .Z(n16628) );
  NAND U16837 ( .A(x[193]), .B(y[170]), .Z(n16480) );
  XOR U16838 ( .A(n16628), .B(n16480), .Z(n16541) );
  XNOR U16839 ( .A(n16540), .B(n16541), .Z(n16561) );
  XOR U16840 ( .A(n16562), .B(n16561), .Z(n16564) );
  XOR U16841 ( .A(n16563), .B(n16564), .Z(n16515) );
  XOR U16842 ( .A(n16516), .B(n16515), .Z(n16501) );
  XNOR U16843 ( .A(n16502), .B(n16501), .Z(n16503) );
  XOR U16844 ( .A(n16504), .B(n16503), .Z(n16520) );
  XNOR U16845 ( .A(n16519), .B(n16520), .Z(n16522) );
  NANDN U16846 ( .A(n16482), .B(n16481), .Z(n16486) );
  NANDN U16847 ( .A(n16484), .B(n16483), .Z(n16485) );
  AND U16848 ( .A(n16486), .B(n16485), .Z(n16526) );
  XNOR U16849 ( .A(n16526), .B(n16525), .Z(n16528) );
  NAND U16850 ( .A(y[48]), .B(x[171]), .Z(n16585) );
  NAND U16851 ( .A(y[11]), .B(x[160]), .Z(n16583) );
  NAND U16852 ( .A(y[129]), .B(x[186]), .Z(n16584) );
  XNOR U16853 ( .A(n16583), .B(n16584), .Z(n16586) );
  XOR U16854 ( .A(n16585), .B(n16586), .Z(n16551) );
  NAND U16855 ( .A(y[51]), .B(x[168]), .Z(n16547) );
  NAND U16856 ( .A(y[49]), .B(x[170]), .Z(n16545) );
  NAND U16857 ( .A(y[128]), .B(x[187]), .Z(n16546) );
  XNOR U16858 ( .A(n16545), .B(n16546), .Z(n16548) );
  XOR U16859 ( .A(n16547), .B(n16548), .Z(n16549) );
  AND U16860 ( .A(y[50]), .B(x[169]), .Z(n16550) );
  XOR U16861 ( .A(n16549), .B(n16550), .Z(n16552) );
  XOR U16862 ( .A(n16551), .B(n16552), .Z(n16527) );
  XOR U16863 ( .A(n16528), .B(n16527), .Z(n16508) );
  NAND U16864 ( .A(n16490), .B(n16489), .Z(n16494) );
  NAND U16865 ( .A(n16492), .B(n16491), .Z(n16493) );
  AND U16866 ( .A(n16494), .B(n16493), .Z(n16507) );
  XNOR U16867 ( .A(n16508), .B(n16507), .Z(n16510) );
  NANDN U16868 ( .A(n16496), .B(n16495), .Z(n16500) );
  OR U16869 ( .A(n16498), .B(n16497), .Z(n16499) );
  AND U16870 ( .A(n16500), .B(n16499), .Z(n16509) );
  XNOR U16871 ( .A(n16510), .B(n16509), .Z(n16521) );
  XOR U16872 ( .A(n16522), .B(n16521), .Z(o[171]) );
  NANDN U16873 ( .A(n16502), .B(n16501), .Z(n16506) );
  NANDN U16874 ( .A(n16504), .B(n16503), .Z(n16505) );
  AND U16875 ( .A(n16506), .B(n16505), .Z(n16595) );
  NANDN U16876 ( .A(n16508), .B(n16507), .Z(n16512) );
  NAND U16877 ( .A(n16510), .B(n16509), .Z(n16511) );
  NAND U16878 ( .A(n16512), .B(n16511), .Z(n16593) );
  NAND U16879 ( .A(n16514), .B(n16513), .Z(n16518) );
  NAND U16880 ( .A(n16516), .B(n16515), .Z(n16517) );
  AND U16881 ( .A(n16518), .B(n16517), .Z(n16594) );
  XOR U16882 ( .A(n16593), .B(n16594), .Z(n16596) );
  XOR U16883 ( .A(n16595), .B(n16596), .Z(n16587) );
  NANDN U16884 ( .A(n16520), .B(n16519), .Z(n16524) );
  NAND U16885 ( .A(n16522), .B(n16521), .Z(n16523) );
  NAND U16886 ( .A(n16524), .B(n16523), .Z(n16588) );
  XNOR U16887 ( .A(n16587), .B(n16588), .Z(n16590) );
  NANDN U16888 ( .A(n16526), .B(n16525), .Z(n16530) );
  NAND U16889 ( .A(n16528), .B(n16527), .Z(n16529) );
  AND U16890 ( .A(n16530), .B(n16529), .Z(n16600) );
  AND U16891 ( .A(x[171]), .B(y[49]), .Z(n16532) );
  NAND U16892 ( .A(x[168]), .B(y[52]), .Z(n16531) );
  XNOR U16893 ( .A(n16532), .B(n16531), .Z(n16659) );
  AND U16894 ( .A(y[50]), .B(x[170]), .Z(n16658) );
  XOR U16895 ( .A(n16659), .B(n16658), .Z(n16667) );
  AND U16896 ( .A(y[51]), .B(x[169]), .Z(n16666) );
  XOR U16897 ( .A(n16667), .B(n16666), .Z(n16669) );
  AND U16898 ( .A(y[128]), .B(x[188]), .Z(n16621) );
  AND U16899 ( .A(y[11]), .B(x[161]), .Z(n16620) );
  XOR U16900 ( .A(n16621), .B(n16620), .Z(n16623) );
  AND U16901 ( .A(y[12]), .B(x[160]), .Z(n16622) );
  XOR U16902 ( .A(n16623), .B(n16622), .Z(n16668) );
  XOR U16903 ( .A(n16669), .B(n16668), .Z(n16665) );
  NANDN U16904 ( .A(n16534), .B(n16533), .Z(n16538) );
  OR U16905 ( .A(n16536), .B(n16535), .Z(n16537) );
  NAND U16906 ( .A(n16538), .B(n16537), .Z(n16662) );
  AND U16907 ( .A(y[171]), .B(x[195]), .Z(n16903) );
  NANDN U16908 ( .A(n16539), .B(n16903), .Z(n16543) );
  NANDN U16909 ( .A(n16541), .B(n16540), .Z(n16542) );
  AND U16910 ( .A(n16543), .B(n16542), .Z(n16663) );
  XOR U16911 ( .A(n16662), .B(n16663), .Z(n16664) );
  XNOR U16912 ( .A(n16665), .B(n16664), .Z(n16689) );
  AND U16913 ( .A(y[8]), .B(x[164]), .Z(n16642) );
  AND U16914 ( .A(y[130]), .B(x[186]), .Z(n16640) );
  NAND U16915 ( .A(y[92]), .B(x[176]), .Z(n16639) );
  XNOR U16916 ( .A(n16640), .B(n16639), .Z(n16641) );
  XNOR U16917 ( .A(n16642), .B(n16641), .Z(n16606) );
  AND U16918 ( .A(x[194]), .B(y[170]), .Z(n16569) );
  NAND U16919 ( .A(n16569), .B(n16544), .Z(n16637) );
  NAND U16920 ( .A(y[88]), .B(x[180]), .Z(n16748) );
  NAND U16921 ( .A(y[172]), .B(x[192]), .Z(n16782) );
  XNOR U16922 ( .A(n16748), .B(n16782), .Z(n16638) );
  XOR U16923 ( .A(n16637), .B(n16638), .Z(n16605) );
  XNOR U16924 ( .A(n16606), .B(n16605), .Z(n16608) );
  XOR U16925 ( .A(n16608), .B(n16607), .Z(n16687) );
  NAND U16926 ( .A(n16550), .B(n16549), .Z(n16554) );
  NAND U16927 ( .A(n16552), .B(n16551), .Z(n16553) );
  AND U16928 ( .A(n16554), .B(n16553), .Z(n16686) );
  XNOR U16929 ( .A(n16689), .B(n16688), .Z(n16599) );
  XNOR U16930 ( .A(n16600), .B(n16599), .Z(n16602) );
  NANDN U16931 ( .A(n16556), .B(n16555), .Z(n16560) );
  NANDN U16932 ( .A(n16558), .B(n16557), .Z(n16559) );
  AND U16933 ( .A(n16560), .B(n16559), .Z(n16675) );
  NANDN U16934 ( .A(n16562), .B(n16561), .Z(n16566) );
  OR U16935 ( .A(n16564), .B(n16563), .Z(n16565) );
  NAND U16936 ( .A(n16566), .B(n16565), .Z(n16674) );
  NAND U16937 ( .A(y[10]), .B(x[162]), .Z(n16653) );
  NAND U16938 ( .A(y[129]), .B(x[187]), .Z(n16652) );
  NAND U16939 ( .A(y[9]), .B(x[163]), .Z(n16651) );
  XOR U16940 ( .A(n16652), .B(n16651), .Z(n16654) );
  XOR U16941 ( .A(n16653), .B(n16654), .Z(n16614) );
  AND U16942 ( .A(x[196]), .B(y[168]), .Z(n16568) );
  NAND U16943 ( .A(x[193]), .B(y[171]), .Z(n16567) );
  XNOR U16944 ( .A(n16568), .B(n16567), .Z(n16633) );
  AND U16945 ( .A(y[169]), .B(x[195]), .Z(n16753) );
  XNOR U16946 ( .A(n16753), .B(n16569), .Z(n16634) );
  XNOR U16947 ( .A(n16633), .B(n16634), .Z(n16612) );
  NANDN U16948 ( .A(n16571), .B(n16570), .Z(n16575) );
  OR U16949 ( .A(n16573), .B(n16572), .Z(n16574) );
  AND U16950 ( .A(n16575), .B(n16574), .Z(n16611) );
  XOR U16951 ( .A(n16612), .B(n16611), .Z(n16613) );
  XNOR U16952 ( .A(n16614), .B(n16613), .Z(n16683) );
  AND U16953 ( .A(y[89]), .B(x[179]), .Z(n16582) );
  NAND U16954 ( .A(n16576), .B(n16582), .Z(n16580) );
  NANDN U16955 ( .A(n16578), .B(n16577), .Z(n16579) );
  AND U16956 ( .A(n16580), .B(n16579), .Z(n16681) );
  AND U16957 ( .A(y[48]), .B(x[172]), .Z(n16625) );
  AND U16958 ( .A(y[132]), .B(x[184]), .Z(n16624) );
  XOR U16959 ( .A(n16625), .B(n16624), .Z(n16627) );
  AND U16960 ( .A(y[131]), .B(x[185]), .Z(n16626) );
  XOR U16961 ( .A(n16627), .B(n16626), .Z(n16671) );
  NAND U16962 ( .A(x[178]), .B(y[90]), .Z(n16581) );
  XNOR U16963 ( .A(n16582), .B(n16581), .Z(n16617) );
  AND U16964 ( .A(y[91]), .B(x[177]), .Z(n16616) );
  XOR U16965 ( .A(n16617), .B(n16616), .Z(n16670) );
  XOR U16966 ( .A(n16671), .B(n16670), .Z(n16673) );
  XOR U16967 ( .A(n16673), .B(n16672), .Z(n16680) );
  XOR U16968 ( .A(n16683), .B(n16682), .Z(n16676) );
  XOR U16969 ( .A(n16677), .B(n16676), .Z(n16601) );
  XNOR U16970 ( .A(n16602), .B(n16601), .Z(n16589) );
  XNOR U16971 ( .A(n16590), .B(n16589), .Z(o[172]) );
  NANDN U16972 ( .A(n16588), .B(n16587), .Z(n16592) );
  NAND U16973 ( .A(n16590), .B(n16589), .Z(n16591) );
  AND U16974 ( .A(n16592), .B(n16591), .Z(n16826) );
  NAND U16975 ( .A(n16594), .B(n16593), .Z(n16598) );
  NAND U16976 ( .A(n16596), .B(n16595), .Z(n16597) );
  NAND U16977 ( .A(n16598), .B(n16597), .Z(n16827) );
  XNOR U16978 ( .A(n16826), .B(n16827), .Z(n16829) );
  NANDN U16979 ( .A(n16600), .B(n16599), .Z(n16604) );
  NAND U16980 ( .A(n16602), .B(n16601), .Z(n16603) );
  AND U16981 ( .A(n16604), .B(n16603), .Z(n16693) );
  NANDN U16982 ( .A(n16606), .B(n16605), .Z(n16610) );
  NAND U16983 ( .A(n16608), .B(n16607), .Z(n16609) );
  NAND U16984 ( .A(n16610), .B(n16609), .Z(n16696) );
  XOR U16985 ( .A(n16696), .B(n16697), .Z(n16700) );
  AND U16986 ( .A(y[90]), .B(x[179]), .Z(n16750) );
  NAND U16987 ( .A(n16615), .B(n16750), .Z(n16619) );
  NAND U16988 ( .A(n16617), .B(n16616), .Z(n16618) );
  NAND U16989 ( .A(n16619), .B(n16618), .Z(n16755) );
  AND U16990 ( .A(y[48]), .B(x[173]), .Z(n16739) );
  AND U16991 ( .A(y[91]), .B(x[178]), .Z(n16738) );
  XOR U16992 ( .A(n16739), .B(n16738), .Z(n16740) );
  AND U16993 ( .A(y[133]), .B(x[184]), .Z(n16884) );
  XOR U16994 ( .A(n16740), .B(n16884), .Z(n16716) );
  AND U16995 ( .A(y[129]), .B(x[188]), .Z(n16744) );
  AND U16996 ( .A(y[8]), .B(x[165]), .Z(n16743) );
  XOR U16997 ( .A(n16744), .B(n16743), .Z(n16745) );
  AND U16998 ( .A(y[9]), .B(x[164]), .Z(n16854) );
  XNOR U16999 ( .A(n16745), .B(n16854), .Z(n16717) );
  XNOR U17000 ( .A(n16716), .B(n16717), .Z(n16718) );
  XNOR U17001 ( .A(n16719), .B(n16718), .Z(n16756) );
  XOR U17002 ( .A(n16755), .B(n16756), .Z(n16758) );
  AND U17003 ( .A(y[170]), .B(x[195]), .Z(n16629) );
  AND U17004 ( .A(n16629), .B(n16628), .Z(n16784) );
  AND U17005 ( .A(x[192]), .B(y[173]), .Z(n16631) );
  AND U17006 ( .A(x[193]), .B(y[172]), .Z(n16630) );
  XOR U17007 ( .A(n16631), .B(n16630), .Z(n16783) );
  XOR U17008 ( .A(n16784), .B(n16783), .Z(n16796) );
  AND U17009 ( .A(y[53]), .B(x[168]), .Z(n16804) );
  AND U17010 ( .A(y[12]), .B(x[161]), .Z(n16803) );
  XOR U17011 ( .A(n16804), .B(n16803), .Z(n16806) );
  AND U17012 ( .A(y[49]), .B(x[172]), .Z(n16805) );
  XOR U17013 ( .A(n16806), .B(n16805), .Z(n16795) );
  XOR U17014 ( .A(n16796), .B(n16795), .Z(n16798) );
  XOR U17015 ( .A(n16797), .B(n16798), .Z(n16757) );
  XOR U17016 ( .A(n16758), .B(n16757), .Z(n16699) );
  XOR U17017 ( .A(n16700), .B(n16699), .Z(n16823) );
  AND U17018 ( .A(y[171]), .B(x[196]), .Z(n16963) );
  NAND U17019 ( .A(n16963), .B(n16632), .Z(n16636) );
  NANDN U17020 ( .A(n16634), .B(n16633), .Z(n16635) );
  NAND U17021 ( .A(n16636), .B(n16635), .Z(n16712) );
  XOR U17022 ( .A(n16712), .B(n16713), .Z(n16715) );
  NANDN U17023 ( .A(n16640), .B(n16639), .Z(n16644) );
  NANDN U17024 ( .A(n16642), .B(n16641), .Z(n16643) );
  AND U17025 ( .A(n16644), .B(n16643), .Z(n16707) );
  AND U17026 ( .A(x[170]), .B(y[51]), .Z(n16646) );
  NAND U17027 ( .A(x[171]), .B(y[50]), .Z(n16645) );
  XNOR U17028 ( .A(n16646), .B(n16645), .Z(n16734) );
  AND U17029 ( .A(y[52]), .B(x[169]), .Z(n16733) );
  XOR U17030 ( .A(n16734), .B(n16733), .Z(n16705) );
  AND U17031 ( .A(y[171]), .B(x[194]), .Z(n16723) );
  AND U17032 ( .A(y[168]), .B(x[197]), .Z(n16722) );
  XOR U17033 ( .A(n16723), .B(n16722), .Z(n16725) );
  AND U17034 ( .A(x[196]), .B(y[169]), .Z(n16648) );
  NAND U17035 ( .A(x[195]), .B(y[170]), .Z(n16647) );
  XNOR U17036 ( .A(n16648), .B(n16647), .Z(n16724) );
  XOR U17037 ( .A(n16725), .B(n16724), .Z(n16704) );
  XOR U17038 ( .A(n16705), .B(n16704), .Z(n16706) );
  XOR U17039 ( .A(n16707), .B(n16706), .Z(n16714) );
  XOR U17040 ( .A(n16715), .B(n16714), .Z(n16768) );
  AND U17041 ( .A(y[89]), .B(x[180]), .Z(n16650) );
  AND U17042 ( .A(x[181]), .B(y[88]), .Z(n16649) );
  XOR U17043 ( .A(n16650), .B(n16649), .Z(n16749) );
  XOR U17044 ( .A(n16750), .B(n16749), .Z(n16772) );
  AND U17045 ( .A(y[128]), .B(x[189]), .Z(n16729) );
  AND U17046 ( .A(y[10]), .B(x[163]), .Z(n16728) );
  XOR U17047 ( .A(n16729), .B(n16728), .Z(n16731) );
  AND U17048 ( .A(y[11]), .B(x[162]), .Z(n16730) );
  XOR U17049 ( .A(n16731), .B(n16730), .Z(n16771) );
  XOR U17050 ( .A(n16772), .B(n16771), .Z(n16774) );
  NAND U17051 ( .A(n16652), .B(n16651), .Z(n16656) );
  NAND U17052 ( .A(n16654), .B(n16653), .Z(n16655) );
  AND U17053 ( .A(n16656), .B(n16655), .Z(n16773) );
  XOR U17054 ( .A(n16774), .B(n16773), .Z(n16766) );
  AND U17055 ( .A(y[52]), .B(x[171]), .Z(n16962) );
  NAND U17056 ( .A(n16962), .B(n16657), .Z(n16661) );
  IV U17057 ( .A(n16658), .Z(n16732) );
  NANDN U17058 ( .A(n16732), .B(n16659), .Z(n16660) );
  NAND U17059 ( .A(n16661), .B(n16660), .Z(n16710) );
  AND U17060 ( .A(y[130]), .B(x[187]), .Z(n16777) );
  AND U17061 ( .A(y[92]), .B(x[177]), .Z(n16867) );
  XOR U17062 ( .A(n16777), .B(n16867), .Z(n16779) );
  AND U17063 ( .A(y[93]), .B(x[176]), .Z(n16778) );
  XOR U17064 ( .A(n16779), .B(n16778), .Z(n16709) );
  AND U17065 ( .A(y[13]), .B(x[160]), .Z(n16788) );
  AND U17066 ( .A(y[132]), .B(x[185]), .Z(n16787) );
  XOR U17067 ( .A(n16788), .B(n16787), .Z(n16790) );
  AND U17068 ( .A(y[131]), .B(x[186]), .Z(n16789) );
  XOR U17069 ( .A(n16790), .B(n16789), .Z(n16708) );
  XOR U17070 ( .A(n16709), .B(n16708), .Z(n16711) );
  XOR U17071 ( .A(n16710), .B(n16711), .Z(n16765) );
  XOR U17072 ( .A(n16766), .B(n16765), .Z(n16767) );
  XOR U17073 ( .A(n16768), .B(n16767), .Z(n16820) );
  XNOR U17074 ( .A(n16761), .B(n16762), .Z(n16764) );
  XNOR U17075 ( .A(n16763), .B(n16764), .Z(n16821) );
  XOR U17076 ( .A(n16820), .B(n16821), .Z(n16822) );
  XOR U17077 ( .A(n16823), .B(n16822), .Z(n16692) );
  XNOR U17078 ( .A(n16693), .B(n16692), .Z(n16695) );
  NANDN U17079 ( .A(n16675), .B(n16674), .Z(n16679) );
  NAND U17080 ( .A(n16677), .B(n16676), .Z(n16678) );
  AND U17081 ( .A(n16679), .B(n16678), .Z(n16817) );
  NANDN U17082 ( .A(n16681), .B(n16680), .Z(n16685) );
  NAND U17083 ( .A(n16683), .B(n16682), .Z(n16684) );
  AND U17084 ( .A(n16685), .B(n16684), .Z(n16815) );
  NANDN U17085 ( .A(n16687), .B(n16686), .Z(n16691) );
  NAND U17086 ( .A(n16689), .B(n16688), .Z(n16690) );
  AND U17087 ( .A(n16691), .B(n16690), .Z(n16814) );
  XOR U17088 ( .A(n16695), .B(n16694), .Z(n16828) );
  XOR U17089 ( .A(n16829), .B(n16828), .Z(o[173]) );
  IV U17090 ( .A(n16696), .Z(n16698) );
  NANDN U17091 ( .A(n16698), .B(n16697), .Z(n16703) );
  IV U17092 ( .A(n16699), .Z(n16701) );
  NANDN U17093 ( .A(n16701), .B(n16700), .Z(n16702) );
  NAND U17094 ( .A(n16703), .B(n16702), .Z(n16832) );
  XOR U17095 ( .A(n16839), .B(n16838), .Z(n16836) );
  XOR U17096 ( .A(n16837), .B(n16836), .Z(n16835) );
  IV U17097 ( .A(n16835), .Z(n16754) );
  NANDN U17098 ( .A(n16717), .B(n16716), .Z(n16721) );
  NANDN U17099 ( .A(n16719), .B(n16718), .Z(n16720) );
  NAND U17100 ( .A(n16721), .B(n16720), .Z(n16842) );
  NAND U17101 ( .A(n16723), .B(n16722), .Z(n16727) );
  NAND U17102 ( .A(n16725), .B(n16724), .Z(n16726) );
  NAND U17103 ( .A(n16727), .B(n16726), .Z(n17041) );
  AND U17104 ( .A(x[171]), .B(y[51]), .Z(n16802) );
  NANDN U17105 ( .A(n16732), .B(n16802), .Z(n16736) );
  NAND U17106 ( .A(n16734), .B(n16733), .Z(n16735) );
  AND U17107 ( .A(n16736), .B(n16735), .Z(n16847) );
  AND U17108 ( .A(y[131]), .B(x[187]), .Z(n16860) );
  AND U17109 ( .A(y[91]), .B(x[179]), .Z(n16859) );
  XOR U17110 ( .A(n16860), .B(n16859), .Z(n16858) );
  AND U17111 ( .A(y[11]), .B(x[163]), .Z(n16857) );
  XOR U17112 ( .A(n16858), .B(n16857), .Z(n16849) );
  IV U17113 ( .A(n16849), .Z(n16737) );
  AND U17114 ( .A(y[132]), .B(x[186]), .Z(n16881) );
  AND U17115 ( .A(y[90]), .B(x[180]), .Z(n16880) );
  XOR U17116 ( .A(n16881), .B(n16880), .Z(n16879) );
  AND U17117 ( .A(y[12]), .B(x[162]), .Z(n16878) );
  XNOR U17118 ( .A(n16879), .B(n16878), .Z(n16848) );
  XOR U17119 ( .A(n16737), .B(n16848), .Z(n16846) );
  XNOR U17120 ( .A(n16847), .B(n16846), .Z(n17043) );
  XOR U17121 ( .A(n17044), .B(n17043), .Z(n17042) );
  XOR U17122 ( .A(n17041), .B(n17042), .Z(n16843) );
  XOR U17123 ( .A(n16842), .B(n16843), .Z(n16841) );
  NAND U17124 ( .A(n16739), .B(n16738), .Z(n16742) );
  NAND U17125 ( .A(n16740), .B(n16884), .Z(n16741) );
  NAND U17126 ( .A(n16742), .B(n16741), .Z(n17002) );
  NAND U17127 ( .A(n16744), .B(n16743), .Z(n16747) );
  NAND U17128 ( .A(n16745), .B(n16854), .Z(n16746) );
  NAND U17129 ( .A(n16747), .B(n16746), .Z(n17001) );
  XOR U17130 ( .A(n17002), .B(n17001), .Z(n17000) );
  AND U17131 ( .A(y[89]), .B(x[181]), .Z(n16871) );
  AND U17132 ( .A(x[165]), .B(y[9]), .Z(n16752) );
  NAND U17133 ( .A(x[164]), .B(y[10]), .Z(n16751) );
  XNOR U17134 ( .A(n16752), .B(n16751), .Z(n16853) );
  AND U17135 ( .A(y[128]), .B(x[190]), .Z(n16852) );
  XOR U17136 ( .A(n16853), .B(n16852), .Z(n17030) );
  AND U17137 ( .A(y[173]), .B(x[193]), .Z(n16909) );
  AND U17138 ( .A(y[170]), .B(x[196]), .Z(n16794) );
  AND U17139 ( .A(n16753), .B(n16794), .Z(n16907) );
  AND U17140 ( .A(y[172]), .B(x[194]), .Z(n16906) );
  XOR U17141 ( .A(n16907), .B(n16906), .Z(n16908) );
  XNOR U17142 ( .A(n16909), .B(n16908), .Z(n17029) );
  XNOR U17143 ( .A(n17028), .B(n17027), .Z(n16999) );
  XOR U17144 ( .A(n17000), .B(n16999), .Z(n16840) );
  XOR U17145 ( .A(n16841), .B(n16840), .Z(n16834) );
  XOR U17146 ( .A(n16754), .B(n16834), .Z(n16833) );
  XOR U17147 ( .A(n16832), .B(n16833), .Z(n17080) );
  NAND U17148 ( .A(n16756), .B(n16755), .Z(n16760) );
  NAND U17149 ( .A(n16758), .B(n16757), .Z(n16759) );
  AND U17150 ( .A(n16760), .B(n16759), .Z(n17079) );
  OR U17151 ( .A(n16766), .B(n16765), .Z(n16770) );
  NANDN U17152 ( .A(n16768), .B(n16767), .Z(n16769) );
  NAND U17153 ( .A(n16770), .B(n16769), .Z(n17059) );
  NAND U17154 ( .A(n16772), .B(n16771), .Z(n16776) );
  NAND U17155 ( .A(n16774), .B(n16773), .Z(n16775) );
  AND U17156 ( .A(n16776), .B(n16775), .Z(n17064) );
  NAND U17157 ( .A(n16777), .B(n16867), .Z(n16781) );
  NAND U17158 ( .A(n16779), .B(n16778), .Z(n16780) );
  NAND U17159 ( .A(n16781), .B(n16780), .Z(n16992) );
  NANDN U17160 ( .A(n16782), .B(n16909), .Z(n16786) );
  NAND U17161 ( .A(n16784), .B(n16783), .Z(n16785) );
  NAND U17162 ( .A(n16786), .B(n16785), .Z(n16996) );
  NAND U17163 ( .A(n16788), .B(n16787), .Z(n16792) );
  NAND U17164 ( .A(n16790), .B(n16789), .Z(n16791) );
  AND U17165 ( .A(n16792), .B(n16791), .Z(n17022) );
  AND U17166 ( .A(y[13]), .B(x[161]), .Z(n16913) );
  AND U17167 ( .A(y[48]), .B(x[174]), .Z(n16912) );
  XOR U17168 ( .A(n16913), .B(n16912), .Z(n16911) );
  AND U17169 ( .A(y[54]), .B(x[168]), .Z(n16910) );
  XOR U17170 ( .A(n16911), .B(n16910), .Z(n17024) );
  NAND U17171 ( .A(x[197]), .B(y[169]), .Z(n16793) );
  XNOR U17172 ( .A(n16794), .B(n16793), .Z(n16905) );
  AND U17173 ( .A(y[168]), .B(x[198]), .Z(n16904) );
  XOR U17174 ( .A(n16905), .B(n16904), .Z(n16902) );
  XNOR U17175 ( .A(n16903), .B(n16902), .Z(n17023) );
  XNOR U17176 ( .A(n17022), .B(n17021), .Z(n16995) );
  XOR U17177 ( .A(n16996), .B(n16995), .Z(n16993) );
  XOR U17178 ( .A(n16992), .B(n16993), .Z(n17063) );
  NAND U17179 ( .A(n16796), .B(n16795), .Z(n16800) );
  NAND U17180 ( .A(n16798), .B(n16797), .Z(n16799) );
  AND U17181 ( .A(n16800), .B(n16799), .Z(n17015) );
  AND U17182 ( .A(y[94]), .B(x[176]), .Z(n16877) );
  AND U17183 ( .A(y[8]), .B(x[166]), .Z(n16876) );
  XOR U17184 ( .A(n16877), .B(n16876), .Z(n16875) );
  AND U17185 ( .A(y[129]), .B(x[189]), .Z(n16874) );
  XOR U17186 ( .A(n16875), .B(n16874), .Z(n17038) );
  AND U17187 ( .A(y[49]), .B(x[173]), .Z(n16888) );
  AND U17188 ( .A(y[52]), .B(x[170]), .Z(n16887) );
  XOR U17189 ( .A(n16888), .B(n16887), .Z(n16886) );
  AND U17190 ( .A(y[53]), .B(x[169]), .Z(n16885) );
  XOR U17191 ( .A(n16886), .B(n16885), .Z(n16894) );
  NAND U17192 ( .A(x[172]), .B(y[50]), .Z(n16801) );
  XNOR U17193 ( .A(n16802), .B(n16801), .Z(n16893) );
  XOR U17194 ( .A(n16894), .B(n16893), .Z(n17037) );
  XOR U17195 ( .A(n17038), .B(n17037), .Z(n17036) );
  AND U17196 ( .A(y[174]), .B(x[192]), .Z(n16870) );
  XOR U17197 ( .A(n16871), .B(n16870), .Z(n16869) );
  AND U17198 ( .A(y[88]), .B(x[182]), .Z(n16868) );
  XOR U17199 ( .A(n16869), .B(n16868), .Z(n17035) );
  XOR U17200 ( .A(n17036), .B(n17035), .Z(n17018) );
  IV U17201 ( .A(n17018), .Z(n16813) );
  NAND U17202 ( .A(n16804), .B(n16803), .Z(n16808) );
  NAND U17203 ( .A(n16806), .B(n16805), .Z(n16807) );
  AND U17204 ( .A(n16808), .B(n16807), .Z(n16899) );
  AND U17205 ( .A(y[130]), .B(x[188]), .Z(n16866) );
  AND U17206 ( .A(x[177]), .B(y[93]), .Z(n16810) );
  AND U17207 ( .A(x[178]), .B(y[92]), .Z(n16809) );
  XOR U17208 ( .A(n16810), .B(n16809), .Z(n16865) );
  XOR U17209 ( .A(n16866), .B(n16865), .Z(n16901) );
  AND U17210 ( .A(y[14]), .B(x[160]), .Z(n16883) );
  AND U17211 ( .A(x[184]), .B(y[134]), .Z(n16812) );
  NAND U17212 ( .A(x[185]), .B(y[133]), .Z(n16811) );
  XNOR U17213 ( .A(n16812), .B(n16811), .Z(n16882) );
  XNOR U17214 ( .A(n16883), .B(n16882), .Z(n16900) );
  XOR U17215 ( .A(n16899), .B(n16898), .Z(n17017) );
  XNOR U17216 ( .A(n16813), .B(n17017), .Z(n17016) );
  XNOR U17217 ( .A(n17015), .B(n17016), .Z(n17065) );
  XOR U17218 ( .A(n17066), .B(n17065), .Z(n17060) );
  XNOR U17219 ( .A(n17059), .B(n17060), .Z(n17058) );
  XNOR U17220 ( .A(n17057), .B(n17058), .Z(n17077) );
  XOR U17221 ( .A(n17078), .B(n17077), .Z(n17084) );
  NANDN U17222 ( .A(n16815), .B(n16814), .Z(n16819) );
  NANDN U17223 ( .A(n16817), .B(n16816), .Z(n16818) );
  AND U17224 ( .A(n16819), .B(n16818), .Z(n17086) );
  NAND U17225 ( .A(n16821), .B(n16820), .Z(n16825) );
  NAND U17226 ( .A(n16823), .B(n16822), .Z(n16824) );
  NAND U17227 ( .A(n16825), .B(n16824), .Z(n17085) );
  NANDN U17228 ( .A(n16827), .B(n16826), .Z(n16831) );
  NAND U17229 ( .A(n16829), .B(n16828), .Z(n16830) );
  NAND U17230 ( .A(n16831), .B(n16830), .Z(n17071) );
  XOR U17231 ( .A(n17072), .B(n17071), .Z(o[174]) );
  NAND U17232 ( .A(n16841), .B(n16840), .Z(n16845) );
  NAND U17233 ( .A(n16843), .B(n16842), .Z(n16844) );
  AND U17234 ( .A(n16845), .B(n16844), .Z(n17056) );
  NAND U17235 ( .A(n16847), .B(n16846), .Z(n16851) );
  NANDN U17236 ( .A(n16849), .B(n16848), .Z(n16850) );
  AND U17237 ( .A(n16851), .B(n16850), .Z(n17014) );
  NAND U17238 ( .A(n16853), .B(n16852), .Z(n16856) );
  AND U17239 ( .A(y[10]), .B(x[165]), .Z(n16961) );
  NAND U17240 ( .A(n16854), .B(n16961), .Z(n16855) );
  AND U17241 ( .A(n16856), .B(n16855), .Z(n16864) );
  NAND U17242 ( .A(n16858), .B(n16857), .Z(n16862) );
  NAND U17243 ( .A(n16860), .B(n16859), .Z(n16861) );
  NAND U17244 ( .A(n16862), .B(n16861), .Z(n16863) );
  XNOR U17245 ( .A(n16864), .B(n16863), .Z(n16873) );
  AND U17246 ( .A(y[93]), .B(x[178]), .Z(n16967) );
  XOR U17247 ( .A(n16873), .B(n16872), .Z(n16892) );
  AND U17248 ( .A(y[134]), .B(x[185]), .Z(n16966) );
  XNOR U17249 ( .A(n16890), .B(n16889), .Z(n16891) );
  XNOR U17250 ( .A(n16892), .B(n16891), .Z(n17012) );
  NAND U17251 ( .A(n16894), .B(n16893), .Z(n16897) );
  AND U17252 ( .A(y[50]), .B(x[171]), .Z(n16895) );
  AND U17253 ( .A(y[51]), .B(x[172]), .Z(n16960) );
  NAND U17254 ( .A(n16895), .B(n16960), .Z(n16896) );
  AND U17255 ( .A(n16897), .B(n16896), .Z(n17010) );
  AND U17256 ( .A(x[169]), .B(y[54]), .Z(n16915) );
  NAND U17257 ( .A(x[170]), .B(y[53]), .Z(n16914) );
  XNOR U17258 ( .A(n16915), .B(n16914), .Z(n16921) );
  AND U17259 ( .A(x[184]), .B(y[135]), .Z(n16919) );
  NAND U17260 ( .A(y[169]), .B(x[196]), .Z(n16916) );
  AND U17261 ( .A(x[197]), .B(n16916), .Z(n16917) );
  NAND U17262 ( .A(n16917), .B(y[170]), .Z(n16918) );
  XNOR U17263 ( .A(n16919), .B(n16918), .Z(n16920) );
  XOR U17264 ( .A(n16921), .B(n16920), .Z(n16929) );
  AND U17265 ( .A(x[160]), .B(y[15]), .Z(n16923) );
  NAND U17266 ( .A(x[186]), .B(y[133]), .Z(n16922) );
  XNOR U17267 ( .A(n16923), .B(n16922), .Z(n16927) );
  AND U17268 ( .A(x[175]), .B(y[48]), .Z(n16925) );
  NAND U17269 ( .A(x[173]), .B(y[50]), .Z(n16924) );
  XNOR U17270 ( .A(n16925), .B(n16924), .Z(n16926) );
  XNOR U17271 ( .A(n16927), .B(n16926), .Z(n16928) );
  AND U17272 ( .A(x[188]), .B(y[131]), .Z(n16931) );
  NAND U17273 ( .A(x[167]), .B(y[8]), .Z(n16930) );
  XNOR U17274 ( .A(n16931), .B(n16930), .Z(n16935) );
  AND U17275 ( .A(x[163]), .B(y[12]), .Z(n16933) );
  NAND U17276 ( .A(x[174]), .B(y[49]), .Z(n16932) );
  XNOR U17277 ( .A(n16933), .B(n16932), .Z(n16934) );
  XOR U17278 ( .A(n16935), .B(n16934), .Z(n16943) );
  AND U17279 ( .A(x[179]), .B(y[92]), .Z(n16937) );
  NAND U17280 ( .A(x[199]), .B(y[168]), .Z(n16936) );
  XNOR U17281 ( .A(n16937), .B(n16936), .Z(n16941) );
  AND U17282 ( .A(x[177]), .B(y[94]), .Z(n16939) );
  NAND U17283 ( .A(x[198]), .B(y[169]), .Z(n16938) );
  XNOR U17284 ( .A(n16939), .B(n16938), .Z(n16940) );
  XNOR U17285 ( .A(n16941), .B(n16940), .Z(n16942) );
  XNOR U17286 ( .A(n16943), .B(n16942), .Z(n16959) );
  AND U17287 ( .A(x[193]), .B(y[174]), .Z(n16945) );
  NAND U17288 ( .A(x[180]), .B(y[91]), .Z(n16944) );
  XNOR U17289 ( .A(n16945), .B(n16944), .Z(n16949) );
  AND U17290 ( .A(x[161]), .B(y[14]), .Z(n16947) );
  NAND U17291 ( .A(x[181]), .B(y[90]), .Z(n16946) );
  XNOR U17292 ( .A(n16947), .B(n16946), .Z(n16948) );
  XOR U17293 ( .A(n16949), .B(n16948), .Z(n16957) );
  AND U17294 ( .A(x[164]), .B(y[11]), .Z(n16951) );
  NAND U17295 ( .A(x[189]), .B(y[130]), .Z(n16950) );
  XNOR U17296 ( .A(n16951), .B(n16950), .Z(n16955) );
  AND U17297 ( .A(x[194]), .B(y[173]), .Z(n16953) );
  NAND U17298 ( .A(x[195]), .B(y[172]), .Z(n16952) );
  XNOR U17299 ( .A(n16953), .B(n16952), .Z(n16954) );
  XNOR U17300 ( .A(n16955), .B(n16954), .Z(n16956) );
  XNOR U17301 ( .A(n16957), .B(n16956), .Z(n16958) );
  XOR U17302 ( .A(n16959), .B(n16958), .Z(n16991) );
  XOR U17303 ( .A(n16961), .B(n16960), .Z(n16965) );
  XNOR U17304 ( .A(n16963), .B(n16962), .Z(n16964) );
  XNOR U17305 ( .A(n16965), .B(n16964), .Z(n16989) );
  AND U17306 ( .A(x[176]), .B(y[95]), .Z(n16987) );
  AND U17307 ( .A(x[168]), .B(y[55]), .Z(n16969) );
  XNOR U17308 ( .A(n16967), .B(n16966), .Z(n16968) );
  XNOR U17309 ( .A(n16969), .B(n16968), .Z(n16985) );
  AND U17310 ( .A(x[166]), .B(y[9]), .Z(n16971) );
  NAND U17311 ( .A(x[182]), .B(y[89]), .Z(n16970) );
  XNOR U17312 ( .A(n16971), .B(n16970), .Z(n16975) );
  AND U17313 ( .A(x[187]), .B(y[132]), .Z(n16973) );
  NAND U17314 ( .A(x[162]), .B(y[13]), .Z(n16972) );
  XNOR U17315 ( .A(n16973), .B(n16972), .Z(n16974) );
  XOR U17316 ( .A(n16975), .B(n16974), .Z(n16983) );
  AND U17317 ( .A(x[192]), .B(y[175]), .Z(n16977) );
  NAND U17318 ( .A(x[183]), .B(y[88]), .Z(n16976) );
  XNOR U17319 ( .A(n16977), .B(n16976), .Z(n16981) );
  AND U17320 ( .A(x[190]), .B(y[129]), .Z(n16979) );
  NAND U17321 ( .A(x[191]), .B(y[128]), .Z(n16978) );
  XNOR U17322 ( .A(n16979), .B(n16978), .Z(n16980) );
  XNOR U17323 ( .A(n16981), .B(n16980), .Z(n16982) );
  XNOR U17324 ( .A(n16983), .B(n16982), .Z(n16984) );
  XNOR U17325 ( .A(n16985), .B(n16984), .Z(n16986) );
  XNOR U17326 ( .A(n16987), .B(n16986), .Z(n16988) );
  XNOR U17327 ( .A(n16989), .B(n16988), .Z(n16990) );
  IV U17328 ( .A(n16992), .Z(n16994) );
  NANDN U17329 ( .A(n16994), .B(n16993), .Z(n16998) );
  NAND U17330 ( .A(n16996), .B(n16995), .Z(n16997) );
  AND U17331 ( .A(n16998), .B(n16997), .Z(n17006) );
  NAND U17332 ( .A(n17000), .B(n16999), .Z(n17004) );
  NAND U17333 ( .A(n17002), .B(n17001), .Z(n17003) );
  NAND U17334 ( .A(n17004), .B(n17003), .Z(n17005) );
  XNOR U17335 ( .A(n17006), .B(n17005), .Z(n17007) );
  XNOR U17336 ( .A(n17008), .B(n17007), .Z(n17009) );
  XNOR U17337 ( .A(n17010), .B(n17009), .Z(n17011) );
  XNOR U17338 ( .A(n17012), .B(n17011), .Z(n17013) );
  XNOR U17339 ( .A(n17014), .B(n17013), .Z(n17054) );
  NANDN U17340 ( .A(n17016), .B(n17015), .Z(n17020) );
  NANDN U17341 ( .A(n17018), .B(n17017), .Z(n17019) );
  AND U17342 ( .A(n17020), .B(n17019), .Z(n17052) );
  NAND U17343 ( .A(n17022), .B(n17021), .Z(n17026) );
  NANDN U17344 ( .A(n17024), .B(n17023), .Z(n17025) );
  AND U17345 ( .A(n17026), .B(n17025), .Z(n17034) );
  NAND U17346 ( .A(n17028), .B(n17027), .Z(n17032) );
  NANDN U17347 ( .A(n17030), .B(n17029), .Z(n17031) );
  NAND U17348 ( .A(n17032), .B(n17031), .Z(n17033) );
  XNOR U17349 ( .A(n17034), .B(n17033), .Z(n17050) );
  NAND U17350 ( .A(n17036), .B(n17035), .Z(n17040) );
  NAND U17351 ( .A(n17038), .B(n17037), .Z(n17039) );
  AND U17352 ( .A(n17040), .B(n17039), .Z(n17048) );
  NAND U17353 ( .A(n17042), .B(n17041), .Z(n17046) );
  NAND U17354 ( .A(n17044), .B(n17043), .Z(n17045) );
  NAND U17355 ( .A(n17046), .B(n17045), .Z(n17047) );
  XNOR U17356 ( .A(n17048), .B(n17047), .Z(n17049) );
  XNOR U17357 ( .A(n17050), .B(n17049), .Z(n17051) );
  XNOR U17358 ( .A(n17052), .B(n17051), .Z(n17053) );
  XNOR U17359 ( .A(n17054), .B(n17053), .Z(n17055) );
  NANDN U17360 ( .A(n17058), .B(n17057), .Z(n17062) );
  AND U17361 ( .A(n17060), .B(n17059), .Z(n17061) );
  ANDN U17362 ( .B(n17062), .A(n17061), .Z(n17070) );
  ANDN U17363 ( .B(n17064), .A(n17063), .Z(n17068) );
  AND U17364 ( .A(n17066), .B(n17065), .Z(n17067) );
  OR U17365 ( .A(n17068), .B(n17067), .Z(n17069) );
  NAND U17366 ( .A(n17072), .B(n17071), .Z(n17076) );
  NANDN U17367 ( .A(n17074), .B(n17073), .Z(n17075) );
  NAND U17368 ( .A(n17078), .B(n17077), .Z(n17082) );
  NANDN U17369 ( .A(n17080), .B(n17079), .Z(n17081) );
  NAND U17370 ( .A(y[176]), .B(x[192]), .Z(n17222) );
  NAND U17371 ( .A(y[56]), .B(x[168]), .Z(n17089) );
  XOR U17372 ( .A(n17222), .B(n17089), .Z(n17090) );
  AND U17373 ( .A(y[16]), .B(x[160]), .Z(n17097) );
  AND U17374 ( .A(y[96]), .B(x[176]), .Z(n17094) );
  XOR U17375 ( .A(n17097), .B(n17094), .Z(n17093) );
  AND U17376 ( .A(y[136]), .B(x[184]), .Z(n17092) );
  XNOR U17377 ( .A(n17093), .B(n17092), .Z(n17091) );
  XNOR U17378 ( .A(n17090), .B(n17091), .Z(o[176]) );
  AND U17379 ( .A(x[161]), .B(y[16]), .Z(n17088) );
  NAND U17380 ( .A(x[160]), .B(y[17]), .Z(n17087) );
  XNOR U17381 ( .A(n17088), .B(n17087), .Z(n17098) );
  NAND U17382 ( .A(y[56]), .B(x[169]), .Z(n17099) );
  XOR U17383 ( .A(n17098), .B(n17099), .Z(n17115) );
  AND U17384 ( .A(y[176]), .B(x[193]), .Z(n17323) );
  NAND U17385 ( .A(y[97]), .B(x[176]), .Z(n17102) );
  XNOR U17386 ( .A(n17323), .B(n17102), .Z(n17103) );
  AND U17387 ( .A(y[177]), .B(x[192]), .Z(n17127) );
  NAND U17388 ( .A(y[96]), .B(x[177]), .Z(n17126) );
  XOR U17389 ( .A(n17127), .B(n17126), .Z(n17104) );
  XOR U17390 ( .A(n17103), .B(n17104), .Z(n17114) );
  AND U17391 ( .A(y[57]), .B(x[168]), .Z(n17346) );
  AND U17392 ( .A(y[137]), .B(x[184]), .Z(n17119) );
  XOR U17393 ( .A(n17346), .B(n17119), .Z(n17121) );
  AND U17394 ( .A(y[136]), .B(x[185]), .Z(n17120) );
  XNOR U17395 ( .A(n17121), .B(n17120), .Z(n17113) );
  XOR U17396 ( .A(n17114), .B(n17113), .Z(n17116) );
  XOR U17397 ( .A(n17115), .B(n17116), .Z(n17110) );
  NAND U17398 ( .A(n17093), .B(n17092), .Z(n17096) );
  AND U17399 ( .A(n17097), .B(n17094), .Z(n17095) );
  ANDN U17400 ( .B(n17096), .A(n17095), .Z(n17107) );
  XNOR U17401 ( .A(n17108), .B(n17107), .Z(n17109) );
  XNOR U17402 ( .A(n17110), .B(n17109), .Z(o[177]) );
  AND U17403 ( .A(y[17]), .B(x[161]), .Z(n17149) );
  NAND U17404 ( .A(n17149), .B(n17097), .Z(n17101) );
  NANDN U17405 ( .A(n17099), .B(n17098), .Z(n17100) );
  NAND U17406 ( .A(n17101), .B(n17100), .Z(n17170) );
  NANDN U17407 ( .A(n17102), .B(n17323), .Z(n17106) );
  NANDN U17408 ( .A(n17104), .B(n17103), .Z(n17105) );
  NAND U17409 ( .A(n17106), .B(n17105), .Z(n17168) );
  AND U17410 ( .A(y[138]), .B(x[184]), .Z(n17174) );
  NAND U17411 ( .A(y[18]), .B(x[160]), .Z(n17175) );
  XNOR U17412 ( .A(n17174), .B(n17175), .Z(n17177) );
  AND U17413 ( .A(y[56]), .B(x[170]), .Z(n17176) );
  XOR U17414 ( .A(n17177), .B(n17176), .Z(n17169) );
  XOR U17415 ( .A(n17168), .B(n17169), .Z(n17171) );
  XNOR U17416 ( .A(n17170), .B(n17171), .Z(n17129) );
  NANDN U17417 ( .A(n17108), .B(n17107), .Z(n17112) );
  NAND U17418 ( .A(n17110), .B(n17109), .Z(n17111) );
  NAND U17419 ( .A(n17112), .B(n17111), .Z(n17128) );
  XOR U17420 ( .A(n17129), .B(n17128), .Z(n17131) );
  NAND U17421 ( .A(n17114), .B(n17113), .Z(n17118) );
  NAND U17422 ( .A(n17116), .B(n17115), .Z(n17117) );
  AND U17423 ( .A(n17118), .B(n17117), .Z(n17137) );
  AND U17424 ( .A(y[16]), .B(x[162]), .Z(n17147) );
  AND U17425 ( .A(y[98]), .B(x[176]), .Z(n17146) );
  XOR U17426 ( .A(n17147), .B(n17146), .Z(n17148) );
  XOR U17427 ( .A(n17149), .B(n17148), .Z(n17183) );
  AND U17428 ( .A(y[136]), .B(x[186]), .Z(n17182) );
  XOR U17429 ( .A(n17183), .B(n17182), .Z(n17185) );
  AND U17430 ( .A(y[96]), .B(x[178]), .Z(n17252) );
  AND U17431 ( .A(y[178]), .B(x[192]), .Z(n17160) );
  XOR U17432 ( .A(n17252), .B(n17160), .Z(n17162) );
  AND U17433 ( .A(y[97]), .B(x[177]), .Z(n17161) );
  XOR U17434 ( .A(n17162), .B(n17161), .Z(n17184) );
  XOR U17435 ( .A(n17185), .B(n17184), .Z(n17134) );
  AND U17436 ( .A(n17346), .B(n17119), .Z(n17123) );
  NAND U17437 ( .A(n17121), .B(n17120), .Z(n17122) );
  NANDN U17438 ( .A(n17123), .B(n17122), .Z(n17142) );
  AND U17439 ( .A(x[194]), .B(y[176]), .Z(n17125) );
  NAND U17440 ( .A(x[193]), .B(y[177]), .Z(n17124) );
  XNOR U17441 ( .A(n17125), .B(n17124), .Z(n17181) );
  ANDN U17442 ( .B(n17127), .A(n17126), .Z(n17180) );
  XOR U17443 ( .A(n17181), .B(n17180), .Z(n17141) );
  AND U17444 ( .A(y[137]), .B(x[185]), .Z(n17152) );
  NAND U17445 ( .A(y[57]), .B(x[169]), .Z(n17153) );
  XNOR U17446 ( .A(n17152), .B(n17153), .Z(n17154) );
  NAND U17447 ( .A(y[58]), .B(x[168]), .Z(n17155) );
  XNOR U17448 ( .A(n17154), .B(n17155), .Z(n17140) );
  XOR U17449 ( .A(n17141), .B(n17140), .Z(n17143) );
  XOR U17450 ( .A(n17142), .B(n17143), .Z(n17135) );
  XOR U17451 ( .A(n17134), .B(n17135), .Z(n17136) );
  XNOR U17452 ( .A(n17137), .B(n17136), .Z(n17130) );
  XNOR U17453 ( .A(n17131), .B(n17130), .Z(o[178]) );
  NAND U17454 ( .A(n17129), .B(n17128), .Z(n17133) );
  NAND U17455 ( .A(n17131), .B(n17130), .Z(n17132) );
  AND U17456 ( .A(n17133), .B(n17132), .Z(n17189) );
  NAND U17457 ( .A(n17135), .B(n17134), .Z(n17139) );
  NAND U17458 ( .A(n17137), .B(n17136), .Z(n17138) );
  NAND U17459 ( .A(n17139), .B(n17138), .Z(n17194) );
  NAND U17460 ( .A(n17141), .B(n17140), .Z(n17145) );
  NAND U17461 ( .A(n17143), .B(n17142), .Z(n17144) );
  NAND U17462 ( .A(n17145), .B(n17144), .Z(n17192) );
  NAND U17463 ( .A(n17147), .B(n17146), .Z(n17151) );
  NAND U17464 ( .A(n17149), .B(n17148), .Z(n17150) );
  NAND U17465 ( .A(n17151), .B(n17150), .Z(n17204) );
  NANDN U17466 ( .A(n17153), .B(n17152), .Z(n17157) );
  NANDN U17467 ( .A(n17155), .B(n17154), .Z(n17156) );
  AND U17468 ( .A(n17157), .B(n17156), .Z(n17243) );
  AND U17469 ( .A(y[139]), .B(x[184]), .Z(n17270) );
  AND U17470 ( .A(y[99]), .B(x[176]), .Z(n17269) );
  NAND U17471 ( .A(y[16]), .B(x[163]), .Z(n17268) );
  XOR U17472 ( .A(n17269), .B(n17268), .Z(n17271) );
  XOR U17473 ( .A(n17270), .B(n17271), .Z(n17241) );
  AND U17474 ( .A(x[179]), .B(y[96]), .Z(n17159) );
  NAND U17475 ( .A(x[178]), .B(y[97]), .Z(n17158) );
  XNOR U17476 ( .A(n17159), .B(n17158), .Z(n17253) );
  NAND U17477 ( .A(y[98]), .B(x[177]), .Z(n17254) );
  XNOR U17478 ( .A(n17253), .B(n17254), .Z(n17240) );
  XNOR U17479 ( .A(n17241), .B(n17240), .Z(n17242) );
  XNOR U17480 ( .A(n17243), .B(n17242), .Z(n17205) );
  XOR U17481 ( .A(n17204), .B(n17205), .Z(n17207) );
  NAND U17482 ( .A(n17252), .B(n17160), .Z(n17164) );
  AND U17483 ( .A(n17162), .B(n17161), .Z(n17163) );
  ANDN U17484 ( .B(n17164), .A(n17163), .Z(n17248) );
  AND U17485 ( .A(y[18]), .B(x[161]), .Z(n17218) );
  AND U17486 ( .A(y[17]), .B(x[162]), .Z(n17217) );
  NAND U17487 ( .A(y[138]), .B(x[185]), .Z(n17216) );
  XOR U17488 ( .A(n17217), .B(n17216), .Z(n17219) );
  XOR U17489 ( .A(n17218), .B(n17219), .Z(n17247) );
  AND U17490 ( .A(x[195]), .B(y[176]), .Z(n17166) );
  NAND U17491 ( .A(x[192]), .B(y[179]), .Z(n17165) );
  XNOR U17492 ( .A(n17166), .B(n17165), .Z(n17223) );
  AND U17493 ( .A(y[177]), .B(x[194]), .Z(n17320) );
  NAND U17494 ( .A(x[193]), .B(y[178]), .Z(n17167) );
  XOR U17495 ( .A(n17320), .B(n17167), .Z(n17224) );
  XNOR U17496 ( .A(n17223), .B(n17224), .Z(n17246) );
  XOR U17497 ( .A(n17247), .B(n17246), .Z(n17249) );
  XOR U17498 ( .A(n17248), .B(n17249), .Z(n17206) );
  XOR U17499 ( .A(n17207), .B(n17206), .Z(n17193) );
  XOR U17500 ( .A(n17192), .B(n17193), .Z(n17195) );
  XOR U17501 ( .A(n17194), .B(n17195), .Z(n17188) );
  XOR U17502 ( .A(n17189), .B(n17188), .Z(n17191) );
  NAND U17503 ( .A(n17169), .B(n17168), .Z(n17173) );
  NAND U17504 ( .A(n17171), .B(n17170), .Z(n17172) );
  AND U17505 ( .A(n17173), .B(n17172), .Z(n17201) );
  NANDN U17506 ( .A(n17175), .B(n17174), .Z(n17179) );
  NAND U17507 ( .A(n17177), .B(n17176), .Z(n17178) );
  AND U17508 ( .A(n17179), .B(n17178), .Z(n17211) );
  XNOR U17509 ( .A(n17211), .B(n17210), .Z(n17213) );
  NAND U17510 ( .A(y[56]), .B(x[171]), .Z(n17262) );
  NAND U17511 ( .A(y[19]), .B(x[160]), .Z(n17260) );
  NAND U17512 ( .A(y[137]), .B(x[186]), .Z(n17259) );
  XOR U17513 ( .A(n17260), .B(n17259), .Z(n17261) );
  XNOR U17514 ( .A(n17262), .B(n17261), .Z(n17237) );
  NAND U17515 ( .A(y[59]), .B(x[168]), .Z(n17231) );
  NAND U17516 ( .A(y[57]), .B(x[170]), .Z(n17229) );
  NAND U17517 ( .A(y[136]), .B(x[187]), .Z(n17228) );
  XOR U17518 ( .A(n17229), .B(n17228), .Z(n17230) );
  XNOR U17519 ( .A(n17231), .B(n17230), .Z(n17235) );
  AND U17520 ( .A(y[58]), .B(x[169]), .Z(n17234) );
  XOR U17521 ( .A(n17235), .B(n17234), .Z(n17236) );
  XOR U17522 ( .A(n17237), .B(n17236), .Z(n17212) );
  XNOR U17523 ( .A(n17213), .B(n17212), .Z(n17199) );
  NAND U17524 ( .A(n17183), .B(n17182), .Z(n17187) );
  NAND U17525 ( .A(n17185), .B(n17184), .Z(n17186) );
  AND U17526 ( .A(n17187), .B(n17186), .Z(n17198) );
  XOR U17527 ( .A(n17199), .B(n17198), .Z(n17200) );
  XNOR U17528 ( .A(n17201), .B(n17200), .Z(n17190) );
  XOR U17529 ( .A(n17191), .B(n17190), .Z(o[179]) );
  NAND U17530 ( .A(n17193), .B(n17192), .Z(n17197) );
  NAND U17531 ( .A(n17195), .B(n17194), .Z(n17196) );
  AND U17532 ( .A(n17197), .B(n17196), .Z(n17280) );
  NAND U17533 ( .A(n17199), .B(n17198), .Z(n17203) );
  NAND U17534 ( .A(n17201), .B(n17200), .Z(n17202) );
  NAND U17535 ( .A(n17203), .B(n17202), .Z(n17278) );
  NAND U17536 ( .A(n17205), .B(n17204), .Z(n17209) );
  NAND U17537 ( .A(n17207), .B(n17206), .Z(n17208) );
  AND U17538 ( .A(n17209), .B(n17208), .Z(n17279) );
  XOR U17539 ( .A(n17278), .B(n17279), .Z(n17281) );
  XOR U17540 ( .A(n17280), .B(n17281), .Z(n17274) );
  XOR U17541 ( .A(n17275), .B(n17274), .Z(n17277) );
  AND U17542 ( .A(x[168]), .B(y[60]), .Z(n17215) );
  NAND U17543 ( .A(x[171]), .B(y[57]), .Z(n17214) );
  XNOR U17544 ( .A(n17215), .B(n17214), .Z(n17347) );
  NAND U17545 ( .A(y[58]), .B(x[170]), .Z(n17407) );
  NAND U17546 ( .A(y[59]), .B(x[169]), .Z(n17357) );
  AND U17547 ( .A(y[136]), .B(x[188]), .Z(n17307) );
  NAND U17548 ( .A(y[19]), .B(x[161]), .Z(n17308) );
  NAND U17549 ( .A(y[20]), .B(x[160]), .Z(n17310) );
  XOR U17550 ( .A(n17359), .B(n17358), .Z(n17353) );
  NANDN U17551 ( .A(n17217), .B(n17216), .Z(n17221) );
  OR U17552 ( .A(n17219), .B(n17218), .Z(n17220) );
  AND U17553 ( .A(n17221), .B(n17220), .Z(n17351) );
  AND U17554 ( .A(y[179]), .B(x[195]), .Z(n17647) );
  NANDN U17555 ( .A(n17222), .B(n17647), .Z(n17226) );
  NANDN U17556 ( .A(n17224), .B(n17223), .Z(n17225) );
  AND U17557 ( .A(n17226), .B(n17225), .Z(n17350) );
  NAND U17558 ( .A(y[16]), .B(x[164]), .Z(n17332) );
  NAND U17559 ( .A(y[138]), .B(x[186]), .Z(n17331) );
  NAND U17560 ( .A(y[100]), .B(x[176]), .Z(n17330) );
  XNOR U17561 ( .A(n17331), .B(n17330), .Z(n17333) );
  AND U17562 ( .A(y[178]), .B(x[194]), .Z(n17267) );
  AND U17563 ( .A(y[177]), .B(x[193]), .Z(n17227) );
  NAND U17564 ( .A(n17267), .B(n17227), .Z(n17328) );
  NAND U17565 ( .A(y[180]), .B(x[192]), .Z(n17502) );
  NAND U17566 ( .A(y[96]), .B(x[180]), .Z(n17428) );
  XNOR U17567 ( .A(n17502), .B(n17428), .Z(n17329) );
  XOR U17568 ( .A(n17328), .B(n17329), .Z(n17290) );
  XOR U17569 ( .A(n17291), .B(n17290), .Z(n17293) );
  NAND U17570 ( .A(n17229), .B(n17228), .Z(n17233) );
  NAND U17571 ( .A(n17231), .B(n17230), .Z(n17232) );
  AND U17572 ( .A(n17233), .B(n17232), .Z(n17292) );
  XOR U17573 ( .A(n17293), .B(n17292), .Z(n17377) );
  NAND U17574 ( .A(n17235), .B(n17234), .Z(n17239) );
  NAND U17575 ( .A(n17237), .B(n17236), .Z(n17238) );
  AND U17576 ( .A(n17239), .B(n17238), .Z(n17376) );
  XNOR U17577 ( .A(n17377), .B(n17376), .Z(n17378) );
  XNOR U17578 ( .A(n17379), .B(n17378), .Z(n17284) );
  XNOR U17579 ( .A(n17285), .B(n17284), .Z(n17287) );
  NANDN U17580 ( .A(n17241), .B(n17240), .Z(n17245) );
  NANDN U17581 ( .A(n17243), .B(n17242), .Z(n17244) );
  AND U17582 ( .A(n17245), .B(n17244), .Z(n17369) );
  NANDN U17583 ( .A(n17247), .B(n17246), .Z(n17251) );
  OR U17584 ( .A(n17249), .B(n17248), .Z(n17250) );
  NAND U17585 ( .A(n17251), .B(n17250), .Z(n17368) );
  XNOR U17586 ( .A(n17369), .B(n17368), .Z(n17371) );
  AND U17587 ( .A(x[179]), .B(y[97]), .Z(n17258) );
  NAND U17588 ( .A(n17252), .B(n17258), .Z(n17256) );
  NANDN U17589 ( .A(n17254), .B(n17253), .Z(n17255) );
  AND U17590 ( .A(n17256), .B(n17255), .Z(n17373) );
  AND U17591 ( .A(y[56]), .B(x[172]), .Z(n17313) );
  NAND U17592 ( .A(y[140]), .B(x[184]), .Z(n17314) );
  NAND U17593 ( .A(y[139]), .B(x[185]), .Z(n17316) );
  NAND U17594 ( .A(x[178]), .B(y[98]), .Z(n17257) );
  XNOR U17595 ( .A(n17258), .B(n17257), .Z(n17303) );
  NAND U17596 ( .A(y[99]), .B(x[177]), .Z(n17304) );
  XOR U17597 ( .A(n17363), .B(n17362), .Z(n17364) );
  NAND U17598 ( .A(n17260), .B(n17259), .Z(n17264) );
  NAND U17599 ( .A(n17262), .B(n17261), .Z(n17263) );
  NAND U17600 ( .A(n17264), .B(n17263), .Z(n17365) );
  XNOR U17601 ( .A(n17373), .B(n17372), .Z(n17375) );
  NAND U17602 ( .A(y[18]), .B(x[162]), .Z(n17342) );
  NAND U17603 ( .A(y[137]), .B(x[187]), .Z(n17341) );
  NAND U17604 ( .A(y[17]), .B(x[163]), .Z(n17340) );
  XNOR U17605 ( .A(n17341), .B(n17340), .Z(n17343) );
  AND U17606 ( .A(x[196]), .B(y[176]), .Z(n17266) );
  NAND U17607 ( .A(x[193]), .B(y[179]), .Z(n17265) );
  XNOR U17608 ( .A(n17266), .B(n17265), .Z(n17325) );
  AND U17609 ( .A(y[177]), .B(x[195]), .Z(n17436) );
  XOR U17610 ( .A(n17436), .B(n17267), .Z(n17324) );
  XOR U17611 ( .A(n17325), .B(n17324), .Z(n17297) );
  XOR U17612 ( .A(n17296), .B(n17297), .Z(n17298) );
  NANDN U17613 ( .A(n17269), .B(n17268), .Z(n17273) );
  OR U17614 ( .A(n17271), .B(n17270), .Z(n17272) );
  NAND U17615 ( .A(n17273), .B(n17272), .Z(n17299) );
  XOR U17616 ( .A(n17375), .B(n17374), .Z(n17370) );
  XOR U17617 ( .A(n17371), .B(n17370), .Z(n17286) );
  XNOR U17618 ( .A(n17287), .B(n17286), .Z(n17276) );
  XNOR U17619 ( .A(n17277), .B(n17276), .Z(o[180]) );
  NAND U17620 ( .A(n17279), .B(n17278), .Z(n17283) );
  NAND U17621 ( .A(n17281), .B(n17280), .Z(n17282) );
  NAND U17622 ( .A(n17283), .B(n17282), .Z(n17527) );
  XNOR U17623 ( .A(n17526), .B(n17527), .Z(n17529) );
  NANDN U17624 ( .A(n17285), .B(n17284), .Z(n17289) );
  NAND U17625 ( .A(n17287), .B(n17286), .Z(n17288) );
  AND U17626 ( .A(n17289), .B(n17288), .Z(n17383) );
  NAND U17627 ( .A(n17291), .B(n17290), .Z(n17295) );
  NAND U17628 ( .A(n17293), .B(n17292), .Z(n17294) );
  AND U17629 ( .A(n17295), .B(n17294), .Z(n17438) );
  NAND U17630 ( .A(n17297), .B(n17296), .Z(n17301) );
  NANDN U17631 ( .A(n17299), .B(n17298), .Z(n17300) );
  NAND U17632 ( .A(n17301), .B(n17300), .Z(n17437) );
  AND U17633 ( .A(y[97]), .B(x[178]), .Z(n17302) );
  AND U17634 ( .A(y[98]), .B(x[179]), .Z(n17429) );
  NAND U17635 ( .A(n17302), .B(n17429), .Z(n17306) );
  NANDN U17636 ( .A(n17304), .B(n17303), .Z(n17305) );
  AND U17637 ( .A(n17306), .B(n17305), .Z(n17389) );
  NANDN U17638 ( .A(n17308), .B(n17307), .Z(n17312) );
  NANDN U17639 ( .A(n17310), .B(n17309), .Z(n17311) );
  NAND U17640 ( .A(n17312), .B(n17311), .Z(n17414) );
  AND U17641 ( .A(y[141]), .B(x[184]), .Z(n17715) );
  AND U17642 ( .A(y[56]), .B(x[173]), .Z(n17419) );
  AND U17643 ( .A(y[99]), .B(x[178]), .Z(n17418) );
  XOR U17644 ( .A(n17419), .B(n17418), .Z(n17420) );
  XOR U17645 ( .A(n17715), .B(n17420), .Z(n17413) );
  AND U17646 ( .A(y[137]), .B(x[188]), .Z(n17424) );
  AND U17647 ( .A(y[16]), .B(x[165]), .Z(n17423) );
  XOR U17648 ( .A(n17424), .B(n17423), .Z(n17425) );
  AND U17649 ( .A(y[17]), .B(x[164]), .Z(n17669) );
  XOR U17650 ( .A(n17425), .B(n17669), .Z(n17412) );
  XOR U17651 ( .A(n17413), .B(n17412), .Z(n17415) );
  XOR U17652 ( .A(n17414), .B(n17415), .Z(n17388) );
  NANDN U17653 ( .A(n17314), .B(n17313), .Z(n17318) );
  NANDN U17654 ( .A(n17316), .B(n17315), .Z(n17317) );
  NAND U17655 ( .A(n17318), .B(n17317), .Z(n17493) );
  AND U17656 ( .A(y[178]), .B(x[195]), .Z(n17319) );
  AND U17657 ( .A(n17320), .B(n17319), .Z(n17504) );
  AND U17658 ( .A(x[192]), .B(y[181]), .Z(n17322) );
  AND U17659 ( .A(x[193]), .B(y[180]), .Z(n17321) );
  XOR U17660 ( .A(n17322), .B(n17321), .Z(n17503) );
  XOR U17661 ( .A(n17504), .B(n17503), .Z(n17492) );
  AND U17662 ( .A(y[57]), .B(x[172]), .Z(n17484) );
  AND U17663 ( .A(y[61]), .B(x[168]), .Z(n17482) );
  AND U17664 ( .A(y[20]), .B(x[161]), .Z(n17481) );
  XOR U17665 ( .A(n17482), .B(n17481), .Z(n17483) );
  XOR U17666 ( .A(n17484), .B(n17483), .Z(n17491) );
  XOR U17667 ( .A(n17492), .B(n17491), .Z(n17494) );
  XOR U17668 ( .A(n17493), .B(n17494), .Z(n17390) );
  XOR U17669 ( .A(n17391), .B(n17390), .Z(n17439) );
  XOR U17670 ( .A(n17440), .B(n17439), .Z(n17524) );
  AND U17671 ( .A(y[179]), .B(x[196]), .Z(n17729) );
  NAND U17672 ( .A(n17729), .B(n17323), .Z(n17327) );
  NAND U17673 ( .A(n17325), .B(n17324), .Z(n17326) );
  AND U17674 ( .A(n17327), .B(n17326), .Z(n17450) );
  NAND U17675 ( .A(n17331), .B(n17330), .Z(n17335) );
  NANDN U17676 ( .A(n17333), .B(n17332), .Z(n17334) );
  AND U17677 ( .A(n17335), .B(n17334), .Z(n17458) );
  AND U17678 ( .A(y[60]), .B(x[169]), .Z(n17408) );
  AND U17679 ( .A(y[58]), .B(x[171]), .Z(n17577) );
  NAND U17680 ( .A(x[170]), .B(y[59]), .Z(n17336) );
  XOR U17681 ( .A(n17577), .B(n17336), .Z(n17409) );
  AND U17682 ( .A(y[177]), .B(x[196]), .Z(n17711) );
  NAND U17683 ( .A(x[195]), .B(y[178]), .Z(n17337) );
  XNOR U17684 ( .A(n17711), .B(n17337), .Z(n17397) );
  AND U17685 ( .A(y[176]), .B(x[197]), .Z(n17394) );
  NAND U17686 ( .A(y[179]), .B(x[194]), .Z(n17395) );
  XOR U17687 ( .A(n17397), .B(n17396), .Z(n17455) );
  XOR U17688 ( .A(n17456), .B(n17455), .Z(n17457) );
  XOR U17689 ( .A(n17458), .B(n17457), .Z(n17451) );
  XOR U17690 ( .A(n17452), .B(n17451), .Z(n17470) );
  AND U17691 ( .A(x[181]), .B(y[96]), .Z(n17339) );
  NAND U17692 ( .A(x[180]), .B(y[97]), .Z(n17338) );
  XOR U17693 ( .A(n17339), .B(n17338), .Z(n17430) );
  AND U17694 ( .A(y[136]), .B(x[189]), .Z(n17400) );
  NAND U17695 ( .A(y[18]), .B(x[163]), .Z(n17401) );
  AND U17696 ( .A(y[19]), .B(x[162]), .Z(n17402) );
  XOR U17697 ( .A(n17403), .B(n17402), .Z(n17473) );
  XOR U17698 ( .A(n17474), .B(n17473), .Z(n17476) );
  NAND U17699 ( .A(n17341), .B(n17340), .Z(n17345) );
  NANDN U17700 ( .A(n17343), .B(n17342), .Z(n17344) );
  AND U17701 ( .A(n17345), .B(n17344), .Z(n17475) );
  XOR U17702 ( .A(n17476), .B(n17475), .Z(n17468) );
  AND U17703 ( .A(y[60]), .B(x[171]), .Z(n17728) );
  NAND U17704 ( .A(n17728), .B(n17346), .Z(n17349) );
  NANDN U17705 ( .A(n17407), .B(n17347), .Z(n17348) );
  AND U17706 ( .A(n17349), .B(n17348), .Z(n17446) );
  AND U17707 ( .A(y[138]), .B(x[187]), .Z(n17497) );
  AND U17708 ( .A(y[100]), .B(x[177]), .Z(n17697) );
  XOR U17709 ( .A(n17497), .B(n17697), .Z(n17499) );
  AND U17710 ( .A(y[101]), .B(x[176]), .Z(n17498) );
  XOR U17711 ( .A(n17499), .B(n17498), .Z(n17444) );
  AND U17712 ( .A(y[21]), .B(x[160]), .Z(n17508) );
  AND U17713 ( .A(y[140]), .B(x[185]), .Z(n17507) );
  XOR U17714 ( .A(n17508), .B(n17507), .Z(n17510) );
  AND U17715 ( .A(y[139]), .B(x[186]), .Z(n17509) );
  XOR U17716 ( .A(n17510), .B(n17509), .Z(n17443) );
  XOR U17717 ( .A(n17444), .B(n17443), .Z(n17445) );
  XOR U17718 ( .A(n17446), .B(n17445), .Z(n17467) );
  NANDN U17719 ( .A(n17351), .B(n17350), .Z(n17355) );
  NANDN U17720 ( .A(n17353), .B(n17352), .Z(n17354) );
  AND U17721 ( .A(n17355), .B(n17354), .Z(n17464) );
  NANDN U17722 ( .A(n17357), .B(n17356), .Z(n17361) );
  NAND U17723 ( .A(n17359), .B(n17358), .Z(n17360) );
  AND U17724 ( .A(n17361), .B(n17360), .Z(n17462) );
  NAND U17725 ( .A(n17363), .B(n17362), .Z(n17367) );
  NANDN U17726 ( .A(n17365), .B(n17364), .Z(n17366) );
  NAND U17727 ( .A(n17367), .B(n17366), .Z(n17461) );
  XOR U17728 ( .A(n17464), .B(n17463), .Z(n17521) );
  XOR U17729 ( .A(n17522), .B(n17521), .Z(n17523) );
  XOR U17730 ( .A(n17524), .B(n17523), .Z(n17382) );
  XNOR U17731 ( .A(n17383), .B(n17382), .Z(n17384) );
  NANDN U17732 ( .A(n17377), .B(n17376), .Z(n17381) );
  NAND U17733 ( .A(n17379), .B(n17378), .Z(n17380) );
  AND U17734 ( .A(n17381), .B(n17380), .Z(n17515) );
  XNOR U17735 ( .A(n17516), .B(n17515), .Z(n17517) );
  XOR U17736 ( .A(n17518), .B(n17517), .Z(n17385) );
  XNOR U17737 ( .A(n17384), .B(n17385), .Z(n17528) );
  XOR U17738 ( .A(n17529), .B(n17528), .Z(o[181]) );
  NANDN U17739 ( .A(n17383), .B(n17382), .Z(n17387) );
  NANDN U17740 ( .A(n17385), .B(n17384), .Z(n17386) );
  AND U17741 ( .A(n17387), .B(n17386), .Z(n17813) );
  NANDN U17742 ( .A(n17389), .B(n17388), .Z(n17393) );
  NAND U17743 ( .A(n17391), .B(n17390), .Z(n17392) );
  AND U17744 ( .A(n17393), .B(n17392), .Z(n17818) );
  NANDN U17745 ( .A(n17395), .B(n17394), .Z(n17399) );
  NAND U17746 ( .A(n17397), .B(n17396), .Z(n17398) );
  NAND U17747 ( .A(n17399), .B(n17398), .Z(n17563) );
  NANDN U17748 ( .A(n17401), .B(n17400), .Z(n17405) );
  NAND U17749 ( .A(n17403), .B(n17402), .Z(n17404) );
  NAND U17750 ( .A(n17405), .B(n17404), .Z(n17566) );
  AND U17751 ( .A(y[59]), .B(x[171]), .Z(n17406) );
  NANDN U17752 ( .A(n17407), .B(n17406), .Z(n17411) );
  NANDN U17753 ( .A(n17409), .B(n17408), .Z(n17410) );
  AND U17754 ( .A(n17411), .B(n17410), .Z(n17641) );
  AND U17755 ( .A(y[139]), .B(x[187]), .Z(n17743) );
  AND U17756 ( .A(y[99]), .B(x[179]), .Z(n17742) );
  XOR U17757 ( .A(n17743), .B(n17742), .Z(n17741) );
  AND U17758 ( .A(y[19]), .B(x[163]), .Z(n17740) );
  XOR U17759 ( .A(n17741), .B(n17740), .Z(n17643) );
  AND U17760 ( .A(y[140]), .B(x[186]), .Z(n17757) );
  AND U17761 ( .A(y[98]), .B(x[180]), .Z(n17756) );
  XOR U17762 ( .A(n17757), .B(n17756), .Z(n17755) );
  AND U17763 ( .A(y[20]), .B(x[162]), .Z(n17754) );
  XNOR U17764 ( .A(n17755), .B(n17754), .Z(n17642) );
  XNOR U17765 ( .A(n17641), .B(n17640), .Z(n17565) );
  XOR U17766 ( .A(n17566), .B(n17565), .Z(n17564) );
  XOR U17767 ( .A(n17563), .B(n17564), .Z(n17542) );
  NAND U17768 ( .A(n17413), .B(n17412), .Z(n17417) );
  NAND U17769 ( .A(n17415), .B(n17414), .Z(n17416) );
  NAND U17770 ( .A(n17417), .B(n17416), .Z(n17541) );
  XOR U17771 ( .A(n17542), .B(n17541), .Z(n17540) );
  NAND U17772 ( .A(n17419), .B(n17418), .Z(n17422) );
  NAND U17773 ( .A(n17715), .B(n17420), .Z(n17421) );
  NAND U17774 ( .A(n17422), .B(n17421), .Z(n17685) );
  NAND U17775 ( .A(n17424), .B(n17423), .Z(n17427) );
  NAND U17776 ( .A(n17425), .B(n17669), .Z(n17426) );
  NAND U17777 ( .A(n17427), .B(n17426), .Z(n17684) );
  XOR U17778 ( .A(n17685), .B(n17684), .Z(n17683) );
  AND U17779 ( .A(y[97]), .B(x[181]), .Z(n17663) );
  NANDN U17780 ( .A(n17428), .B(n17663), .Z(n17432) );
  NANDN U17781 ( .A(n17430), .B(n17429), .Z(n17431) );
  AND U17782 ( .A(n17432), .B(n17431), .Z(n17689) );
  AND U17783 ( .A(x[164]), .B(y[18]), .Z(n17434) );
  NAND U17784 ( .A(x[165]), .B(y[17]), .Z(n17433) );
  XNOR U17785 ( .A(n17434), .B(n17433), .Z(n17667) );
  AND U17786 ( .A(y[136]), .B(x[190]), .Z(n17666) );
  XOR U17787 ( .A(n17667), .B(n17666), .Z(n17691) );
  AND U17788 ( .A(y[181]), .B(x[193]), .Z(n17655) );
  AND U17789 ( .A(y[178]), .B(x[196]), .Z(n17435) );
  AND U17790 ( .A(n17436), .B(n17435), .Z(n17653) );
  AND U17791 ( .A(y[180]), .B(x[194]), .Z(n17652) );
  XOR U17792 ( .A(n17653), .B(n17652), .Z(n17654) );
  XNOR U17793 ( .A(n17655), .B(n17654), .Z(n17690) );
  XNOR U17794 ( .A(n17689), .B(n17688), .Z(n17682) );
  XOR U17795 ( .A(n17683), .B(n17682), .Z(n17539) );
  XOR U17796 ( .A(n17540), .B(n17539), .Z(n17538) );
  NANDN U17797 ( .A(n17438), .B(n17437), .Z(n17442) );
  NAND U17798 ( .A(n17440), .B(n17439), .Z(n17441) );
  AND U17799 ( .A(n17442), .B(n17441), .Z(n17537) );
  NAND U17800 ( .A(n17444), .B(n17443), .Z(n17448) );
  NANDN U17801 ( .A(n17446), .B(n17445), .Z(n17447) );
  AND U17802 ( .A(n17448), .B(n17447), .Z(n17546) );
  NANDN U17803 ( .A(n17450), .B(n17449), .Z(n17454) );
  NAND U17804 ( .A(n17452), .B(n17451), .Z(n17453) );
  AND U17805 ( .A(n17454), .B(n17453), .Z(n17545) );
  XOR U17806 ( .A(n17546), .B(n17545), .Z(n17544) );
  NAND U17807 ( .A(n17456), .B(n17455), .Z(n17460) );
  NAND U17808 ( .A(n17458), .B(n17457), .Z(n17459) );
  AND U17809 ( .A(n17460), .B(n17459), .Z(n17543) );
  XOR U17810 ( .A(n17544), .B(n17543), .Z(n17535) );
  XOR U17811 ( .A(n17536), .B(n17535), .Z(n17817) );
  XOR U17812 ( .A(n17818), .B(n17817), .Z(n17820) );
  NANDN U17813 ( .A(n17462), .B(n17461), .Z(n17466) );
  NAND U17814 ( .A(n17464), .B(n17463), .Z(n17465) );
  AND U17815 ( .A(n17466), .B(n17465), .Z(n17797) );
  NANDN U17816 ( .A(n17468), .B(n17467), .Z(n17472) );
  NANDN U17817 ( .A(n17470), .B(n17469), .Z(n17471) );
  NAND U17818 ( .A(n17472), .B(n17471), .Z(n17798) );
  NAND U17819 ( .A(n17474), .B(n17473), .Z(n17478) );
  NAND U17820 ( .A(n17476), .B(n17475), .Z(n17477) );
  AND U17821 ( .A(n17478), .B(n17477), .Z(n17803) );
  AND U17822 ( .A(y[102]), .B(x[176]), .Z(n17703) );
  AND U17823 ( .A(y[16]), .B(x[166]), .Z(n17702) );
  XOR U17824 ( .A(n17703), .B(n17702), .Z(n17701) );
  AND U17825 ( .A(y[137]), .B(x[189]), .Z(n17700) );
  XOR U17826 ( .A(n17701), .B(n17700), .Z(n17572) );
  AND U17827 ( .A(y[57]), .B(x[173]), .Z(n17751) );
  AND U17828 ( .A(y[60]), .B(x[170]), .Z(n17750) );
  XOR U17829 ( .A(n17751), .B(n17750), .Z(n17749) );
  AND U17830 ( .A(y[61]), .B(x[169]), .Z(n17748) );
  XOR U17831 ( .A(n17749), .B(n17748), .Z(n17576) );
  AND U17832 ( .A(x[172]), .B(y[58]), .Z(n17480) );
  NAND U17833 ( .A(x[171]), .B(y[59]), .Z(n17479) );
  XNOR U17834 ( .A(n17480), .B(n17479), .Z(n17575) );
  XOR U17835 ( .A(n17576), .B(n17575), .Z(n17571) );
  XOR U17836 ( .A(n17572), .B(n17571), .Z(n17570) );
  AND U17837 ( .A(y[182]), .B(x[192]), .Z(n17662) );
  XOR U17838 ( .A(n17663), .B(n17662), .Z(n17661) );
  AND U17839 ( .A(y[96]), .B(x[182]), .Z(n17660) );
  XOR U17840 ( .A(n17661), .B(n17660), .Z(n17569) );
  XOR U17841 ( .A(n17570), .B(n17569), .Z(n17555) );
  NAND U17842 ( .A(n17482), .B(n17481), .Z(n17486) );
  NAND U17843 ( .A(n17484), .B(n17483), .Z(n17485) );
  AND U17844 ( .A(n17486), .B(n17485), .Z(n17779) );
  AND U17845 ( .A(y[138]), .B(x[188]), .Z(n17695) );
  AND U17846 ( .A(x[177]), .B(y[101]), .Z(n17488) );
  AND U17847 ( .A(x[178]), .B(y[100]), .Z(n17487) );
  XOR U17848 ( .A(n17488), .B(n17487), .Z(n17694) );
  XNOR U17849 ( .A(n17695), .B(n17694), .Z(n17777) );
  AND U17850 ( .A(y[22]), .B(x[160]), .Z(n17713) );
  AND U17851 ( .A(y[142]), .B(x[184]), .Z(n17490) );
  AND U17852 ( .A(x[185]), .B(y[141]), .Z(n17489) );
  XOR U17853 ( .A(n17490), .B(n17489), .Z(n17712) );
  XOR U17854 ( .A(n17713), .B(n17712), .Z(n17776) );
  XNOR U17855 ( .A(n17779), .B(n17778), .Z(n17556) );
  NAND U17856 ( .A(n17492), .B(n17491), .Z(n17496) );
  NAND U17857 ( .A(n17494), .B(n17493), .Z(n17495) );
  AND U17858 ( .A(n17496), .B(n17495), .Z(n17557) );
  XOR U17859 ( .A(n17558), .B(n17557), .Z(n17802) );
  XOR U17860 ( .A(n17803), .B(n17802), .Z(n17805) );
  NAND U17861 ( .A(n17497), .B(n17697), .Z(n17501) );
  NAND U17862 ( .A(n17499), .B(n17498), .Z(n17500) );
  NAND U17863 ( .A(n17501), .B(n17500), .Z(n17549) );
  NANDN U17864 ( .A(n17502), .B(n17655), .Z(n17506) );
  NAND U17865 ( .A(n17504), .B(n17503), .Z(n17505) );
  NAND U17866 ( .A(n17506), .B(n17505), .Z(n17552) );
  NAND U17867 ( .A(n17508), .B(n17507), .Z(n17512) );
  NAND U17868 ( .A(n17510), .B(n17509), .Z(n17511) );
  AND U17869 ( .A(n17512), .B(n17511), .Z(n17771) );
  AND U17870 ( .A(y[21]), .B(x[161]), .Z(n17737) );
  AND U17871 ( .A(y[56]), .B(x[174]), .Z(n17736) );
  XOR U17872 ( .A(n17737), .B(n17736), .Z(n17735) );
  AND U17873 ( .A(y[62]), .B(x[168]), .Z(n17734) );
  XOR U17874 ( .A(n17735), .B(n17734), .Z(n17772) );
  AND U17875 ( .A(x[197]), .B(y[177]), .Z(n17514) );
  NAND U17876 ( .A(x[196]), .B(y[178]), .Z(n17513) );
  XNOR U17877 ( .A(n17514), .B(n17513), .Z(n17649) );
  AND U17878 ( .A(y[176]), .B(x[198]), .Z(n17648) );
  XOR U17879 ( .A(n17649), .B(n17648), .Z(n17646) );
  XNOR U17880 ( .A(n17647), .B(n17646), .Z(n17773) );
  XNOR U17881 ( .A(n17771), .B(n17770), .Z(n17551) );
  XOR U17882 ( .A(n17552), .B(n17551), .Z(n17550) );
  XOR U17883 ( .A(n17549), .B(n17550), .Z(n17804) );
  XOR U17884 ( .A(n17798), .B(n17799), .Z(n17796) );
  XOR U17885 ( .A(n17797), .B(n17796), .Z(n17819) );
  XOR U17886 ( .A(n17820), .B(n17819), .Z(n17534) );
  NANDN U17887 ( .A(n17516), .B(n17515), .Z(n17520) );
  NANDN U17888 ( .A(n17518), .B(n17517), .Z(n17519) );
  AND U17889 ( .A(n17520), .B(n17519), .Z(n17533) );
  XOR U17890 ( .A(n17533), .B(n17532), .Z(n17525) );
  XOR U17891 ( .A(n17534), .B(n17525), .Z(n17814) );
  NANDN U17892 ( .A(n17527), .B(n17526), .Z(n17531) );
  NAND U17893 ( .A(n17529), .B(n17528), .Z(n17530) );
  NAND U17894 ( .A(n17531), .B(n17530), .Z(n17811) );
  XOR U17895 ( .A(n17812), .B(n17811), .Z(o[182]) );
  NAND U17896 ( .A(n17544), .B(n17543), .Z(n17548) );
  NAND U17897 ( .A(n17546), .B(n17545), .Z(n17547) );
  AND U17898 ( .A(n17548), .B(n17547), .Z(n17795) );
  NAND U17899 ( .A(n17550), .B(n17549), .Z(n17554) );
  AND U17900 ( .A(n17552), .B(n17551), .Z(n17553) );
  ANDN U17901 ( .B(n17554), .A(n17553), .Z(n17562) );
  ANDN U17902 ( .B(n17556), .A(n17555), .Z(n17560) );
  AND U17903 ( .A(n17558), .B(n17557), .Z(n17559) );
  OR U17904 ( .A(n17560), .B(n17559), .Z(n17561) );
  XNOR U17905 ( .A(n17562), .B(n17561), .Z(n17793) );
  NAND U17906 ( .A(n17564), .B(n17563), .Z(n17568) );
  NAND U17907 ( .A(n17566), .B(n17565), .Z(n17567) );
  AND U17908 ( .A(n17568), .B(n17567), .Z(n17791) );
  NAND U17909 ( .A(n17570), .B(n17569), .Z(n17574) );
  NAND U17910 ( .A(n17572), .B(n17571), .Z(n17573) );
  AND U17911 ( .A(n17574), .B(n17573), .Z(n17681) );
  NAND U17912 ( .A(n17576), .B(n17575), .Z(n17579) );
  AND U17913 ( .A(y[59]), .B(x[172]), .Z(n17629) );
  NAND U17914 ( .A(n17577), .B(n17629), .Z(n17578) );
  AND U17915 ( .A(n17579), .B(n17578), .Z(n17639) );
  AND U17916 ( .A(x[189]), .B(y[138]), .Z(n17581) );
  NAND U17917 ( .A(x[194]), .B(y[181]), .Z(n17580) );
  XNOR U17918 ( .A(n17581), .B(n17580), .Z(n17585) );
  AND U17919 ( .A(x[161]), .B(y[22]), .Z(n17583) );
  NAND U17920 ( .A(x[181]), .B(y[98]), .Z(n17582) );
  XNOR U17921 ( .A(n17583), .B(n17582), .Z(n17584) );
  XOR U17922 ( .A(n17585), .B(n17584), .Z(n17593) );
  AND U17923 ( .A(x[177]), .B(y[102]), .Z(n17587) );
  NAND U17924 ( .A(x[179]), .B(y[100]), .Z(n17586) );
  XNOR U17925 ( .A(n17587), .B(n17586), .Z(n17591) );
  AND U17926 ( .A(x[195]), .B(y[180]), .Z(n17589) );
  NAND U17927 ( .A(x[164]), .B(y[19]), .Z(n17588) );
  XNOR U17928 ( .A(n17589), .B(n17588), .Z(n17590) );
  XNOR U17929 ( .A(n17591), .B(n17590), .Z(n17592) );
  XNOR U17930 ( .A(n17593), .B(n17592), .Z(n17637) );
  AND U17931 ( .A(x[186]), .B(y[141]), .Z(n17598) );
  AND U17932 ( .A(y[178]), .B(x[197]), .Z(n17710) );
  AND U17933 ( .A(x[173]), .B(y[58]), .Z(n17595) );
  NAND U17934 ( .A(x[170]), .B(y[61]), .Z(n17594) );
  XNOR U17935 ( .A(n17595), .B(n17594), .Z(n17596) );
  XNOR U17936 ( .A(n17710), .B(n17596), .Z(n17597) );
  XNOR U17937 ( .A(n17598), .B(n17597), .Z(n17614) );
  AND U17938 ( .A(x[168]), .B(y[63]), .Z(n17600) );
  NAND U17939 ( .A(x[180]), .B(y[99]), .Z(n17599) );
  XNOR U17940 ( .A(n17600), .B(n17599), .Z(n17604) );
  AND U17941 ( .A(x[176]), .B(y[103]), .Z(n17602) );
  NAND U17942 ( .A(x[191]), .B(y[136]), .Z(n17601) );
  XNOR U17943 ( .A(n17602), .B(n17601), .Z(n17603) );
  XOR U17944 ( .A(n17604), .B(n17603), .Z(n17612) );
  AND U17945 ( .A(x[184]), .B(y[143]), .Z(n17606) );
  NAND U17946 ( .A(x[187]), .B(y[140]), .Z(n17605) );
  XNOR U17947 ( .A(n17606), .B(n17605), .Z(n17610) );
  AND U17948 ( .A(x[169]), .B(y[62]), .Z(n17608) );
  NAND U17949 ( .A(x[175]), .B(y[56]), .Z(n17607) );
  XNOR U17950 ( .A(n17608), .B(n17607), .Z(n17609) );
  XNOR U17951 ( .A(n17610), .B(n17609), .Z(n17611) );
  XNOR U17952 ( .A(n17612), .B(n17611), .Z(n17613) );
  XOR U17953 ( .A(n17614), .B(n17613), .Z(n17635) );
  AND U17954 ( .A(x[192]), .B(y[183]), .Z(n17616) );
  NAND U17955 ( .A(x[183]), .B(y[96]), .Z(n17615) );
  XNOR U17956 ( .A(n17616), .B(n17615), .Z(n17620) );
  AND U17957 ( .A(x[160]), .B(y[23]), .Z(n17618) );
  NAND U17958 ( .A(x[193]), .B(y[182]), .Z(n17617) );
  XNOR U17959 ( .A(n17618), .B(n17617), .Z(n17619) );
  XOR U17960 ( .A(n17620), .B(n17619), .Z(n17628) );
  AND U17961 ( .A(x[166]), .B(y[17]), .Z(n17622) );
  NAND U17962 ( .A(x[182]), .B(y[97]), .Z(n17621) );
  XNOR U17963 ( .A(n17622), .B(n17621), .Z(n17626) );
  AND U17964 ( .A(x[188]), .B(y[139]), .Z(n17624) );
  NAND U17965 ( .A(x[167]), .B(y[16]), .Z(n17623) );
  XNOR U17966 ( .A(n17624), .B(n17623), .Z(n17625) );
  XNOR U17967 ( .A(n17626), .B(n17625), .Z(n17627) );
  XNOR U17968 ( .A(n17628), .B(n17627), .Z(n17633) );
  AND U17969 ( .A(y[101]), .B(x[178]), .Z(n17696) );
  AND U17970 ( .A(y[142]), .B(x[185]), .Z(n17714) );
  XOR U17971 ( .A(n17696), .B(n17714), .Z(n17631) );
  AND U17972 ( .A(y[18]), .B(x[165]), .Z(n17668) );
  XNOR U17973 ( .A(n17668), .B(n17629), .Z(n17630) );
  XNOR U17974 ( .A(n17631), .B(n17630), .Z(n17632) );
  XNOR U17975 ( .A(n17633), .B(n17632), .Z(n17634) );
  XNOR U17976 ( .A(n17635), .B(n17634), .Z(n17636) );
  XNOR U17977 ( .A(n17637), .B(n17636), .Z(n17638) );
  XNOR U17978 ( .A(n17639), .B(n17638), .Z(n17679) );
  NAND U17979 ( .A(n17641), .B(n17640), .Z(n17645) );
  NANDN U17980 ( .A(n17643), .B(n17642), .Z(n17644) );
  AND U17981 ( .A(n17645), .B(n17644), .Z(n17677) );
  NAND U17982 ( .A(n17647), .B(n17646), .Z(n17651) );
  AND U17983 ( .A(n17649), .B(n17648), .Z(n17650) );
  ANDN U17984 ( .B(n17651), .A(n17650), .Z(n17659) );
  AND U17985 ( .A(n17653), .B(n17652), .Z(n17657) );
  AND U17986 ( .A(n17655), .B(n17654), .Z(n17656) );
  OR U17987 ( .A(n17657), .B(n17656), .Z(n17658) );
  XNOR U17988 ( .A(n17659), .B(n17658), .Z(n17675) );
  NAND U17989 ( .A(n17661), .B(n17660), .Z(n17665) );
  NAND U17990 ( .A(n17663), .B(n17662), .Z(n17664) );
  AND U17991 ( .A(n17665), .B(n17664), .Z(n17673) );
  NAND U17992 ( .A(n17667), .B(n17666), .Z(n17671) );
  NAND U17993 ( .A(n17669), .B(n17668), .Z(n17670) );
  NAND U17994 ( .A(n17671), .B(n17670), .Z(n17672) );
  XNOR U17995 ( .A(n17673), .B(n17672), .Z(n17674) );
  XNOR U17996 ( .A(n17675), .B(n17674), .Z(n17676) );
  XNOR U17997 ( .A(n17677), .B(n17676), .Z(n17678) );
  XNOR U17998 ( .A(n17679), .B(n17678), .Z(n17680) );
  XNOR U17999 ( .A(n17681), .B(n17680), .Z(n17789) );
  NAND U18000 ( .A(n17683), .B(n17682), .Z(n17687) );
  NAND U18001 ( .A(n17685), .B(n17684), .Z(n17686) );
  AND U18002 ( .A(n17687), .B(n17686), .Z(n17787) );
  NAND U18003 ( .A(n17689), .B(n17688), .Z(n17693) );
  NANDN U18004 ( .A(n17691), .B(n17690), .Z(n17692) );
  AND U18005 ( .A(n17693), .B(n17692), .Z(n17769) );
  NAND U18006 ( .A(n17695), .B(n17694), .Z(n17699) );
  NAND U18007 ( .A(n17697), .B(n17696), .Z(n17698) );
  AND U18008 ( .A(n17699), .B(n17698), .Z(n17707) );
  NAND U18009 ( .A(n17701), .B(n17700), .Z(n17705) );
  NAND U18010 ( .A(n17703), .B(n17702), .Z(n17704) );
  NAND U18011 ( .A(n17705), .B(n17704), .Z(n17706) );
  XNOR U18012 ( .A(n17707), .B(n17706), .Z(n17767) );
  AND U18013 ( .A(x[162]), .B(y[21]), .Z(n17709) );
  NAND U18014 ( .A(x[190]), .B(y[137]), .Z(n17708) );
  XNOR U18015 ( .A(n17709), .B(n17708), .Z(n17733) );
  AND U18016 ( .A(n17711), .B(n17710), .Z(n17727) );
  NAND U18017 ( .A(n17713), .B(n17712), .Z(n17717) );
  NAND U18018 ( .A(n17715), .B(n17714), .Z(n17716) );
  AND U18019 ( .A(n17717), .B(n17716), .Z(n17725) );
  AND U18020 ( .A(x[174]), .B(y[57]), .Z(n17719) );
  NAND U18021 ( .A(x[163]), .B(y[20]), .Z(n17718) );
  XNOR U18022 ( .A(n17719), .B(n17718), .Z(n17723) );
  AND U18023 ( .A(x[199]), .B(y[176]), .Z(n17721) );
  NAND U18024 ( .A(x[198]), .B(y[177]), .Z(n17720) );
  XNOR U18025 ( .A(n17721), .B(n17720), .Z(n17722) );
  XNOR U18026 ( .A(n17723), .B(n17722), .Z(n17724) );
  XNOR U18027 ( .A(n17725), .B(n17724), .Z(n17726) );
  XOR U18028 ( .A(n17727), .B(n17726), .Z(n17731) );
  XNOR U18029 ( .A(n17729), .B(n17728), .Z(n17730) );
  XNOR U18030 ( .A(n17731), .B(n17730), .Z(n17732) );
  XOR U18031 ( .A(n17733), .B(n17732), .Z(n17765) );
  NAND U18032 ( .A(n17735), .B(n17734), .Z(n17739) );
  NAND U18033 ( .A(n17737), .B(n17736), .Z(n17738) );
  AND U18034 ( .A(n17739), .B(n17738), .Z(n17747) );
  NAND U18035 ( .A(n17741), .B(n17740), .Z(n17745) );
  NAND U18036 ( .A(n17743), .B(n17742), .Z(n17744) );
  NAND U18037 ( .A(n17745), .B(n17744), .Z(n17746) );
  XNOR U18038 ( .A(n17747), .B(n17746), .Z(n17763) );
  NAND U18039 ( .A(n17749), .B(n17748), .Z(n17753) );
  NAND U18040 ( .A(n17751), .B(n17750), .Z(n17752) );
  AND U18041 ( .A(n17753), .B(n17752), .Z(n17761) );
  NAND U18042 ( .A(n17755), .B(n17754), .Z(n17759) );
  NAND U18043 ( .A(n17757), .B(n17756), .Z(n17758) );
  NAND U18044 ( .A(n17759), .B(n17758), .Z(n17760) );
  XNOR U18045 ( .A(n17761), .B(n17760), .Z(n17762) );
  XNOR U18046 ( .A(n17763), .B(n17762), .Z(n17764) );
  XNOR U18047 ( .A(n17765), .B(n17764), .Z(n17766) );
  XNOR U18048 ( .A(n17767), .B(n17766), .Z(n17768) );
  XNOR U18049 ( .A(n17769), .B(n17768), .Z(n17785) );
  NAND U18050 ( .A(n17771), .B(n17770), .Z(n17775) );
  ANDN U18051 ( .B(n17773), .A(n17772), .Z(n17774) );
  ANDN U18052 ( .B(n17775), .A(n17774), .Z(n17783) );
  ANDN U18053 ( .B(n17777), .A(n17776), .Z(n17781) );
  ANDN U18054 ( .B(n17779), .A(n17778), .Z(n17780) );
  OR U18055 ( .A(n17781), .B(n17780), .Z(n17782) );
  XNOR U18056 ( .A(n17783), .B(n17782), .Z(n17784) );
  XNOR U18057 ( .A(n17785), .B(n17784), .Z(n17786) );
  XNOR U18058 ( .A(n17787), .B(n17786), .Z(n17788) );
  XNOR U18059 ( .A(n17789), .B(n17788), .Z(n17790) );
  XNOR U18060 ( .A(n17791), .B(n17790), .Z(n17792) );
  XNOR U18061 ( .A(n17793), .B(n17792), .Z(n17794) );
  NAND U18062 ( .A(n17797), .B(n17796), .Z(n17801) );
  AND U18063 ( .A(n17799), .B(n17798), .Z(n17800) );
  ANDN U18064 ( .B(n17801), .A(n17800), .Z(n17809) );
  AND U18065 ( .A(n17803), .B(n17802), .Z(n17807) );
  ANDN U18066 ( .B(n17805), .A(n17804), .Z(n17806) );
  OR U18067 ( .A(n17807), .B(n17806), .Z(n17808) );
  XNOR U18068 ( .A(n17809), .B(n17808), .Z(n17810) );
  NAND U18069 ( .A(n17812), .B(n17811), .Z(n17816) );
  ANDN U18070 ( .B(n17814), .A(n17813), .Z(n17815) );
  AND U18071 ( .A(n17818), .B(n17817), .Z(n17822) );
  AND U18072 ( .A(n17820), .B(n17819), .Z(n17821) );
  NAND U18073 ( .A(y[184]), .B(x[192]), .Z(n17970) );
  NAND U18074 ( .A(y[64]), .B(x[168]), .Z(n17825) );
  XOR U18075 ( .A(n17970), .B(n17825), .Z(n17826) );
  AND U18076 ( .A(y[24]), .B(x[160]), .Z(n17833) );
  AND U18077 ( .A(y[104]), .B(x[176]), .Z(n17830) );
  XOR U18078 ( .A(n17833), .B(n17830), .Z(n17829) );
  AND U18079 ( .A(y[144]), .B(x[184]), .Z(n17828) );
  XNOR U18080 ( .A(n17829), .B(n17828), .Z(n17827) );
  XNOR U18081 ( .A(n17826), .B(n17827), .Z(o[184]) );
  AND U18082 ( .A(x[161]), .B(y[24]), .Z(n17824) );
  NAND U18083 ( .A(x[160]), .B(y[25]), .Z(n17823) );
  XNOR U18084 ( .A(n17824), .B(n17823), .Z(n17834) );
  NAND U18085 ( .A(y[64]), .B(x[169]), .Z(n17835) );
  XOR U18086 ( .A(n17834), .B(n17835), .Z(n17851) );
  AND U18087 ( .A(y[184]), .B(x[193]), .Z(n18059) );
  NAND U18088 ( .A(y[105]), .B(x[176]), .Z(n17838) );
  XNOR U18089 ( .A(n18059), .B(n17838), .Z(n17839) );
  AND U18090 ( .A(y[185]), .B(x[192]), .Z(n17862) );
  NAND U18091 ( .A(y[104]), .B(x[177]), .Z(n17861) );
  XOR U18092 ( .A(n17862), .B(n17861), .Z(n17840) );
  XOR U18093 ( .A(n17839), .B(n17840), .Z(n17850) );
  AND U18094 ( .A(y[65]), .B(x[168]), .Z(n18085) );
  AND U18095 ( .A(y[145]), .B(x[184]), .Z(n17855) );
  XOR U18096 ( .A(n18085), .B(n17855), .Z(n17857) );
  AND U18097 ( .A(y[144]), .B(x[185]), .Z(n17856) );
  XNOR U18098 ( .A(n17857), .B(n17856), .Z(n17849) );
  XOR U18099 ( .A(n17850), .B(n17849), .Z(n17852) );
  XOR U18100 ( .A(n17851), .B(n17852), .Z(n17846) );
  NAND U18101 ( .A(n17829), .B(n17828), .Z(n17832) );
  AND U18102 ( .A(n17833), .B(n17830), .Z(n17831) );
  ANDN U18103 ( .B(n17832), .A(n17831), .Z(n17843) );
  XNOR U18104 ( .A(n17844), .B(n17843), .Z(n17845) );
  XNOR U18105 ( .A(n17846), .B(n17845), .Z(o[185]) );
  AND U18106 ( .A(y[25]), .B(x[161]), .Z(n17892) );
  NAND U18107 ( .A(n17892), .B(n17833), .Z(n17837) );
  NANDN U18108 ( .A(n17835), .B(n17834), .Z(n17836) );
  NAND U18109 ( .A(n17837), .B(n17836), .Z(n17904) );
  NANDN U18110 ( .A(n17838), .B(n18059), .Z(n17842) );
  NANDN U18111 ( .A(n17840), .B(n17839), .Z(n17841) );
  NAND U18112 ( .A(n17842), .B(n17841), .Z(n17902) );
  AND U18113 ( .A(y[146]), .B(x[184]), .Z(n17908) );
  NAND U18114 ( .A(y[26]), .B(x[160]), .Z(n17909) );
  XNOR U18115 ( .A(n17908), .B(n17909), .Z(n17911) );
  AND U18116 ( .A(y[64]), .B(x[170]), .Z(n17910) );
  XOR U18117 ( .A(n17911), .B(n17910), .Z(n17903) );
  XOR U18118 ( .A(n17902), .B(n17903), .Z(n17905) );
  XNOR U18119 ( .A(n17904), .B(n17905), .Z(n17864) );
  NANDN U18120 ( .A(n17844), .B(n17843), .Z(n17848) );
  NAND U18121 ( .A(n17846), .B(n17845), .Z(n17847) );
  NAND U18122 ( .A(n17848), .B(n17847), .Z(n17863) );
  XOR U18123 ( .A(n17864), .B(n17863), .Z(n17866) );
  NAND U18124 ( .A(n17850), .B(n17849), .Z(n17854) );
  NAND U18125 ( .A(n17852), .B(n17851), .Z(n17853) );
  AND U18126 ( .A(n17854), .B(n17853), .Z(n17872) );
  AND U18127 ( .A(y[24]), .B(x[162]), .Z(n17890) );
  AND U18128 ( .A(y[106]), .B(x[176]), .Z(n17889) );
  XOR U18129 ( .A(n17890), .B(n17889), .Z(n17891) );
  XOR U18130 ( .A(n17892), .B(n17891), .Z(n17917) );
  AND U18131 ( .A(y[144]), .B(x[186]), .Z(n17916) );
  XOR U18132 ( .A(n17917), .B(n17916), .Z(n17919) );
  AND U18133 ( .A(y[104]), .B(x[178]), .Z(n17987) );
  AND U18134 ( .A(y[186]), .B(x[192]), .Z(n17881) );
  XOR U18135 ( .A(n17987), .B(n17881), .Z(n17883) );
  AND U18136 ( .A(y[105]), .B(x[177]), .Z(n17882) );
  XOR U18137 ( .A(n17883), .B(n17882), .Z(n17918) );
  XOR U18138 ( .A(n17919), .B(n17918), .Z(n17869) );
  AND U18139 ( .A(n18085), .B(n17855), .Z(n17859) );
  NAND U18140 ( .A(n17857), .B(n17856), .Z(n17858) );
  NANDN U18141 ( .A(n17859), .B(n17858), .Z(n17877) );
  AND U18142 ( .A(x[193]), .B(y[185]), .Z(n17949) );
  NAND U18143 ( .A(x[194]), .B(y[184]), .Z(n17860) );
  XNOR U18144 ( .A(n17949), .B(n17860), .Z(n17915) );
  ANDN U18145 ( .B(n17862), .A(n17861), .Z(n17914) );
  XOR U18146 ( .A(n17915), .B(n17914), .Z(n17876) );
  AND U18147 ( .A(y[145]), .B(x[185]), .Z(n17895) );
  NAND U18148 ( .A(y[65]), .B(x[169]), .Z(n17896) );
  XNOR U18149 ( .A(n17895), .B(n17896), .Z(n17897) );
  NAND U18150 ( .A(y[66]), .B(x[168]), .Z(n17898) );
  XNOR U18151 ( .A(n17897), .B(n17898), .Z(n17875) );
  XOR U18152 ( .A(n17876), .B(n17875), .Z(n17878) );
  XOR U18153 ( .A(n17877), .B(n17878), .Z(n17870) );
  XOR U18154 ( .A(n17869), .B(n17870), .Z(n17871) );
  XNOR U18155 ( .A(n17872), .B(n17871), .Z(n17865) );
  XNOR U18156 ( .A(n17866), .B(n17865), .Z(o[186]) );
  NAND U18157 ( .A(n17864), .B(n17863), .Z(n17868) );
  NAND U18158 ( .A(n17866), .B(n17865), .Z(n17867) );
  AND U18159 ( .A(n17868), .B(n17867), .Z(n17923) );
  NAND U18160 ( .A(n17870), .B(n17869), .Z(n17874) );
  NAND U18161 ( .A(n17872), .B(n17871), .Z(n17873) );
  NAND U18162 ( .A(n17874), .B(n17873), .Z(n17928) );
  NAND U18163 ( .A(n17876), .B(n17875), .Z(n17880) );
  NAND U18164 ( .A(n17878), .B(n17877), .Z(n17879) );
  NAND U18165 ( .A(n17880), .B(n17879), .Z(n17926) );
  AND U18166 ( .A(y[26]), .B(x[161]), .Z(n17966) );
  AND U18167 ( .A(y[25]), .B(x[162]), .Z(n17965) );
  NAND U18168 ( .A(y[146]), .B(x[185]), .Z(n17964) );
  XOR U18169 ( .A(n17965), .B(n17964), .Z(n17967) );
  XOR U18170 ( .A(n17966), .B(n17967), .Z(n17984) );
  NAND U18171 ( .A(n17987), .B(n17881), .Z(n17885) );
  AND U18172 ( .A(n17883), .B(n17882), .Z(n17884) );
  ANDN U18173 ( .B(n17885), .A(n17884), .Z(n17982) );
  AND U18174 ( .A(x[195]), .B(y[184]), .Z(n17887) );
  NAND U18175 ( .A(x[192]), .B(y[187]), .Z(n17886) );
  XNOR U18176 ( .A(n17887), .B(n17886), .Z(n17971) );
  AND U18177 ( .A(x[194]), .B(y[185]), .Z(n18055) );
  NAND U18178 ( .A(x[193]), .B(y[186]), .Z(n17888) );
  XOR U18179 ( .A(n18055), .B(n17888), .Z(n17972) );
  XNOR U18180 ( .A(n17971), .B(n17972), .Z(n17981) );
  XNOR U18181 ( .A(n17982), .B(n17981), .Z(n17983) );
  XNOR U18182 ( .A(n17984), .B(n17983), .Z(n17940) );
  NAND U18183 ( .A(n17890), .B(n17889), .Z(n17894) );
  NAND U18184 ( .A(n17892), .B(n17891), .Z(n17893) );
  NAND U18185 ( .A(n17894), .B(n17893), .Z(n17938) );
  NANDN U18186 ( .A(n17896), .B(n17895), .Z(n17900) );
  NANDN U18187 ( .A(n17898), .B(n17897), .Z(n17899) );
  AND U18188 ( .A(n17900), .B(n17899), .Z(n17977) );
  AND U18189 ( .A(y[147]), .B(x[184]), .Z(n18006) );
  AND U18190 ( .A(y[107]), .B(x[176]), .Z(n18005) );
  NAND U18191 ( .A(y[24]), .B(x[163]), .Z(n18004) );
  XOR U18192 ( .A(n18005), .B(n18004), .Z(n18007) );
  XOR U18193 ( .A(n18006), .B(n18007), .Z(n17976) );
  AND U18194 ( .A(x[178]), .B(y[105]), .Z(n18038) );
  NAND U18195 ( .A(x[179]), .B(y[104]), .Z(n17901) );
  XNOR U18196 ( .A(n18038), .B(n17901), .Z(n17989) );
  NAND U18197 ( .A(y[106]), .B(x[177]), .Z(n17990) );
  XOR U18198 ( .A(n17976), .B(n17975), .Z(n17978) );
  XOR U18199 ( .A(n17977), .B(n17978), .Z(n17939) );
  XOR U18200 ( .A(n17938), .B(n17939), .Z(n17941) );
  XOR U18201 ( .A(n17940), .B(n17941), .Z(n17927) );
  XOR U18202 ( .A(n17926), .B(n17927), .Z(n17929) );
  XOR U18203 ( .A(n17928), .B(n17929), .Z(n17922) );
  XOR U18204 ( .A(n17923), .B(n17922), .Z(n17925) );
  NAND U18205 ( .A(n17903), .B(n17902), .Z(n17907) );
  NAND U18206 ( .A(n17905), .B(n17904), .Z(n17906) );
  AND U18207 ( .A(n17907), .B(n17906), .Z(n17935) );
  NANDN U18208 ( .A(n17909), .B(n17908), .Z(n17913) );
  NAND U18209 ( .A(n17911), .B(n17910), .Z(n17912) );
  AND U18210 ( .A(n17913), .B(n17912), .Z(n17945) );
  XNOR U18211 ( .A(n17945), .B(n17944), .Z(n17947) );
  AND U18212 ( .A(y[64]), .B(x[171]), .Z(n17997) );
  AND U18213 ( .A(y[27]), .B(x[160]), .Z(n17996) );
  NAND U18214 ( .A(y[145]), .B(x[186]), .Z(n17995) );
  XOR U18215 ( .A(n17996), .B(n17995), .Z(n17998) );
  XOR U18216 ( .A(n17997), .B(n17998), .Z(n17959) );
  AND U18217 ( .A(y[67]), .B(x[168]), .Z(n17952) );
  AND U18218 ( .A(y[65]), .B(x[170]), .Z(n17951) );
  NAND U18219 ( .A(y[144]), .B(x[187]), .Z(n17950) );
  XOR U18220 ( .A(n17951), .B(n17950), .Z(n17953) );
  XOR U18221 ( .A(n17952), .B(n17953), .Z(n17957) );
  AND U18222 ( .A(y[66]), .B(x[169]), .Z(n17956) );
  XNOR U18223 ( .A(n17947), .B(n17946), .Z(n17933) );
  NAND U18224 ( .A(n17917), .B(n17916), .Z(n17921) );
  NAND U18225 ( .A(n17919), .B(n17918), .Z(n17920) );
  AND U18226 ( .A(n17921), .B(n17920), .Z(n17932) );
  XOR U18227 ( .A(n17933), .B(n17932), .Z(n17934) );
  XNOR U18228 ( .A(n17935), .B(n17934), .Z(n17924) );
  XOR U18229 ( .A(n17925), .B(n17924), .Z(o[187]) );
  NAND U18230 ( .A(n17927), .B(n17926), .Z(n17931) );
  NAND U18231 ( .A(n17929), .B(n17928), .Z(n17930) );
  AND U18232 ( .A(n17931), .B(n17930), .Z(n18016) );
  NAND U18233 ( .A(n17933), .B(n17932), .Z(n17937) );
  NAND U18234 ( .A(n17935), .B(n17934), .Z(n17936) );
  NAND U18235 ( .A(n17937), .B(n17936), .Z(n18014) );
  NAND U18236 ( .A(n17939), .B(n17938), .Z(n17943) );
  NAND U18237 ( .A(n17941), .B(n17940), .Z(n17942) );
  AND U18238 ( .A(n17943), .B(n17942), .Z(n18015) );
  XOR U18239 ( .A(n18014), .B(n18015), .Z(n18017) );
  XOR U18240 ( .A(n18016), .B(n18017), .Z(n18010) );
  XOR U18241 ( .A(n18011), .B(n18010), .Z(n18013) );
  AND U18242 ( .A(y[24]), .B(x[164]), .Z(n18073) );
  AND U18243 ( .A(y[146]), .B(x[186]), .Z(n18072) );
  NAND U18244 ( .A(y[108]), .B(x[176]), .Z(n18071) );
  XOR U18245 ( .A(n18072), .B(n18071), .Z(n18074) );
  XOR U18246 ( .A(n18073), .B(n18074), .Z(n18027) );
  AND U18247 ( .A(y[186]), .B(x[194]), .Z(n17948) );
  AND U18248 ( .A(n17949), .B(n17948), .Z(n18066) );
  NAND U18249 ( .A(y[104]), .B(x[180]), .Z(n18193) );
  IV U18250 ( .A(n18193), .Z(n18064) );
  NAND U18251 ( .A(y[188]), .B(x[192]), .Z(n18233) );
  XNOR U18252 ( .A(n18064), .B(n18233), .Z(n18065) );
  XOR U18253 ( .A(n18066), .B(n18065), .Z(n18026) );
  XNOR U18254 ( .A(n18027), .B(n18026), .Z(n18029) );
  NANDN U18255 ( .A(n17951), .B(n17950), .Z(n17955) );
  OR U18256 ( .A(n17953), .B(n17952), .Z(n17954) );
  AND U18257 ( .A(n17955), .B(n17954), .Z(n18028) );
  XOR U18258 ( .A(n18029), .B(n18028), .Z(n18120) );
  NANDN U18259 ( .A(n17957), .B(n17956), .Z(n17961) );
  NANDN U18260 ( .A(n17959), .B(n17958), .Z(n17960) );
  AND U18261 ( .A(n17961), .B(n17960), .Z(n18119) );
  AND U18262 ( .A(y[66]), .B(x[170]), .Z(n18178) );
  AND U18263 ( .A(x[168]), .B(y[68]), .Z(n17963) );
  NAND U18264 ( .A(x[171]), .B(y[65]), .Z(n17962) );
  XOR U18265 ( .A(n17963), .B(n17962), .Z(n18086) );
  XNOR U18266 ( .A(n18178), .B(n18086), .Z(n18089) );
  NAND U18267 ( .A(y[67]), .B(x[169]), .Z(n18090) );
  XNOR U18268 ( .A(n18089), .B(n18090), .Z(n18092) );
  AND U18269 ( .A(y[144]), .B(x[188]), .Z(n18043) );
  NAND U18270 ( .A(y[27]), .B(x[161]), .Z(n18044) );
  XNOR U18271 ( .A(n18043), .B(n18044), .Z(n18045) );
  NAND U18272 ( .A(y[28]), .B(x[160]), .Z(n18046) );
  XNOR U18273 ( .A(n18045), .B(n18046), .Z(n18091) );
  XOR U18274 ( .A(n18092), .B(n18091), .Z(n18104) );
  NANDN U18275 ( .A(n17965), .B(n17964), .Z(n17969) );
  OR U18276 ( .A(n17967), .B(n17966), .Z(n17968) );
  AND U18277 ( .A(n17969), .B(n17968), .Z(n18102) );
  AND U18278 ( .A(y[187]), .B(x[195]), .Z(n18313) );
  NANDN U18279 ( .A(n17970), .B(n18313), .Z(n17974) );
  NANDN U18280 ( .A(n17972), .B(n17971), .Z(n17973) );
  AND U18281 ( .A(n17974), .B(n17973), .Z(n18101) );
  XNOR U18282 ( .A(n18102), .B(n18101), .Z(n18103) );
  XNOR U18283 ( .A(n18104), .B(n18103), .Z(n18121) );
  XNOR U18284 ( .A(n18122), .B(n18121), .Z(n18020) );
  XNOR U18285 ( .A(n18021), .B(n18020), .Z(n18023) );
  NANDN U18286 ( .A(n17976), .B(n17975), .Z(n17980) );
  OR U18287 ( .A(n17978), .B(n17977), .Z(n17979) );
  AND U18288 ( .A(n17980), .B(n17979), .Z(n18108) );
  NANDN U18289 ( .A(n17982), .B(n17981), .Z(n17986) );
  NANDN U18290 ( .A(n17984), .B(n17983), .Z(n17985) );
  NAND U18291 ( .A(n17986), .B(n17985), .Z(n18107) );
  AND U18292 ( .A(y[105]), .B(x[179]), .Z(n17988) );
  NAND U18293 ( .A(n17988), .B(n17987), .Z(n17992) );
  NANDN U18294 ( .A(n17990), .B(n17989), .Z(n17991) );
  AND U18295 ( .A(n17992), .B(n17991), .Z(n18114) );
  AND U18296 ( .A(y[64]), .B(x[172]), .Z(n18049) );
  NAND U18297 ( .A(y[148]), .B(x[184]), .Z(n18050) );
  XNOR U18298 ( .A(n18049), .B(n18050), .Z(n18051) );
  NAND U18299 ( .A(y[147]), .B(x[185]), .Z(n18052) );
  XNOR U18300 ( .A(n18051), .B(n18052), .Z(n18095) );
  AND U18301 ( .A(x[178]), .B(y[106]), .Z(n17994) );
  NAND U18302 ( .A(x[179]), .B(y[105]), .Z(n17993) );
  XNOR U18303 ( .A(n17994), .B(n17993), .Z(n18039) );
  NAND U18304 ( .A(y[107]), .B(x[177]), .Z(n18040) );
  XOR U18305 ( .A(n18039), .B(n18040), .Z(n18096) );
  XNOR U18306 ( .A(n18095), .B(n18096), .Z(n18097) );
  NANDN U18307 ( .A(n17996), .B(n17995), .Z(n18000) );
  OR U18308 ( .A(n17998), .B(n17997), .Z(n17999) );
  NAND U18309 ( .A(n18000), .B(n17999), .Z(n18098) );
  XNOR U18310 ( .A(n18097), .B(n18098), .Z(n18113) );
  NAND U18311 ( .A(y[26]), .B(x[162]), .Z(n18081) );
  NAND U18312 ( .A(y[145]), .B(x[187]), .Z(n18080) );
  NAND U18313 ( .A(y[25]), .B(x[163]), .Z(n18079) );
  XNOR U18314 ( .A(n18080), .B(n18079), .Z(n18082) );
  AND U18315 ( .A(x[196]), .B(y[184]), .Z(n18002) );
  NAND U18316 ( .A(x[193]), .B(y[187]), .Z(n18001) );
  XNOR U18317 ( .A(n18002), .B(n18001), .Z(n18060) );
  AND U18318 ( .A(y[185]), .B(x[195]), .Z(n18201) );
  NAND U18319 ( .A(x[194]), .B(y[186]), .Z(n18003) );
  XOR U18320 ( .A(n18201), .B(n18003), .Z(n18061) );
  XNOR U18321 ( .A(n18060), .B(n18061), .Z(n18032) );
  XOR U18322 ( .A(n18033), .B(n18032), .Z(n18034) );
  NANDN U18323 ( .A(n18005), .B(n18004), .Z(n18009) );
  OR U18324 ( .A(n18007), .B(n18006), .Z(n18008) );
  NAND U18325 ( .A(n18009), .B(n18008), .Z(n18035) );
  XOR U18326 ( .A(n18034), .B(n18035), .Z(n18116) );
  XOR U18327 ( .A(n18110), .B(n18109), .Z(n18022) );
  XNOR U18328 ( .A(n18023), .B(n18022), .Z(n18012) );
  XNOR U18329 ( .A(n18013), .B(n18012), .Z(o[188]) );
  NAND U18330 ( .A(n18015), .B(n18014), .Z(n18019) );
  NAND U18331 ( .A(n18017), .B(n18016), .Z(n18018) );
  NAND U18332 ( .A(n18019), .B(n18018), .Z(n18263) );
  XNOR U18333 ( .A(n18262), .B(n18263), .Z(n18265) );
  NANDN U18334 ( .A(n18021), .B(n18020), .Z(n18025) );
  NAND U18335 ( .A(n18023), .B(n18022), .Z(n18024) );
  AND U18336 ( .A(n18025), .B(n18024), .Z(n18126) );
  NANDN U18337 ( .A(n18027), .B(n18026), .Z(n18031) );
  NAND U18338 ( .A(n18029), .B(n18028), .Z(n18030) );
  AND U18339 ( .A(n18031), .B(n18030), .Z(n18142) );
  NAND U18340 ( .A(n18033), .B(n18032), .Z(n18037) );
  NANDN U18341 ( .A(n18035), .B(n18034), .Z(n18036) );
  NAND U18342 ( .A(n18037), .B(n18036), .Z(n18141) );
  XNOR U18343 ( .A(n18142), .B(n18141), .Z(n18144) );
  AND U18344 ( .A(y[106]), .B(x[179]), .Z(n18194) );
  NAND U18345 ( .A(n18038), .B(n18194), .Z(n18042) );
  NANDN U18346 ( .A(n18040), .B(n18039), .Z(n18041) );
  NAND U18347 ( .A(n18042), .B(n18041), .Z(n18202) );
  NANDN U18348 ( .A(n18044), .B(n18043), .Z(n18048) );
  NANDN U18349 ( .A(n18046), .B(n18045), .Z(n18047) );
  AND U18350 ( .A(n18048), .B(n18047), .Z(n18162) );
  AND U18351 ( .A(y[149]), .B(x[184]), .Z(n18488) );
  AND U18352 ( .A(y[64]), .B(x[173]), .Z(n18184) );
  AND U18353 ( .A(y[107]), .B(x[178]), .Z(n18183) );
  XOR U18354 ( .A(n18184), .B(n18183), .Z(n18185) );
  XOR U18355 ( .A(n18488), .B(n18185), .Z(n18159) );
  AND U18356 ( .A(y[25]), .B(x[164]), .Z(n18452) );
  AND U18357 ( .A(y[145]), .B(x[188]), .Z(n18189) );
  AND U18358 ( .A(y[24]), .B(x[165]), .Z(n18188) );
  XOR U18359 ( .A(n18189), .B(n18188), .Z(n18190) );
  XNOR U18360 ( .A(n18452), .B(n18190), .Z(n18160) );
  XNOR U18361 ( .A(n18159), .B(n18160), .Z(n18161) );
  XNOR U18362 ( .A(n18162), .B(n18161), .Z(n18203) );
  XOR U18363 ( .A(n18202), .B(n18203), .Z(n18204) );
  NANDN U18364 ( .A(n18050), .B(n18049), .Z(n18054) );
  NANDN U18365 ( .A(n18052), .B(n18051), .Z(n18053) );
  NAND U18366 ( .A(n18054), .B(n18053), .Z(n18258) );
  AND U18367 ( .A(y[186]), .B(x[195]), .Z(n18056) );
  AND U18368 ( .A(n18056), .B(n18055), .Z(n18235) );
  AND U18369 ( .A(x[192]), .B(y[189]), .Z(n18058) );
  AND U18370 ( .A(x[193]), .B(y[188]), .Z(n18057) );
  XOR U18371 ( .A(n18058), .B(n18057), .Z(n18234) );
  XOR U18372 ( .A(n18235), .B(n18234), .Z(n18257) );
  AND U18373 ( .A(y[69]), .B(x[168]), .Z(n18247) );
  AND U18374 ( .A(y[28]), .B(x[161]), .Z(n18246) );
  XOR U18375 ( .A(n18247), .B(n18246), .Z(n18249) );
  AND U18376 ( .A(y[65]), .B(x[172]), .Z(n18248) );
  XOR U18377 ( .A(n18249), .B(n18248), .Z(n18256) );
  XOR U18378 ( .A(n18257), .B(n18256), .Z(n18259) );
  XNOR U18379 ( .A(n18258), .B(n18259), .Z(n18205) );
  XOR U18380 ( .A(n18144), .B(n18143), .Z(n18132) );
  AND U18381 ( .A(y[187]), .B(x[196]), .Z(n18466) );
  NAND U18382 ( .A(n18466), .B(n18059), .Z(n18063) );
  NANDN U18383 ( .A(n18061), .B(n18060), .Z(n18062) );
  AND U18384 ( .A(n18063), .B(n18062), .Z(n18154) );
  NANDN U18385 ( .A(n18064), .B(n18233), .Z(n18068) );
  NANDN U18386 ( .A(n18066), .B(n18065), .Z(n18067) );
  AND U18387 ( .A(n18068), .B(n18067), .Z(n18153) );
  XNOR U18388 ( .A(n18154), .B(n18153), .Z(n18156) );
  AND U18389 ( .A(y[187]), .B(x[194]), .Z(n18165) );
  NAND U18390 ( .A(y[184]), .B(x[197]), .Z(n18166) );
  AND U18391 ( .A(y[185]), .B(x[196]), .Z(n18448) );
  NAND U18392 ( .A(x[195]), .B(y[186]), .Z(n18069) );
  XOR U18393 ( .A(n18448), .B(n18069), .Z(n18168) );
  AND U18394 ( .A(y[66]), .B(x[171]), .Z(n18386) );
  NAND U18395 ( .A(x[170]), .B(y[67]), .Z(n18070) );
  XNOR U18396 ( .A(n18386), .B(n18070), .Z(n18179) );
  NAND U18397 ( .A(y[68]), .B(x[169]), .Z(n18180) );
  XOR U18398 ( .A(n18146), .B(n18145), .Z(n18147) );
  NANDN U18399 ( .A(n18072), .B(n18071), .Z(n18076) );
  OR U18400 ( .A(n18074), .B(n18073), .Z(n18075) );
  NAND U18401 ( .A(n18076), .B(n18075), .Z(n18148) );
  XNOR U18402 ( .A(n18147), .B(n18148), .Z(n18155) );
  XOR U18403 ( .A(n18156), .B(n18155), .Z(n18216) );
  AND U18404 ( .A(x[180]), .B(y[105]), .Z(n18078) );
  NAND U18405 ( .A(x[181]), .B(y[104]), .Z(n18077) );
  XOR U18406 ( .A(n18078), .B(n18077), .Z(n18195) );
  XNOR U18407 ( .A(n18194), .B(n18195), .Z(n18238) );
  AND U18408 ( .A(y[144]), .B(x[189]), .Z(n18171) );
  NAND U18409 ( .A(y[26]), .B(x[163]), .Z(n18172) );
  XNOR U18410 ( .A(n18171), .B(n18172), .Z(n18173) );
  NAND U18411 ( .A(y[27]), .B(x[162]), .Z(n18174) );
  XOR U18412 ( .A(n18173), .B(n18174), .Z(n18239) );
  NAND U18413 ( .A(n18080), .B(n18079), .Z(n18084) );
  NANDN U18414 ( .A(n18082), .B(n18081), .Z(n18083) );
  AND U18415 ( .A(n18084), .B(n18083), .Z(n18240) );
  XOR U18416 ( .A(n18241), .B(n18240), .Z(n18215) );
  AND U18417 ( .A(y[68]), .B(x[171]), .Z(n18465) );
  NAND U18418 ( .A(n18465), .B(n18085), .Z(n18088) );
  NANDN U18419 ( .A(n18086), .B(n18178), .Z(n18087) );
  AND U18420 ( .A(n18088), .B(n18087), .Z(n18152) );
  AND U18421 ( .A(y[146]), .B(x[187]), .Z(n18220) );
  AND U18422 ( .A(y[108]), .B(x[177]), .Z(n18434) );
  XOR U18423 ( .A(n18220), .B(n18434), .Z(n18222) );
  AND U18424 ( .A(y[109]), .B(x[176]), .Z(n18221) );
  XOR U18425 ( .A(n18222), .B(n18221), .Z(n18150) );
  AND U18426 ( .A(y[29]), .B(x[160]), .Z(n18226) );
  AND U18427 ( .A(y[148]), .B(x[185]), .Z(n18225) );
  XOR U18428 ( .A(n18226), .B(n18225), .Z(n18228) );
  AND U18429 ( .A(y[147]), .B(x[186]), .Z(n18227) );
  XOR U18430 ( .A(n18228), .B(n18227), .Z(n18149) );
  XOR U18431 ( .A(n18150), .B(n18149), .Z(n18151) );
  XOR U18432 ( .A(n18152), .B(n18151), .Z(n18214) );
  XOR U18433 ( .A(n18215), .B(n18214), .Z(n18217) );
  XOR U18434 ( .A(n18216), .B(n18217), .Z(n18130) );
  NANDN U18435 ( .A(n18090), .B(n18089), .Z(n18094) );
  NAND U18436 ( .A(n18092), .B(n18091), .Z(n18093) );
  AND U18437 ( .A(n18094), .B(n18093), .Z(n18209) );
  NANDN U18438 ( .A(n18096), .B(n18095), .Z(n18100) );
  NANDN U18439 ( .A(n18098), .B(n18097), .Z(n18099) );
  NAND U18440 ( .A(n18100), .B(n18099), .Z(n18208) );
  XNOR U18441 ( .A(n18209), .B(n18208), .Z(n18210) );
  NANDN U18442 ( .A(n18102), .B(n18101), .Z(n18106) );
  NANDN U18443 ( .A(n18104), .B(n18103), .Z(n18105) );
  NAND U18444 ( .A(n18106), .B(n18105), .Z(n18211) );
  XNOR U18445 ( .A(n18210), .B(n18211), .Z(n18129) );
  XOR U18446 ( .A(n18132), .B(n18131), .Z(n18125) );
  XNOR U18447 ( .A(n18126), .B(n18125), .Z(n18128) );
  NANDN U18448 ( .A(n18108), .B(n18107), .Z(n18112) );
  NAND U18449 ( .A(n18110), .B(n18109), .Z(n18111) );
  AND U18450 ( .A(n18112), .B(n18111), .Z(n18138) );
  NANDN U18451 ( .A(n18114), .B(n18113), .Z(n18118) );
  NANDN U18452 ( .A(n18116), .B(n18115), .Z(n18117) );
  AND U18453 ( .A(n18118), .B(n18117), .Z(n18136) );
  NANDN U18454 ( .A(n18120), .B(n18119), .Z(n18124) );
  NAND U18455 ( .A(n18122), .B(n18121), .Z(n18123) );
  AND U18456 ( .A(n18124), .B(n18123), .Z(n18135) );
  XOR U18457 ( .A(n18128), .B(n18127), .Z(n18264) );
  XOR U18458 ( .A(n18265), .B(n18264), .Z(o[189]) );
  NANDN U18459 ( .A(n18130), .B(n18129), .Z(n18134) );
  NAND U18460 ( .A(n18132), .B(n18131), .Z(n18133) );
  AND U18461 ( .A(n18134), .B(n18133), .Z(n18559) );
  NANDN U18462 ( .A(n18136), .B(n18135), .Z(n18140) );
  NANDN U18463 ( .A(n18138), .B(n18137), .Z(n18139) );
  NAND U18464 ( .A(n18140), .B(n18139), .Z(n18560) );
  NANDN U18465 ( .A(n18154), .B(n18153), .Z(n18158) );
  NAND U18466 ( .A(n18156), .B(n18155), .Z(n18157) );
  AND U18467 ( .A(n18158), .B(n18157), .Z(n18276) );
  XOR U18468 ( .A(n18277), .B(n18276), .Z(n18274) );
  XOR U18469 ( .A(n18275), .B(n18274), .Z(n18271) );
  NANDN U18470 ( .A(n18160), .B(n18159), .Z(n18164) );
  NANDN U18471 ( .A(n18162), .B(n18161), .Z(n18163) );
  NAND U18472 ( .A(n18164), .B(n18163), .Z(n18282) );
  NANDN U18473 ( .A(n18166), .B(n18165), .Z(n18170) );
  NANDN U18474 ( .A(n18168), .B(n18167), .Z(n18169) );
  NAND U18475 ( .A(n18170), .B(n18169), .Z(n18300) );
  NANDN U18476 ( .A(n18172), .B(n18171), .Z(n18176) );
  NANDN U18477 ( .A(n18174), .B(n18173), .Z(n18175) );
  NAND U18478 ( .A(n18176), .B(n18175), .Z(n18303) );
  AND U18479 ( .A(y[67]), .B(x[171]), .Z(n18177) );
  NAND U18480 ( .A(n18178), .B(n18177), .Z(n18182) );
  NANDN U18481 ( .A(n18180), .B(n18179), .Z(n18181) );
  AND U18482 ( .A(n18182), .B(n18181), .Z(n18514) );
  AND U18483 ( .A(y[147]), .B(x[187]), .Z(n18406) );
  AND U18484 ( .A(y[107]), .B(x[179]), .Z(n18405) );
  XOR U18485 ( .A(n18406), .B(n18405), .Z(n18404) );
  AND U18486 ( .A(y[27]), .B(x[163]), .Z(n18403) );
  XOR U18487 ( .A(n18404), .B(n18403), .Z(n18516) );
  AND U18488 ( .A(y[148]), .B(x[186]), .Z(n18480) );
  AND U18489 ( .A(y[106]), .B(x[180]), .Z(n18479) );
  XOR U18490 ( .A(n18480), .B(n18479), .Z(n18478) );
  AND U18491 ( .A(y[28]), .B(x[162]), .Z(n18477) );
  XNOR U18492 ( .A(n18478), .B(n18477), .Z(n18515) );
  XNOR U18493 ( .A(n18514), .B(n18513), .Z(n18302) );
  XOR U18494 ( .A(n18303), .B(n18302), .Z(n18301) );
  XOR U18495 ( .A(n18300), .B(n18301), .Z(n18283) );
  XOR U18496 ( .A(n18282), .B(n18283), .Z(n18281) );
  NAND U18497 ( .A(n18184), .B(n18183), .Z(n18187) );
  NAND U18498 ( .A(n18488), .B(n18185), .Z(n18186) );
  NAND U18499 ( .A(n18187), .B(n18186), .Z(n18422) );
  NAND U18500 ( .A(n18189), .B(n18188), .Z(n18192) );
  NAND U18501 ( .A(n18452), .B(n18190), .Z(n18191) );
  NAND U18502 ( .A(n18192), .B(n18191), .Z(n18421) );
  XOR U18503 ( .A(n18422), .B(n18421), .Z(n18420) );
  AND U18504 ( .A(y[105]), .B(x[181]), .Z(n18440) );
  NANDN U18505 ( .A(n18193), .B(n18440), .Z(n18197) );
  NANDN U18506 ( .A(n18195), .B(n18194), .Z(n18196) );
  AND U18507 ( .A(n18197), .B(n18196), .Z(n18426) );
  AND U18508 ( .A(x[165]), .B(y[25]), .Z(n18199) );
  NAND U18509 ( .A(x[164]), .B(y[26]), .Z(n18198) );
  XNOR U18510 ( .A(n18199), .B(n18198), .Z(n18450) );
  AND U18511 ( .A(y[144]), .B(x[190]), .Z(n18449) );
  XOR U18512 ( .A(n18450), .B(n18449), .Z(n18428) );
  AND U18513 ( .A(y[189]), .B(x[193]), .Z(n18390) );
  AND U18514 ( .A(y[186]), .B(x[196]), .Z(n18200) );
  AND U18515 ( .A(n18201), .B(n18200), .Z(n18392) );
  AND U18516 ( .A(y[188]), .B(x[194]), .Z(n18391) );
  XOR U18517 ( .A(n18392), .B(n18391), .Z(n18389) );
  XNOR U18518 ( .A(n18390), .B(n18389), .Z(n18427) );
  XNOR U18519 ( .A(n18426), .B(n18425), .Z(n18419) );
  XOR U18520 ( .A(n18420), .B(n18419), .Z(n18280) );
  XOR U18521 ( .A(n18281), .B(n18280), .Z(n18270) );
  XOR U18522 ( .A(n18269), .B(n18268), .Z(n18569) );
  NAND U18523 ( .A(n18203), .B(n18202), .Z(n18207) );
  NANDN U18524 ( .A(n18205), .B(n18204), .Z(n18206) );
  AND U18525 ( .A(n18207), .B(n18206), .Z(n18570) );
  XOR U18526 ( .A(n18569), .B(n18570), .Z(n18572) );
  NANDN U18527 ( .A(n18209), .B(n18208), .Z(n18213) );
  NANDN U18528 ( .A(n18211), .B(n18210), .Z(n18212) );
  AND U18529 ( .A(n18213), .B(n18212), .Z(n18534) );
  NANDN U18530 ( .A(n18215), .B(n18214), .Z(n18219) );
  OR U18531 ( .A(n18217), .B(n18216), .Z(n18218) );
  AND U18532 ( .A(n18219), .B(n18218), .Z(n18536) );
  NAND U18533 ( .A(n18220), .B(n18434), .Z(n18224) );
  NAND U18534 ( .A(n18222), .B(n18221), .Z(n18223) );
  AND U18535 ( .A(n18224), .B(n18223), .Z(n18293) );
  NAND U18536 ( .A(n18226), .B(n18225), .Z(n18230) );
  NAND U18537 ( .A(n18228), .B(n18227), .Z(n18229) );
  AND U18538 ( .A(n18230), .B(n18229), .Z(n18508) );
  AND U18539 ( .A(y[29]), .B(x[161]), .Z(n18474) );
  AND U18540 ( .A(y[64]), .B(x[174]), .Z(n18473) );
  XOR U18541 ( .A(n18474), .B(n18473), .Z(n18472) );
  AND U18542 ( .A(y[70]), .B(x[168]), .Z(n18471) );
  XOR U18543 ( .A(n18472), .B(n18471), .Z(n18510) );
  AND U18544 ( .A(x[197]), .B(y[185]), .Z(n18232) );
  NAND U18545 ( .A(x[196]), .B(y[186]), .Z(n18231) );
  XNOR U18546 ( .A(n18232), .B(n18231), .Z(n18315) );
  AND U18547 ( .A(y[184]), .B(x[198]), .Z(n18314) );
  XOR U18548 ( .A(n18315), .B(n18314), .Z(n18312) );
  XNOR U18549 ( .A(n18313), .B(n18312), .Z(n18509) );
  XOR U18550 ( .A(n18508), .B(n18507), .Z(n18295) );
  NANDN U18551 ( .A(n18233), .B(n18390), .Z(n18237) );
  NAND U18552 ( .A(n18235), .B(n18234), .Z(n18236) );
  NAND U18553 ( .A(n18237), .B(n18236), .Z(n18294) );
  XOR U18554 ( .A(n18293), .B(n18292), .Z(n18539) );
  NANDN U18555 ( .A(n18239), .B(n18238), .Z(n18243) );
  NAND U18556 ( .A(n18241), .B(n18240), .Z(n18242) );
  AND U18557 ( .A(n18243), .B(n18242), .Z(n18541) );
  AND U18558 ( .A(y[190]), .B(x[192]), .Z(n18439) );
  XOR U18559 ( .A(n18440), .B(n18439), .Z(n18438) );
  AND U18560 ( .A(y[104]), .B(x[182]), .Z(n18437) );
  XOR U18561 ( .A(n18438), .B(n18437), .Z(n18307) );
  AND U18562 ( .A(y[110]), .B(x[176]), .Z(n18400) );
  AND U18563 ( .A(y[24]), .B(x[166]), .Z(n18399) );
  XOR U18564 ( .A(n18400), .B(n18399), .Z(n18398) );
  AND U18565 ( .A(y[145]), .B(x[189]), .Z(n18397) );
  XOR U18566 ( .A(n18398), .B(n18397), .Z(n18309) );
  AND U18567 ( .A(y[65]), .B(x[173]), .Z(n18494) );
  AND U18568 ( .A(y[68]), .B(x[170]), .Z(n18493) );
  XOR U18569 ( .A(n18494), .B(n18493), .Z(n18492) );
  AND U18570 ( .A(y[69]), .B(x[169]), .Z(n18491) );
  XOR U18571 ( .A(n18492), .B(n18491), .Z(n18384) );
  AND U18572 ( .A(x[172]), .B(y[66]), .Z(n18245) );
  NAND U18573 ( .A(x[171]), .B(y[67]), .Z(n18244) );
  XNOR U18574 ( .A(n18245), .B(n18244), .Z(n18383) );
  XOR U18575 ( .A(n18384), .B(n18383), .Z(n18308) );
  XOR U18576 ( .A(n18309), .B(n18308), .Z(n18306) );
  XOR U18577 ( .A(n18307), .B(n18306), .Z(n18289) );
  NAND U18578 ( .A(n18247), .B(n18246), .Z(n18251) );
  NAND U18579 ( .A(n18249), .B(n18248), .Z(n18250) );
  AND U18580 ( .A(n18251), .B(n18250), .Z(n18377) );
  AND U18581 ( .A(y[146]), .B(x[188]), .Z(n18432) );
  AND U18582 ( .A(x[177]), .B(y[109]), .Z(n18253) );
  AND U18583 ( .A(x[178]), .B(y[108]), .Z(n18252) );
  XOR U18584 ( .A(n18253), .B(n18252), .Z(n18431) );
  XOR U18585 ( .A(n18432), .B(n18431), .Z(n18380) );
  AND U18586 ( .A(y[30]), .B(x[160]), .Z(n18486) );
  AND U18587 ( .A(y[150]), .B(x[184]), .Z(n18255) );
  AND U18588 ( .A(x[185]), .B(y[149]), .Z(n18254) );
  XOR U18589 ( .A(n18255), .B(n18254), .Z(n18485) );
  XNOR U18590 ( .A(n18486), .B(n18485), .Z(n18379) );
  XNOR U18591 ( .A(n18377), .B(n18378), .Z(n18288) );
  NAND U18592 ( .A(n18257), .B(n18256), .Z(n18261) );
  NAND U18593 ( .A(n18259), .B(n18258), .Z(n18260) );
  NAND U18594 ( .A(n18261), .B(n18260), .Z(n18287) );
  XOR U18595 ( .A(n18286), .B(n18287), .Z(n18542) );
  XOR U18596 ( .A(n18539), .B(n18540), .Z(n18535) );
  XOR U18597 ( .A(n18534), .B(n18533), .Z(n18571) );
  XOR U18598 ( .A(n18572), .B(n18571), .Z(n18557) );
  XNOR U18599 ( .A(n18558), .B(n18557), .Z(n18553) );
  NANDN U18600 ( .A(n18263), .B(n18262), .Z(n18267) );
  NAND U18601 ( .A(n18265), .B(n18264), .Z(n18266) );
  NAND U18602 ( .A(n18267), .B(n18266), .Z(n18551) );
  XOR U18603 ( .A(n18552), .B(n18551), .Z(o[190]) );
  NANDN U18604 ( .A(n18269), .B(n18268), .Z(n18273) );
  NANDN U18605 ( .A(n18271), .B(n18270), .Z(n18272) );
  AND U18606 ( .A(n18273), .B(n18272), .Z(n18568) );
  NAND U18607 ( .A(n18275), .B(n18274), .Z(n18279) );
  NAND U18608 ( .A(n18277), .B(n18276), .Z(n18278) );
  AND U18609 ( .A(n18279), .B(n18278), .Z(n18550) );
  NAND U18610 ( .A(n18281), .B(n18280), .Z(n18285) );
  NAND U18611 ( .A(n18283), .B(n18282), .Z(n18284) );
  AND U18612 ( .A(n18285), .B(n18284), .Z(n18532) );
  NANDN U18613 ( .A(n18287), .B(n18286), .Z(n18291) );
  NANDN U18614 ( .A(n18289), .B(n18288), .Z(n18290) );
  AND U18615 ( .A(n18291), .B(n18290), .Z(n18299) );
  NANDN U18616 ( .A(n18293), .B(n18292), .Z(n18297) );
  NANDN U18617 ( .A(n18295), .B(n18294), .Z(n18296) );
  NAND U18618 ( .A(n18297), .B(n18296), .Z(n18298) );
  XNOR U18619 ( .A(n18299), .B(n18298), .Z(n18530) );
  NAND U18620 ( .A(n18301), .B(n18300), .Z(n18305) );
  NAND U18621 ( .A(n18303), .B(n18302), .Z(n18304) );
  AND U18622 ( .A(n18305), .B(n18304), .Z(n18528) );
  NAND U18623 ( .A(n18307), .B(n18306), .Z(n18311) );
  NAND U18624 ( .A(n18309), .B(n18308), .Z(n18310) );
  AND U18625 ( .A(n18311), .B(n18310), .Z(n18418) );
  NAND U18626 ( .A(n18313), .B(n18312), .Z(n18317) );
  NAND U18627 ( .A(n18315), .B(n18314), .Z(n18316) );
  AND U18628 ( .A(n18317), .B(n18316), .Z(n18376) );
  AND U18629 ( .A(x[164]), .B(y[27]), .Z(n18319) );
  NAND U18630 ( .A(x[187]), .B(y[148]), .Z(n18318) );
  XNOR U18631 ( .A(n18319), .B(n18318), .Z(n18323) );
  AND U18632 ( .A(x[176]), .B(y[111]), .Z(n18321) );
  NAND U18633 ( .A(x[194]), .B(y[189]), .Z(n18320) );
  XNOR U18634 ( .A(n18321), .B(n18320), .Z(n18322) );
  XOR U18635 ( .A(n18323), .B(n18322), .Z(n18331) );
  AND U18636 ( .A(x[177]), .B(y[110]), .Z(n18325) );
  NAND U18637 ( .A(x[162]), .B(y[29]), .Z(n18324) );
  XNOR U18638 ( .A(n18325), .B(n18324), .Z(n18329) );
  AND U18639 ( .A(x[163]), .B(y[28]), .Z(n18327) );
  NAND U18640 ( .A(x[174]), .B(y[65]), .Z(n18326) );
  XNOR U18641 ( .A(n18327), .B(n18326), .Z(n18328) );
  XNOR U18642 ( .A(n18329), .B(n18328), .Z(n18330) );
  XNOR U18643 ( .A(n18331), .B(n18330), .Z(n18374) );
  AND U18644 ( .A(x[173]), .B(y[66]), .Z(n18336) );
  AND U18645 ( .A(y[150]), .B(x[185]), .Z(n18487) );
  AND U18646 ( .A(x[170]), .B(y[69]), .Z(n18333) );
  NAND U18647 ( .A(x[186]), .B(y[149]), .Z(n18332) );
  XNOR U18648 ( .A(n18333), .B(n18332), .Z(n18334) );
  XNOR U18649 ( .A(n18487), .B(n18334), .Z(n18335) );
  XNOR U18650 ( .A(n18336), .B(n18335), .Z(n18352) );
  AND U18651 ( .A(x[199]), .B(y[184]), .Z(n18338) );
  NAND U18652 ( .A(x[190]), .B(y[145]), .Z(n18337) );
  XNOR U18653 ( .A(n18338), .B(n18337), .Z(n18342) );
  AND U18654 ( .A(x[198]), .B(y[185]), .Z(n18340) );
  NAND U18655 ( .A(x[180]), .B(y[107]), .Z(n18339) );
  XNOR U18656 ( .A(n18340), .B(n18339), .Z(n18341) );
  XOR U18657 ( .A(n18342), .B(n18341), .Z(n18350) );
  AND U18658 ( .A(x[184]), .B(y[151]), .Z(n18344) );
  NAND U18659 ( .A(x[179]), .B(y[108]), .Z(n18343) );
  XNOR U18660 ( .A(n18344), .B(n18343), .Z(n18348) );
  AND U18661 ( .A(x[169]), .B(y[70]), .Z(n18346) );
  NAND U18662 ( .A(x[175]), .B(y[64]), .Z(n18345) );
  XNOR U18663 ( .A(n18346), .B(n18345), .Z(n18347) );
  XNOR U18664 ( .A(n18348), .B(n18347), .Z(n18349) );
  XNOR U18665 ( .A(n18350), .B(n18349), .Z(n18351) );
  XOR U18666 ( .A(n18352), .B(n18351), .Z(n18372) );
  AND U18667 ( .A(x[191]), .B(y[144]), .Z(n18354) );
  NAND U18668 ( .A(x[188]), .B(y[147]), .Z(n18353) );
  XNOR U18669 ( .A(n18354), .B(n18353), .Z(n18358) );
  AND U18670 ( .A(x[160]), .B(y[31]), .Z(n18356) );
  NAND U18671 ( .A(x[167]), .B(y[24]), .Z(n18355) );
  XNOR U18672 ( .A(n18356), .B(n18355), .Z(n18357) );
  XOR U18673 ( .A(n18358), .B(n18357), .Z(n18366) );
  AND U18674 ( .A(x[161]), .B(y[30]), .Z(n18360) );
  NAND U18675 ( .A(x[181]), .B(y[106]), .Z(n18359) );
  XNOR U18676 ( .A(n18360), .B(n18359), .Z(n18364) );
  AND U18677 ( .A(x[168]), .B(y[71]), .Z(n18362) );
  NAND U18678 ( .A(x[195]), .B(y[188]), .Z(n18361) );
  XNOR U18679 ( .A(n18362), .B(n18361), .Z(n18363) );
  XNOR U18680 ( .A(n18364), .B(n18363), .Z(n18365) );
  XNOR U18681 ( .A(n18366), .B(n18365), .Z(n18370) );
  AND U18682 ( .A(y[67]), .B(x[172]), .Z(n18385) );
  AND U18683 ( .A(y[109]), .B(x[178]), .Z(n18433) );
  XOR U18684 ( .A(n18385), .B(n18433), .Z(n18368) );
  AND U18685 ( .A(y[26]), .B(x[165]), .Z(n18451) );
  AND U18686 ( .A(y[186]), .B(x[197]), .Z(n18447) );
  XNOR U18687 ( .A(n18451), .B(n18447), .Z(n18367) );
  XNOR U18688 ( .A(n18368), .B(n18367), .Z(n18369) );
  XNOR U18689 ( .A(n18370), .B(n18369), .Z(n18371) );
  XNOR U18690 ( .A(n18372), .B(n18371), .Z(n18373) );
  XNOR U18691 ( .A(n18374), .B(n18373), .Z(n18375) );
  XNOR U18692 ( .A(n18376), .B(n18375), .Z(n18416) );
  NANDN U18693 ( .A(n18378), .B(n18377), .Z(n18382) );
  NANDN U18694 ( .A(n18380), .B(n18379), .Z(n18381) );
  AND U18695 ( .A(n18382), .B(n18381), .Z(n18414) );
  NAND U18696 ( .A(n18384), .B(n18383), .Z(n18388) );
  NAND U18697 ( .A(n18386), .B(n18385), .Z(n18387) );
  AND U18698 ( .A(n18388), .B(n18387), .Z(n18396) );
  NAND U18699 ( .A(n18390), .B(n18389), .Z(n18394) );
  NAND U18700 ( .A(n18392), .B(n18391), .Z(n18393) );
  NAND U18701 ( .A(n18394), .B(n18393), .Z(n18395) );
  XNOR U18702 ( .A(n18396), .B(n18395), .Z(n18412) );
  NAND U18703 ( .A(n18398), .B(n18397), .Z(n18402) );
  NAND U18704 ( .A(n18400), .B(n18399), .Z(n18401) );
  AND U18705 ( .A(n18402), .B(n18401), .Z(n18410) );
  NAND U18706 ( .A(n18404), .B(n18403), .Z(n18408) );
  NAND U18707 ( .A(n18406), .B(n18405), .Z(n18407) );
  NAND U18708 ( .A(n18408), .B(n18407), .Z(n18409) );
  XNOR U18709 ( .A(n18410), .B(n18409), .Z(n18411) );
  XNOR U18710 ( .A(n18412), .B(n18411), .Z(n18413) );
  XNOR U18711 ( .A(n18414), .B(n18413), .Z(n18415) );
  XNOR U18712 ( .A(n18416), .B(n18415), .Z(n18417) );
  XNOR U18713 ( .A(n18418), .B(n18417), .Z(n18526) );
  NAND U18714 ( .A(n18420), .B(n18419), .Z(n18424) );
  NAND U18715 ( .A(n18422), .B(n18421), .Z(n18423) );
  AND U18716 ( .A(n18424), .B(n18423), .Z(n18524) );
  NAND U18717 ( .A(n18426), .B(n18425), .Z(n18430) );
  NANDN U18718 ( .A(n18428), .B(n18427), .Z(n18429) );
  AND U18719 ( .A(n18430), .B(n18429), .Z(n18506) );
  NAND U18720 ( .A(n18432), .B(n18431), .Z(n18436) );
  NAND U18721 ( .A(n18434), .B(n18433), .Z(n18435) );
  AND U18722 ( .A(n18436), .B(n18435), .Z(n18444) );
  NAND U18723 ( .A(n18438), .B(n18437), .Z(n18442) );
  NAND U18724 ( .A(n18440), .B(n18439), .Z(n18441) );
  NAND U18725 ( .A(n18442), .B(n18441), .Z(n18443) );
  XNOR U18726 ( .A(n18444), .B(n18443), .Z(n18504) );
  AND U18727 ( .A(x[189]), .B(y[146]), .Z(n18446) );
  NAND U18728 ( .A(x[183]), .B(y[104]), .Z(n18445) );
  XNOR U18729 ( .A(n18446), .B(n18445), .Z(n18470) );
  AND U18730 ( .A(n18448), .B(n18447), .Z(n18464) );
  NAND U18731 ( .A(n18450), .B(n18449), .Z(n18454) );
  NAND U18732 ( .A(n18452), .B(n18451), .Z(n18453) );
  AND U18733 ( .A(n18454), .B(n18453), .Z(n18462) );
  AND U18734 ( .A(x[192]), .B(y[191]), .Z(n18456) );
  NAND U18735 ( .A(x[182]), .B(y[105]), .Z(n18455) );
  XNOR U18736 ( .A(n18456), .B(n18455), .Z(n18460) );
  AND U18737 ( .A(x[193]), .B(y[190]), .Z(n18458) );
  NAND U18738 ( .A(x[166]), .B(y[25]), .Z(n18457) );
  XNOR U18739 ( .A(n18458), .B(n18457), .Z(n18459) );
  XNOR U18740 ( .A(n18460), .B(n18459), .Z(n18461) );
  XNOR U18741 ( .A(n18462), .B(n18461), .Z(n18463) );
  XOR U18742 ( .A(n18464), .B(n18463), .Z(n18468) );
  XNOR U18743 ( .A(n18466), .B(n18465), .Z(n18467) );
  XNOR U18744 ( .A(n18468), .B(n18467), .Z(n18469) );
  XOR U18745 ( .A(n18470), .B(n18469), .Z(n18502) );
  NAND U18746 ( .A(n18472), .B(n18471), .Z(n18476) );
  NAND U18747 ( .A(n18474), .B(n18473), .Z(n18475) );
  AND U18748 ( .A(n18476), .B(n18475), .Z(n18484) );
  NAND U18749 ( .A(n18478), .B(n18477), .Z(n18482) );
  NAND U18750 ( .A(n18480), .B(n18479), .Z(n18481) );
  NAND U18751 ( .A(n18482), .B(n18481), .Z(n18483) );
  XNOR U18752 ( .A(n18484), .B(n18483), .Z(n18500) );
  NAND U18753 ( .A(n18486), .B(n18485), .Z(n18490) );
  NAND U18754 ( .A(n18488), .B(n18487), .Z(n18489) );
  AND U18755 ( .A(n18490), .B(n18489), .Z(n18498) );
  NAND U18756 ( .A(n18492), .B(n18491), .Z(n18496) );
  NAND U18757 ( .A(n18494), .B(n18493), .Z(n18495) );
  NAND U18758 ( .A(n18496), .B(n18495), .Z(n18497) );
  XNOR U18759 ( .A(n18498), .B(n18497), .Z(n18499) );
  XNOR U18760 ( .A(n18500), .B(n18499), .Z(n18501) );
  XNOR U18761 ( .A(n18502), .B(n18501), .Z(n18503) );
  XNOR U18762 ( .A(n18504), .B(n18503), .Z(n18505) );
  XNOR U18763 ( .A(n18506), .B(n18505), .Z(n18522) );
  NAND U18764 ( .A(n18508), .B(n18507), .Z(n18512) );
  NANDN U18765 ( .A(n18510), .B(n18509), .Z(n18511) );
  AND U18766 ( .A(n18512), .B(n18511), .Z(n18520) );
  NAND U18767 ( .A(n18514), .B(n18513), .Z(n18518) );
  NANDN U18768 ( .A(n18516), .B(n18515), .Z(n18517) );
  NAND U18769 ( .A(n18518), .B(n18517), .Z(n18519) );
  XNOR U18770 ( .A(n18520), .B(n18519), .Z(n18521) );
  XNOR U18771 ( .A(n18522), .B(n18521), .Z(n18523) );
  XNOR U18772 ( .A(n18524), .B(n18523), .Z(n18525) );
  XNOR U18773 ( .A(n18526), .B(n18525), .Z(n18527) );
  XNOR U18774 ( .A(n18528), .B(n18527), .Z(n18529) );
  XNOR U18775 ( .A(n18530), .B(n18529), .Z(n18531) );
  XNOR U18776 ( .A(n18532), .B(n18531), .Z(n18548) );
  NAND U18777 ( .A(n18534), .B(n18533), .Z(n18538) );
  NANDN U18778 ( .A(n18536), .B(n18535), .Z(n18537) );
  AND U18779 ( .A(n18538), .B(n18537), .Z(n18546) );
  NAND U18780 ( .A(n18540), .B(n18539), .Z(n18544) );
  NANDN U18781 ( .A(n18542), .B(n18541), .Z(n18543) );
  NAND U18782 ( .A(n18544), .B(n18543), .Z(n18545) );
  XNOR U18783 ( .A(n18546), .B(n18545), .Z(n18547) );
  XNOR U18784 ( .A(n18548), .B(n18547), .Z(n18549) );
  XNOR U18785 ( .A(n18550), .B(n18549), .Z(n18566) );
  NAND U18786 ( .A(n18552), .B(n18551), .Z(n18556) );
  NANDN U18787 ( .A(n18554), .B(n18553), .Z(n18555) );
  AND U18788 ( .A(n18556), .B(n18555), .Z(n18564) );
  NAND U18789 ( .A(n18558), .B(n18557), .Z(n18562) );
  NANDN U18790 ( .A(n18560), .B(n18559), .Z(n18561) );
  NAND U18791 ( .A(n18562), .B(n18561), .Z(n18563) );
  XNOR U18792 ( .A(n18564), .B(n18563), .Z(n18565) );
  XNOR U18793 ( .A(n18566), .B(n18565), .Z(n18567) );
  XNOR U18794 ( .A(n18568), .B(n18567), .Z(n18576) );
  AND U18795 ( .A(n18570), .B(n18569), .Z(n18574) );
  AND U18796 ( .A(n18572), .B(n18571), .Z(n18573) );
  NOR U18797 ( .A(n18574), .B(n18573), .Z(n18575) );
  XNOR U18798 ( .A(n18576), .B(n18575), .Z(o[191]) );
  NAND U18799 ( .A(y[192]), .B(x[192]), .Z(n18715) );
  NAND U18800 ( .A(y[72]), .B(x[168]), .Z(n18579) );
  XOR U18801 ( .A(n18715), .B(n18579), .Z(n18580) );
  AND U18802 ( .A(y[32]), .B(x[160]), .Z(n18587) );
  AND U18803 ( .A(y[112]), .B(x[176]), .Z(n18584) );
  XOR U18804 ( .A(n18587), .B(n18584), .Z(n18583) );
  AND U18805 ( .A(y[152]), .B(x[184]), .Z(n18582) );
  XNOR U18806 ( .A(n18583), .B(n18582), .Z(n18581) );
  XNOR U18807 ( .A(n18580), .B(n18581), .Z(o[192]) );
  AND U18808 ( .A(x[161]), .B(y[32]), .Z(n18578) );
  NAND U18809 ( .A(x[160]), .B(y[33]), .Z(n18577) );
  XNOR U18810 ( .A(n18578), .B(n18577), .Z(n18589) );
  AND U18811 ( .A(y[72]), .B(x[169]), .Z(n18588) );
  XOR U18812 ( .A(n18589), .B(n18588), .Z(n18606) );
  AND U18813 ( .A(y[192]), .B(x[193]), .Z(n18818) );
  AND U18814 ( .A(y[113]), .B(x[176]), .Z(n18592) );
  XOR U18815 ( .A(n18818), .B(n18592), .Z(n18594) );
  AND U18816 ( .A(y[193]), .B(x[192]), .Z(n18616) );
  NAND U18817 ( .A(y[112]), .B(x[177]), .Z(n18615) );
  XNOR U18818 ( .A(n18616), .B(n18615), .Z(n18593) );
  XOR U18819 ( .A(n18594), .B(n18593), .Z(n18604) );
  AND U18820 ( .A(y[73]), .B(x[168]), .Z(n18842) );
  AND U18821 ( .A(y[153]), .B(x[184]), .Z(n18609) );
  XOR U18822 ( .A(n18842), .B(n18609), .Z(n18611) );
  AND U18823 ( .A(y[152]), .B(x[185]), .Z(n18610) );
  XNOR U18824 ( .A(n18611), .B(n18610), .Z(n18603) );
  XNOR U18825 ( .A(n18604), .B(n18603), .Z(n18605) );
  XNOR U18826 ( .A(n18606), .B(n18605), .Z(n18600) );
  NAND U18827 ( .A(n18583), .B(n18582), .Z(n18586) );
  AND U18828 ( .A(n18587), .B(n18584), .Z(n18585) );
  ANDN U18829 ( .B(n18586), .A(n18585), .Z(n18597) );
  XNOR U18830 ( .A(n18598), .B(n18597), .Z(n18599) );
  XNOR U18831 ( .A(n18600), .B(n18599), .Z(o[193]) );
  NAND U18832 ( .A(y[33]), .B(x[161]), .Z(n18638) );
  NANDN U18833 ( .A(n18638), .B(n18587), .Z(n18591) );
  NAND U18834 ( .A(n18589), .B(n18588), .Z(n18590) );
  AND U18835 ( .A(n18591), .B(n18590), .Z(n18673) );
  NAND U18836 ( .A(n18818), .B(n18592), .Z(n18596) );
  NAND U18837 ( .A(n18594), .B(n18593), .Z(n18595) );
  AND U18838 ( .A(n18596), .B(n18595), .Z(n18672) );
  AND U18839 ( .A(y[154]), .B(x[184]), .Z(n18657) );
  NAND U18840 ( .A(y[34]), .B(x[160]), .Z(n18658) );
  XNOR U18841 ( .A(n18657), .B(n18658), .Z(n18659) );
  NAND U18842 ( .A(y[72]), .B(x[170]), .Z(n18660) );
  XNOR U18843 ( .A(n18659), .B(n18660), .Z(n18671) );
  XOR U18844 ( .A(n18672), .B(n18671), .Z(n18674) );
  XOR U18845 ( .A(n18673), .B(n18674), .Z(n18618) );
  NANDN U18846 ( .A(n18598), .B(n18597), .Z(n18602) );
  NAND U18847 ( .A(n18600), .B(n18599), .Z(n18601) );
  NAND U18848 ( .A(n18602), .B(n18601), .Z(n18617) );
  XNOR U18849 ( .A(n18618), .B(n18617), .Z(n18620) );
  NANDN U18850 ( .A(n18604), .B(n18603), .Z(n18608) );
  NANDN U18851 ( .A(n18606), .B(n18605), .Z(n18607) );
  AND U18852 ( .A(n18608), .B(n18607), .Z(n18626) );
  AND U18853 ( .A(y[32]), .B(x[162]), .Z(n18635) );
  NAND U18854 ( .A(y[114]), .B(x[176]), .Z(n18636) );
  XNOR U18855 ( .A(n18635), .B(n18636), .Z(n18637) );
  AND U18856 ( .A(y[152]), .B(x[186]), .Z(n18665) );
  XOR U18857 ( .A(n18666), .B(n18665), .Z(n18668) );
  AND U18858 ( .A(y[112]), .B(x[178]), .Z(n18746) );
  AND U18859 ( .A(y[194]), .B(x[192]), .Z(n18648) );
  XOR U18860 ( .A(n18746), .B(n18648), .Z(n18650) );
  AND U18861 ( .A(y[113]), .B(x[177]), .Z(n18649) );
  XOR U18862 ( .A(n18650), .B(n18649), .Z(n18667) );
  XOR U18863 ( .A(n18668), .B(n18667), .Z(n18623) );
  NAND U18864 ( .A(n18842), .B(n18609), .Z(n18613) );
  AND U18865 ( .A(n18611), .B(n18610), .Z(n18612) );
  ANDN U18866 ( .B(n18613), .A(n18612), .Z(n18632) );
  AND U18867 ( .A(y[193]), .B(x[193]), .Z(n18720) );
  NAND U18868 ( .A(x[194]), .B(y[192]), .Z(n18614) );
  XNOR U18869 ( .A(n18720), .B(n18614), .Z(n18664) );
  ANDN U18870 ( .B(n18616), .A(n18615), .Z(n18663) );
  XOR U18871 ( .A(n18664), .B(n18663), .Z(n18629) );
  AND U18872 ( .A(y[153]), .B(x[185]), .Z(n18641) );
  NAND U18873 ( .A(y[73]), .B(x[169]), .Z(n18642) );
  XNOR U18874 ( .A(n18641), .B(n18642), .Z(n18643) );
  NAND U18875 ( .A(y[74]), .B(x[168]), .Z(n18644) );
  XOR U18876 ( .A(n18643), .B(n18644), .Z(n18630) );
  XNOR U18877 ( .A(n18629), .B(n18630), .Z(n18631) );
  XOR U18878 ( .A(n18632), .B(n18631), .Z(n18624) );
  XNOR U18879 ( .A(n18623), .B(n18624), .Z(n18625) );
  XNOR U18880 ( .A(n18626), .B(n18625), .Z(n18619) );
  XNOR U18881 ( .A(n18620), .B(n18619), .Z(o[194]) );
  NANDN U18882 ( .A(n18618), .B(n18617), .Z(n18622) );
  NAND U18883 ( .A(n18620), .B(n18619), .Z(n18621) );
  AND U18884 ( .A(n18622), .B(n18621), .Z(n18695) );
  NANDN U18885 ( .A(n18624), .B(n18623), .Z(n18628) );
  NAND U18886 ( .A(n18626), .B(n18625), .Z(n18627) );
  AND U18887 ( .A(n18628), .B(n18627), .Z(n18680) );
  NANDN U18888 ( .A(n18630), .B(n18629), .Z(n18634) );
  NANDN U18889 ( .A(n18632), .B(n18631), .Z(n18633) );
  AND U18890 ( .A(n18634), .B(n18633), .Z(n18678) );
  NANDN U18891 ( .A(n18636), .B(n18635), .Z(n18640) );
  NANDN U18892 ( .A(n18638), .B(n18637), .Z(n18639) );
  NAND U18893 ( .A(n18640), .B(n18639), .Z(n18689) );
  NANDN U18894 ( .A(n18642), .B(n18641), .Z(n18646) );
  NANDN U18895 ( .A(n18644), .B(n18643), .Z(n18645) );
  AND U18896 ( .A(n18646), .B(n18645), .Z(n18736) );
  AND U18897 ( .A(y[155]), .B(x[184]), .Z(n18764) );
  AND U18898 ( .A(y[115]), .B(x[176]), .Z(n18763) );
  NAND U18899 ( .A(y[32]), .B(x[163]), .Z(n18762) );
  XOR U18900 ( .A(n18763), .B(n18762), .Z(n18765) );
  XOR U18901 ( .A(n18764), .B(n18765), .Z(n18734) );
  AND U18902 ( .A(y[113]), .B(x[178]), .Z(n18798) );
  NAND U18903 ( .A(x[179]), .B(y[112]), .Z(n18647) );
  XNOR U18904 ( .A(n18798), .B(n18647), .Z(n18748) );
  AND U18905 ( .A(y[114]), .B(x[177]), .Z(n18747) );
  XOR U18906 ( .A(n18748), .B(n18747), .Z(n18733) );
  XNOR U18907 ( .A(n18734), .B(n18733), .Z(n18735) );
  XNOR U18908 ( .A(n18736), .B(n18735), .Z(n18690) );
  XOR U18909 ( .A(n18689), .B(n18690), .Z(n18692) );
  NAND U18910 ( .A(n18746), .B(n18648), .Z(n18652) );
  AND U18911 ( .A(n18650), .B(n18649), .Z(n18651) );
  ANDN U18912 ( .B(n18652), .A(n18651), .Z(n18741) );
  AND U18913 ( .A(y[34]), .B(x[161]), .Z(n18711) );
  AND U18914 ( .A(y[33]), .B(x[162]), .Z(n18710) );
  NAND U18915 ( .A(y[154]), .B(x[185]), .Z(n18709) );
  XOR U18916 ( .A(n18710), .B(n18709), .Z(n18712) );
  XOR U18917 ( .A(n18711), .B(n18712), .Z(n18740) );
  AND U18918 ( .A(x[195]), .B(y[192]), .Z(n18654) );
  NAND U18919 ( .A(x[192]), .B(y[195]), .Z(n18653) );
  XNOR U18920 ( .A(n18654), .B(n18653), .Z(n18716) );
  AND U18921 ( .A(x[193]), .B(y[194]), .Z(n18656) );
  NAND U18922 ( .A(x[194]), .B(y[193]), .Z(n18655) );
  XOR U18923 ( .A(n18656), .B(n18655), .Z(n18717) );
  XNOR U18924 ( .A(n18716), .B(n18717), .Z(n18739) );
  XOR U18925 ( .A(n18740), .B(n18739), .Z(n18742) );
  XOR U18926 ( .A(n18741), .B(n18742), .Z(n18691) );
  XOR U18927 ( .A(n18692), .B(n18691), .Z(n18677) );
  XNOR U18928 ( .A(n18678), .B(n18677), .Z(n18679) );
  XOR U18929 ( .A(n18680), .B(n18679), .Z(n18696) );
  XNOR U18930 ( .A(n18695), .B(n18696), .Z(n18698) );
  NANDN U18931 ( .A(n18658), .B(n18657), .Z(n18662) );
  NANDN U18932 ( .A(n18660), .B(n18659), .Z(n18661) );
  AND U18933 ( .A(n18662), .B(n18661), .Z(n18702) );
  AND U18934 ( .A(y[193]), .B(x[194]), .Z(n18815) );
  XNOR U18935 ( .A(n18702), .B(n18701), .Z(n18704) );
  AND U18936 ( .A(y[72]), .B(x[171]), .Z(n18756) );
  AND U18937 ( .A(y[35]), .B(x[160]), .Z(n18754) );
  NAND U18938 ( .A(y[153]), .B(x[186]), .Z(n18753) );
  XNOR U18939 ( .A(n18754), .B(n18753), .Z(n18755) );
  XOR U18940 ( .A(n18756), .B(n18755), .Z(n18729) );
  AND U18941 ( .A(y[75]), .B(x[168]), .Z(n18724) );
  AND U18942 ( .A(y[73]), .B(x[170]), .Z(n18722) );
  NAND U18943 ( .A(y[152]), .B(x[187]), .Z(n18721) );
  XNOR U18944 ( .A(n18722), .B(n18721), .Z(n18723) );
  XOR U18945 ( .A(n18724), .B(n18723), .Z(n18727) );
  AND U18946 ( .A(y[74]), .B(x[169]), .Z(n18728) );
  XOR U18947 ( .A(n18727), .B(n18728), .Z(n18730) );
  XOR U18948 ( .A(n18729), .B(n18730), .Z(n18703) );
  XOR U18949 ( .A(n18704), .B(n18703), .Z(n18684) );
  NAND U18950 ( .A(n18666), .B(n18665), .Z(n18670) );
  NAND U18951 ( .A(n18668), .B(n18667), .Z(n18669) );
  AND U18952 ( .A(n18670), .B(n18669), .Z(n18683) );
  XNOR U18953 ( .A(n18684), .B(n18683), .Z(n18686) );
  NANDN U18954 ( .A(n18672), .B(n18671), .Z(n18676) );
  OR U18955 ( .A(n18674), .B(n18673), .Z(n18675) );
  AND U18956 ( .A(n18676), .B(n18675), .Z(n18685) );
  XNOR U18957 ( .A(n18686), .B(n18685), .Z(n18697) );
  XOR U18958 ( .A(n18698), .B(n18697), .Z(o[195]) );
  NANDN U18959 ( .A(n18678), .B(n18677), .Z(n18682) );
  NANDN U18960 ( .A(n18680), .B(n18679), .Z(n18681) );
  AND U18961 ( .A(n18682), .B(n18681), .Z(n18776) );
  NANDN U18962 ( .A(n18684), .B(n18683), .Z(n18688) );
  NAND U18963 ( .A(n18686), .B(n18685), .Z(n18687) );
  NAND U18964 ( .A(n18688), .B(n18687), .Z(n18774) );
  NAND U18965 ( .A(n18690), .B(n18689), .Z(n18694) );
  NAND U18966 ( .A(n18692), .B(n18691), .Z(n18693) );
  AND U18967 ( .A(n18694), .B(n18693), .Z(n18775) );
  XOR U18968 ( .A(n18774), .B(n18775), .Z(n18777) );
  XOR U18969 ( .A(n18776), .B(n18777), .Z(n18768) );
  NANDN U18970 ( .A(n18696), .B(n18695), .Z(n18700) );
  NAND U18971 ( .A(n18698), .B(n18697), .Z(n18699) );
  NAND U18972 ( .A(n18700), .B(n18699), .Z(n18769) );
  XNOR U18973 ( .A(n18768), .B(n18769), .Z(n18771) );
  NANDN U18974 ( .A(n18702), .B(n18701), .Z(n18706) );
  NAND U18975 ( .A(n18704), .B(n18703), .Z(n18705) );
  AND U18976 ( .A(n18706), .B(n18705), .Z(n18781) );
  AND U18977 ( .A(x[168]), .B(y[76]), .Z(n18708) );
  NAND U18978 ( .A(x[171]), .B(y[73]), .Z(n18707) );
  XNOR U18979 ( .A(n18708), .B(n18707), .Z(n18843) );
  NAND U18980 ( .A(y[74]), .B(x[170]), .Z(n18899) );
  NAND U18981 ( .A(y[75]), .B(x[169]), .Z(n18847) );
  XNOR U18982 ( .A(n18846), .B(n18847), .Z(n18849) );
  AND U18983 ( .A(y[152]), .B(x[188]), .Z(n18803) );
  NAND U18984 ( .A(y[35]), .B(x[161]), .Z(n18804) );
  XNOR U18985 ( .A(n18803), .B(n18804), .Z(n18805) );
  NAND U18986 ( .A(y[36]), .B(x[160]), .Z(n18806) );
  XNOR U18987 ( .A(n18805), .B(n18806), .Z(n18848) );
  XOR U18988 ( .A(n18849), .B(n18848), .Z(n18861) );
  NANDN U18989 ( .A(n18710), .B(n18709), .Z(n18714) );
  OR U18990 ( .A(n18712), .B(n18711), .Z(n18713) );
  AND U18991 ( .A(n18714), .B(n18713), .Z(n18859) );
  AND U18992 ( .A(y[195]), .B(x[195]), .Z(n19247) );
  NANDN U18993 ( .A(n18715), .B(n19247), .Z(n18719) );
  NANDN U18994 ( .A(n18717), .B(n18716), .Z(n18718) );
  AND U18995 ( .A(n18719), .B(n18718), .Z(n18858) );
  XNOR U18996 ( .A(n18859), .B(n18858), .Z(n18860) );
  XNOR U18997 ( .A(n18861), .B(n18860), .Z(n18879) );
  NAND U18998 ( .A(y[32]), .B(x[164]), .Z(n18827) );
  NAND U18999 ( .A(y[154]), .B(x[186]), .Z(n18826) );
  NAND U19000 ( .A(y[116]), .B(x[176]), .Z(n18825) );
  XNOR U19001 ( .A(n18826), .B(n18825), .Z(n18828) );
  AND U19002 ( .A(y[194]), .B(x[194]), .Z(n18761) );
  NAND U19003 ( .A(n18761), .B(n18720), .Z(n18823) );
  NAND U19004 ( .A(y[196]), .B(x[192]), .Z(n18999) );
  NAND U19005 ( .A(y[112]), .B(x[180]), .Z(n18916) );
  XNOR U19006 ( .A(n18999), .B(n18916), .Z(n18824) );
  XOR U19007 ( .A(n18823), .B(n18824), .Z(n18786) );
  XOR U19008 ( .A(n18787), .B(n18786), .Z(n18788) );
  NANDN U19009 ( .A(n18722), .B(n18721), .Z(n18726) );
  NANDN U19010 ( .A(n18724), .B(n18723), .Z(n18725) );
  NAND U19011 ( .A(n18726), .B(n18725), .Z(n18789) );
  XOR U19012 ( .A(n18788), .B(n18789), .Z(n18876) );
  NAND U19013 ( .A(n18728), .B(n18727), .Z(n18732) );
  NAND U19014 ( .A(n18730), .B(n18729), .Z(n18731) );
  AND U19015 ( .A(n18732), .B(n18731), .Z(n18877) );
  XOR U19016 ( .A(n18876), .B(n18877), .Z(n18878) );
  XNOR U19017 ( .A(n18879), .B(n18878), .Z(n18780) );
  XNOR U19018 ( .A(n18781), .B(n18780), .Z(n18783) );
  NANDN U19019 ( .A(n18734), .B(n18733), .Z(n18738) );
  NANDN U19020 ( .A(n18736), .B(n18735), .Z(n18737) );
  NAND U19021 ( .A(n18738), .B(n18737), .Z(n18865) );
  NANDN U19022 ( .A(n18740), .B(n18739), .Z(n18744) );
  OR U19023 ( .A(n18742), .B(n18741), .Z(n18743) );
  NAND U19024 ( .A(n18744), .B(n18743), .Z(n18864) );
  XOR U19025 ( .A(n18865), .B(n18864), .Z(n18867) );
  AND U19026 ( .A(y[113]), .B(x[179]), .Z(n18745) );
  NAND U19027 ( .A(n18746), .B(n18745), .Z(n18750) );
  NAND U19028 ( .A(n18748), .B(n18747), .Z(n18749) );
  NAND U19029 ( .A(n18750), .B(n18749), .Z(n18870) );
  AND U19030 ( .A(y[72]), .B(x[172]), .Z(n18809) );
  NAND U19031 ( .A(y[156]), .B(x[184]), .Z(n18810) );
  XNOR U19032 ( .A(n18809), .B(n18810), .Z(n18811) );
  NAND U19033 ( .A(y[155]), .B(x[185]), .Z(n18812) );
  XNOR U19034 ( .A(n18811), .B(n18812), .Z(n18852) );
  AND U19035 ( .A(x[178]), .B(y[114]), .Z(n18752) );
  NAND U19036 ( .A(x[179]), .B(y[113]), .Z(n18751) );
  XNOR U19037 ( .A(n18752), .B(n18751), .Z(n18799) );
  NAND U19038 ( .A(y[115]), .B(x[177]), .Z(n18800) );
  XOR U19039 ( .A(n18799), .B(n18800), .Z(n18853) );
  XNOR U19040 ( .A(n18852), .B(n18853), .Z(n18854) );
  NANDN U19041 ( .A(n18754), .B(n18753), .Z(n18758) );
  NANDN U19042 ( .A(n18756), .B(n18755), .Z(n18757) );
  NAND U19043 ( .A(n18758), .B(n18757), .Z(n18855) );
  XNOR U19044 ( .A(n18854), .B(n18855), .Z(n18871) );
  XOR U19045 ( .A(n18870), .B(n18871), .Z(n18873) );
  NAND U19046 ( .A(y[34]), .B(x[162]), .Z(n18838) );
  NAND U19047 ( .A(y[153]), .B(x[187]), .Z(n18837) );
  NAND U19048 ( .A(y[33]), .B(x[163]), .Z(n18836) );
  XNOR U19049 ( .A(n18837), .B(n18836), .Z(n18839) );
  AND U19050 ( .A(x[196]), .B(y[192]), .Z(n18760) );
  NAND U19051 ( .A(x[193]), .B(y[195]), .Z(n18759) );
  XNOR U19052 ( .A(n18760), .B(n18759), .Z(n18820) );
  AND U19053 ( .A(y[193]), .B(x[195]), .Z(n18923) );
  XOR U19054 ( .A(n18761), .B(n18923), .Z(n18819) );
  XOR U19055 ( .A(n18820), .B(n18819), .Z(n18792) );
  XOR U19056 ( .A(n18793), .B(n18792), .Z(n18794) );
  NANDN U19057 ( .A(n18763), .B(n18762), .Z(n18767) );
  OR U19058 ( .A(n18765), .B(n18764), .Z(n18766) );
  NAND U19059 ( .A(n18767), .B(n18766), .Z(n18795) );
  XNOR U19060 ( .A(n18794), .B(n18795), .Z(n18872) );
  XOR U19061 ( .A(n18873), .B(n18872), .Z(n18866) );
  XOR U19062 ( .A(n18867), .B(n18866), .Z(n18782) );
  XNOR U19063 ( .A(n18783), .B(n18782), .Z(n18770) );
  XNOR U19064 ( .A(n18771), .B(n18770), .Z(o[196]) );
  NANDN U19065 ( .A(n18769), .B(n18768), .Z(n18773) );
  NAND U19066 ( .A(n18771), .B(n18770), .Z(n18772) );
  AND U19067 ( .A(n18773), .B(n18772), .Z(n19025) );
  NAND U19068 ( .A(n18775), .B(n18774), .Z(n18779) );
  NAND U19069 ( .A(n18777), .B(n18776), .Z(n18778) );
  NAND U19070 ( .A(n18779), .B(n18778), .Z(n19026) );
  XNOR U19071 ( .A(n19025), .B(n19026), .Z(n19028) );
  NANDN U19072 ( .A(n18781), .B(n18780), .Z(n18785) );
  NAND U19073 ( .A(n18783), .B(n18782), .Z(n18784) );
  AND U19074 ( .A(n18785), .B(n18784), .Z(n18883) );
  NAND U19075 ( .A(n18787), .B(n18786), .Z(n18791) );
  NANDN U19076 ( .A(n18789), .B(n18788), .Z(n18790) );
  AND U19077 ( .A(n18791), .B(n18790), .Z(n18935) );
  NAND U19078 ( .A(n18793), .B(n18792), .Z(n18797) );
  NANDN U19079 ( .A(n18795), .B(n18794), .Z(n18796) );
  NAND U19080 ( .A(n18797), .B(n18796), .Z(n18934) );
  AND U19081 ( .A(y[114]), .B(x[179]), .Z(n18917) );
  NAND U19082 ( .A(n18798), .B(n18917), .Z(n18802) );
  NANDN U19083 ( .A(n18800), .B(n18799), .Z(n18801) );
  AND U19084 ( .A(n18802), .B(n18801), .Z(n18887) );
  NANDN U19085 ( .A(n18804), .B(n18803), .Z(n18808) );
  NANDN U19086 ( .A(n18806), .B(n18805), .Z(n18807) );
  NAND U19087 ( .A(n18808), .B(n18807), .Z(n18912) );
  AND U19088 ( .A(y[157]), .B(x[184]), .Z(n19121) );
  AND U19089 ( .A(y[72]), .B(x[173]), .Z(n18930) );
  AND U19090 ( .A(y[115]), .B(x[178]), .Z(n18929) );
  XOR U19091 ( .A(n18930), .B(n18929), .Z(n18931) );
  XOR U19092 ( .A(n19121), .B(n18931), .Z(n18911) );
  AND U19093 ( .A(y[153]), .B(x[188]), .Z(n18925) );
  AND U19094 ( .A(y[32]), .B(x[165]), .Z(n18924) );
  XOR U19095 ( .A(n18925), .B(n18924), .Z(n18926) );
  AND U19096 ( .A(y[33]), .B(x[164]), .Z(n19089) );
  XOR U19097 ( .A(n18926), .B(n19089), .Z(n18910) );
  XOR U19098 ( .A(n18911), .B(n18910), .Z(n18913) );
  XOR U19099 ( .A(n18912), .B(n18913), .Z(n18886) );
  NANDN U19100 ( .A(n18810), .B(n18809), .Z(n18814) );
  NANDN U19101 ( .A(n18812), .B(n18811), .Z(n18813) );
  NAND U19102 ( .A(n18814), .B(n18813), .Z(n18990) );
  AND U19103 ( .A(x[195]), .B(y[194]), .Z(n18833) );
  AND U19104 ( .A(n18815), .B(n18833), .Z(n19001) );
  AND U19105 ( .A(x[192]), .B(y[197]), .Z(n18817) );
  AND U19106 ( .A(x[193]), .B(y[196]), .Z(n18816) );
  XOR U19107 ( .A(n18817), .B(n18816), .Z(n19000) );
  XOR U19108 ( .A(n19001), .B(n19000), .Z(n18989) );
  AND U19109 ( .A(y[73]), .B(x[172]), .Z(n18981) );
  AND U19110 ( .A(y[77]), .B(x[168]), .Z(n18979) );
  AND U19111 ( .A(y[36]), .B(x[161]), .Z(n18978) );
  XOR U19112 ( .A(n18979), .B(n18978), .Z(n18980) );
  XOR U19113 ( .A(n18981), .B(n18980), .Z(n18988) );
  XOR U19114 ( .A(n18989), .B(n18988), .Z(n18991) );
  XOR U19115 ( .A(n18990), .B(n18991), .Z(n18888) );
  XOR U19116 ( .A(n18889), .B(n18888), .Z(n18936) );
  XOR U19117 ( .A(n18937), .B(n18936), .Z(n19020) );
  AND U19118 ( .A(y[195]), .B(x[196]), .Z(n19114) );
  NAND U19119 ( .A(n19114), .B(n18818), .Z(n18822) );
  NAND U19120 ( .A(n18820), .B(n18819), .Z(n18821) );
  AND U19121 ( .A(n18822), .B(n18821), .Z(n18947) );
  NAND U19122 ( .A(n18826), .B(n18825), .Z(n18830) );
  NANDN U19123 ( .A(n18828), .B(n18827), .Z(n18829) );
  AND U19124 ( .A(n18830), .B(n18829), .Z(n18955) );
  AND U19125 ( .A(y[76]), .B(x[169]), .Z(n18900) );
  AND U19126 ( .A(y[74]), .B(x[171]), .Z(n19179) );
  NAND U19127 ( .A(x[170]), .B(y[75]), .Z(n18831) );
  XOR U19128 ( .A(n19179), .B(n18831), .Z(n18901) );
  NAND U19129 ( .A(x[196]), .B(y[193]), .Z(n18832) );
  XNOR U19130 ( .A(n18833), .B(n18832), .Z(n18895) );
  AND U19131 ( .A(y[192]), .B(x[197]), .Z(n18892) );
  NAND U19132 ( .A(y[195]), .B(x[194]), .Z(n18893) );
  XOR U19133 ( .A(n18895), .B(n18894), .Z(n18952) );
  XOR U19134 ( .A(n18953), .B(n18952), .Z(n18954) );
  XOR U19135 ( .A(n18955), .B(n18954), .Z(n18948) );
  XOR U19136 ( .A(n18949), .B(n18948), .Z(n18967) );
  AND U19137 ( .A(x[180]), .B(y[113]), .Z(n18835) );
  NAND U19138 ( .A(x[181]), .B(y[112]), .Z(n18834) );
  XOR U19139 ( .A(n18835), .B(n18834), .Z(n18918) );
  AND U19140 ( .A(y[152]), .B(x[189]), .Z(n18904) );
  NAND U19141 ( .A(y[34]), .B(x[163]), .Z(n18905) );
  AND U19142 ( .A(y[35]), .B(x[162]), .Z(n18906) );
  XOR U19143 ( .A(n18907), .B(n18906), .Z(n18970) );
  XOR U19144 ( .A(n18971), .B(n18970), .Z(n18973) );
  NAND U19145 ( .A(n18837), .B(n18836), .Z(n18841) );
  NANDN U19146 ( .A(n18839), .B(n18838), .Z(n18840) );
  AND U19147 ( .A(n18841), .B(n18840), .Z(n18972) );
  XOR U19148 ( .A(n18973), .B(n18972), .Z(n18965) );
  AND U19149 ( .A(y[76]), .B(x[171]), .Z(n19113) );
  NAND U19150 ( .A(n19113), .B(n18842), .Z(n18845) );
  NANDN U19151 ( .A(n18899), .B(n18843), .Z(n18844) );
  AND U19152 ( .A(n18845), .B(n18844), .Z(n18943) );
  AND U19153 ( .A(y[154]), .B(x[187]), .Z(n18994) );
  AND U19154 ( .A(y[116]), .B(x[177]), .Z(n19126) );
  XOR U19155 ( .A(n18994), .B(n19126), .Z(n18996) );
  AND U19156 ( .A(y[117]), .B(x[176]), .Z(n18995) );
  XOR U19157 ( .A(n18996), .B(n18995), .Z(n18941) );
  AND U19158 ( .A(y[37]), .B(x[160]), .Z(n19005) );
  AND U19159 ( .A(y[156]), .B(x[185]), .Z(n19004) );
  XOR U19160 ( .A(n19005), .B(n19004), .Z(n19007) );
  AND U19161 ( .A(y[155]), .B(x[186]), .Z(n19006) );
  XOR U19162 ( .A(n19007), .B(n19006), .Z(n18940) );
  XOR U19163 ( .A(n18941), .B(n18940), .Z(n18942) );
  XOR U19164 ( .A(n18943), .B(n18942), .Z(n18964) );
  NANDN U19165 ( .A(n18847), .B(n18846), .Z(n18851) );
  NAND U19166 ( .A(n18849), .B(n18848), .Z(n18850) );
  NAND U19167 ( .A(n18851), .B(n18850), .Z(n18959) );
  NANDN U19168 ( .A(n18853), .B(n18852), .Z(n18857) );
  NANDN U19169 ( .A(n18855), .B(n18854), .Z(n18856) );
  NAND U19170 ( .A(n18857), .B(n18856), .Z(n18958) );
  XOR U19171 ( .A(n18959), .B(n18958), .Z(n18961) );
  NANDN U19172 ( .A(n18859), .B(n18858), .Z(n18863) );
  NANDN U19173 ( .A(n18861), .B(n18860), .Z(n18862) );
  AND U19174 ( .A(n18863), .B(n18862), .Z(n18960) );
  XOR U19175 ( .A(n18961), .B(n18960), .Z(n19018) );
  XNOR U19176 ( .A(n19020), .B(n19021), .Z(n18882) );
  XNOR U19177 ( .A(n18883), .B(n18882), .Z(n18885) );
  NAND U19178 ( .A(n18865), .B(n18864), .Z(n18869) );
  NAND U19179 ( .A(n18867), .B(n18866), .Z(n18868) );
  NAND U19180 ( .A(n18869), .B(n18868), .Z(n19014) );
  NAND U19181 ( .A(n18871), .B(n18870), .Z(n18875) );
  NAND U19182 ( .A(n18873), .B(n18872), .Z(n18874) );
  NAND U19183 ( .A(n18875), .B(n18874), .Z(n19012) );
  NAND U19184 ( .A(n18877), .B(n18876), .Z(n18881) );
  NAND U19185 ( .A(n18879), .B(n18878), .Z(n18880) );
  AND U19186 ( .A(n18881), .B(n18880), .Z(n19013) );
  XOR U19187 ( .A(n19012), .B(n19013), .Z(n19015) );
  XOR U19188 ( .A(n19014), .B(n19015), .Z(n18884) );
  XOR U19189 ( .A(n18885), .B(n18884), .Z(n19027) );
  XOR U19190 ( .A(n19028), .B(n19027), .Z(o[197]) );
  NANDN U19191 ( .A(n18887), .B(n18886), .Z(n18891) );
  NAND U19192 ( .A(n18889), .B(n18888), .Z(n18890) );
  AND U19193 ( .A(n18891), .B(n18890), .Z(n19036) );
  NANDN U19194 ( .A(n18893), .B(n18892), .Z(n18897) );
  NAND U19195 ( .A(n18895), .B(n18894), .Z(n18896) );
  NAND U19196 ( .A(n18897), .B(n18896), .Z(n19069) );
  AND U19197 ( .A(y[75]), .B(x[171]), .Z(n18898) );
  NANDN U19198 ( .A(n18899), .B(n18898), .Z(n18903) );
  NANDN U19199 ( .A(n18901), .B(n18900), .Z(n18902) );
  AND U19200 ( .A(n18903), .B(n18902), .Z(n19282) );
  AND U19201 ( .A(y[155]), .B(x[187]), .Z(n19140) );
  AND U19202 ( .A(y[115]), .B(x[179]), .Z(n19139) );
  XOR U19203 ( .A(n19140), .B(n19139), .Z(n19138) );
  AND U19204 ( .A(y[35]), .B(x[163]), .Z(n19137) );
  XOR U19205 ( .A(n19138), .B(n19137), .Z(n19281) );
  AND U19206 ( .A(y[156]), .B(x[186]), .Z(n19100) );
  AND U19207 ( .A(y[114]), .B(x[180]), .Z(n19099) );
  XOR U19208 ( .A(n19100), .B(n19099), .Z(n19098) );
  AND U19209 ( .A(y[36]), .B(x[162]), .Z(n19097) );
  XNOR U19210 ( .A(n19098), .B(n19097), .Z(n19280) );
  XNOR U19211 ( .A(n19282), .B(n19283), .Z(n19072) );
  NANDN U19212 ( .A(n18905), .B(n18904), .Z(n18909) );
  NAND U19213 ( .A(n18907), .B(n18906), .Z(n18908) );
  NAND U19214 ( .A(n18909), .B(n18908), .Z(n19071) );
  XOR U19215 ( .A(n19069), .B(n19070), .Z(n19046) );
  NAND U19216 ( .A(n18911), .B(n18910), .Z(n18915) );
  NAND U19217 ( .A(n18913), .B(n18912), .Z(n18914) );
  NAND U19218 ( .A(n18915), .B(n18914), .Z(n19045) );
  XOR U19219 ( .A(n19046), .B(n19045), .Z(n19043) );
  AND U19220 ( .A(y[113]), .B(x[181]), .Z(n19084) );
  NANDN U19221 ( .A(n18916), .B(n19084), .Z(n18920) );
  NANDN U19222 ( .A(n18918), .B(n18917), .Z(n18919) );
  AND U19223 ( .A(n18920), .B(n18919), .Z(n19075) );
  AND U19224 ( .A(x[165]), .B(y[33]), .Z(n18922) );
  NAND U19225 ( .A(x[164]), .B(y[34]), .Z(n18921) );
  XNOR U19226 ( .A(n18922), .B(n18921), .Z(n19088) );
  AND U19227 ( .A(y[152]), .B(x[190]), .Z(n19087) );
  XOR U19228 ( .A(n19088), .B(n19087), .Z(n19078) );
  AND U19229 ( .A(y[197]), .B(x[193]), .Z(n19255) );
  AND U19230 ( .A(x[196]), .B(y[194]), .Z(n19011) );
  AND U19231 ( .A(n18923), .B(n19011), .Z(n19253) );
  AND U19232 ( .A(y[196]), .B(x[194]), .Z(n19252) );
  XOR U19233 ( .A(n19253), .B(n19252), .Z(n19254) );
  XNOR U19234 ( .A(n19255), .B(n19254), .Z(n19077) );
  XOR U19235 ( .A(n19075), .B(n19076), .Z(n19171) );
  NAND U19236 ( .A(n18925), .B(n18924), .Z(n18928) );
  NAND U19237 ( .A(n18926), .B(n19089), .Z(n18927) );
  NAND U19238 ( .A(n18928), .B(n18927), .Z(n19174) );
  NAND U19239 ( .A(n18930), .B(n18929), .Z(n18933) );
  NAND U19240 ( .A(n19121), .B(n18931), .Z(n18932) );
  NAND U19241 ( .A(n18933), .B(n18932), .Z(n19173) );
  XNOR U19242 ( .A(n19174), .B(n19173), .Z(n19172) );
  XNOR U19243 ( .A(n19043), .B(n19044), .Z(n19313) );
  NANDN U19244 ( .A(n18935), .B(n18934), .Z(n18939) );
  NAND U19245 ( .A(n18937), .B(n18936), .Z(n18938) );
  AND U19246 ( .A(n18939), .B(n18938), .Z(n19312) );
  NAND U19247 ( .A(n18941), .B(n18940), .Z(n18945) );
  NANDN U19248 ( .A(n18943), .B(n18942), .Z(n18944) );
  AND U19249 ( .A(n18945), .B(n18944), .Z(n19058) );
  NANDN U19250 ( .A(n18947), .B(n18946), .Z(n18951) );
  NAND U19251 ( .A(n18949), .B(n18948), .Z(n18950) );
  AND U19252 ( .A(n18951), .B(n18950), .Z(n19057) );
  XOR U19253 ( .A(n19058), .B(n19057), .Z(n19056) );
  NAND U19254 ( .A(n18953), .B(n18952), .Z(n18957) );
  NAND U19255 ( .A(n18955), .B(n18954), .Z(n18956) );
  AND U19256 ( .A(n18957), .B(n18956), .Z(n19055) );
  XOR U19257 ( .A(n19056), .B(n19055), .Z(n19310) );
  XOR U19258 ( .A(n19311), .B(n19310), .Z(n19035) );
  XOR U19259 ( .A(n19036), .B(n19035), .Z(n19038) );
  NAND U19260 ( .A(n18959), .B(n18958), .Z(n18963) );
  NAND U19261 ( .A(n18961), .B(n18960), .Z(n18962) );
  AND U19262 ( .A(n18963), .B(n18962), .Z(n19304) );
  NANDN U19263 ( .A(n18965), .B(n18964), .Z(n18969) );
  NANDN U19264 ( .A(n18967), .B(n18966), .Z(n18968) );
  NAND U19265 ( .A(n18969), .B(n18968), .Z(n19306) );
  NAND U19266 ( .A(n18971), .B(n18970), .Z(n18975) );
  NAND U19267 ( .A(n18973), .B(n18972), .Z(n18974) );
  AND U19268 ( .A(n18975), .B(n18974), .Z(n19042) );
  AND U19269 ( .A(y[118]), .B(x[176]), .Z(n19134) );
  AND U19270 ( .A(y[32]), .B(x[166]), .Z(n19133) );
  XOR U19271 ( .A(n19134), .B(n19133), .Z(n19132) );
  AND U19272 ( .A(y[153]), .B(x[189]), .Z(n19131) );
  XOR U19273 ( .A(n19132), .B(n19131), .Z(n19162) );
  AND U19274 ( .A(y[73]), .B(x[173]), .Z(n19267) );
  AND U19275 ( .A(y[76]), .B(x[170]), .Z(n19266) );
  XOR U19276 ( .A(n19267), .B(n19266), .Z(n19269) );
  AND U19277 ( .A(y[77]), .B(x[169]), .Z(n19268) );
  XOR U19278 ( .A(n19269), .B(n19268), .Z(n19178) );
  AND U19279 ( .A(x[172]), .B(y[74]), .Z(n18977) );
  NAND U19280 ( .A(x[171]), .B(y[75]), .Z(n18976) );
  XNOR U19281 ( .A(n18977), .B(n18976), .Z(n19177) );
  XOR U19282 ( .A(n19178), .B(n19177), .Z(n19161) );
  XOR U19283 ( .A(n19162), .B(n19161), .Z(n19160) );
  AND U19284 ( .A(y[198]), .B(x[192]), .Z(n19083) );
  XOR U19285 ( .A(n19084), .B(n19083), .Z(n19082) );
  AND U19286 ( .A(y[112]), .B(x[182]), .Z(n19081) );
  XOR U19287 ( .A(n19082), .B(n19081), .Z(n19159) );
  XOR U19288 ( .A(n19160), .B(n19159), .Z(n19065) );
  NAND U19289 ( .A(n18979), .B(n18978), .Z(n18983) );
  NAND U19290 ( .A(n18981), .B(n18980), .Z(n18982) );
  AND U19291 ( .A(n18983), .B(n18982), .Z(n19153) );
  AND U19292 ( .A(y[154]), .B(x[188]), .Z(n19125) );
  AND U19293 ( .A(x[177]), .B(y[117]), .Z(n18985) );
  AND U19294 ( .A(x[178]), .B(y[116]), .Z(n18984) );
  XOR U19295 ( .A(n18985), .B(n18984), .Z(n19124) );
  XOR U19296 ( .A(n19125), .B(n19124), .Z(n19156) );
  AND U19297 ( .A(y[38]), .B(x[160]), .Z(n19120) );
  AND U19298 ( .A(y[158]), .B(x[184]), .Z(n18987) );
  AND U19299 ( .A(x[185]), .B(y[157]), .Z(n18986) );
  XOR U19300 ( .A(n18987), .B(n18986), .Z(n19119) );
  XNOR U19301 ( .A(n19120), .B(n19119), .Z(n19155) );
  XNOR U19302 ( .A(n19153), .B(n19154), .Z(n19066) );
  NAND U19303 ( .A(n18989), .B(n18988), .Z(n18993) );
  NAND U19304 ( .A(n18991), .B(n18990), .Z(n18992) );
  AND U19305 ( .A(n18993), .B(n18992), .Z(n19063) );
  XOR U19306 ( .A(n19064), .B(n19063), .Z(n19041) );
  XOR U19307 ( .A(n19042), .B(n19041), .Z(n19040) );
  NAND U19308 ( .A(n18994), .B(n19126), .Z(n18998) );
  NAND U19309 ( .A(n18996), .B(n18995), .Z(n18997) );
  NAND U19310 ( .A(n18998), .B(n18997), .Z(n19049) );
  NANDN U19311 ( .A(n18999), .B(n19255), .Z(n19003) );
  NAND U19312 ( .A(n19001), .B(n19000), .Z(n19002) );
  NAND U19313 ( .A(n19003), .B(n19002), .Z(n19051) );
  NAND U19314 ( .A(n19005), .B(n19004), .Z(n19009) );
  NAND U19315 ( .A(n19007), .B(n19006), .Z(n19008) );
  AND U19316 ( .A(n19009), .B(n19008), .Z(n19277) );
  AND U19317 ( .A(y[37]), .B(x[161]), .Z(n19261) );
  AND U19318 ( .A(y[72]), .B(x[174]), .Z(n19260) );
  XOR U19319 ( .A(n19261), .B(n19260), .Z(n19263) );
  AND U19320 ( .A(y[78]), .B(x[168]), .Z(n19262) );
  XNOR U19321 ( .A(n19263), .B(n19262), .Z(n19275) );
  NAND U19322 ( .A(x[197]), .B(y[193]), .Z(n19010) );
  XNOR U19323 ( .A(n19011), .B(n19010), .Z(n19249) );
  AND U19324 ( .A(y[192]), .B(x[198]), .Z(n19248) );
  XOR U19325 ( .A(n19249), .B(n19248), .Z(n19246) );
  XOR U19326 ( .A(n19247), .B(n19246), .Z(n19274) );
  XNOR U19327 ( .A(n19277), .B(n19276), .Z(n19052) );
  XOR U19328 ( .A(n19049), .B(n19050), .Z(n19039) );
  XOR U19329 ( .A(n19040), .B(n19039), .Z(n19307) );
  XNOR U19330 ( .A(n19306), .B(n19307), .Z(n19305) );
  XOR U19331 ( .A(n19038), .B(n19037), .Z(n19320) );
  NAND U19332 ( .A(n19013), .B(n19012), .Z(n19017) );
  NAND U19333 ( .A(n19015), .B(n19014), .Z(n19016) );
  AND U19334 ( .A(n19017), .B(n19016), .Z(n19319) );
  NANDN U19335 ( .A(n19019), .B(n19018), .Z(n19023) );
  NANDN U19336 ( .A(n19021), .B(n19020), .Z(n19022) );
  AND U19337 ( .A(n19023), .B(n19022), .Z(n19318) );
  XNOR U19338 ( .A(n19319), .B(n19318), .Z(n19024) );
  XOR U19339 ( .A(n19320), .B(n19024), .Z(n19034) );
  NANDN U19340 ( .A(n19026), .B(n19025), .Z(n19030) );
  NAND U19341 ( .A(n19028), .B(n19027), .Z(n19029) );
  NAND U19342 ( .A(n19030), .B(n19029), .Z(n19031) );
  XOR U19343 ( .A(n19032), .B(n19031), .Z(o[198]) );
  NANDN U19344 ( .A(n19044), .B(n19043), .Z(n19048) );
  NAND U19345 ( .A(n19046), .B(n19045), .Z(n19047) );
  AND U19346 ( .A(n19048), .B(n19047), .Z(n19303) );
  NANDN U19347 ( .A(n19050), .B(n19049), .Z(n19054) );
  NANDN U19348 ( .A(n19052), .B(n19051), .Z(n19053) );
  AND U19349 ( .A(n19054), .B(n19053), .Z(n19062) );
  NAND U19350 ( .A(n19056), .B(n19055), .Z(n19060) );
  NAND U19351 ( .A(n19058), .B(n19057), .Z(n19059) );
  NAND U19352 ( .A(n19060), .B(n19059), .Z(n19061) );
  XNOR U19353 ( .A(n19062), .B(n19061), .Z(n19301) );
  NAND U19354 ( .A(n19064), .B(n19063), .Z(n19068) );
  ANDN U19355 ( .B(n19066), .A(n19065), .Z(n19067) );
  ANDN U19356 ( .B(n19068), .A(n19067), .Z(n19299) );
  NAND U19357 ( .A(n19070), .B(n19069), .Z(n19074) );
  NANDN U19358 ( .A(n19072), .B(n19071), .Z(n19073) );
  AND U19359 ( .A(n19074), .B(n19073), .Z(n19170) );
  NANDN U19360 ( .A(n19076), .B(n19075), .Z(n19080) );
  NANDN U19361 ( .A(n19078), .B(n19077), .Z(n19079) );
  AND U19362 ( .A(n19080), .B(n19079), .Z(n19152) );
  NAND U19363 ( .A(n19082), .B(n19081), .Z(n19086) );
  NAND U19364 ( .A(n19084), .B(n19083), .Z(n19085) );
  AND U19365 ( .A(n19086), .B(n19085), .Z(n19093) );
  NAND U19366 ( .A(n19088), .B(n19087), .Z(n19091) );
  AND U19367 ( .A(y[34]), .B(x[165]), .Z(n19235) );
  NAND U19368 ( .A(n19089), .B(n19235), .Z(n19090) );
  NAND U19369 ( .A(n19091), .B(n19090), .Z(n19092) );
  XNOR U19370 ( .A(n19093), .B(n19092), .Z(n19150) );
  AND U19371 ( .A(x[160]), .B(y[39]), .Z(n19095) );
  NAND U19372 ( .A(x[193]), .B(y[198]), .Z(n19094) );
  XNOR U19373 ( .A(n19095), .B(n19094), .Z(n19118) );
  AND U19374 ( .A(y[193]), .B(x[196]), .Z(n19096) );
  AND U19375 ( .A(y[194]), .B(x[197]), .Z(n19199) );
  AND U19376 ( .A(n19096), .B(n19199), .Z(n19112) );
  NAND U19377 ( .A(n19098), .B(n19097), .Z(n19102) );
  NAND U19378 ( .A(n19100), .B(n19099), .Z(n19101) );
  AND U19379 ( .A(n19102), .B(n19101), .Z(n19110) );
  AND U19380 ( .A(x[192]), .B(y[199]), .Z(n19104) );
  NAND U19381 ( .A(x[183]), .B(y[112]), .Z(n19103) );
  XNOR U19382 ( .A(n19104), .B(n19103), .Z(n19108) );
  AND U19383 ( .A(x[189]), .B(y[154]), .Z(n19106) );
  NAND U19384 ( .A(x[181]), .B(y[114]), .Z(n19105) );
  XNOR U19385 ( .A(n19106), .B(n19105), .Z(n19107) );
  XNOR U19386 ( .A(n19108), .B(n19107), .Z(n19109) );
  XNOR U19387 ( .A(n19110), .B(n19109), .Z(n19111) );
  XOR U19388 ( .A(n19112), .B(n19111), .Z(n19116) );
  XNOR U19389 ( .A(n19114), .B(n19113), .Z(n19115) );
  XNOR U19390 ( .A(n19116), .B(n19115), .Z(n19117) );
  XOR U19391 ( .A(n19118), .B(n19117), .Z(n19148) );
  NAND U19392 ( .A(n19120), .B(n19119), .Z(n19123) );
  AND U19393 ( .A(y[158]), .B(x[185]), .Z(n19232) );
  NAND U19394 ( .A(n19121), .B(n19232), .Z(n19122) );
  AND U19395 ( .A(n19123), .B(n19122), .Z(n19130) );
  NAND U19396 ( .A(n19125), .B(n19124), .Z(n19128) );
  AND U19397 ( .A(y[117]), .B(x[178]), .Z(n19233) );
  NAND U19398 ( .A(n19126), .B(n19233), .Z(n19127) );
  NAND U19399 ( .A(n19128), .B(n19127), .Z(n19129) );
  XNOR U19400 ( .A(n19130), .B(n19129), .Z(n19146) );
  NAND U19401 ( .A(n19132), .B(n19131), .Z(n19136) );
  NAND U19402 ( .A(n19134), .B(n19133), .Z(n19135) );
  AND U19403 ( .A(n19136), .B(n19135), .Z(n19144) );
  NAND U19404 ( .A(n19138), .B(n19137), .Z(n19142) );
  NAND U19405 ( .A(n19140), .B(n19139), .Z(n19141) );
  NAND U19406 ( .A(n19142), .B(n19141), .Z(n19143) );
  XNOR U19407 ( .A(n19144), .B(n19143), .Z(n19145) );
  XNOR U19408 ( .A(n19146), .B(n19145), .Z(n19147) );
  XNOR U19409 ( .A(n19148), .B(n19147), .Z(n19149) );
  XNOR U19410 ( .A(n19150), .B(n19149), .Z(n19151) );
  XNOR U19411 ( .A(n19152), .B(n19151), .Z(n19168) );
  NANDN U19412 ( .A(n19154), .B(n19153), .Z(n19158) );
  NANDN U19413 ( .A(n19156), .B(n19155), .Z(n19157) );
  AND U19414 ( .A(n19158), .B(n19157), .Z(n19166) );
  NAND U19415 ( .A(n19160), .B(n19159), .Z(n19164) );
  NAND U19416 ( .A(n19162), .B(n19161), .Z(n19163) );
  NAND U19417 ( .A(n19164), .B(n19163), .Z(n19165) );
  XNOR U19418 ( .A(n19166), .B(n19165), .Z(n19167) );
  XNOR U19419 ( .A(n19168), .B(n19167), .Z(n19169) );
  XNOR U19420 ( .A(n19170), .B(n19169), .Z(n19297) );
  NANDN U19421 ( .A(n19172), .B(n19171), .Z(n19176) );
  AND U19422 ( .A(n19174), .B(n19173), .Z(n19175) );
  ANDN U19423 ( .B(n19176), .A(n19175), .Z(n19295) );
  NAND U19424 ( .A(n19178), .B(n19177), .Z(n19181) );
  AND U19425 ( .A(y[75]), .B(x[172]), .Z(n19234) );
  NAND U19426 ( .A(n19179), .B(n19234), .Z(n19180) );
  AND U19427 ( .A(n19181), .B(n19180), .Z(n19245) );
  AND U19428 ( .A(x[167]), .B(y[32]), .Z(n19183) );
  NAND U19429 ( .A(x[199]), .B(y[192]), .Z(n19182) );
  XNOR U19430 ( .A(n19183), .B(n19182), .Z(n19187) );
  AND U19431 ( .A(x[162]), .B(y[37]), .Z(n19185) );
  NAND U19432 ( .A(x[198]), .B(y[193]), .Z(n19184) );
  XNOR U19433 ( .A(n19185), .B(n19184), .Z(n19186) );
  XOR U19434 ( .A(n19187), .B(n19186), .Z(n19195) );
  AND U19435 ( .A(x[195]), .B(y[196]), .Z(n19189) );
  NAND U19436 ( .A(x[166]), .B(y[33]), .Z(n19188) );
  XNOR U19437 ( .A(n19189), .B(n19188), .Z(n19193) );
  AND U19438 ( .A(x[188]), .B(y[155]), .Z(n19191) );
  NAND U19439 ( .A(x[182]), .B(y[113]), .Z(n19190) );
  XNOR U19440 ( .A(n19191), .B(n19190), .Z(n19192) );
  XNOR U19441 ( .A(n19193), .B(n19192), .Z(n19194) );
  XNOR U19442 ( .A(n19195), .B(n19194), .Z(n19243) );
  AND U19443 ( .A(x[186]), .B(y[157]), .Z(n19201) );
  AND U19444 ( .A(x[184]), .B(y[159]), .Z(n19197) );
  NAND U19445 ( .A(x[169]), .B(y[78]), .Z(n19196) );
  XNOR U19446 ( .A(n19197), .B(n19196), .Z(n19198) );
  XNOR U19447 ( .A(n19199), .B(n19198), .Z(n19200) );
  XNOR U19448 ( .A(n19201), .B(n19200), .Z(n19217) );
  AND U19449 ( .A(x[194]), .B(y[197]), .Z(n19203) );
  NAND U19450 ( .A(x[164]), .B(y[35]), .Z(n19202) );
  XNOR U19451 ( .A(n19203), .B(n19202), .Z(n19207) );
  AND U19452 ( .A(x[177]), .B(y[118]), .Z(n19205) );
  NAND U19453 ( .A(x[191]), .B(y[152]), .Z(n19204) );
  XNOR U19454 ( .A(n19205), .B(n19204), .Z(n19206) );
  XOR U19455 ( .A(n19207), .B(n19206), .Z(n19215) );
  AND U19456 ( .A(x[168]), .B(y[79]), .Z(n19209) );
  NAND U19457 ( .A(x[170]), .B(y[77]), .Z(n19208) );
  XNOR U19458 ( .A(n19209), .B(n19208), .Z(n19213) );
  AND U19459 ( .A(x[173]), .B(y[74]), .Z(n19211) );
  NAND U19460 ( .A(x[175]), .B(y[72]), .Z(n19210) );
  XNOR U19461 ( .A(n19211), .B(n19210), .Z(n19212) );
  XNOR U19462 ( .A(n19213), .B(n19212), .Z(n19214) );
  XNOR U19463 ( .A(n19215), .B(n19214), .Z(n19216) );
  XOR U19464 ( .A(n19217), .B(n19216), .Z(n19241) );
  AND U19465 ( .A(x[179]), .B(y[116]), .Z(n19219) );
  NAND U19466 ( .A(x[187]), .B(y[156]), .Z(n19218) );
  XNOR U19467 ( .A(n19219), .B(n19218), .Z(n19223) );
  AND U19468 ( .A(x[161]), .B(y[38]), .Z(n19221) );
  NAND U19469 ( .A(x[180]), .B(y[115]), .Z(n19220) );
  XNOR U19470 ( .A(n19221), .B(n19220), .Z(n19222) );
  XOR U19471 ( .A(n19223), .B(n19222), .Z(n19231) );
  AND U19472 ( .A(x[163]), .B(y[36]), .Z(n19225) );
  NAND U19473 ( .A(x[190]), .B(y[153]), .Z(n19224) );
  XNOR U19474 ( .A(n19225), .B(n19224), .Z(n19229) );
  AND U19475 ( .A(x[176]), .B(y[119]), .Z(n19227) );
  NAND U19476 ( .A(x[174]), .B(y[73]), .Z(n19226) );
  XNOR U19477 ( .A(n19227), .B(n19226), .Z(n19228) );
  XNOR U19478 ( .A(n19229), .B(n19228), .Z(n19230) );
  XNOR U19479 ( .A(n19231), .B(n19230), .Z(n19239) );
  XOR U19480 ( .A(n19233), .B(n19232), .Z(n19237) );
  XNOR U19481 ( .A(n19235), .B(n19234), .Z(n19236) );
  XNOR U19482 ( .A(n19237), .B(n19236), .Z(n19238) );
  XNOR U19483 ( .A(n19239), .B(n19238), .Z(n19240) );
  XNOR U19484 ( .A(n19241), .B(n19240), .Z(n19242) );
  XNOR U19485 ( .A(n19243), .B(n19242), .Z(n19244) );
  XNOR U19486 ( .A(n19245), .B(n19244), .Z(n19293) );
  NAND U19487 ( .A(n19247), .B(n19246), .Z(n19251) );
  AND U19488 ( .A(n19249), .B(n19248), .Z(n19250) );
  ANDN U19489 ( .B(n19251), .A(n19250), .Z(n19259) );
  AND U19490 ( .A(n19253), .B(n19252), .Z(n19257) );
  AND U19491 ( .A(n19255), .B(n19254), .Z(n19256) );
  OR U19492 ( .A(n19257), .B(n19256), .Z(n19258) );
  XNOR U19493 ( .A(n19259), .B(n19258), .Z(n19291) );
  AND U19494 ( .A(n19261), .B(n19260), .Z(n19265) );
  AND U19495 ( .A(n19263), .B(n19262), .Z(n19264) );
  NOR U19496 ( .A(n19265), .B(n19264), .Z(n19273) );
  NAND U19497 ( .A(n19267), .B(n19266), .Z(n19271) );
  NAND U19498 ( .A(n19269), .B(n19268), .Z(n19270) );
  AND U19499 ( .A(n19271), .B(n19270), .Z(n19272) );
  XNOR U19500 ( .A(n19273), .B(n19272), .Z(n19289) );
  ANDN U19501 ( .B(n19275), .A(n19274), .Z(n19279) );
  ANDN U19502 ( .B(n19277), .A(n19276), .Z(n19278) );
  NOR U19503 ( .A(n19279), .B(n19278), .Z(n19287) );
  NANDN U19504 ( .A(n19281), .B(n19280), .Z(n19285) );
  NANDN U19505 ( .A(n19283), .B(n19282), .Z(n19284) );
  AND U19506 ( .A(n19285), .B(n19284), .Z(n19286) );
  XNOR U19507 ( .A(n19287), .B(n19286), .Z(n19288) );
  XNOR U19508 ( .A(n19289), .B(n19288), .Z(n19290) );
  XNOR U19509 ( .A(n19291), .B(n19290), .Z(n19292) );
  XNOR U19510 ( .A(n19293), .B(n19292), .Z(n19294) );
  XNOR U19511 ( .A(n19295), .B(n19294), .Z(n19296) );
  XNOR U19512 ( .A(n19297), .B(n19296), .Z(n19298) );
  XNOR U19513 ( .A(n19299), .B(n19298), .Z(n19300) );
  XNOR U19514 ( .A(n19301), .B(n19300), .Z(n19302) );
  NANDN U19515 ( .A(n19305), .B(n19304), .Z(n19309) );
  NAND U19516 ( .A(n19307), .B(n19306), .Z(n19308) );
  AND U19517 ( .A(n19309), .B(n19308), .Z(n19317) );
  NAND U19518 ( .A(n19311), .B(n19310), .Z(n19315) );
  NANDN U19519 ( .A(n19313), .B(n19312), .Z(n19314) );
  NAND U19520 ( .A(n19315), .B(n19314), .Z(n19316) );
endmodule

