
module sum_N16384_CC256 ( clk, rst, a, b, c );
  input [63:0] a;
  input [63:0] b;
  output [63:0] c;
  input clk, rst;
  wire   carry_on, carry_on_d, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318;

  DFF carry_on_reg ( .D(carry_on_d), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        carry_on) );
  XOR U4 ( .A(n2), .B(n3), .Z(carry_on_d) );
  ANDN U5 ( .B(n4), .A(n5), .Z(n2) );
  XOR U6 ( .A(b[63]), .B(n3), .Z(n4) );
  XNOR U7 ( .A(b[9]), .B(n6), .Z(c[9]) );
  XNOR U8 ( .A(b[8]), .B(n7), .Z(c[8]) );
  XNOR U9 ( .A(b[7]), .B(n8), .Z(c[7]) );
  XNOR U10 ( .A(b[6]), .B(n9), .Z(c[6]) );
  XNOR U11 ( .A(b[63]), .B(n5), .Z(c[63]) );
  XNOR U12 ( .A(a[63]), .B(n3), .Z(n5) );
  XNOR U13 ( .A(n10), .B(n11), .Z(n3) );
  ANDN U14 ( .B(n12), .A(n13), .Z(n10) );
  XNOR U15 ( .A(b[62]), .B(n11), .Z(n12) );
  XNOR U16 ( .A(b[62]), .B(n13), .Z(c[62]) );
  XNOR U17 ( .A(a[62]), .B(n14), .Z(n13) );
  IV U18 ( .A(n11), .Z(n14) );
  XOR U19 ( .A(n15), .B(n16), .Z(n11) );
  ANDN U20 ( .B(n17), .A(n18), .Z(n15) );
  XNOR U21 ( .A(b[61]), .B(n16), .Z(n17) );
  XNOR U22 ( .A(b[61]), .B(n18), .Z(c[61]) );
  XNOR U23 ( .A(a[61]), .B(n19), .Z(n18) );
  IV U24 ( .A(n16), .Z(n19) );
  XOR U25 ( .A(n20), .B(n21), .Z(n16) );
  ANDN U26 ( .B(n22), .A(n23), .Z(n20) );
  XNOR U27 ( .A(b[60]), .B(n21), .Z(n22) );
  XNOR U28 ( .A(b[60]), .B(n23), .Z(c[60]) );
  XNOR U29 ( .A(a[60]), .B(n24), .Z(n23) );
  IV U30 ( .A(n21), .Z(n24) );
  XOR U31 ( .A(n25), .B(n26), .Z(n21) );
  ANDN U32 ( .B(n27), .A(n28), .Z(n25) );
  XNOR U33 ( .A(b[59]), .B(n26), .Z(n27) );
  XNOR U34 ( .A(b[5]), .B(n29), .Z(c[5]) );
  XNOR U35 ( .A(b[59]), .B(n28), .Z(c[59]) );
  XNOR U36 ( .A(a[59]), .B(n30), .Z(n28) );
  IV U37 ( .A(n26), .Z(n30) );
  XOR U38 ( .A(n31), .B(n32), .Z(n26) );
  ANDN U39 ( .B(n33), .A(n34), .Z(n31) );
  XNOR U40 ( .A(b[58]), .B(n32), .Z(n33) );
  XNOR U41 ( .A(b[58]), .B(n34), .Z(c[58]) );
  XNOR U42 ( .A(a[58]), .B(n35), .Z(n34) );
  IV U43 ( .A(n32), .Z(n35) );
  XOR U44 ( .A(n36), .B(n37), .Z(n32) );
  ANDN U45 ( .B(n38), .A(n39), .Z(n36) );
  XNOR U46 ( .A(b[57]), .B(n37), .Z(n38) );
  XNOR U47 ( .A(b[57]), .B(n39), .Z(c[57]) );
  XNOR U48 ( .A(a[57]), .B(n40), .Z(n39) );
  IV U49 ( .A(n37), .Z(n40) );
  XOR U50 ( .A(n41), .B(n42), .Z(n37) );
  ANDN U51 ( .B(n43), .A(n44), .Z(n41) );
  XNOR U52 ( .A(b[56]), .B(n42), .Z(n43) );
  XNOR U53 ( .A(b[56]), .B(n44), .Z(c[56]) );
  XNOR U54 ( .A(a[56]), .B(n45), .Z(n44) );
  IV U55 ( .A(n42), .Z(n45) );
  XOR U56 ( .A(n46), .B(n47), .Z(n42) );
  ANDN U57 ( .B(n48), .A(n49), .Z(n46) );
  XNOR U58 ( .A(b[55]), .B(n47), .Z(n48) );
  XNOR U59 ( .A(b[55]), .B(n49), .Z(c[55]) );
  XNOR U60 ( .A(a[55]), .B(n50), .Z(n49) );
  IV U61 ( .A(n47), .Z(n50) );
  XOR U62 ( .A(n51), .B(n52), .Z(n47) );
  ANDN U63 ( .B(n53), .A(n54), .Z(n51) );
  XNOR U64 ( .A(b[54]), .B(n52), .Z(n53) );
  XNOR U65 ( .A(b[54]), .B(n54), .Z(c[54]) );
  XNOR U66 ( .A(a[54]), .B(n55), .Z(n54) );
  IV U67 ( .A(n52), .Z(n55) );
  XOR U68 ( .A(n56), .B(n57), .Z(n52) );
  ANDN U69 ( .B(n58), .A(n59), .Z(n56) );
  XNOR U70 ( .A(b[53]), .B(n57), .Z(n58) );
  XNOR U71 ( .A(b[53]), .B(n59), .Z(c[53]) );
  XNOR U72 ( .A(a[53]), .B(n60), .Z(n59) );
  IV U73 ( .A(n57), .Z(n60) );
  XOR U74 ( .A(n61), .B(n62), .Z(n57) );
  ANDN U75 ( .B(n63), .A(n64), .Z(n61) );
  XNOR U76 ( .A(b[52]), .B(n62), .Z(n63) );
  XNOR U77 ( .A(b[52]), .B(n64), .Z(c[52]) );
  XNOR U78 ( .A(a[52]), .B(n65), .Z(n64) );
  IV U79 ( .A(n62), .Z(n65) );
  XOR U80 ( .A(n66), .B(n67), .Z(n62) );
  ANDN U81 ( .B(n68), .A(n69), .Z(n66) );
  XNOR U82 ( .A(b[51]), .B(n67), .Z(n68) );
  XNOR U83 ( .A(b[51]), .B(n69), .Z(c[51]) );
  XNOR U84 ( .A(a[51]), .B(n70), .Z(n69) );
  IV U85 ( .A(n67), .Z(n70) );
  XOR U86 ( .A(n71), .B(n72), .Z(n67) );
  ANDN U87 ( .B(n73), .A(n74), .Z(n71) );
  XNOR U88 ( .A(b[50]), .B(n72), .Z(n73) );
  XNOR U89 ( .A(b[50]), .B(n74), .Z(c[50]) );
  XNOR U90 ( .A(a[50]), .B(n75), .Z(n74) );
  IV U91 ( .A(n72), .Z(n75) );
  XOR U92 ( .A(n76), .B(n77), .Z(n72) );
  ANDN U93 ( .B(n78), .A(n79), .Z(n76) );
  XNOR U94 ( .A(b[49]), .B(n77), .Z(n78) );
  XNOR U95 ( .A(b[4]), .B(n80), .Z(c[4]) );
  XNOR U96 ( .A(b[49]), .B(n79), .Z(c[49]) );
  XNOR U97 ( .A(a[49]), .B(n81), .Z(n79) );
  IV U98 ( .A(n77), .Z(n81) );
  XOR U99 ( .A(n82), .B(n83), .Z(n77) );
  ANDN U100 ( .B(n84), .A(n85), .Z(n82) );
  XNOR U101 ( .A(b[48]), .B(n83), .Z(n84) );
  XNOR U102 ( .A(b[48]), .B(n85), .Z(c[48]) );
  XNOR U103 ( .A(a[48]), .B(n86), .Z(n85) );
  IV U104 ( .A(n83), .Z(n86) );
  XOR U105 ( .A(n87), .B(n88), .Z(n83) );
  ANDN U106 ( .B(n89), .A(n90), .Z(n87) );
  XNOR U107 ( .A(b[47]), .B(n88), .Z(n89) );
  XNOR U108 ( .A(b[47]), .B(n90), .Z(c[47]) );
  XNOR U109 ( .A(a[47]), .B(n91), .Z(n90) );
  IV U110 ( .A(n88), .Z(n91) );
  XOR U111 ( .A(n92), .B(n93), .Z(n88) );
  ANDN U112 ( .B(n94), .A(n95), .Z(n92) );
  XNOR U113 ( .A(b[46]), .B(n93), .Z(n94) );
  XNOR U114 ( .A(b[46]), .B(n95), .Z(c[46]) );
  XNOR U115 ( .A(a[46]), .B(n96), .Z(n95) );
  IV U116 ( .A(n93), .Z(n96) );
  XOR U117 ( .A(n97), .B(n98), .Z(n93) );
  ANDN U118 ( .B(n99), .A(n100), .Z(n97) );
  XNOR U119 ( .A(b[45]), .B(n98), .Z(n99) );
  XNOR U120 ( .A(b[45]), .B(n100), .Z(c[45]) );
  XNOR U121 ( .A(a[45]), .B(n101), .Z(n100) );
  IV U122 ( .A(n98), .Z(n101) );
  XOR U123 ( .A(n102), .B(n103), .Z(n98) );
  ANDN U124 ( .B(n104), .A(n105), .Z(n102) );
  XNOR U125 ( .A(b[44]), .B(n103), .Z(n104) );
  XNOR U126 ( .A(b[44]), .B(n105), .Z(c[44]) );
  XNOR U127 ( .A(a[44]), .B(n106), .Z(n105) );
  IV U128 ( .A(n103), .Z(n106) );
  XOR U129 ( .A(n107), .B(n108), .Z(n103) );
  ANDN U130 ( .B(n109), .A(n110), .Z(n107) );
  XNOR U131 ( .A(b[43]), .B(n108), .Z(n109) );
  XNOR U132 ( .A(b[43]), .B(n110), .Z(c[43]) );
  XNOR U133 ( .A(a[43]), .B(n111), .Z(n110) );
  IV U134 ( .A(n108), .Z(n111) );
  XOR U135 ( .A(n112), .B(n113), .Z(n108) );
  ANDN U136 ( .B(n114), .A(n115), .Z(n112) );
  XNOR U137 ( .A(b[42]), .B(n113), .Z(n114) );
  XNOR U138 ( .A(b[42]), .B(n115), .Z(c[42]) );
  XNOR U139 ( .A(a[42]), .B(n116), .Z(n115) );
  IV U140 ( .A(n113), .Z(n116) );
  XOR U141 ( .A(n117), .B(n118), .Z(n113) );
  ANDN U142 ( .B(n119), .A(n120), .Z(n117) );
  XNOR U143 ( .A(b[41]), .B(n118), .Z(n119) );
  XNOR U144 ( .A(b[41]), .B(n120), .Z(c[41]) );
  XNOR U145 ( .A(a[41]), .B(n121), .Z(n120) );
  IV U146 ( .A(n118), .Z(n121) );
  XOR U147 ( .A(n122), .B(n123), .Z(n118) );
  ANDN U148 ( .B(n124), .A(n125), .Z(n122) );
  XNOR U149 ( .A(b[40]), .B(n123), .Z(n124) );
  XNOR U150 ( .A(b[40]), .B(n125), .Z(c[40]) );
  XNOR U151 ( .A(a[40]), .B(n126), .Z(n125) );
  IV U152 ( .A(n123), .Z(n126) );
  XOR U153 ( .A(n127), .B(n128), .Z(n123) );
  ANDN U154 ( .B(n129), .A(n130), .Z(n127) );
  XNOR U155 ( .A(b[39]), .B(n128), .Z(n129) );
  XNOR U156 ( .A(b[3]), .B(n131), .Z(c[3]) );
  XNOR U157 ( .A(b[39]), .B(n130), .Z(c[39]) );
  XNOR U158 ( .A(a[39]), .B(n132), .Z(n130) );
  IV U159 ( .A(n128), .Z(n132) );
  XOR U160 ( .A(n133), .B(n134), .Z(n128) );
  ANDN U161 ( .B(n135), .A(n136), .Z(n133) );
  XNOR U162 ( .A(b[38]), .B(n134), .Z(n135) );
  XNOR U163 ( .A(b[38]), .B(n136), .Z(c[38]) );
  XNOR U164 ( .A(a[38]), .B(n137), .Z(n136) );
  IV U165 ( .A(n134), .Z(n137) );
  XOR U166 ( .A(n138), .B(n139), .Z(n134) );
  ANDN U167 ( .B(n140), .A(n141), .Z(n138) );
  XNOR U168 ( .A(b[37]), .B(n139), .Z(n140) );
  XNOR U169 ( .A(b[37]), .B(n141), .Z(c[37]) );
  XNOR U170 ( .A(a[37]), .B(n142), .Z(n141) );
  IV U171 ( .A(n139), .Z(n142) );
  XOR U172 ( .A(n143), .B(n144), .Z(n139) );
  ANDN U173 ( .B(n145), .A(n146), .Z(n143) );
  XNOR U174 ( .A(b[36]), .B(n144), .Z(n145) );
  XNOR U175 ( .A(b[36]), .B(n146), .Z(c[36]) );
  XNOR U176 ( .A(a[36]), .B(n147), .Z(n146) );
  IV U177 ( .A(n144), .Z(n147) );
  XOR U178 ( .A(n148), .B(n149), .Z(n144) );
  ANDN U179 ( .B(n150), .A(n151), .Z(n148) );
  XNOR U180 ( .A(b[35]), .B(n149), .Z(n150) );
  XNOR U181 ( .A(b[35]), .B(n151), .Z(c[35]) );
  XNOR U182 ( .A(a[35]), .B(n152), .Z(n151) );
  IV U183 ( .A(n149), .Z(n152) );
  XOR U184 ( .A(n153), .B(n154), .Z(n149) );
  ANDN U185 ( .B(n155), .A(n156), .Z(n153) );
  XNOR U186 ( .A(b[34]), .B(n154), .Z(n155) );
  XNOR U187 ( .A(b[34]), .B(n156), .Z(c[34]) );
  XNOR U188 ( .A(a[34]), .B(n157), .Z(n156) );
  IV U189 ( .A(n154), .Z(n157) );
  XOR U190 ( .A(n158), .B(n159), .Z(n154) );
  ANDN U191 ( .B(n160), .A(n161), .Z(n158) );
  XNOR U192 ( .A(b[33]), .B(n159), .Z(n160) );
  XNOR U193 ( .A(b[33]), .B(n161), .Z(c[33]) );
  XNOR U194 ( .A(a[33]), .B(n162), .Z(n161) );
  IV U195 ( .A(n159), .Z(n162) );
  XOR U196 ( .A(n163), .B(n164), .Z(n159) );
  ANDN U197 ( .B(n165), .A(n166), .Z(n163) );
  XNOR U198 ( .A(b[32]), .B(n164), .Z(n165) );
  XNOR U199 ( .A(b[32]), .B(n166), .Z(c[32]) );
  XNOR U200 ( .A(a[32]), .B(n167), .Z(n166) );
  IV U201 ( .A(n164), .Z(n167) );
  XOR U202 ( .A(n168), .B(n169), .Z(n164) );
  ANDN U203 ( .B(n170), .A(n171), .Z(n168) );
  XNOR U204 ( .A(b[31]), .B(n169), .Z(n170) );
  XNOR U205 ( .A(b[31]), .B(n171), .Z(c[31]) );
  XNOR U206 ( .A(a[31]), .B(n172), .Z(n171) );
  IV U207 ( .A(n169), .Z(n172) );
  XOR U208 ( .A(n173), .B(n174), .Z(n169) );
  ANDN U209 ( .B(n175), .A(n176), .Z(n173) );
  XNOR U210 ( .A(b[30]), .B(n174), .Z(n175) );
  XNOR U211 ( .A(b[30]), .B(n176), .Z(c[30]) );
  XNOR U212 ( .A(a[30]), .B(n177), .Z(n176) );
  IV U213 ( .A(n174), .Z(n177) );
  XOR U214 ( .A(n178), .B(n179), .Z(n174) );
  ANDN U215 ( .B(n180), .A(n181), .Z(n178) );
  XNOR U216 ( .A(b[29]), .B(n179), .Z(n180) );
  XNOR U217 ( .A(b[2]), .B(n182), .Z(c[2]) );
  XNOR U218 ( .A(b[29]), .B(n181), .Z(c[29]) );
  XNOR U219 ( .A(a[29]), .B(n183), .Z(n181) );
  IV U220 ( .A(n179), .Z(n183) );
  XOR U221 ( .A(n184), .B(n185), .Z(n179) );
  ANDN U222 ( .B(n186), .A(n187), .Z(n184) );
  XNOR U223 ( .A(b[28]), .B(n185), .Z(n186) );
  XNOR U224 ( .A(b[28]), .B(n187), .Z(c[28]) );
  XNOR U225 ( .A(a[28]), .B(n188), .Z(n187) );
  IV U226 ( .A(n185), .Z(n188) );
  XOR U227 ( .A(n189), .B(n190), .Z(n185) );
  ANDN U228 ( .B(n191), .A(n192), .Z(n189) );
  XNOR U229 ( .A(b[27]), .B(n190), .Z(n191) );
  XNOR U230 ( .A(b[27]), .B(n192), .Z(c[27]) );
  XNOR U231 ( .A(a[27]), .B(n193), .Z(n192) );
  IV U232 ( .A(n190), .Z(n193) );
  XOR U233 ( .A(n194), .B(n195), .Z(n190) );
  ANDN U234 ( .B(n196), .A(n197), .Z(n194) );
  XNOR U235 ( .A(b[26]), .B(n195), .Z(n196) );
  XNOR U236 ( .A(b[26]), .B(n197), .Z(c[26]) );
  XNOR U237 ( .A(a[26]), .B(n198), .Z(n197) );
  IV U238 ( .A(n195), .Z(n198) );
  XOR U239 ( .A(n199), .B(n200), .Z(n195) );
  ANDN U240 ( .B(n201), .A(n202), .Z(n199) );
  XNOR U241 ( .A(b[25]), .B(n200), .Z(n201) );
  XNOR U242 ( .A(b[25]), .B(n202), .Z(c[25]) );
  XNOR U243 ( .A(a[25]), .B(n203), .Z(n202) );
  IV U244 ( .A(n200), .Z(n203) );
  XOR U245 ( .A(n204), .B(n205), .Z(n200) );
  ANDN U246 ( .B(n206), .A(n207), .Z(n204) );
  XNOR U247 ( .A(b[24]), .B(n205), .Z(n206) );
  XNOR U248 ( .A(b[24]), .B(n207), .Z(c[24]) );
  XNOR U249 ( .A(a[24]), .B(n208), .Z(n207) );
  IV U250 ( .A(n205), .Z(n208) );
  XOR U251 ( .A(n209), .B(n210), .Z(n205) );
  ANDN U252 ( .B(n211), .A(n212), .Z(n209) );
  XNOR U253 ( .A(b[23]), .B(n210), .Z(n211) );
  XNOR U254 ( .A(b[23]), .B(n212), .Z(c[23]) );
  XNOR U255 ( .A(a[23]), .B(n213), .Z(n212) );
  IV U256 ( .A(n210), .Z(n213) );
  XOR U257 ( .A(n214), .B(n215), .Z(n210) );
  ANDN U258 ( .B(n216), .A(n217), .Z(n214) );
  XNOR U259 ( .A(b[22]), .B(n215), .Z(n216) );
  XNOR U260 ( .A(b[22]), .B(n217), .Z(c[22]) );
  XNOR U261 ( .A(a[22]), .B(n218), .Z(n217) );
  IV U262 ( .A(n215), .Z(n218) );
  XOR U263 ( .A(n219), .B(n220), .Z(n215) );
  ANDN U264 ( .B(n221), .A(n222), .Z(n219) );
  XNOR U265 ( .A(b[21]), .B(n220), .Z(n221) );
  XNOR U266 ( .A(b[21]), .B(n222), .Z(c[21]) );
  XNOR U267 ( .A(a[21]), .B(n223), .Z(n222) );
  IV U268 ( .A(n220), .Z(n223) );
  XOR U269 ( .A(n224), .B(n225), .Z(n220) );
  ANDN U270 ( .B(n226), .A(n227), .Z(n224) );
  XNOR U271 ( .A(b[20]), .B(n225), .Z(n226) );
  XNOR U272 ( .A(b[20]), .B(n227), .Z(c[20]) );
  XNOR U273 ( .A(a[20]), .B(n228), .Z(n227) );
  IV U274 ( .A(n225), .Z(n228) );
  XOR U275 ( .A(n229), .B(n230), .Z(n225) );
  ANDN U276 ( .B(n231), .A(n232), .Z(n229) );
  XNOR U277 ( .A(b[19]), .B(n230), .Z(n231) );
  XNOR U278 ( .A(b[1]), .B(n233), .Z(c[1]) );
  XNOR U279 ( .A(b[19]), .B(n232), .Z(c[19]) );
  XNOR U280 ( .A(a[19]), .B(n234), .Z(n232) );
  IV U281 ( .A(n230), .Z(n234) );
  XOR U282 ( .A(n235), .B(n236), .Z(n230) );
  ANDN U283 ( .B(n237), .A(n238), .Z(n235) );
  XNOR U284 ( .A(b[18]), .B(n236), .Z(n237) );
  XNOR U285 ( .A(b[18]), .B(n238), .Z(c[18]) );
  XNOR U286 ( .A(a[18]), .B(n239), .Z(n238) );
  IV U287 ( .A(n236), .Z(n239) );
  XOR U288 ( .A(n240), .B(n241), .Z(n236) );
  ANDN U289 ( .B(n242), .A(n243), .Z(n240) );
  XNOR U290 ( .A(b[17]), .B(n241), .Z(n242) );
  XNOR U291 ( .A(b[17]), .B(n243), .Z(c[17]) );
  XNOR U292 ( .A(a[17]), .B(n244), .Z(n243) );
  IV U293 ( .A(n241), .Z(n244) );
  XOR U294 ( .A(n245), .B(n246), .Z(n241) );
  ANDN U295 ( .B(n247), .A(n248), .Z(n245) );
  XNOR U296 ( .A(b[16]), .B(n246), .Z(n247) );
  XNOR U297 ( .A(b[16]), .B(n248), .Z(c[16]) );
  XNOR U298 ( .A(a[16]), .B(n249), .Z(n248) );
  IV U299 ( .A(n246), .Z(n249) );
  XOR U300 ( .A(n250), .B(n251), .Z(n246) );
  ANDN U301 ( .B(n252), .A(n253), .Z(n250) );
  XNOR U302 ( .A(b[15]), .B(n251), .Z(n252) );
  XNOR U303 ( .A(b[15]), .B(n253), .Z(c[15]) );
  XNOR U304 ( .A(a[15]), .B(n254), .Z(n253) );
  IV U305 ( .A(n251), .Z(n254) );
  XOR U306 ( .A(n255), .B(n256), .Z(n251) );
  ANDN U307 ( .B(n257), .A(n258), .Z(n255) );
  XNOR U308 ( .A(b[14]), .B(n256), .Z(n257) );
  XNOR U309 ( .A(b[14]), .B(n258), .Z(c[14]) );
  XNOR U310 ( .A(a[14]), .B(n259), .Z(n258) );
  IV U311 ( .A(n256), .Z(n259) );
  XOR U312 ( .A(n260), .B(n261), .Z(n256) );
  ANDN U313 ( .B(n262), .A(n263), .Z(n260) );
  XNOR U314 ( .A(b[13]), .B(n261), .Z(n262) );
  XNOR U315 ( .A(b[13]), .B(n263), .Z(c[13]) );
  XNOR U316 ( .A(a[13]), .B(n264), .Z(n263) );
  IV U317 ( .A(n261), .Z(n264) );
  XOR U318 ( .A(n265), .B(n266), .Z(n261) );
  ANDN U319 ( .B(n267), .A(n268), .Z(n265) );
  XNOR U320 ( .A(b[12]), .B(n266), .Z(n267) );
  XNOR U321 ( .A(b[12]), .B(n268), .Z(c[12]) );
  XNOR U322 ( .A(a[12]), .B(n269), .Z(n268) );
  IV U323 ( .A(n266), .Z(n269) );
  XOR U324 ( .A(n270), .B(n271), .Z(n266) );
  ANDN U325 ( .B(n272), .A(n273), .Z(n270) );
  XNOR U326 ( .A(b[11]), .B(n271), .Z(n272) );
  XNOR U327 ( .A(b[11]), .B(n273), .Z(c[11]) );
  XNOR U328 ( .A(a[11]), .B(n274), .Z(n273) );
  IV U329 ( .A(n271), .Z(n274) );
  XOR U330 ( .A(n275), .B(n276), .Z(n271) );
  ANDN U331 ( .B(n277), .A(n278), .Z(n275) );
  XNOR U332 ( .A(b[10]), .B(n276), .Z(n277) );
  XNOR U333 ( .A(b[10]), .B(n278), .Z(c[10]) );
  XNOR U334 ( .A(a[10]), .B(n279), .Z(n278) );
  IV U335 ( .A(n276), .Z(n279) );
  XOR U336 ( .A(n280), .B(n281), .Z(n276) );
  ANDN U337 ( .B(n282), .A(n6), .Z(n280) );
  XNOR U338 ( .A(a[9]), .B(n283), .Z(n6) );
  IV U339 ( .A(n281), .Z(n283) );
  XNOR U340 ( .A(b[9]), .B(n281), .Z(n282) );
  XOR U341 ( .A(n284), .B(n285), .Z(n281) );
  ANDN U342 ( .B(n286), .A(n7), .Z(n284) );
  XNOR U343 ( .A(a[8]), .B(n287), .Z(n7) );
  IV U344 ( .A(n285), .Z(n287) );
  XNOR U345 ( .A(b[8]), .B(n285), .Z(n286) );
  XOR U346 ( .A(n288), .B(n289), .Z(n285) );
  ANDN U347 ( .B(n290), .A(n8), .Z(n288) );
  XNOR U348 ( .A(a[7]), .B(n291), .Z(n8) );
  IV U349 ( .A(n289), .Z(n291) );
  XNOR U350 ( .A(b[7]), .B(n289), .Z(n290) );
  XOR U351 ( .A(n292), .B(n293), .Z(n289) );
  ANDN U352 ( .B(n294), .A(n9), .Z(n292) );
  XNOR U353 ( .A(a[6]), .B(n295), .Z(n9) );
  IV U354 ( .A(n293), .Z(n295) );
  XNOR U355 ( .A(b[6]), .B(n293), .Z(n294) );
  XOR U356 ( .A(n296), .B(n297), .Z(n293) );
  ANDN U357 ( .B(n298), .A(n29), .Z(n296) );
  XNOR U358 ( .A(a[5]), .B(n299), .Z(n29) );
  IV U359 ( .A(n297), .Z(n299) );
  XNOR U360 ( .A(b[5]), .B(n297), .Z(n298) );
  XOR U361 ( .A(n300), .B(n301), .Z(n297) );
  ANDN U362 ( .B(n302), .A(n80), .Z(n300) );
  XNOR U363 ( .A(a[4]), .B(n303), .Z(n80) );
  IV U364 ( .A(n301), .Z(n303) );
  XNOR U365 ( .A(b[4]), .B(n301), .Z(n302) );
  XOR U366 ( .A(n304), .B(n305), .Z(n301) );
  ANDN U367 ( .B(n306), .A(n131), .Z(n304) );
  XNOR U368 ( .A(a[3]), .B(n307), .Z(n131) );
  IV U369 ( .A(n305), .Z(n307) );
  XNOR U370 ( .A(b[3]), .B(n305), .Z(n306) );
  XOR U371 ( .A(n308), .B(n309), .Z(n305) );
  ANDN U372 ( .B(n310), .A(n182), .Z(n308) );
  XNOR U373 ( .A(a[2]), .B(n311), .Z(n182) );
  IV U374 ( .A(n309), .Z(n311) );
  XNOR U375 ( .A(b[2]), .B(n309), .Z(n310) );
  XOR U376 ( .A(n312), .B(n313), .Z(n309) );
  ANDN U377 ( .B(n314), .A(n233), .Z(n312) );
  XNOR U378 ( .A(a[1]), .B(n315), .Z(n233) );
  IV U379 ( .A(n313), .Z(n315) );
  XNOR U380 ( .A(b[1]), .B(n313), .Z(n314) );
  XOR U381 ( .A(carry_on), .B(n316), .Z(n313) );
  NANDN U382 ( .A(n317), .B(n318), .Z(n316) );
  XOR U383 ( .A(carry_on), .B(b[0]), .Z(n318) );
  XNOR U384 ( .A(b[0]), .B(n317), .Z(c[0]) );
  XNOR U385 ( .A(a[0]), .B(carry_on), .Z(n317) );
endmodule

