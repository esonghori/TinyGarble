
module hamming ( x, y, o );
  input [159:0] x;
  input [159:0] y;
  output [7:0] o;
  wire   n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079;

  IV U4045 ( .A(n4166), .Z(n2802) );
  NOR U4046 ( .A(n4165), .B(n2802), .Z(n2803) );
  NOR U4047 ( .A(n4167), .B(n2803), .Z(n2804) );
  NOR U4048 ( .A(n4164), .B(n4163), .Z(n2805) );
  NOR U4049 ( .A(n2805), .B(n2804), .Z(n4658) );
  XOR U4050 ( .A(n4605), .B(n4602), .Z(n2806) );
  NOR U4051 ( .A(n4603), .B(n2806), .Z(n2807) );
  NOR U4052 ( .A(n4604), .B(n4605), .Z(n2808) );
  NOR U4053 ( .A(n2807), .B(n4606), .Z(n2809) );
  IV U4054 ( .A(n2809), .Z(n2810) );
  NOR U4055 ( .A(n2808), .B(n2810), .Z(n2811) );
  NOR U4056 ( .A(n4608), .B(n4607), .Z(n2812) );
  NOR U4057 ( .A(n4609), .B(n2812), .Z(n2813) );
  NOR U4058 ( .A(n2811), .B(n2813), .Z(n5120) );
  XOR U4059 ( .A(x[159]), .B(y[159]), .Z(n2814) );
  IV U4060 ( .A(n2814), .Z(n2820) );
  XOR U4061 ( .A(x[158]), .B(y[158]), .Z(n2816) );
  XOR U4062 ( .A(x[157]), .B(y[157]), .Z(n2821) );
  XOR U4063 ( .A(x[156]), .B(y[156]), .Z(n2824) );
  XOR U4064 ( .A(x[155]), .B(y[155]), .Z(n3432) );
  XOR U4065 ( .A(x[154]), .B(y[154]), .Z(n3429) );
  XOR U4066 ( .A(x[153]), .B(y[153]), .Z(n3426) );
  XOR U4067 ( .A(x[152]), .B(y[152]), .Z(n3423) );
  XOR U4068 ( .A(x[151]), .B(y[151]), .Z(n2830) );
  XOR U4069 ( .A(x[150]), .B(y[150]), .Z(n2827) );
  XOR U4070 ( .A(x[149]), .B(y[149]), .Z(n2836) );
  XOR U4071 ( .A(x[148]), .B(y[148]), .Z(n2833) );
  XOR U4072 ( .A(x[147]), .B(y[147]), .Z(n2842) );
  XOR U4073 ( .A(x[146]), .B(y[146]), .Z(n2839) );
  XOR U4074 ( .A(x[145]), .B(y[145]), .Z(n3418) );
  XOR U4075 ( .A(x[144]), .B(y[144]), .Z(n3415) );
  XOR U4076 ( .A(x[143]), .B(y[143]), .Z(n2845) );
  XOR U4077 ( .A(x[142]), .B(y[142]), .Z(n2849) );
  XOR U4078 ( .A(x[141]), .B(y[141]), .Z(n3408) );
  XOR U4079 ( .A(x[140]), .B(y[140]), .Z(n2852) );
  XOR U4080 ( .A(x[139]), .B(y[139]), .Z(n2858) );
  XOR U4081 ( .A(x[138]), .B(y[138]), .Z(n2855) );
  XOR U4082 ( .A(x[137]), .B(y[137]), .Z(n2864) );
  XOR U4083 ( .A(x[136]), .B(y[136]), .Z(n2861) );
  XOR U4084 ( .A(x[135]), .B(y[135]), .Z(n2867) );
  XOR U4085 ( .A(x[134]), .B(y[134]), .Z(n3400) );
  XOR U4086 ( .A(x[133]), .B(y[133]), .Z(n3397) );
  XOR U4087 ( .A(x[132]), .B(y[132]), .Z(n2873) );
  XOR U4088 ( .A(x[131]), .B(y[131]), .Z(n2870) );
  XOR U4089 ( .A(x[130]), .B(y[130]), .Z(n2876) );
  XOR U4090 ( .A(x[129]), .B(y[129]), .Z(n3390) );
  XOR U4091 ( .A(x[128]), .B(y[128]), .Z(n2879) );
  XOR U4092 ( .A(x[127]), .B(y[127]), .Z(n3384) );
  XOR U4093 ( .A(x[126]), .B(y[126]), .Z(n3381) );
  XOR U4094 ( .A(x[125]), .B(y[125]), .Z(n2885) );
  XOR U4095 ( .A(x[124]), .B(y[124]), .Z(n2882) );
  XOR U4096 ( .A(x[123]), .B(y[123]), .Z(n2891) );
  XOR U4097 ( .A(x[122]), .B(y[122]), .Z(n2888) );
  XOR U4098 ( .A(x[121]), .B(y[121]), .Z(n3375) );
  XOR U4099 ( .A(x[120]), .B(y[120]), .Z(n3372) );
  XOR U4100 ( .A(x[119]), .B(y[119]), .Z(n2897) );
  XOR U4101 ( .A(x[118]), .B(y[118]), .Z(n2894) );
  XOR U4102 ( .A(x[117]), .B(y[117]), .Z(n2903) );
  XOR U4103 ( .A(x[116]), .B(y[116]), .Z(n2900) );
  XOR U4104 ( .A(x[115]), .B(y[115]), .Z(n3366) );
  XOR U4105 ( .A(x[114]), .B(y[114]), .Z(n3363) );
  XOR U4106 ( .A(x[113]), .B(y[113]), .Z(n3359) );
  XOR U4107 ( .A(x[112]), .B(y[112]), .Z(n3356) );
  XOR U4108 ( .A(x[111]), .B(y[111]), .Z(n3352) );
  XOR U4109 ( .A(x[110]), .B(y[110]), .Z(n3349) );
  XOR U4110 ( .A(x[109]), .B(y[109]), .Z(n3345) );
  XOR U4111 ( .A(x[108]), .B(y[108]), .Z(n3342) );
  XOR U4112 ( .A(x[107]), .B(y[107]), .Z(n3338) );
  XOR U4113 ( .A(x[106]), .B(y[106]), .Z(n3335) );
  XOR U4114 ( .A(x[105]), .B(y[105]), .Z(n2909) );
  XOR U4115 ( .A(x[104]), .B(y[104]), .Z(n2906) );
  XOR U4116 ( .A(x[103]), .B(y[103]), .Z(n3330) );
  XOR U4117 ( .A(x[102]), .B(y[102]), .Z(n3327) );
  XOR U4118 ( .A(x[101]), .B(y[101]), .Z(n2915) );
  XOR U4119 ( .A(x[100]), .B(y[100]), .Z(n2912) );
  XOR U4120 ( .A(x[99]), .B(y[99]), .Z(n2918) );
  XOR U4121 ( .A(x[98]), .B(y[98]), .Z(n3321) );
  XOR U4122 ( .A(x[97]), .B(y[97]), .Z(n3318) );
  XOR U4123 ( .A(x[96]), .B(y[96]), .Z(n2921) );
  XOR U4124 ( .A(x[95]), .B(y[95]), .Z(n2925) );
  XOR U4125 ( .A(x[94]), .B(y[94]), .Z(n2928) );
  XOR U4126 ( .A(x[93]), .B(y[93]), .Z(n3306) );
  XOR U4127 ( .A(x[92]), .B(y[92]), .Z(n2931) );
  XOR U4128 ( .A(x[91]), .B(y[91]), .Z(n2937) );
  XOR U4129 ( .A(x[90]), .B(y[90]), .Z(n2934) );
  XOR U4130 ( .A(x[89]), .B(y[89]), .Z(n2943) );
  XOR U4131 ( .A(x[88]), .B(y[88]), .Z(n2940) );
  XOR U4132 ( .A(x[87]), .B(y[87]), .Z(n2946) );
  XOR U4133 ( .A(x[86]), .B(y[86]), .Z(n2952) );
  XOR U4134 ( .A(x[85]), .B(y[85]), .Z(n2949) );
  XOR U4135 ( .A(x[84]), .B(y[84]), .Z(n2958) );
  XOR U4136 ( .A(x[83]), .B(y[83]), .Z(n2955) );
  XOR U4137 ( .A(x[82]), .B(y[82]), .Z(n3297) );
  XOR U4138 ( .A(x[81]), .B(y[81]), .Z(n3294) );
  XOR U4139 ( .A(x[80]), .B(y[80]), .Z(n2964) );
  XOR U4140 ( .A(x[79]), .B(y[79]), .Z(n2961) );
  XOR U4141 ( .A(x[78]), .B(y[78]), .Z(n2967) );
  XOR U4142 ( .A(x[77]), .B(y[77]), .Z(n3289) );
  XOR U4143 ( .A(x[76]), .B(y[76]), .Z(n3286) );
  XOR U4144 ( .A(x[75]), .B(y[75]), .Z(n2970) );
  XOR U4145 ( .A(x[74]), .B(y[74]), .Z(n2977) );
  XOR U4146 ( .A(x[73]), .B(y[73]), .Z(n2974) );
  XOR U4147 ( .A(x[72]), .B(y[72]), .Z(n3281) );
  XOR U4148 ( .A(x[71]), .B(y[71]), .Z(n3278) );
  XOR U4149 ( .A(x[70]), .B(y[70]), .Z(n2980) );
  XOR U4150 ( .A(x[69]), .B(y[69]), .Z(n3271) );
  XOR U4151 ( .A(x[68]), .B(y[68]), .Z(n2983) );
  XOR U4152 ( .A(x[67]), .B(y[67]), .Z(n3265) );
  XOR U4153 ( .A(x[66]), .B(y[66]), .Z(n3262) );
  XOR U4154 ( .A(x[65]), .B(y[65]), .Z(n3258) );
  XOR U4155 ( .A(x[64]), .B(y[64]), .Z(n3255) );
  XOR U4156 ( .A(x[63]), .B(y[63]), .Z(n3251) );
  XOR U4157 ( .A(x[62]), .B(y[62]), .Z(n3248) );
  XOR U4158 ( .A(x[61]), .B(y[61]), .Z(n2986) );
  XOR U4159 ( .A(x[60]), .B(y[60]), .Z(n2992) );
  XOR U4160 ( .A(x[59]), .B(y[59]), .Z(n2989) );
  XOR U4161 ( .A(x[58]), .B(y[58]), .Z(n3231) );
  XOR U4162 ( .A(x[57]), .B(y[57]), .Z(n3234) );
  XOR U4163 ( .A(x[56]), .B(y[56]), .Z(n2995) );
  XOR U4164 ( .A(x[55]), .B(y[55]), .Z(n2998) );
  XOR U4165 ( .A(x[54]), .B(y[54]), .Z(n3215) );
  XOR U4166 ( .A(x[53]), .B(y[53]), .Z(n3001) );
  XOR U4167 ( .A(x[52]), .B(y[52]), .Z(n3205) );
  XOR U4168 ( .A(x[51]), .B(y[51]), .Z(n3202) );
  XOR U4169 ( .A(x[50]), .B(y[50]), .Z(n3198) );
  XOR U4170 ( .A(x[49]), .B(y[49]), .Z(n3195) );
  XOR U4171 ( .A(x[48]), .B(y[48]), .Z(n3007) );
  XOR U4172 ( .A(x[47]), .B(y[47]), .Z(n3004) );
  XOR U4173 ( .A(x[46]), .B(y[46]), .Z(n3190) );
  XOR U4174 ( .A(x[45]), .B(y[45]), .Z(n3187) );
  XOR U4175 ( .A(x[44]), .B(y[44]), .Z(n3013) );
  XOR U4176 ( .A(x[43]), .B(y[43]), .Z(n3010) );
  XOR U4177 ( .A(x[42]), .B(y[42]), .Z(n3182) );
  XOR U4178 ( .A(x[41]), .B(y[41]), .Z(n3179) );
  XOR U4179 ( .A(x[40]), .B(y[40]), .Z(n3019) );
  XOR U4180 ( .A(x[39]), .B(y[39]), .Z(n3016) );
  XOR U4181 ( .A(x[38]), .B(y[38]), .Z(n3167) );
  XOR U4182 ( .A(x[37]), .B(y[37]), .Z(n3163) );
  XOR U4183 ( .A(x[36]), .B(y[36]), .Z(n3170) );
  XOR U4184 ( .A(x[35]), .B(y[35]), .Z(n3158) );
  XOR U4185 ( .A(x[34]), .B(y[34]), .Z(n3155) );
  XOR U4186 ( .A(x[33]), .B(y[33]), .Z(n3022) );
  XOR U4187 ( .A(x[32]), .B(y[32]), .Z(n3151) );
  XOR U4188 ( .A(x[31]), .B(y[31]), .Z(n3148) );
  XOR U4189 ( .A(x[30]), .B(y[30]), .Z(n3144) );
  XOR U4190 ( .A(x[29]), .B(y[29]), .Z(n3141) );
  XOR U4191 ( .A(x[28]), .B(y[28]), .Z(n3028) );
  XOR U4192 ( .A(x[27]), .B(y[27]), .Z(n3025) );
  XOR U4193 ( .A(x[26]), .B(y[26]), .Z(n3031) );
  XOR U4194 ( .A(x[25]), .B(y[25]), .Z(n3133) );
  XOR U4195 ( .A(x[24]), .B(y[24]), .Z(n3034) );
  XOR U4196 ( .A(x[23]), .B(y[23]), .Z(n3037) );
  XOR U4197 ( .A(x[22]), .B(y[22]), .Z(n3127) );
  XOR U4198 ( .A(x[21]), .B(y[21]), .Z(n3124) );
  XOR U4199 ( .A(x[20]), .B(y[20]), .Z(n3120) );
  XOR U4200 ( .A(x[19]), .B(y[19]), .Z(n3117) );
  XOR U4201 ( .A(x[18]), .B(y[18]), .Z(n3113) );
  XOR U4202 ( .A(x[17]), .B(y[17]), .Z(n3110) );
  XOR U4203 ( .A(x[16]), .B(y[16]), .Z(n3043) );
  XOR U4204 ( .A(x[15]), .B(y[15]), .Z(n3040) );
  XOR U4205 ( .A(x[14]), .B(y[14]), .Z(n3105) );
  XOR U4206 ( .A(x[13]), .B(y[13]), .Z(n3102) );
  XOR U4207 ( .A(x[12]), .B(y[12]), .Z(n3098) );
  XOR U4208 ( .A(x[11]), .B(y[11]), .Z(n3095) );
  XOR U4209 ( .A(x[10]), .B(y[10]), .Z(n3091) );
  XOR U4210 ( .A(x[9]), .B(y[9]), .Z(n3088) );
  XOR U4211 ( .A(x[8]), .B(y[8]), .Z(n3046) );
  XOR U4212 ( .A(x[7]), .B(y[7]), .Z(n3082) );
  XOR U4213 ( .A(x[6]), .B(y[6]), .Z(n3049) );
  XOR U4214 ( .A(x[5]), .B(y[5]), .Z(n3076) );
  XOR U4215 ( .A(x[4]), .B(y[4]), .Z(n3064) );
  XOR U4216 ( .A(x[3]), .B(y[3]), .Z(n3058) );
  XOR U4217 ( .A(x[2]), .B(y[2]), .Z(n3055) );
  XOR U4218 ( .A(x[1]), .B(y[1]), .Z(n2815) );
  IV U4219 ( .A(n2815), .Z(n3054) );
  XOR U4220 ( .A(x[0]), .B(y[0]), .Z(n3052) );
  XOR U4221 ( .A(n3054), .B(n3052), .Z(n3056) );
  XOR U4222 ( .A(n3055), .B(n3056), .Z(n3059) );
  XOR U4223 ( .A(n3058), .B(n3059), .Z(n3066) );
  XOR U4224 ( .A(n3064), .B(n3066), .Z(n3078) );
  XOR U4225 ( .A(n3076), .B(n3078), .Z(n3051) );
  XOR U4226 ( .A(n3049), .B(n3051), .Z(n3084) );
  XOR U4227 ( .A(n3082), .B(n3084), .Z(n3048) );
  XOR U4228 ( .A(n3046), .B(n3048), .Z(n3090) );
  XOR U4229 ( .A(n3088), .B(n3090), .Z(n3093) );
  XOR U4230 ( .A(n3091), .B(n3093), .Z(n3097) );
  XOR U4231 ( .A(n3095), .B(n3097), .Z(n3100) );
  XOR U4232 ( .A(n3098), .B(n3100), .Z(n3103) );
  XOR U4233 ( .A(n3102), .B(n3103), .Z(n3106) );
  XOR U4234 ( .A(n3105), .B(n3106), .Z(n3041) );
  XOR U4235 ( .A(n3040), .B(n3041), .Z(n3045) );
  XOR U4236 ( .A(n3043), .B(n3045), .Z(n3112) );
  XOR U4237 ( .A(n3110), .B(n3112), .Z(n3114) );
  XOR U4238 ( .A(n3113), .B(n3114), .Z(n3118) );
  XOR U4239 ( .A(n3117), .B(n3118), .Z(n3121) );
  XOR U4240 ( .A(n3120), .B(n3121), .Z(n3125) );
  XOR U4241 ( .A(n3124), .B(n3125), .Z(n3128) );
  XOR U4242 ( .A(n3127), .B(n3128), .Z(n3038) );
  XOR U4243 ( .A(n3037), .B(n3038), .Z(n3035) );
  XOR U4244 ( .A(n3034), .B(n3035), .Z(n3135) );
  XOR U4245 ( .A(n3133), .B(n3135), .Z(n3032) );
  XOR U4246 ( .A(n3031), .B(n3032), .Z(n3027) );
  XOR U4247 ( .A(n3025), .B(n3027), .Z(n3029) );
  XOR U4248 ( .A(n3028), .B(n3029), .Z(n3142) );
  XOR U4249 ( .A(n3141), .B(n3142), .Z(n3146) );
  XOR U4250 ( .A(n3144), .B(n3146), .Z(n3150) );
  XOR U4251 ( .A(n3148), .B(n3150), .Z(n3153) );
  XOR U4252 ( .A(n3151), .B(n3153), .Z(n3024) );
  XOR U4253 ( .A(n3022), .B(n3024), .Z(n3156) );
  XOR U4254 ( .A(n3155), .B(n3156), .Z(n3159) );
  XOR U4255 ( .A(n3158), .B(n3159), .Z(n3171) );
  XOR U4256 ( .A(n3170), .B(n3171), .Z(n3164) );
  XOR U4257 ( .A(n3163), .B(n3164), .Z(n3169) );
  XOR U4258 ( .A(n3167), .B(n3169), .Z(n3018) );
  XOR U4259 ( .A(n3016), .B(n3018), .Z(n3020) );
  XOR U4260 ( .A(n3019), .B(n3020), .Z(n3180) );
  XOR U4261 ( .A(n3179), .B(n3180), .Z(n3184) );
  XOR U4262 ( .A(n3182), .B(n3184), .Z(n3012) );
  XOR U4263 ( .A(n3010), .B(n3012), .Z(n3015) );
  XOR U4264 ( .A(n3013), .B(n3015), .Z(n3188) );
  XOR U4265 ( .A(n3187), .B(n3188), .Z(n3191) );
  XOR U4266 ( .A(n3190), .B(n3191), .Z(n3006) );
  XOR U4267 ( .A(n3004), .B(n3006), .Z(n3009) );
  XOR U4268 ( .A(n3007), .B(n3009), .Z(n3197) );
  XOR U4269 ( .A(n3195), .B(n3197), .Z(n3199) );
  XOR U4270 ( .A(n3198), .B(n3199), .Z(n3203) );
  XOR U4271 ( .A(n3202), .B(n3203), .Z(n3206) );
  XOR U4272 ( .A(n3205), .B(n3206), .Z(n3003) );
  XOR U4273 ( .A(n3001), .B(n3003), .Z(n3217) );
  XOR U4274 ( .A(n3215), .B(n3217), .Z(n3000) );
  XOR U4275 ( .A(n2998), .B(n3000), .Z(n2996) );
  XOR U4276 ( .A(n2995), .B(n2996), .Z(n3236) );
  XOR U4277 ( .A(n3234), .B(n3236), .Z(n3232) );
  XOR U4278 ( .A(n3231), .B(n3232), .Z(n2991) );
  XOR U4279 ( .A(n2989), .B(n2991), .Z(n2993) );
  XOR U4280 ( .A(n2992), .B(n2993), .Z(n2987) );
  XOR U4281 ( .A(n2986), .B(n2987), .Z(n3249) );
  XOR U4282 ( .A(n3248), .B(n3249), .Z(n3252) );
  XOR U4283 ( .A(n3251), .B(n3252), .Z(n3256) );
  XOR U4284 ( .A(n3255), .B(n3256), .Z(n3259) );
  XOR U4285 ( .A(n3258), .B(n3259), .Z(n3263) );
  XOR U4286 ( .A(n3262), .B(n3263), .Z(n3266) );
  XOR U4287 ( .A(n3265), .B(n3266), .Z(n2985) );
  XOR U4288 ( .A(n2983), .B(n2985), .Z(n3273) );
  XOR U4289 ( .A(n3271), .B(n3273), .Z(n2981) );
  XOR U4290 ( .A(n2980), .B(n2981), .Z(n3279) );
  XOR U4291 ( .A(n3278), .B(n3279), .Z(n3283) );
  XOR U4292 ( .A(n3281), .B(n3283), .Z(n2976) );
  XOR U4293 ( .A(n2974), .B(n2976), .Z(n2978) );
  XOR U4294 ( .A(n2977), .B(n2978), .Z(n2971) );
  XOR U4295 ( .A(n2970), .B(n2971), .Z(n3288) );
  XOR U4296 ( .A(n3286), .B(n3288), .Z(n3291) );
  XOR U4297 ( .A(n3289), .B(n3291), .Z(n2968) );
  XOR U4298 ( .A(n2967), .B(n2968), .Z(n2962) );
  XOR U4299 ( .A(n2961), .B(n2962), .Z(n2965) );
  XOR U4300 ( .A(n2964), .B(n2965), .Z(n3295) );
  XOR U4301 ( .A(n3294), .B(n3295), .Z(n3298) );
  XOR U4302 ( .A(n3297), .B(n3298), .Z(n2956) );
  XOR U4303 ( .A(n2955), .B(n2956), .Z(n2960) );
  XOR U4304 ( .A(n2958), .B(n2960), .Z(n2950) );
  XOR U4305 ( .A(n2949), .B(n2950), .Z(n2953) );
  XOR U4306 ( .A(n2952), .B(n2953), .Z(n2948) );
  XOR U4307 ( .A(n2946), .B(n2948), .Z(n2941) );
  XOR U4308 ( .A(n2940), .B(n2941), .Z(n2944) );
  XOR U4309 ( .A(n2943), .B(n2944), .Z(n2935) );
  XOR U4310 ( .A(n2934), .B(n2935), .Z(n2938) );
  XOR U4311 ( .A(n2937), .B(n2938), .Z(n2932) );
  XOR U4312 ( .A(n2931), .B(n2932), .Z(n3307) );
  XOR U4313 ( .A(n3306), .B(n3307), .Z(n2929) );
  XOR U4314 ( .A(n2928), .B(n2929), .Z(n2926) );
  XOR U4315 ( .A(n2925), .B(n2926), .Z(n2922) );
  XOR U4316 ( .A(n2921), .B(n2922), .Z(n3320) );
  XOR U4317 ( .A(n3318), .B(n3320), .Z(n3322) );
  XOR U4318 ( .A(n3321), .B(n3322), .Z(n2920) );
  XOR U4319 ( .A(n2918), .B(n2920), .Z(n2914) );
  XOR U4320 ( .A(n2912), .B(n2914), .Z(n2917) );
  XOR U4321 ( .A(n2915), .B(n2917), .Z(n3328) );
  XOR U4322 ( .A(n3327), .B(n3328), .Z(n3331) );
  XOR U4323 ( .A(n3330), .B(n3331), .Z(n2908) );
  XOR U4324 ( .A(n2906), .B(n2908), .Z(n2911) );
  XOR U4325 ( .A(n2909), .B(n2911), .Z(n3336) );
  XOR U4326 ( .A(n3335), .B(n3336), .Z(n3339) );
  XOR U4327 ( .A(n3338), .B(n3339), .Z(n3343) );
  XOR U4328 ( .A(n3342), .B(n3343), .Z(n3346) );
  XOR U4329 ( .A(n3345), .B(n3346), .Z(n3350) );
  XOR U4330 ( .A(n3349), .B(n3350), .Z(n3354) );
  XOR U4331 ( .A(n3352), .B(n3354), .Z(n3358) );
  XOR U4332 ( .A(n3356), .B(n3358), .Z(n3361) );
  XOR U4333 ( .A(n3359), .B(n3361), .Z(n3364) );
  XOR U4334 ( .A(n3363), .B(n3364), .Z(n3367) );
  XOR U4335 ( .A(n3366), .B(n3367), .Z(n2902) );
  XOR U4336 ( .A(n2900), .B(n2902), .Z(n2905) );
  XOR U4337 ( .A(n2903), .B(n2905), .Z(n2895) );
  XOR U4338 ( .A(n2894), .B(n2895), .Z(n2899) );
  XOR U4339 ( .A(n2897), .B(n2899), .Z(n3374) );
  XOR U4340 ( .A(n3372), .B(n3374), .Z(n3377) );
  XOR U4341 ( .A(n3375), .B(n3377), .Z(n2889) );
  XOR U4342 ( .A(n2888), .B(n2889), .Z(n2892) );
  XOR U4343 ( .A(n2891), .B(n2892), .Z(n2884) );
  XOR U4344 ( .A(n2882), .B(n2884), .Z(n2887) );
  XOR U4345 ( .A(n2885), .B(n2887), .Z(n3382) );
  XOR U4346 ( .A(n3381), .B(n3382), .Z(n3385) );
  XOR U4347 ( .A(n3384), .B(n3385), .Z(n2880) );
  XOR U4348 ( .A(n2879), .B(n2880), .Z(n3391) );
  XOR U4349 ( .A(n3390), .B(n3391), .Z(n2877) );
  XOR U4350 ( .A(n2876), .B(n2877), .Z(n2871) );
  XOR U4351 ( .A(n2870), .B(n2871), .Z(n2875) );
  XOR U4352 ( .A(n2873), .B(n2875), .Z(n3399) );
  XOR U4353 ( .A(n3397), .B(n3399), .Z(n3401) );
  XOR U4354 ( .A(n3400), .B(n3401), .Z(n2868) );
  XOR U4355 ( .A(n2867), .B(n2868), .Z(n2863) );
  XOR U4356 ( .A(n2861), .B(n2863), .Z(n2866) );
  XOR U4357 ( .A(n2864), .B(n2866), .Z(n2856) );
  XOR U4358 ( .A(n2855), .B(n2856), .Z(n2859) );
  XOR U4359 ( .A(n2858), .B(n2859), .Z(n2854) );
  XOR U4360 ( .A(n2852), .B(n2854), .Z(n3410) );
  XOR U4361 ( .A(n3408), .B(n3410), .Z(n2850) );
  XOR U4362 ( .A(n2849), .B(n2850), .Z(n2847) );
  XOR U4363 ( .A(n2845), .B(n2847), .Z(n3417) );
  XOR U4364 ( .A(n3415), .B(n3417), .Z(n3420) );
  XOR U4365 ( .A(n3418), .B(n3420), .Z(n2841) );
  XOR U4366 ( .A(n2839), .B(n2841), .Z(n2844) );
  XOR U4367 ( .A(n2842), .B(n2844), .Z(n2834) );
  XOR U4368 ( .A(n2833), .B(n2834), .Z(n2837) );
  XOR U4369 ( .A(n2836), .B(n2837), .Z(n2828) );
  XOR U4370 ( .A(n2827), .B(n2828), .Z(n2831) );
  XOR U4371 ( .A(n2830), .B(n2831), .Z(n3424) );
  XOR U4372 ( .A(n3423), .B(n3424), .Z(n3427) );
  XOR U4373 ( .A(n3426), .B(n3427), .Z(n3430) );
  XOR U4374 ( .A(n3429), .B(n3430), .Z(n3433) );
  XOR U4375 ( .A(n3432), .B(n3433), .Z(n2825) );
  XOR U4376 ( .A(n2824), .B(n2825), .Z(n2822) );
  XOR U4377 ( .A(n2821), .B(n2822), .Z(n2817) );
  XOR U4378 ( .A(n2816), .B(n2817), .Z(n2819) );
  XOR U4379 ( .A(n2820), .B(n2819), .Z(o[0]) );
  IV U4380 ( .A(n2816), .Z(n2818) );
  NOR U4381 ( .A(n2818), .B(n2817), .Z(n3436) );
  NOR U4382 ( .A(n2820), .B(n2819), .Z(n3908) );
  NOR U4383 ( .A(n3436), .B(n3908), .Z(n3435) );
  IV U4384 ( .A(n2821), .Z(n2823) );
  NOR U4385 ( .A(n2823), .B(n2822), .Z(n3905) );
  IV U4386 ( .A(n2824), .Z(n2826) );
  NOR U4387 ( .A(n2826), .B(n2825), .Z(n3900) );
  IV U4388 ( .A(n2827), .Z(n2829) );
  NOR U4389 ( .A(n2829), .B(n2828), .Z(n4422) );
  IV U4390 ( .A(n2830), .Z(n2832) );
  NOR U4391 ( .A(n2832), .B(n2831), .Z(n4420) );
  NOR U4392 ( .A(n4422), .B(n4420), .Z(n3893) );
  IV U4393 ( .A(n2833), .Z(n2835) );
  NOR U4394 ( .A(n2835), .B(n2834), .Z(n4890) );
  IV U4395 ( .A(n2836), .Z(n2838) );
  NOR U4396 ( .A(n2838), .B(n2837), .Z(n4885) );
  NOR U4397 ( .A(n4890), .B(n4885), .Z(n4856) );
  IV U4398 ( .A(n2839), .Z(n2840) );
  NOR U4399 ( .A(n2841), .B(n2840), .Z(n3883) );
  IV U4400 ( .A(n2842), .Z(n2843) );
  NOR U4401 ( .A(n2844), .B(n2843), .Z(n3439) );
  NOR U4402 ( .A(n3883), .B(n3439), .Z(n3422) );
  IV U4403 ( .A(n2845), .Z(n2846) );
  NOR U4404 ( .A(n2847), .B(n2846), .Z(n2848) );
  IV U4405 ( .A(n2848), .Z(n3447) );
  IV U4406 ( .A(n2849), .Z(n2851) );
  NOR U4407 ( .A(n2851), .B(n2850), .Z(n3413) );
  IV U4408 ( .A(n3413), .Z(n3407) );
  IV U4409 ( .A(n2852), .Z(n2853) );
  NOR U4410 ( .A(n2854), .B(n2853), .Z(n3875) );
  IV U4411 ( .A(n2855), .Z(n2857) );
  NOR U4412 ( .A(n2857), .B(n2856), .Z(n3953) );
  IV U4413 ( .A(n2858), .Z(n2860) );
  NOR U4414 ( .A(n2860), .B(n2859), .Z(n3948) );
  NOR U4415 ( .A(n3953), .B(n3948), .Z(n3874) );
  IV U4416 ( .A(n2861), .Z(n2862) );
  NOR U4417 ( .A(n2863), .B(n2862), .Z(n3453) );
  IV U4418 ( .A(n2864), .Z(n2865) );
  NOR U4419 ( .A(n2866), .B(n2865), .Z(n3448) );
  NOR U4420 ( .A(n3453), .B(n3448), .Z(n3405) );
  IV U4421 ( .A(n2867), .Z(n2869) );
  NOR U4422 ( .A(n2869), .B(n2868), .Z(n3451) );
  IV U4423 ( .A(n2870), .Z(n2872) );
  NOR U4424 ( .A(n2872), .B(n2871), .Z(n3974) );
  IV U4425 ( .A(n2873), .Z(n2874) );
  NOR U4426 ( .A(n2875), .B(n2874), .Z(n3970) );
  NOR U4427 ( .A(n3974), .B(n3970), .Z(n3863) );
  IV U4428 ( .A(n2876), .Z(n2878) );
  NOR U4429 ( .A(n2878), .B(n2877), .Z(n3395) );
  IV U4430 ( .A(n3395), .Z(n3389) );
  IV U4431 ( .A(n2879), .Z(n2881) );
  NOR U4432 ( .A(n2881), .B(n2880), .Z(n3459) );
  IV U4433 ( .A(n2882), .Z(n2883) );
  NOR U4434 ( .A(n2884), .B(n2883), .Z(n3859) );
  IV U4435 ( .A(n2885), .Z(n2886) );
  NOR U4436 ( .A(n2887), .B(n2886), .Z(n3853) );
  NOR U4437 ( .A(n3859), .B(n3853), .Z(n3380) );
  IV U4438 ( .A(n2888), .Z(n2890) );
  NOR U4439 ( .A(n2890), .B(n2889), .Z(n3842) );
  IV U4440 ( .A(n2891), .Z(n2893) );
  NOR U4441 ( .A(n2893), .B(n2892), .Z(n3467) );
  NOR U4442 ( .A(n3842), .B(n3467), .Z(n3379) );
  IV U4443 ( .A(n2894), .Z(n2896) );
  NOR U4444 ( .A(n2896), .B(n2895), .Z(n3834) );
  IV U4445 ( .A(n2897), .Z(n2898) );
  NOR U4446 ( .A(n2899), .B(n2898), .Z(n3471) );
  NOR U4447 ( .A(n3834), .B(n3471), .Z(n3371) );
  IV U4448 ( .A(n2900), .Z(n2901) );
  NOR U4449 ( .A(n2902), .B(n2901), .Z(n3478) );
  IV U4450 ( .A(n2903), .Z(n2904) );
  NOR U4451 ( .A(n2905), .B(n2904), .Z(n3475) );
  NOR U4452 ( .A(n3478), .B(n3475), .Z(n3370) );
  IV U4453 ( .A(n2906), .Z(n2907) );
  NOR U4454 ( .A(n2908), .B(n2907), .Z(n3497) );
  IV U4455 ( .A(n2909), .Z(n2910) );
  NOR U4456 ( .A(n2911), .B(n2910), .Z(n3495) );
  NOR U4457 ( .A(n3497), .B(n3495), .Z(n3334) );
  IV U4458 ( .A(n2912), .Z(n2913) );
  NOR U4459 ( .A(n2914), .B(n2913), .Z(n3503) );
  IV U4460 ( .A(n2915), .Z(n2916) );
  NOR U4461 ( .A(n2917), .B(n2916), .Z(n3807) );
  NOR U4462 ( .A(n3503), .B(n3807), .Z(n3326) );
  IV U4463 ( .A(n2918), .Z(n2919) );
  NOR U4464 ( .A(n2920), .B(n2919), .Z(n3505) );
  IV U4465 ( .A(n2921), .Z(n2923) );
  NOR U4466 ( .A(n2923), .B(n2922), .Z(n2924) );
  IV U4467 ( .A(n2924), .Z(n3513) );
  IV U4468 ( .A(n2925), .Z(n2927) );
  NOR U4469 ( .A(n2927), .B(n2926), .Z(n3313) );
  IV U4470 ( .A(n2928), .Z(n2930) );
  NOR U4471 ( .A(n2930), .B(n2929), .Z(n3310) );
  IV U4472 ( .A(n3310), .Z(n3305) );
  IV U4473 ( .A(n2931), .Z(n2933) );
  NOR U4474 ( .A(n2933), .B(n2932), .Z(n3516) );
  IV U4475 ( .A(n2934), .Z(n2936) );
  NOR U4476 ( .A(n2936), .B(n2935), .Z(n4310) );
  IV U4477 ( .A(n2937), .Z(n2939) );
  NOR U4478 ( .A(n2939), .B(n2938), .Z(n4054) );
  NOR U4479 ( .A(n4310), .B(n4054), .Z(n3521) );
  IV U4480 ( .A(n2940), .Z(n2942) );
  NOR U4481 ( .A(n2942), .B(n2941), .Z(n3526) );
  IV U4482 ( .A(n2943), .Z(n2945) );
  NOR U4483 ( .A(n2945), .B(n2944), .Z(n3522) );
  NOR U4484 ( .A(n3526), .B(n3522), .Z(n3303) );
  IV U4485 ( .A(n2946), .Z(n2947) );
  NOR U4486 ( .A(n2948), .B(n2947), .Z(n4308) );
  IV U4487 ( .A(n2949), .Z(n2951) );
  NOR U4488 ( .A(n2951), .B(n2950), .Z(n3792) );
  IV U4489 ( .A(n2952), .Z(n2954) );
  NOR U4490 ( .A(n2954), .B(n2953), .Z(n3529) );
  NOR U4491 ( .A(n3792), .B(n3529), .Z(n3302) );
  IV U4492 ( .A(n2955), .Z(n2957) );
  NOR U4493 ( .A(n2957), .B(n2956), .Z(n3534) );
  IV U4494 ( .A(n2958), .Z(n2959) );
  NOR U4495 ( .A(n2960), .B(n2959), .Z(n3795) );
  NOR U4496 ( .A(n3534), .B(n3795), .Z(n3301) );
  IV U4497 ( .A(n2961), .Z(n2963) );
  NOR U4498 ( .A(n2963), .B(n2962), .Z(n4067) );
  IV U4499 ( .A(n2964), .Z(n2966) );
  NOR U4500 ( .A(n2966), .B(n2965), .Z(n4061) );
  NOR U4501 ( .A(n4067), .B(n4061), .Z(n3789) );
  IV U4502 ( .A(n2967), .Z(n2969) );
  NOR U4503 ( .A(n2969), .B(n2968), .Z(n3787) );
  IV U4504 ( .A(n2970), .Z(n2972) );
  NOR U4505 ( .A(n2972), .B(n2971), .Z(n2973) );
  IV U4506 ( .A(n2973), .Z(n3778) );
  IV U4507 ( .A(n2974), .Z(n2975) );
  NOR U4508 ( .A(n2976), .B(n2975), .Z(n3544) );
  IV U4509 ( .A(n2977), .Z(n2979) );
  NOR U4510 ( .A(n2979), .B(n2978), .Z(n3542) );
  NOR U4511 ( .A(n3544), .B(n3542), .Z(n3285) );
  IV U4512 ( .A(n2980), .Z(n2982) );
  NOR U4513 ( .A(n2982), .B(n2981), .Z(n3276) );
  IV U4514 ( .A(n3276), .Z(n3270) );
  IV U4515 ( .A(n2983), .Z(n2984) );
  NOR U4516 ( .A(n2985), .B(n2984), .Z(n3549) );
  IV U4517 ( .A(n2986), .Z(n2988) );
  NOR U4518 ( .A(n2988), .B(n2987), .Z(n3751) );
  IV U4519 ( .A(n2989), .Z(n2990) );
  NOR U4520 ( .A(n2991), .B(n2990), .Z(n3566) );
  IV U4521 ( .A(n2992), .Z(n2994) );
  NOR U4522 ( .A(n2994), .B(n2993), .Z(n3748) );
  NOR U4523 ( .A(n3566), .B(n3748), .Z(n3247) );
  IV U4524 ( .A(n2995), .Z(n2997) );
  NOR U4525 ( .A(n2997), .B(n2996), .Z(n3226) );
  IV U4526 ( .A(n2998), .Z(n2999) );
  NOR U4527 ( .A(n3000), .B(n2999), .Z(n3224) );
  IV U4528 ( .A(n3224), .Z(n3214) );
  IV U4529 ( .A(n3001), .Z(n3002) );
  NOR U4530 ( .A(n3003), .B(n3002), .Z(n3209) );
  IV U4531 ( .A(n3004), .Z(n3005) );
  NOR U4532 ( .A(n3006), .B(n3005), .Z(n3722) );
  IV U4533 ( .A(n3007), .Z(n3008) );
  NOR U4534 ( .A(n3009), .B(n3008), .Z(n3569) );
  NOR U4535 ( .A(n3722), .B(n3569), .Z(n3194) );
  IV U4536 ( .A(n3010), .Z(n3011) );
  NOR U4537 ( .A(n3012), .B(n3011), .Z(n4603) );
  IV U4538 ( .A(n3013), .Z(n3014) );
  NOR U4539 ( .A(n3015), .B(n3014), .Z(n4604) );
  NOR U4540 ( .A(n4603), .B(n4604), .Z(n3713) );
  IV U4541 ( .A(n3016), .Z(n3017) );
  NOR U4542 ( .A(n3018), .B(n3017), .Z(n3577) );
  IV U4543 ( .A(n3019), .Z(n3021) );
  NOR U4544 ( .A(n3021), .B(n3020), .Z(n3705) );
  NOR U4545 ( .A(n3577), .B(n3705), .Z(n3178) );
  IV U4546 ( .A(n3022), .Z(n3023) );
  NOR U4547 ( .A(n3024), .B(n3023), .Z(n3693) );
  IV U4548 ( .A(n3025), .Z(n3026) );
  NOR U4549 ( .A(n3027), .B(n3026), .Z(n3679) );
  IV U4550 ( .A(n3028), .Z(n3030) );
  NOR U4551 ( .A(n3030), .B(n3029), .Z(n3593) );
  NOR U4552 ( .A(n3679), .B(n3593), .Z(n3140) );
  IV U4553 ( .A(n3031), .Z(n3033) );
  NOR U4554 ( .A(n3033), .B(n3032), .Z(n3138) );
  IV U4555 ( .A(n3138), .Z(n3132) );
  IV U4556 ( .A(n3034), .Z(n3036) );
  NOR U4557 ( .A(n3036), .B(n3035), .Z(n3598) );
  IV U4558 ( .A(n3037), .Z(n3039) );
  NOR U4559 ( .A(n3039), .B(n3038), .Z(n3602) );
  IV U4560 ( .A(n3040), .Z(n3042) );
  NOR U4561 ( .A(n3042), .B(n3041), .Z(n3670) );
  IV U4562 ( .A(n3043), .Z(n3044) );
  NOR U4563 ( .A(n3045), .B(n3044), .Z(n3619) );
  NOR U4564 ( .A(n3670), .B(n3619), .Z(n3109) );
  IV U4565 ( .A(n3046), .Z(n3047) );
  NOR U4566 ( .A(n3048), .B(n3047), .Z(n3086) );
  IV U4567 ( .A(n3086), .Z(n3081) );
  IV U4568 ( .A(n3049), .Z(n3050) );
  NOR U4569 ( .A(n3051), .B(n3050), .Z(n3645) );
  IV U4570 ( .A(n3052), .Z(n3053) );
  NOR U4571 ( .A(n3054), .B(n3053), .Z(n3067) );
  IV U4572 ( .A(n3055), .Z(n3057) );
  NOR U4573 ( .A(n3057), .B(n3056), .Z(n3061) );
  IV U4574 ( .A(n3058), .Z(n3060) );
  NOR U4575 ( .A(n3060), .B(n3059), .Z(n3068) );
  NOR U4576 ( .A(n3061), .B(n3068), .Z(n3062) );
  IV U4577 ( .A(n3062), .Z(n3063) );
  NOR U4578 ( .A(n3067), .B(n3063), .Z(n3072) );
  IV U4579 ( .A(n3064), .Z(n3065) );
  NOR U4580 ( .A(n3066), .B(n3065), .Z(n3074) );
  IV U4581 ( .A(n3067), .Z(n3070) );
  IV U4582 ( .A(n3068), .Z(n3069) );
  NOR U4583 ( .A(n3070), .B(n3069), .Z(n3641) );
  NOR U4584 ( .A(n3074), .B(n3641), .Z(n3071) );
  NOR U4585 ( .A(n3072), .B(n3071), .Z(n3652) );
  IV U4586 ( .A(n3072), .Z(n3073) );
  NOR U4587 ( .A(n3074), .B(n3073), .Z(n3075) );
  NOR U4588 ( .A(n3652), .B(n3075), .Z(n3642) );
  IV U4589 ( .A(n3076), .Z(n3077) );
  NOR U4590 ( .A(n3078), .B(n3077), .Z(n3079) );
  IV U4591 ( .A(n3079), .Z(n3644) );
  XOR U4592 ( .A(n3642), .B(n3644), .Z(n3646) );
  XOR U4593 ( .A(n3645), .B(n3646), .Z(n3080) );
  NOR U4594 ( .A(n3081), .B(n3080), .Z(n3637) );
  IV U4595 ( .A(n3082), .Z(n3083) );
  NOR U4596 ( .A(n3084), .B(n3083), .Z(n3638) );
  NOR U4597 ( .A(n3645), .B(n3638), .Z(n3085) );
  XOR U4598 ( .A(n3085), .B(n3646), .Z(n3633) );
  NOR U4599 ( .A(n3086), .B(n3633), .Z(n3087) );
  NOR U4600 ( .A(n3637), .B(n3087), .Z(n3626) );
  IV U4601 ( .A(n3088), .Z(n3089) );
  NOR U4602 ( .A(n3090), .B(n3089), .Z(n3632) );
  IV U4603 ( .A(n3091), .Z(n3092) );
  NOR U4604 ( .A(n3093), .B(n3092), .Z(n3627) );
  NOR U4605 ( .A(n3632), .B(n3627), .Z(n3094) );
  XOR U4606 ( .A(n3626), .B(n3094), .Z(n3662) );
  IV U4607 ( .A(n3095), .Z(n3096) );
  NOR U4608 ( .A(n3097), .B(n3096), .Z(n3624) );
  IV U4609 ( .A(n3098), .Z(n3099) );
  NOR U4610 ( .A(n3100), .B(n3099), .Z(n3660) );
  NOR U4611 ( .A(n3624), .B(n3660), .Z(n3101) );
  XOR U4612 ( .A(n3662), .B(n3101), .Z(n3622) );
  IV U4613 ( .A(n3102), .Z(n3104) );
  NOR U4614 ( .A(n3104), .B(n3103), .Z(n3621) );
  IV U4615 ( .A(n3105), .Z(n3107) );
  NOR U4616 ( .A(n3107), .B(n3106), .Z(n3667) );
  NOR U4617 ( .A(n3621), .B(n3667), .Z(n3108) );
  XOR U4618 ( .A(n3622), .B(n3108), .Z(n3671) );
  XOR U4619 ( .A(n3109), .B(n3671), .Z(n3614) );
  IV U4620 ( .A(n3110), .Z(n3111) );
  NOR U4621 ( .A(n3112), .B(n3111), .Z(n3616) );
  IV U4622 ( .A(n3113), .Z(n3115) );
  NOR U4623 ( .A(n3115), .B(n3114), .Z(n3613) );
  NOR U4624 ( .A(n3616), .B(n3613), .Z(n3116) );
  XOR U4625 ( .A(n3614), .B(n3116), .Z(n3612) );
  IV U4626 ( .A(n3117), .Z(n3119) );
  NOR U4627 ( .A(n3119), .B(n3118), .Z(n3610) );
  IV U4628 ( .A(n3120), .Z(n3122) );
  NOR U4629 ( .A(n3122), .B(n3121), .Z(n3608) );
  NOR U4630 ( .A(n3610), .B(n3608), .Z(n3123) );
  XOR U4631 ( .A(n3612), .B(n3123), .Z(n3606) );
  IV U4632 ( .A(n3124), .Z(n3126) );
  NOR U4633 ( .A(n3126), .B(n3125), .Z(n3674) );
  IV U4634 ( .A(n3127), .Z(n3129) );
  NOR U4635 ( .A(n3129), .B(n3128), .Z(n3605) );
  NOR U4636 ( .A(n3674), .B(n3605), .Z(n3130) );
  XOR U4637 ( .A(n3606), .B(n3130), .Z(n3604) );
  XOR U4638 ( .A(n3602), .B(n3604), .Z(n3599) );
  XOR U4639 ( .A(n3598), .B(n3599), .Z(n3131) );
  NOR U4640 ( .A(n3132), .B(n3131), .Z(n3683) );
  IV U4641 ( .A(n3133), .Z(n3134) );
  NOR U4642 ( .A(n3135), .B(n3134), .Z(n3596) );
  NOR U4643 ( .A(n3598), .B(n3596), .Z(n3136) );
  XOR U4644 ( .A(n3136), .B(n3599), .Z(n3137) );
  NOR U4645 ( .A(n3138), .B(n3137), .Z(n3139) );
  NOR U4646 ( .A(n3683), .B(n3139), .Z(n3594) );
  XOR U4647 ( .A(n3140), .B(n3594), .Z(n3591) );
  IV U4648 ( .A(n3141), .Z(n3143) );
  NOR U4649 ( .A(n3143), .B(n3142), .Z(n3590) );
  IV U4650 ( .A(n3144), .Z(n3145) );
  NOR U4651 ( .A(n3146), .B(n3145), .Z(n3588) );
  NOR U4652 ( .A(n3590), .B(n3588), .Z(n3147) );
  XOR U4653 ( .A(n3591), .B(n3147), .Z(n3582) );
  IV U4654 ( .A(n3148), .Z(n3149) );
  NOR U4655 ( .A(n3150), .B(n3149), .Z(n3585) );
  IV U4656 ( .A(n3151), .Z(n3152) );
  NOR U4657 ( .A(n3153), .B(n3152), .Z(n3583) );
  NOR U4658 ( .A(n3585), .B(n3583), .Z(n3154) );
  XOR U4659 ( .A(n3582), .B(n3154), .Z(n3694) );
  XOR U4660 ( .A(n3693), .B(n3694), .Z(n3701) );
  IV U4661 ( .A(n3701), .Z(n3162) );
  IV U4662 ( .A(n3155), .Z(n3157) );
  NOR U4663 ( .A(n3157), .B(n3156), .Z(n3686) );
  IV U4664 ( .A(n3158), .Z(n3160) );
  NOR U4665 ( .A(n3160), .B(n3159), .Z(n3700) );
  NOR U4666 ( .A(n3686), .B(n3700), .Z(n3161) );
  XOR U4667 ( .A(n3162), .B(n3161), .Z(n3581) );
  IV U4668 ( .A(n3163), .Z(n3165) );
  NOR U4669 ( .A(n3165), .B(n3164), .Z(n3166) );
  IV U4670 ( .A(n3166), .Z(n3174) );
  NOR U4671 ( .A(n3581), .B(n3174), .Z(n4189) );
  IV U4672 ( .A(n3167), .Z(n3168) );
  NOR U4673 ( .A(n3169), .B(n3168), .Z(n3573) );
  IV U4674 ( .A(n3170), .Z(n3172) );
  NOR U4675 ( .A(n3172), .B(n3171), .Z(n3173) );
  IV U4676 ( .A(n3173), .Z(n3580) );
  XOR U4677 ( .A(n3580), .B(n3581), .Z(n3574) );
  XOR U4678 ( .A(n3573), .B(n3574), .Z(n3176) );
  NOR U4679 ( .A(n3574), .B(n3174), .Z(n3175) );
  NOR U4680 ( .A(n3176), .B(n3175), .Z(n3177) );
  NOR U4681 ( .A(n4189), .B(n3177), .Z(n3578) );
  XOR U4682 ( .A(n3178), .B(n3578), .Z(n3710) );
  IV U4683 ( .A(n3179), .Z(n3181) );
  NOR U4684 ( .A(n3181), .B(n3180), .Z(n3708) );
  IV U4685 ( .A(n3182), .Z(n3183) );
  NOR U4686 ( .A(n3184), .B(n3183), .Z(n3571) );
  NOR U4687 ( .A(n3708), .B(n3571), .Z(n3185) );
  XOR U4688 ( .A(n3710), .B(n3185), .Z(n3186) );
  IV U4689 ( .A(n3186), .Z(n4205) );
  XOR U4690 ( .A(n3713), .B(n4205), .Z(n3715) );
  IV U4691 ( .A(n3187), .Z(n3189) );
  NOR U4692 ( .A(n3189), .B(n3188), .Z(n3714) );
  IV U4693 ( .A(n3190), .Z(n3192) );
  NOR U4694 ( .A(n3192), .B(n3191), .Z(n3719) );
  NOR U4695 ( .A(n3714), .B(n3719), .Z(n3193) );
  XOR U4696 ( .A(n3715), .B(n3193), .Z(n3723) );
  XOR U4697 ( .A(n3194), .B(n3723), .Z(n3727) );
  IV U4698 ( .A(n3195), .Z(n3196) );
  NOR U4699 ( .A(n3197), .B(n3196), .Z(n3726) );
  IV U4700 ( .A(n3198), .Z(n3200) );
  NOR U4701 ( .A(n3200), .B(n3199), .Z(n3729) );
  NOR U4702 ( .A(n3726), .B(n3729), .Z(n3201) );
  XOR U4703 ( .A(n3727), .B(n3201), .Z(n3736) );
  IV U4704 ( .A(n3202), .Z(n3204) );
  NOR U4705 ( .A(n3204), .B(n3203), .Z(n3734) );
  IV U4706 ( .A(n3205), .Z(n3207) );
  NOR U4707 ( .A(n3207), .B(n3206), .Z(n3732) );
  NOR U4708 ( .A(n3734), .B(n3732), .Z(n3208) );
  XOR U4709 ( .A(n3736), .B(n3208), .Z(n3220) );
  NOR U4710 ( .A(n3209), .B(n3220), .Z(n3212) );
  IV U4711 ( .A(n3209), .Z(n3211) );
  XOR U4712 ( .A(n3734), .B(n3736), .Z(n3210) );
  NOR U4713 ( .A(n3211), .B(n3210), .Z(n3739) );
  NOR U4714 ( .A(n3212), .B(n3739), .Z(n3218) );
  IV U4715 ( .A(n3218), .Z(n3213) );
  NOR U4716 ( .A(n3214), .B(n3213), .Z(n3568) );
  IV U4717 ( .A(n3215), .Z(n3216) );
  NOR U4718 ( .A(n3217), .B(n3216), .Z(n3219) );
  NOR U4719 ( .A(n3219), .B(n3218), .Z(n3223) );
  IV U4720 ( .A(n3219), .Z(n3222) );
  IV U4721 ( .A(n3220), .Z(n3221) );
  NOR U4722 ( .A(n3222), .B(n3221), .Z(n4095) );
  NOR U4723 ( .A(n3223), .B(n4095), .Z(n3227) );
  NOR U4724 ( .A(n3224), .B(n3227), .Z(n3225) );
  NOR U4725 ( .A(n3568), .B(n3225), .Z(n3237) );
  NOR U4726 ( .A(n3226), .B(n3237), .Z(n3230) );
  IV U4727 ( .A(n3226), .Z(n3229) );
  IV U4728 ( .A(n3227), .Z(n3228) );
  NOR U4729 ( .A(n3229), .B(n3228), .Z(n3744) );
  NOR U4730 ( .A(n3230), .B(n3744), .Z(n3563) );
  IV U4731 ( .A(n3231), .Z(n3233) );
  NOR U4732 ( .A(n3233), .B(n3232), .Z(n3244) );
  IV U4733 ( .A(n3244), .Z(n3565) );
  NOR U4734 ( .A(n3563), .B(n3565), .Z(n3246) );
  IV U4735 ( .A(n3234), .Z(n3235) );
  NOR U4736 ( .A(n3236), .B(n3235), .Z(n3240) );
  IV U4737 ( .A(n3240), .Z(n3239) );
  IV U4738 ( .A(n3237), .Z(n3238) );
  NOR U4739 ( .A(n3239), .B(n3238), .Z(n4244) );
  NOR U4740 ( .A(n3563), .B(n3240), .Z(n3241) );
  NOR U4741 ( .A(n4244), .B(n3241), .Z(n3242) );
  IV U4742 ( .A(n3242), .Z(n3243) );
  NOR U4743 ( .A(n3244), .B(n3243), .Z(n3245) );
  NOR U4744 ( .A(n3246), .B(n3245), .Z(n3749) );
  XOR U4745 ( .A(n3247), .B(n3749), .Z(n3746) );
  XOR U4746 ( .A(n3751), .B(n3746), .Z(n3758) );
  IV U4747 ( .A(n3248), .Z(n3250) );
  NOR U4748 ( .A(n3250), .B(n3249), .Z(n3745) );
  IV U4749 ( .A(n3251), .Z(n3253) );
  NOR U4750 ( .A(n3253), .B(n3252), .Z(n3757) );
  NOR U4751 ( .A(n3745), .B(n3757), .Z(n3254) );
  XOR U4752 ( .A(n3758), .B(n3254), .Z(n3562) );
  IV U4753 ( .A(n3255), .Z(n3257) );
  NOR U4754 ( .A(n3257), .B(n3256), .Z(n3560) );
  IV U4755 ( .A(n3258), .Z(n3260) );
  NOR U4756 ( .A(n3260), .B(n3259), .Z(n3558) );
  NOR U4757 ( .A(n3560), .B(n3558), .Z(n3261) );
  XOR U4758 ( .A(n3562), .B(n3261), .Z(n3553) );
  IV U4759 ( .A(n3262), .Z(n3264) );
  NOR U4760 ( .A(n3264), .B(n3263), .Z(n3555) );
  IV U4761 ( .A(n3265), .Z(n3267) );
  NOR U4762 ( .A(n3267), .B(n3266), .Z(n3552) );
  NOR U4763 ( .A(n3555), .B(n3552), .Z(n3268) );
  XOR U4764 ( .A(n3553), .B(n3268), .Z(n3551) );
  XOR U4765 ( .A(n3549), .B(n3551), .Z(n3269) );
  NOR U4766 ( .A(n3270), .B(n3269), .Z(n4077) );
  IV U4767 ( .A(n3271), .Z(n3272) );
  NOR U4768 ( .A(n3273), .B(n3272), .Z(n3547) );
  NOR U4769 ( .A(n3549), .B(n3547), .Z(n3274) );
  XOR U4770 ( .A(n3551), .B(n3274), .Z(n3275) );
  NOR U4771 ( .A(n3276), .B(n3275), .Z(n3277) );
  NOR U4772 ( .A(n4077), .B(n3277), .Z(n3765) );
  IV U4773 ( .A(n3278), .Z(n3280) );
  NOR U4774 ( .A(n3280), .B(n3279), .Z(n3767) );
  IV U4775 ( .A(n3281), .Z(n3282) );
  NOR U4776 ( .A(n3283), .B(n3282), .Z(n3764) );
  NOR U4777 ( .A(n3767), .B(n3764), .Z(n3284) );
  XOR U4778 ( .A(n3765), .B(n3284), .Z(n3545) );
  XOR U4779 ( .A(n3285), .B(n3545), .Z(n3777) );
  XOR U4780 ( .A(n3778), .B(n3777), .Z(n3540) );
  IV U4781 ( .A(n3286), .Z(n3287) );
  NOR U4782 ( .A(n3288), .B(n3287), .Z(n3780) );
  IV U4783 ( .A(n3289), .Z(n3290) );
  NOR U4784 ( .A(n3291), .B(n3290), .Z(n3539) );
  NOR U4785 ( .A(n3780), .B(n3539), .Z(n3292) );
  XOR U4786 ( .A(n3540), .B(n3292), .Z(n3293) );
  IV U4787 ( .A(n3293), .Z(n4068) );
  XOR U4788 ( .A(n3787), .B(n4068), .Z(n4063) );
  XOR U4789 ( .A(n3789), .B(n4063), .Z(n3532) );
  IV U4790 ( .A(n3294), .Z(n3296) );
  NOR U4791 ( .A(n3296), .B(n3295), .Z(n3536) );
  IV U4792 ( .A(n3297), .Z(n3299) );
  NOR U4793 ( .A(n3299), .B(n3298), .Z(n3531) );
  NOR U4794 ( .A(n3536), .B(n3531), .Z(n3300) );
  XOR U4795 ( .A(n3532), .B(n3300), .Z(n3796) );
  XOR U4796 ( .A(n3301), .B(n3796), .Z(n3528) );
  XOR U4797 ( .A(n3302), .B(n3528), .Z(n4297) );
  XOR U4798 ( .A(n4308), .B(n4297), .Z(n3523) );
  XOR U4799 ( .A(n3303), .B(n3523), .Z(n3520) );
  XOR U4800 ( .A(n3521), .B(n3520), .Z(n3517) );
  XOR U4801 ( .A(n3516), .B(n3517), .Z(n3304) );
  NOR U4802 ( .A(n3305), .B(n3304), .Z(n4318) );
  IV U4803 ( .A(n3306), .Z(n3308) );
  NOR U4804 ( .A(n3308), .B(n3307), .Z(n3514) );
  NOR U4805 ( .A(n3516), .B(n3514), .Z(n3309) );
  XOR U4806 ( .A(n3309), .B(n3517), .Z(n3314) );
  NOR U4807 ( .A(n3310), .B(n3314), .Z(n3311) );
  NOR U4808 ( .A(n4318), .B(n3311), .Z(n3312) );
  NOR U4809 ( .A(n3313), .B(n3312), .Z(n3317) );
  IV U4810 ( .A(n3313), .Z(n3316) );
  IV U4811 ( .A(n3314), .Z(n3315) );
  NOR U4812 ( .A(n3316), .B(n3315), .Z(n4321) );
  NOR U4813 ( .A(n3317), .B(n4321), .Z(n3509) );
  XOR U4814 ( .A(n3513), .B(n3509), .Z(n3802) );
  IV U4815 ( .A(n3318), .Z(n3319) );
  NOR U4816 ( .A(n3320), .B(n3319), .Z(n3508) );
  IV U4817 ( .A(n3321), .Z(n3323) );
  NOR U4818 ( .A(n3323), .B(n3322), .Z(n3801) );
  NOR U4819 ( .A(n3508), .B(n3801), .Z(n3324) );
  XOR U4820 ( .A(n3802), .B(n3324), .Z(n3325) );
  IV U4821 ( .A(n3325), .Z(n3507) );
  XOR U4822 ( .A(n3505), .B(n3507), .Z(n3808) );
  XOR U4823 ( .A(n3326), .B(n3808), .Z(n3500) );
  IV U4824 ( .A(n3327), .Z(n3329) );
  NOR U4825 ( .A(n3329), .B(n3328), .Z(n3804) );
  IV U4826 ( .A(n3330), .Z(n3332) );
  NOR U4827 ( .A(n3332), .B(n3331), .Z(n3501) );
  NOR U4828 ( .A(n3804), .B(n3501), .Z(n3333) );
  XOR U4829 ( .A(n3500), .B(n3333), .Z(n3498) );
  XOR U4830 ( .A(n3334), .B(n3498), .Z(n3490) );
  IV U4831 ( .A(n3335), .Z(n3337) );
  NOR U4832 ( .A(n3337), .B(n3336), .Z(n3492) );
  IV U4833 ( .A(n3338), .Z(n3340) );
  NOR U4834 ( .A(n3340), .B(n3339), .Z(n3489) );
  NOR U4835 ( .A(n3492), .B(n3489), .Z(n3341) );
  XOR U4836 ( .A(n3490), .B(n3341), .Z(n3816) );
  IV U4837 ( .A(n3342), .Z(n3344) );
  NOR U4838 ( .A(n3344), .B(n3343), .Z(n3814) );
  IV U4839 ( .A(n3345), .Z(n3347) );
  NOR U4840 ( .A(n3347), .B(n3346), .Z(n3812) );
  NOR U4841 ( .A(n3814), .B(n3812), .Z(n3348) );
  XOR U4842 ( .A(n3816), .B(n3348), .Z(n3483) );
  IV U4843 ( .A(n3349), .Z(n3351) );
  NOR U4844 ( .A(n3351), .B(n3350), .Z(n3486) );
  IV U4845 ( .A(n3352), .Z(n3353) );
  NOR U4846 ( .A(n3354), .B(n3353), .Z(n3482) );
  NOR U4847 ( .A(n3486), .B(n3482), .Z(n3355) );
  XOR U4848 ( .A(n3483), .B(n3355), .Z(n3823) );
  IV U4849 ( .A(n3356), .Z(n3357) );
  NOR U4850 ( .A(n3358), .B(n3357), .Z(n3819) );
  IV U4851 ( .A(n3359), .Z(n3360) );
  NOR U4852 ( .A(n3361), .B(n3360), .Z(n3821) );
  NOR U4853 ( .A(n3819), .B(n3821), .Z(n3362) );
  XOR U4854 ( .A(n3823), .B(n3362), .Z(n3479) );
  IV U4855 ( .A(n3363), .Z(n3365) );
  NOR U4856 ( .A(n3365), .B(n3364), .Z(n3826) );
  IV U4857 ( .A(n3366), .Z(n3368) );
  NOR U4858 ( .A(n3368), .B(n3367), .Z(n3824) );
  NOR U4859 ( .A(n3826), .B(n3824), .Z(n3369) );
  XOR U4860 ( .A(n3479), .B(n3369), .Z(n3476) );
  XOR U4861 ( .A(n3370), .B(n3476), .Z(n3470) );
  XOR U4862 ( .A(n3371), .B(n3470), .Z(n3838) );
  IV U4863 ( .A(n3372), .Z(n3373) );
  NOR U4864 ( .A(n3374), .B(n3373), .Z(n3832) );
  IV U4865 ( .A(n3375), .Z(n3376) );
  NOR U4866 ( .A(n3377), .B(n3376), .Z(n3837) );
  NOR U4867 ( .A(n3832), .B(n3837), .Z(n3378) );
  XOR U4868 ( .A(n3838), .B(n3378), .Z(n3466) );
  XOR U4869 ( .A(n3379), .B(n3466), .Z(n3858) );
  XOR U4870 ( .A(n3380), .B(n3858), .Z(n3463) );
  IV U4871 ( .A(n3381), .Z(n3383) );
  NOR U4872 ( .A(n3383), .B(n3382), .Z(n3857) );
  IV U4873 ( .A(n3384), .Z(n3386) );
  NOR U4874 ( .A(n3386), .B(n3385), .Z(n3462) );
  NOR U4875 ( .A(n3857), .B(n3462), .Z(n3387) );
  XOR U4876 ( .A(n3463), .B(n3387), .Z(n3461) );
  XOR U4877 ( .A(n3459), .B(n3461), .Z(n3388) );
  NOR U4878 ( .A(n3389), .B(n3388), .Z(n3980) );
  IV U4879 ( .A(n3390), .Z(n3392) );
  NOR U4880 ( .A(n3392), .B(n3391), .Z(n3457) );
  NOR U4881 ( .A(n3459), .B(n3457), .Z(n3393) );
  XOR U4882 ( .A(n3461), .B(n3393), .Z(n3394) );
  NOR U4883 ( .A(n3395), .B(n3394), .Z(n3396) );
  NOR U4884 ( .A(n3980), .B(n3396), .Z(n3862) );
  XOR U4885 ( .A(n3863), .B(n3862), .Z(n3870) );
  IV U4886 ( .A(n3397), .Z(n3398) );
  NOR U4887 ( .A(n3399), .B(n3398), .Z(n3864) );
  IV U4888 ( .A(n3400), .Z(n3402) );
  NOR U4889 ( .A(n3402), .B(n3401), .Z(n3869) );
  NOR U4890 ( .A(n3864), .B(n3869), .Z(n3403) );
  XOR U4891 ( .A(n3870), .B(n3403), .Z(n3404) );
  IV U4892 ( .A(n3404), .Z(n3455) );
  XOR U4893 ( .A(n3451), .B(n3455), .Z(n3449) );
  XOR U4894 ( .A(n3405), .B(n3449), .Z(n3873) );
  XOR U4895 ( .A(n3874), .B(n3873), .Z(n3880) );
  XOR U4896 ( .A(n3875), .B(n3880), .Z(n3406) );
  NOR U4897 ( .A(n3407), .B(n3406), .Z(n3938) );
  IV U4898 ( .A(n3408), .Z(n3409) );
  NOR U4899 ( .A(n3410), .B(n3409), .Z(n3879) );
  NOR U4900 ( .A(n3875), .B(n3879), .Z(n3411) );
  XOR U4901 ( .A(n3411), .B(n3880), .Z(n3412) );
  NOR U4902 ( .A(n3413), .B(n3412), .Z(n3414) );
  NOR U4903 ( .A(n3938), .B(n3414), .Z(n3443) );
  XOR U4904 ( .A(n3447), .B(n3443), .Z(n3887) );
  IV U4905 ( .A(n3415), .Z(n3416) );
  NOR U4906 ( .A(n3417), .B(n3416), .Z(n3442) );
  IV U4907 ( .A(n3418), .Z(n3419) );
  NOR U4908 ( .A(n3420), .B(n3419), .Z(n3886) );
  NOR U4909 ( .A(n3442), .B(n3886), .Z(n3421) );
  XOR U4910 ( .A(n3887), .B(n3421), .Z(n3438) );
  XOR U4911 ( .A(n3422), .B(n3438), .Z(n4850) );
  XOR U4912 ( .A(n4856), .B(n4850), .Z(n3892) );
  XOR U4913 ( .A(n3893), .B(n3892), .Z(n4390) );
  IV U4914 ( .A(n3423), .Z(n3425) );
  NOR U4915 ( .A(n3425), .B(n3424), .Z(n4398) );
  IV U4916 ( .A(n3426), .Z(n3428) );
  NOR U4917 ( .A(n3428), .B(n3427), .Z(n4393) );
  NOR U4918 ( .A(n4398), .B(n4393), .Z(n3890) );
  XOR U4919 ( .A(n4390), .B(n3890), .Z(n3898) );
  IV U4920 ( .A(n3429), .Z(n3431) );
  NOR U4921 ( .A(n3431), .B(n3430), .Z(n3923) );
  IV U4922 ( .A(n3432), .Z(n3434) );
  NOR U4923 ( .A(n3434), .B(n3433), .Z(n3921) );
  NOR U4924 ( .A(n3923), .B(n3921), .Z(n3899) );
  XOR U4925 ( .A(n3898), .B(n3899), .Z(n3902) );
  XOR U4926 ( .A(n3900), .B(n3902), .Z(n3907) );
  XOR U4927 ( .A(n3905), .B(n3907), .Z(n3910) );
  XOR U4928 ( .A(n3435), .B(n3910), .Z(o[1]) );
  IV U4929 ( .A(n3436), .Z(n3437) );
  NOR U4930 ( .A(n3907), .B(n3437), .Z(n3912) );
  NOR U4931 ( .A(n4856), .B(n4850), .Z(n3894) );
  IV U4932 ( .A(n3438), .Z(n3885) );
  IV U4933 ( .A(n3439), .Z(n3440) );
  NOR U4934 ( .A(n3885), .B(n3440), .Z(n3441) );
  IV U4935 ( .A(n3441), .Z(n4428) );
  IV U4936 ( .A(n3442), .Z(n3444) );
  IV U4937 ( .A(n3443), .Z(n3446) );
  NOR U4938 ( .A(n3444), .B(n3446), .Z(n3445) );
  IV U4939 ( .A(n3445), .Z(n3934) );
  NOR U4940 ( .A(n3447), .B(n3446), .Z(n3936) );
  NOR U4941 ( .A(n3938), .B(n3936), .Z(n3882) );
  IV U4942 ( .A(n3448), .Z(n3450) );
  NOR U4943 ( .A(n3450), .B(n3449), .Z(n3959) );
  IV U4944 ( .A(n3451), .Z(n3452) );
  NOR U4945 ( .A(n3455), .B(n3452), .Z(n3964) );
  IV U4946 ( .A(n3453), .Z(n3454) );
  NOR U4947 ( .A(n3455), .B(n3454), .Z(n3956) );
  XOR U4948 ( .A(n3964), .B(n3956), .Z(n3456) );
  NOR U4949 ( .A(n3959), .B(n3456), .Z(n3872) );
  IV U4950 ( .A(n3457), .Z(n3458) );
  NOR U4951 ( .A(n3461), .B(n3458), .Z(n3977) );
  IV U4952 ( .A(n3459), .Z(n3460) );
  NOR U4953 ( .A(n3461), .B(n3460), .Z(n3983) );
  IV U4954 ( .A(n3462), .Z(n3465) );
  IV U4955 ( .A(n3463), .Z(n3464) );
  NOR U4956 ( .A(n3465), .B(n3464), .Z(n4366) );
  IV U4957 ( .A(n3466), .Z(n3844) );
  IV U4958 ( .A(n3467), .Z(n3468) );
  NOR U4959 ( .A(n3844), .B(n3468), .Z(n3469) );
  IV U4960 ( .A(n3469), .Z(n3849) );
  IV U4961 ( .A(n3470), .Z(n3833) );
  IV U4962 ( .A(n3471), .Z(n3472) );
  NOR U4963 ( .A(n3833), .B(n3472), .Z(n3473) );
  IV U4964 ( .A(n3473), .Z(n3995) );
  IV U4965 ( .A(n3834), .Z(n3474) );
  NOR U4966 ( .A(n3833), .B(n3474), .Z(n3999) );
  IV U4967 ( .A(n3475), .Z(n3477) );
  NOR U4968 ( .A(n3477), .B(n3476), .Z(n4001) );
  NOR U4969 ( .A(n3999), .B(n4001), .Z(n3831) );
  IV U4970 ( .A(n3478), .Z(n3481) );
  IV U4971 ( .A(n3479), .Z(n3827) );
  XOR U4972 ( .A(n3826), .B(n3827), .Z(n3480) );
  NOR U4973 ( .A(n3481), .B(n3480), .Z(n4004) );
  IV U4974 ( .A(n3482), .Z(n3485) );
  IV U4975 ( .A(n3483), .Z(n3484) );
  NOR U4976 ( .A(n3485), .B(n3484), .Z(n4016) );
  IV U4977 ( .A(n3486), .Z(n3488) );
  XOR U4978 ( .A(n3814), .B(n3816), .Z(n3487) );
  NOR U4979 ( .A(n3488), .B(n3487), .Z(n4013) );
  IV U4980 ( .A(n3489), .Z(n3491) );
  IV U4981 ( .A(n3490), .Z(n3493) );
  NOR U4982 ( .A(n3491), .B(n3493), .Z(n4024) );
  IV U4983 ( .A(n3492), .Z(n3494) );
  NOR U4984 ( .A(n3494), .B(n3493), .Z(n4030) );
  IV U4985 ( .A(n3495), .Z(n3496) );
  NOR U4986 ( .A(n3496), .B(n3498), .Z(n4027) );
  IV U4987 ( .A(n3497), .Z(n3499) );
  NOR U4988 ( .A(n3499), .B(n3498), .Z(n4036) );
  IV U4989 ( .A(n3500), .Z(n3806) );
  IV U4990 ( .A(n3501), .Z(n3502) );
  NOR U4991 ( .A(n3806), .B(n3502), .Z(n4033) );
  IV U4992 ( .A(n3503), .Z(n3504) );
  NOR U4993 ( .A(n3507), .B(n3504), .Z(n4336) );
  IV U4994 ( .A(n3505), .Z(n3506) );
  NOR U4995 ( .A(n3507), .B(n3506), .Z(n4325) );
  IV U4996 ( .A(n3508), .Z(n3510) );
  IV U4997 ( .A(n3509), .Z(n3512) );
  NOR U4998 ( .A(n3510), .B(n3512), .Z(n3511) );
  IV U4999 ( .A(n3511), .Z(n4330) );
  NOR U5000 ( .A(n3513), .B(n3512), .Z(n4045) );
  NOR U5001 ( .A(n4321), .B(n4045), .Z(n3800) );
  IV U5002 ( .A(n3514), .Z(n3515) );
  NOR U5003 ( .A(n3515), .B(n3517), .Z(n4048) );
  IV U5004 ( .A(n3516), .Z(n3518) );
  NOR U5005 ( .A(n3518), .B(n3517), .Z(n4052) );
  XOR U5006 ( .A(n4048), .B(n4052), .Z(n3519) );
  NOR U5007 ( .A(n4318), .B(n3519), .Z(n3799) );
  IV U5008 ( .A(n3520), .Z(n4055) );
  NOR U5009 ( .A(n4055), .B(n3521), .Z(n3525) );
  IV U5010 ( .A(n3522), .Z(n3524) );
  NOR U5011 ( .A(n3524), .B(n3523), .Z(n4313) );
  NOR U5012 ( .A(n3525), .B(n4313), .Z(n3798) );
  NOR U5013 ( .A(n4308), .B(n3526), .Z(n3527) );
  NOR U5014 ( .A(n3527), .B(n4297), .Z(n4303) );
  IV U5015 ( .A(n3528), .Z(n3794) );
  IV U5016 ( .A(n3529), .Z(n3530) );
  NOR U5017 ( .A(n3794), .B(n3530), .Z(n4295) );
  IV U5018 ( .A(n3531), .Z(n3533) );
  IV U5019 ( .A(n3532), .Z(n3537) );
  NOR U5020 ( .A(n3533), .B(n3537), .Z(n4554) );
  IV U5021 ( .A(n3534), .Z(n3535) );
  NOR U5022 ( .A(n3535), .B(n3796), .Z(n4549) );
  NOR U5023 ( .A(n4554), .B(n4549), .Z(n4289) );
  IV U5024 ( .A(n3536), .Z(n3538) );
  NOR U5025 ( .A(n3538), .B(n3537), .Z(n4058) );
  IV U5026 ( .A(n3539), .Z(n3541) );
  NOR U5027 ( .A(n3541), .B(n3540), .Z(n3785) );
  IV U5028 ( .A(n3785), .Z(n3776) );
  IV U5029 ( .A(n3542), .Z(n3543) );
  NOR U5030 ( .A(n3543), .B(n3545), .Z(n4075) );
  IV U5031 ( .A(n3544), .Z(n3546) );
  NOR U5032 ( .A(n3546), .B(n3545), .Z(n3772) );
  IV U5033 ( .A(n3772), .Z(n3763) );
  IV U5034 ( .A(n3547), .Z(n3548) );
  NOR U5035 ( .A(n3551), .B(n3548), .Z(n4265) );
  IV U5036 ( .A(n3549), .Z(n3550) );
  NOR U5037 ( .A(n3551), .B(n3550), .Z(n4580) );
  IV U5038 ( .A(n3552), .Z(n3554) );
  IV U5039 ( .A(n3553), .Z(n3556) );
  NOR U5040 ( .A(n3554), .B(n3556), .Z(n4756) );
  NOR U5041 ( .A(n4580), .B(n4756), .Z(n4081) );
  IV U5042 ( .A(n3555), .Z(n3557) );
  NOR U5043 ( .A(n3557), .B(n3556), .Z(n4082) );
  IV U5044 ( .A(n3558), .Z(n3559) );
  NOR U5045 ( .A(n3562), .B(n3559), .Z(n4257) );
  NOR U5046 ( .A(n4082), .B(n4257), .Z(n3761) );
  IV U5047 ( .A(n3560), .Z(n3561) );
  NOR U5048 ( .A(n3562), .B(n3561), .Z(n4254) );
  IV U5049 ( .A(n3563), .Z(n3564) );
  NOR U5050 ( .A(n3565), .B(n3564), .Z(n4723) );
  IV U5051 ( .A(n3566), .Z(n3567) );
  NOR U5052 ( .A(n3567), .B(n3749), .Z(n4732) );
  NOR U5053 ( .A(n4723), .B(n4732), .Z(n4247) );
  IV U5054 ( .A(n3568), .Z(n3740) );
  IV U5055 ( .A(n3569), .Z(n3570) );
  NOR U5056 ( .A(n3570), .B(n3723), .Z(n4101) );
  IV U5057 ( .A(n3571), .Z(n3572) );
  NOR U5058 ( .A(n3710), .B(n3572), .Z(n4199) );
  IV U5059 ( .A(n3573), .Z(n3576) );
  IV U5060 ( .A(n3574), .Z(n3575) );
  NOR U5061 ( .A(n3576), .B(n3575), .Z(n4685) );
  IV U5062 ( .A(n3577), .Z(n3579) );
  IV U5063 ( .A(n3578), .Z(n3706) );
  NOR U5064 ( .A(n3579), .B(n3706), .Z(n4693) );
  NOR U5065 ( .A(n4685), .B(n4693), .Z(n4193) );
  NOR U5066 ( .A(n3581), .B(n3580), .Z(n4110) );
  NOR U5067 ( .A(n4110), .B(n4189), .Z(n3704) );
  IV U5068 ( .A(n3582), .Z(n3587) );
  IV U5069 ( .A(n3583), .Z(n3584) );
  NOR U5070 ( .A(n3587), .B(n3584), .Z(n3689) );
  IV U5071 ( .A(n3585), .Z(n3586) );
  NOR U5072 ( .A(n3587), .B(n3586), .Z(n4115) );
  IV U5073 ( .A(n3588), .Z(n3589) );
  NOR U5074 ( .A(n3589), .B(n3591), .Z(n4120) );
  NOR U5075 ( .A(n4115), .B(n4120), .Z(n3685) );
  IV U5076 ( .A(n3590), .Z(n3592) );
  NOR U5077 ( .A(n3592), .B(n3591), .Z(n4117) );
  IV U5078 ( .A(n3593), .Z(n3595) );
  IV U5079 ( .A(n3594), .Z(n3680) );
  NOR U5080 ( .A(n3595), .B(n3680), .Z(n4126) );
  IV U5081 ( .A(n3596), .Z(n3597) );
  NOR U5082 ( .A(n3597), .B(n3599), .Z(n4176) );
  IV U5083 ( .A(n3598), .Z(n3600) );
  NOR U5084 ( .A(n3600), .B(n3599), .Z(n3601) );
  IV U5085 ( .A(n3601), .Z(n4174) );
  IV U5086 ( .A(n3602), .Z(n3603) );
  NOR U5087 ( .A(n3604), .B(n3603), .Z(n4129) );
  IV U5088 ( .A(n3605), .Z(n3607) );
  IV U5089 ( .A(n3606), .Z(n3675) );
  NOR U5090 ( .A(n3607), .B(n3675), .Z(n4170) );
  NOR U5091 ( .A(n4129), .B(n4170), .Z(n3678) );
  IV U5092 ( .A(n3608), .Z(n3609) );
  NOR U5093 ( .A(n3612), .B(n3609), .Z(n4131) );
  IV U5094 ( .A(n3610), .Z(n3611) );
  NOR U5095 ( .A(n3612), .B(n3611), .Z(n4141) );
  IV U5096 ( .A(n3613), .Z(n3615) );
  IV U5097 ( .A(n3614), .Z(n3617) );
  NOR U5098 ( .A(n3615), .B(n3617), .Z(n4138) );
  IV U5099 ( .A(n3616), .Z(n3618) );
  NOR U5100 ( .A(n3618), .B(n3617), .Z(n4149) );
  IV U5101 ( .A(n3619), .Z(n3620) );
  NOR U5102 ( .A(n3620), .B(n3671), .Z(n4146) );
  IV U5103 ( .A(n3621), .Z(n3623) );
  IV U5104 ( .A(n3622), .Z(n3668) );
  NOR U5105 ( .A(n3623), .B(n3668), .Z(n3666) );
  IV U5106 ( .A(n3666), .Z(n3659) );
  IV U5107 ( .A(n3624), .Z(n3625) );
  NOR U5108 ( .A(n3662), .B(n3625), .Z(n3631) );
  IV U5109 ( .A(n3626), .Z(n3629) );
  IV U5110 ( .A(n3627), .Z(n3628) );
  NOR U5111 ( .A(n3629), .B(n3628), .Z(n3630) );
  NOR U5112 ( .A(n3631), .B(n3630), .Z(n4166) );
  IV U5113 ( .A(n3632), .Z(n3635) );
  IV U5114 ( .A(n3633), .Z(n3634) );
  NOR U5115 ( .A(n3635), .B(n3634), .Z(n3636) );
  NOR U5116 ( .A(n3637), .B(n3636), .Z(n3657) );
  IV U5117 ( .A(n3638), .Z(n3639) );
  NOR U5118 ( .A(n3639), .B(n3646), .Z(n3653) );
  IV U5119 ( .A(n3653), .Z(n3640) );
  NOR U5120 ( .A(n3641), .B(n3640), .Z(n3655) );
  IV U5121 ( .A(n3642), .Z(n3643) );
  NOR U5122 ( .A(n3644), .B(n3643), .Z(n3649) );
  IV U5123 ( .A(n3645), .Z(n3647) );
  NOR U5124 ( .A(n3647), .B(n3646), .Z(n3648) );
  NOR U5125 ( .A(n3649), .B(n3648), .Z(n3650) );
  IV U5126 ( .A(n3650), .Z(n3651) );
  NOR U5127 ( .A(n3652), .B(n3651), .Z(n4163) );
  NOR U5128 ( .A(n3653), .B(n4163), .Z(n3654) );
  NOR U5129 ( .A(n3655), .B(n3654), .Z(n3656) );
  XOR U5130 ( .A(n3657), .B(n3656), .Z(n4164) );
  XOR U5131 ( .A(n4166), .B(n4164), .Z(n3658) );
  NOR U5132 ( .A(n3659), .B(n3658), .Z(n4162) );
  IV U5133 ( .A(n4164), .Z(n4167) );
  IV U5134 ( .A(n4166), .Z(n3663) );
  IV U5135 ( .A(n3660), .Z(n3661) );
  NOR U5136 ( .A(n3662), .B(n3661), .Z(n4165) );
  NOR U5137 ( .A(n3663), .B(n4165), .Z(n3664) );
  XOR U5138 ( .A(n4167), .B(n3664), .Z(n3665) );
  NOR U5139 ( .A(n3666), .B(n3665), .Z(n4159) );
  NOR U5140 ( .A(n4162), .B(n4159), .Z(n4155) );
  IV U5141 ( .A(n3667), .Z(n3669) );
  NOR U5142 ( .A(n3669), .B(n3668), .Z(n4158) );
  IV U5143 ( .A(n3670), .Z(n3672) );
  NOR U5144 ( .A(n3672), .B(n3671), .Z(n4154) );
  NOR U5145 ( .A(n4158), .B(n4154), .Z(n3673) );
  XOR U5146 ( .A(n4155), .B(n3673), .Z(n4148) );
  XOR U5147 ( .A(n4146), .B(n4148), .Z(n4151) );
  XOR U5148 ( .A(n4149), .B(n4151), .Z(n4140) );
  XOR U5149 ( .A(n4138), .B(n4140), .Z(n4143) );
  XOR U5150 ( .A(n4141), .B(n4143), .Z(n4132) );
  XOR U5151 ( .A(n4131), .B(n4132), .Z(n4172) );
  IV U5152 ( .A(n3674), .Z(n3676) );
  NOR U5153 ( .A(n3676), .B(n3675), .Z(n4134) );
  XOR U5154 ( .A(n4172), .B(n4134), .Z(n3677) );
  XOR U5155 ( .A(n3678), .B(n3677), .Z(n4173) );
  XOR U5156 ( .A(n4174), .B(n4173), .Z(n4177) );
  XOR U5157 ( .A(n4176), .B(n4177), .Z(n4124) );
  IV U5158 ( .A(n3679), .Z(n3681) );
  NOR U5159 ( .A(n3681), .B(n3680), .Z(n3682) );
  NOR U5160 ( .A(n3683), .B(n3682), .Z(n4125) );
  XOR U5161 ( .A(n4124), .B(n4125), .Z(n3684) );
  IV U5162 ( .A(n3684), .Z(n4127) );
  XOR U5163 ( .A(n4126), .B(n4127), .Z(n4118) );
  XOR U5164 ( .A(n4117), .B(n4118), .Z(n4122) );
  XOR U5165 ( .A(n3685), .B(n4122), .Z(n3690) );
  NOR U5166 ( .A(n3689), .B(n3690), .Z(n4114) );
  IV U5167 ( .A(n3686), .Z(n3687) );
  NOR U5168 ( .A(n3687), .B(n3694), .Z(n3698) );
  IV U5169 ( .A(n3698), .Z(n3688) );
  NOR U5170 ( .A(n4114), .B(n3688), .Z(n4680) );
  IV U5171 ( .A(n3689), .Z(n3692) );
  IV U5172 ( .A(n3690), .Z(n3691) );
  NOR U5173 ( .A(n3692), .B(n3691), .Z(n4621) );
  IV U5174 ( .A(n3693), .Z(n3695) );
  NOR U5175 ( .A(n3695), .B(n3694), .Z(n4112) );
  XOR U5176 ( .A(n4114), .B(n4112), .Z(n3696) );
  NOR U5177 ( .A(n4621), .B(n3696), .Z(n3697) );
  NOR U5178 ( .A(n3698), .B(n3697), .Z(n3699) );
  NOR U5179 ( .A(n4680), .B(n3699), .Z(n4184) );
  IV U5180 ( .A(n3700), .Z(n3702) );
  NOR U5181 ( .A(n3702), .B(n3701), .Z(n3703) );
  IV U5182 ( .A(n3703), .Z(n4185) );
  XOR U5183 ( .A(n4184), .B(n4185), .Z(n4190) );
  XOR U5184 ( .A(n3704), .B(n4190), .Z(n4192) );
  XOR U5185 ( .A(n4193), .B(n4192), .Z(n4202) );
  IV U5186 ( .A(n3705), .Z(n3707) );
  NOR U5187 ( .A(n3707), .B(n3706), .Z(n4197) );
  IV U5188 ( .A(n3708), .Z(n3709) );
  NOR U5189 ( .A(n3710), .B(n3709), .Z(n4201) );
  NOR U5190 ( .A(n4197), .B(n4201), .Z(n3711) );
  XOR U5191 ( .A(n4202), .B(n3711), .Z(n3712) );
  IV U5192 ( .A(n3712), .Z(n4206) );
  XOR U5193 ( .A(n4199), .B(n4206), .Z(n4108) );
  NOR U5194 ( .A(n3713), .B(n4205), .Z(n3717) );
  IV U5195 ( .A(n3714), .Z(n3716) );
  IV U5196 ( .A(n3715), .Z(n3720) );
  NOR U5197 ( .A(n3716), .B(n3720), .Z(n4107) );
  NOR U5198 ( .A(n3717), .B(n4107), .Z(n3718) );
  XOR U5199 ( .A(n4108), .B(n3718), .Z(n4104) );
  IV U5200 ( .A(n3719), .Z(n3721) );
  NOR U5201 ( .A(n3721), .B(n3720), .Z(n4219) );
  IV U5202 ( .A(n3722), .Z(n3724) );
  NOR U5203 ( .A(n3724), .B(n3723), .Z(n4105) );
  NOR U5204 ( .A(n4219), .B(n4105), .Z(n3725) );
  XOR U5205 ( .A(n4104), .B(n3725), .Z(n4102) );
  XOR U5206 ( .A(n4101), .B(n4102), .Z(n4233) );
  IV U5207 ( .A(n3726), .Z(n3728) );
  IV U5208 ( .A(n3727), .Z(n3730) );
  NOR U5209 ( .A(n3728), .B(n3730), .Z(n4231) );
  XOR U5210 ( .A(n4233), .B(n4231), .Z(n4236) );
  IV U5211 ( .A(n3729), .Z(n3731) );
  NOR U5212 ( .A(n3731), .B(n3730), .Z(n4234) );
  XOR U5213 ( .A(n4236), .B(n4234), .Z(n4238) );
  IV U5214 ( .A(n4238), .Z(n3738) );
  IV U5215 ( .A(n3732), .Z(n3733) );
  NOR U5216 ( .A(n3736), .B(n3733), .Z(n4237) );
  IV U5217 ( .A(n3734), .Z(n3735) );
  NOR U5218 ( .A(n3736), .B(n3735), .Z(n4099) );
  NOR U5219 ( .A(n4237), .B(n4099), .Z(n3737) );
  XOR U5220 ( .A(n3738), .B(n3737), .Z(n4240) );
  NOR U5221 ( .A(n3740), .B(n4240), .Z(n4718) );
  IV U5222 ( .A(n3739), .Z(n4241) );
  XOR U5223 ( .A(n4241), .B(n4240), .Z(n4096) );
  XOR U5224 ( .A(n4095), .B(n4096), .Z(n3742) );
  NOR U5225 ( .A(n4096), .B(n3740), .Z(n3741) );
  NOR U5226 ( .A(n3742), .B(n3741), .Z(n3743) );
  NOR U5227 ( .A(n4718), .B(n3743), .Z(n4092) );
  IV U5228 ( .A(n3744), .Z(n4094) );
  XOR U5229 ( .A(n4092), .B(n4094), .Z(n4245) );
  XOR U5230 ( .A(n4244), .B(n4245), .Z(n4725) );
  XOR U5231 ( .A(n4247), .B(n4725), .Z(n4087) );
  IV U5232 ( .A(n3745), .Z(n3747) );
  IV U5233 ( .A(n3746), .Z(n3752) );
  NOR U5234 ( .A(n3747), .B(n3752), .Z(n4088) );
  IV U5235 ( .A(n3748), .Z(n3750) );
  NOR U5236 ( .A(n3750), .B(n3749), .Z(n4251) );
  IV U5237 ( .A(n3751), .Z(n3753) );
  NOR U5238 ( .A(n3753), .B(n3752), .Z(n4090) );
  NOR U5239 ( .A(n4251), .B(n4090), .Z(n3754) );
  IV U5240 ( .A(n3754), .Z(n3755) );
  NOR U5241 ( .A(n4088), .B(n3755), .Z(n3756) );
  XOR U5242 ( .A(n4087), .B(n3756), .Z(n4086) );
  IV U5243 ( .A(n3757), .Z(n3760) );
  IV U5244 ( .A(n3758), .Z(n3759) );
  NOR U5245 ( .A(n3760), .B(n3759), .Z(n4084) );
  XOR U5246 ( .A(n4086), .B(n4084), .Z(n4255) );
  XOR U5247 ( .A(n4254), .B(n4255), .Z(n4259) );
  XOR U5248 ( .A(n3761), .B(n4259), .Z(n4080) );
  XOR U5249 ( .A(n4081), .B(n4080), .Z(n4266) );
  XOR U5250 ( .A(n4265), .B(n4266), .Z(n4263) );
  XOR U5251 ( .A(n4077), .B(n4263), .Z(n3762) );
  NOR U5252 ( .A(n3763), .B(n3762), .Z(n4764) );
  IV U5253 ( .A(n3764), .Z(n3766) );
  IV U5254 ( .A(n3765), .Z(n3768) );
  NOR U5255 ( .A(n3766), .B(n3768), .Z(n4274) );
  IV U5256 ( .A(n3767), .Z(n3769) );
  NOR U5257 ( .A(n3769), .B(n3768), .Z(n4262) );
  NOR U5258 ( .A(n4077), .B(n4262), .Z(n3770) );
  XOR U5259 ( .A(n3770), .B(n4263), .Z(n4275) );
  XOR U5260 ( .A(n4274), .B(n4275), .Z(n3771) );
  NOR U5261 ( .A(n3772), .B(n3771), .Z(n3773) );
  NOR U5262 ( .A(n4764), .B(n3773), .Z(n3774) );
  IV U5263 ( .A(n3774), .Z(n4282) );
  XOR U5264 ( .A(n4075), .B(n4282), .Z(n3775) );
  NOR U5265 ( .A(n3776), .B(n3775), .Z(n4562) );
  IV U5266 ( .A(n3777), .Z(n3781) );
  NOR U5267 ( .A(n3778), .B(n3781), .Z(n4072) );
  NOR U5268 ( .A(n4075), .B(n4072), .Z(n3779) );
  XOR U5269 ( .A(n3779), .B(n4282), .Z(n3783) );
  IV U5270 ( .A(n3780), .Z(n3782) );
  NOR U5271 ( .A(n3782), .B(n3781), .Z(n4280) );
  XOR U5272 ( .A(n3783), .B(n4280), .Z(n3784) );
  NOR U5273 ( .A(n3785), .B(n3784), .Z(n3786) );
  NOR U5274 ( .A(n4562), .B(n3786), .Z(n4062) );
  IV U5275 ( .A(n3787), .Z(n3788) );
  NOR U5276 ( .A(n4068), .B(n3788), .Z(n4283) );
  NOR U5277 ( .A(n3789), .B(n4063), .Z(n3790) );
  NOR U5278 ( .A(n4283), .B(n3790), .Z(n3791) );
  XOR U5279 ( .A(n4062), .B(n3791), .Z(n4060) );
  XOR U5280 ( .A(n4058), .B(n4060), .Z(n4551) );
  XOR U5281 ( .A(n4289), .B(n4551), .Z(n4290) );
  IV U5282 ( .A(n3792), .Z(n3793) );
  NOR U5283 ( .A(n3794), .B(n3793), .Z(n4538) );
  IV U5284 ( .A(n3795), .Z(n3797) );
  NOR U5285 ( .A(n3797), .B(n3796), .Z(n4546) );
  NOR U5286 ( .A(n4538), .B(n4546), .Z(n4291) );
  XOR U5287 ( .A(n4290), .B(n4291), .Z(n4300) );
  XOR U5288 ( .A(n4295), .B(n4300), .Z(n4305) );
  XOR U5289 ( .A(n4303), .B(n4305), .Z(n4315) );
  XOR U5290 ( .A(n3798), .B(n4315), .Z(n4049) );
  XOR U5291 ( .A(n3799), .B(n4049), .Z(n4322) );
  XOR U5292 ( .A(n3800), .B(n4322), .Z(n4328) );
  XOR U5293 ( .A(n4330), .B(n4328), .Z(n4043) );
  IV U5294 ( .A(n3801), .Z(n3803) );
  NOR U5295 ( .A(n3803), .B(n3802), .Z(n4041) );
  XOR U5296 ( .A(n4043), .B(n4041), .Z(n4326) );
  XOR U5297 ( .A(n4325), .B(n4326), .Z(n4337) );
  XOR U5298 ( .A(n4336), .B(n4337), .Z(n4341) );
  IV U5299 ( .A(n3804), .Z(n3805) );
  NOR U5300 ( .A(n3806), .B(n3805), .Z(n4039) );
  IV U5301 ( .A(n3807), .Z(n3809) );
  NOR U5302 ( .A(n3809), .B(n3808), .Z(n4339) );
  NOR U5303 ( .A(n4039), .B(n4339), .Z(n3810) );
  XOR U5304 ( .A(n4341), .B(n3810), .Z(n3811) );
  IV U5305 ( .A(n3811), .Z(n4035) );
  XOR U5306 ( .A(n4033), .B(n4035), .Z(n4037) );
  XOR U5307 ( .A(n4036), .B(n4037), .Z(n4028) );
  XOR U5308 ( .A(n4027), .B(n4028), .Z(n4031) );
  XOR U5309 ( .A(n4030), .B(n4031), .Z(n4026) );
  XOR U5310 ( .A(n4024), .B(n4026), .Z(n4020) );
  IV U5311 ( .A(n4020), .Z(n3818) );
  IV U5312 ( .A(n3812), .Z(n3813) );
  NOR U5313 ( .A(n3816), .B(n3813), .Z(n4019) );
  IV U5314 ( .A(n3814), .Z(n3815) );
  NOR U5315 ( .A(n3816), .B(n3815), .Z(n4022) );
  NOR U5316 ( .A(n4019), .B(n4022), .Z(n3817) );
  XOR U5317 ( .A(n3818), .B(n3817), .Z(n4015) );
  XOR U5318 ( .A(n4013), .B(n4015), .Z(n4017) );
  XOR U5319 ( .A(n4016), .B(n4017), .Z(n4011) );
  IV U5320 ( .A(n3819), .Z(n3820) );
  NOR U5321 ( .A(n3823), .B(n3820), .Z(n4009) );
  XOR U5322 ( .A(n4011), .B(n4009), .Z(n4347) );
  IV U5323 ( .A(n3821), .Z(n3822) );
  NOR U5324 ( .A(n3823), .B(n3822), .Z(n4345) );
  XOR U5325 ( .A(n4347), .B(n4345), .Z(n4349) );
  IV U5326 ( .A(n3824), .Z(n3825) );
  NOR U5327 ( .A(n3825), .B(n3827), .Z(n4007) );
  IV U5328 ( .A(n3826), .Z(n3828) );
  NOR U5329 ( .A(n3828), .B(n3827), .Z(n4348) );
  NOR U5330 ( .A(n4007), .B(n4348), .Z(n3829) );
  XOR U5331 ( .A(n4349), .B(n3829), .Z(n3830) );
  IV U5332 ( .A(n3830), .Z(n4005) );
  XOR U5333 ( .A(n4004), .B(n4005), .Z(n4003) );
  XOR U5334 ( .A(n3831), .B(n4003), .Z(n3993) );
  XOR U5335 ( .A(n3995), .B(n3993), .Z(n3998) );
  IV U5336 ( .A(n3832), .Z(n3836) );
  XOR U5337 ( .A(n3834), .B(n3833), .Z(n3835) );
  NOR U5338 ( .A(n3836), .B(n3835), .Z(n3996) );
  XOR U5339 ( .A(n3998), .B(n3996), .Z(n3992) );
  IV U5340 ( .A(n3837), .Z(n3839) );
  NOR U5341 ( .A(n3839), .B(n3838), .Z(n3840) );
  IV U5342 ( .A(n3840), .Z(n3991) );
  XOR U5343 ( .A(n3992), .B(n3991), .Z(n3850) );
  IV U5344 ( .A(n3850), .Z(n3841) );
  NOR U5345 ( .A(n3849), .B(n3841), .Z(n4358) );
  IV U5346 ( .A(n3842), .Z(n3843) );
  NOR U5347 ( .A(n3844), .B(n3843), .Z(n3847) );
  IV U5348 ( .A(n3847), .Z(n3845) );
  NOR U5349 ( .A(n3845), .B(n3992), .Z(n4354) );
  NOR U5350 ( .A(n4358), .B(n4354), .Z(n3846) );
  IV U5351 ( .A(n3846), .Z(n4353) );
  NOR U5352 ( .A(n3847), .B(n3850), .Z(n3848) );
  NOR U5353 ( .A(n4353), .B(n3848), .Z(n3852) );
  NOR U5354 ( .A(n3850), .B(n3849), .Z(n3851) );
  NOR U5355 ( .A(n3852), .B(n3851), .Z(n4470) );
  IV U5356 ( .A(n4470), .Z(n3856) );
  IV U5357 ( .A(n3853), .Z(n3854) );
  NOR U5358 ( .A(n3854), .B(n3858), .Z(n4468) );
  IV U5359 ( .A(n3859), .Z(n3855) );
  NOR U5360 ( .A(n3855), .B(n3858), .Z(n4473) );
  NOR U5361 ( .A(n4468), .B(n4473), .Z(n3987) );
  XOR U5362 ( .A(n3856), .B(n3987), .Z(n3990) );
  IV U5363 ( .A(n3857), .Z(n3861) );
  XOR U5364 ( .A(n3859), .B(n3858), .Z(n3860) );
  NOR U5365 ( .A(n3861), .B(n3860), .Z(n3988) );
  XOR U5366 ( .A(n3990), .B(n3988), .Z(n4367) );
  XOR U5367 ( .A(n4366), .B(n4367), .Z(n3984) );
  XOR U5368 ( .A(n3983), .B(n3984), .Z(n3978) );
  XOR U5369 ( .A(n3977), .B(n3978), .Z(n3981) );
  XOR U5370 ( .A(n3980), .B(n3981), .Z(n3968) );
  IV U5371 ( .A(n3862), .Z(n3971) );
  NOR U5372 ( .A(n3863), .B(n3971), .Z(n3866) );
  IV U5373 ( .A(n3864), .Z(n3865) );
  NOR U5374 ( .A(n3865), .B(n3870), .Z(n3967) );
  NOR U5375 ( .A(n3866), .B(n3967), .Z(n3867) );
  XOR U5376 ( .A(n3968), .B(n3867), .Z(n3868) );
  IV U5377 ( .A(n3868), .Z(n3963) );
  IV U5378 ( .A(n3869), .Z(n3871) );
  NOR U5379 ( .A(n3871), .B(n3870), .Z(n3961) );
  XOR U5380 ( .A(n3963), .B(n3961), .Z(n3965) );
  XOR U5381 ( .A(n3872), .B(n3965), .Z(n3945) );
  IV U5382 ( .A(n3873), .Z(n3950) );
  NOR U5383 ( .A(n3874), .B(n3950), .Z(n3877) );
  IV U5384 ( .A(n3875), .Z(n3876) );
  NOR U5385 ( .A(n3876), .B(n3880), .Z(n3946) );
  NOR U5386 ( .A(n3877), .B(n3946), .Z(n3878) );
  XOR U5387 ( .A(n3945), .B(n3878), .Z(n3944) );
  IV U5388 ( .A(n3879), .Z(n3881) );
  NOR U5389 ( .A(n3881), .B(n3880), .Z(n3942) );
  XOR U5390 ( .A(n3944), .B(n3942), .Z(n3940) );
  XOR U5391 ( .A(n3882), .B(n3940), .Z(n3933) );
  XOR U5392 ( .A(n3934), .B(n3933), .Z(n4431) );
  IV U5393 ( .A(n3883), .Z(n3884) );
  NOR U5394 ( .A(n3885), .B(n3884), .Z(n3929) );
  IV U5395 ( .A(n3886), .Z(n3888) );
  NOR U5396 ( .A(n3888), .B(n3887), .Z(n3931) );
  NOR U5397 ( .A(n3929), .B(n3931), .Z(n3889) );
  XOR U5398 ( .A(n4431), .B(n3889), .Z(n3926) );
  XOR U5399 ( .A(n4428), .B(n3926), .Z(n4851) );
  XOR U5400 ( .A(n3894), .B(n4851), .Z(n4391) );
  NOR U5401 ( .A(n3890), .B(n4390), .Z(n3896) );
  IV U5402 ( .A(n3896), .Z(n3891) );
  NOR U5403 ( .A(n4391), .B(n3891), .Z(n4388) );
  IV U5404 ( .A(n3892), .Z(n4415) );
  NOR U5405 ( .A(n3893), .B(n4415), .Z(n4385) );
  NOR U5406 ( .A(n3894), .B(n4385), .Z(n3895) );
  XOR U5407 ( .A(n3895), .B(n4851), .Z(n3917) );
  NOR U5408 ( .A(n3896), .B(n3917), .Z(n3897) );
  NOR U5409 ( .A(n4388), .B(n3897), .Z(n4406) );
  IV U5410 ( .A(n3898), .Z(n3919) );
  NOR U5411 ( .A(n3899), .B(n3919), .Z(n3903) );
  IV U5412 ( .A(n3900), .Z(n3901) );
  NOR U5413 ( .A(n3902), .B(n3901), .Z(n4407) );
  NOR U5414 ( .A(n3903), .B(n4407), .Z(n3904) );
  XOR U5415 ( .A(n4406), .B(n3904), .Z(n4412) );
  IV U5416 ( .A(n3905), .Z(n3906) );
  NOR U5417 ( .A(n3907), .B(n3906), .Z(n4410) );
  XOR U5418 ( .A(n4412), .B(n4410), .Z(n3914) );
  XOR U5419 ( .A(n3912), .B(n3914), .Z(n3916) );
  IV U5420 ( .A(n3908), .Z(n3909) );
  NOR U5421 ( .A(n3910), .B(n3909), .Z(n3911) );
  IV U5422 ( .A(n3911), .Z(n3915) );
  XOR U5423 ( .A(n3916), .B(n3915), .Z(o[2]) );
  IV U5424 ( .A(n3912), .Z(n3913) );
  NOR U5425 ( .A(n3914), .B(n3913), .Z(n5795) );
  NOR U5426 ( .A(n3916), .B(n3915), .Z(n5786) );
  NOR U5427 ( .A(n5795), .B(n5786), .Z(n4871) );
  IV U5428 ( .A(n3917), .Z(n3918) );
  NOR U5429 ( .A(n3919), .B(n3918), .Z(n3920) );
  IV U5430 ( .A(n3920), .Z(n3925) );
  IV U5431 ( .A(n3921), .Z(n3922) );
  NOR U5432 ( .A(n3925), .B(n3922), .Z(n4862) );
  IV U5433 ( .A(n3923), .Z(n3924) );
  NOR U5434 ( .A(n3925), .B(n3924), .Z(n4858) );
  IV U5435 ( .A(n4391), .Z(n3928) );
  IV U5436 ( .A(n3926), .Z(n3927) );
  NOR U5437 ( .A(n3928), .B(n3927), .Z(n4384) );
  IV U5438 ( .A(n3929), .Z(n3930) );
  NOR U5439 ( .A(n4431), .B(n3930), .Z(n4425) );
  IV U5440 ( .A(n3931), .Z(n3932) );
  NOR U5441 ( .A(n4431), .B(n3932), .Z(n4436) );
  IV U5442 ( .A(n3933), .Z(n3935) );
  NOR U5443 ( .A(n3935), .B(n3934), .Z(n4434) );
  IV U5444 ( .A(n3936), .Z(n3937) );
  NOR U5445 ( .A(n3940), .B(n3937), .Z(n4844) );
  IV U5446 ( .A(n3938), .Z(n3939) );
  NOR U5447 ( .A(n3940), .B(n3939), .Z(n4842) );
  XOR U5448 ( .A(n4844), .B(n4842), .Z(n3941) );
  NOR U5449 ( .A(n4434), .B(n3941), .Z(n4383) );
  IV U5450 ( .A(n3942), .Z(n3943) );
  NOR U5451 ( .A(n3944), .B(n3943), .Z(n4439) );
  IV U5452 ( .A(n3945), .Z(n3949) );
  IV U5453 ( .A(n3946), .Z(n3947) );
  NOR U5454 ( .A(n3949), .B(n3947), .Z(n4836) );
  NOR U5455 ( .A(n4439), .B(n4836), .Z(n4382) );
  IV U5456 ( .A(n3948), .Z(n3952) );
  NOR U5457 ( .A(n3950), .B(n3949), .Z(n3951) );
  IV U5458 ( .A(n3951), .Z(n3954) );
  NOR U5459 ( .A(n3952), .B(n3954), .Z(n4833) );
  IV U5460 ( .A(n3953), .Z(n3955) );
  NOR U5461 ( .A(n3955), .B(n3954), .Z(n4441) );
  XOR U5462 ( .A(n3964), .B(n3965), .Z(n3958) );
  IV U5463 ( .A(n3956), .Z(n3957) );
  NOR U5464 ( .A(n3958), .B(n3957), .Z(n4448) );
  IV U5465 ( .A(n3959), .Z(n3960) );
  NOR U5466 ( .A(n3960), .B(n3965), .Z(n4446) );
  NOR U5467 ( .A(n4448), .B(n4446), .Z(n4381) );
  IV U5468 ( .A(n3961), .Z(n3962) );
  NOR U5469 ( .A(n3963), .B(n3962), .Z(n4456) );
  IV U5470 ( .A(n3964), .Z(n3966) );
  NOR U5471 ( .A(n3966), .B(n3965), .Z(n4451) );
  NOR U5472 ( .A(n4456), .B(n4451), .Z(n4380) );
  IV U5473 ( .A(n3967), .Z(n3969) );
  NOR U5474 ( .A(n3969), .B(n3968), .Z(n4453) );
  IV U5475 ( .A(n3970), .Z(n3973) );
  NOR U5476 ( .A(n3971), .B(n3981), .Z(n3972) );
  IV U5477 ( .A(n3972), .Z(n3975) );
  NOR U5478 ( .A(n3973), .B(n3975), .Z(n4462) );
  IV U5479 ( .A(n3974), .Z(n3976) );
  NOR U5480 ( .A(n3976), .B(n3975), .Z(n4459) );
  IV U5481 ( .A(n3977), .Z(n3979) );
  NOR U5482 ( .A(n3979), .B(n3978), .Z(n4930) );
  IV U5483 ( .A(n3980), .Z(n3982) );
  NOR U5484 ( .A(n3982), .B(n3981), .Z(n4925) );
  NOR U5485 ( .A(n4930), .B(n4925), .Z(n4465) );
  IV U5486 ( .A(n4465), .Z(n4379) );
  IV U5487 ( .A(n3983), .Z(n3985) );
  NOR U5488 ( .A(n3985), .B(n3984), .Z(n3986) );
  IV U5489 ( .A(n3986), .Z(n4375) );
  NOR U5490 ( .A(n4470), .B(n3987), .Z(n4369) );
  IV U5491 ( .A(n3988), .Z(n3989) );
  NOR U5492 ( .A(n3990), .B(n3989), .Z(n4466) );
  NOR U5493 ( .A(n4369), .B(n4466), .Z(n4364) );
  NOR U5494 ( .A(n3992), .B(n3991), .Z(n4477) );
  IV U5495 ( .A(n3993), .Z(n3994) );
  NOR U5496 ( .A(n3995), .B(n3994), .Z(n4958) );
  IV U5497 ( .A(n3996), .Z(n3997) );
  NOR U5498 ( .A(n3998), .B(n3997), .Z(n4951) );
  NOR U5499 ( .A(n4958), .B(n4951), .Z(n4476) );
  IV U5500 ( .A(n3999), .Z(n4000) );
  NOR U5501 ( .A(n4000), .B(n4003), .Z(n4481) );
  IV U5502 ( .A(n4001), .Z(n4002) );
  NOR U5503 ( .A(n4003), .B(n4002), .Z(n4822) );
  IV U5504 ( .A(n4004), .Z(n4006) );
  NOR U5505 ( .A(n4006), .B(n4005), .Z(n4819) );
  IV U5506 ( .A(n4007), .Z(n4008) );
  NOR U5507 ( .A(n4008), .B(n4349), .Z(n4484) );
  IV U5508 ( .A(n4009), .Z(n4010) );
  NOR U5509 ( .A(n4011), .B(n4010), .Z(n4012) );
  IV U5510 ( .A(n4012), .Z(n4814) );
  IV U5511 ( .A(n4013), .Z(n4014) );
  NOR U5512 ( .A(n4015), .B(n4014), .Z(n4493) );
  IV U5513 ( .A(n4016), .Z(n4018) );
  NOR U5514 ( .A(n4018), .B(n4017), .Z(n4809) );
  NOR U5515 ( .A(n4493), .B(n4809), .Z(n4344) );
  IV U5516 ( .A(n4019), .Z(n4021) );
  NOR U5517 ( .A(n4021), .B(n4020), .Z(n4490) );
  IV U5518 ( .A(n4022), .Z(n4023) );
  NOR U5519 ( .A(n4023), .B(n4026), .Z(n4797) );
  IV U5520 ( .A(n4024), .Z(n4025) );
  NOR U5521 ( .A(n4026), .B(n4025), .Z(n4495) );
  IV U5522 ( .A(n4027), .Z(n4029) );
  NOR U5523 ( .A(n4029), .B(n4028), .Z(n4499) );
  IV U5524 ( .A(n4030), .Z(n4032) );
  NOR U5525 ( .A(n4032), .B(n4031), .Z(n4800) );
  NOR U5526 ( .A(n4499), .B(n4800), .Z(n4343) );
  IV U5527 ( .A(n4033), .Z(n4034) );
  NOR U5528 ( .A(n4035), .B(n4034), .Z(n4509) );
  IV U5529 ( .A(n4036), .Z(n4038) );
  NOR U5530 ( .A(n4038), .B(n4037), .Z(n4502) );
  NOR U5531 ( .A(n4509), .B(n4502), .Z(n4342) );
  IV U5532 ( .A(n4039), .Z(n4040) );
  NOR U5533 ( .A(n4341), .B(n4040), .Z(n4506) );
  IV U5534 ( .A(n4041), .Z(n4042) );
  NOR U5535 ( .A(n4043), .B(n4042), .Z(n4044) );
  IV U5536 ( .A(n4044), .Z(n4332) );
  IV U5537 ( .A(n4045), .Z(n4046) );
  NOR U5538 ( .A(n4046), .B(n4322), .Z(n4047) );
  IV U5539 ( .A(n4047), .Z(n4790) );
  IV U5540 ( .A(n4048), .Z(n4051) );
  IV U5541 ( .A(n4049), .Z(n4320) );
  XOR U5542 ( .A(n4052), .B(n4320), .Z(n4050) );
  NOR U5543 ( .A(n4051), .B(n4050), .Z(n4521) );
  IV U5544 ( .A(n4052), .Z(n4053) );
  NOR U5545 ( .A(n4320), .B(n4053), .Z(n4780) );
  IV U5546 ( .A(n4054), .Z(n4057) );
  NOR U5547 ( .A(n4055), .B(n4315), .Z(n4056) );
  IV U5548 ( .A(n4056), .Z(n4311) );
  NOR U5549 ( .A(n4057), .B(n4311), .Z(n4525) );
  NOR U5550 ( .A(n4780), .B(n4525), .Z(n4317) );
  IV U5551 ( .A(n4058), .Z(n4059) );
  NOR U5552 ( .A(n4060), .B(n4059), .Z(n4557) );
  IV U5553 ( .A(n4061), .Z(n4066) );
  IV U5554 ( .A(n4062), .Z(n4284) );
  NOR U5555 ( .A(n4063), .B(n4284), .Z(n4064) );
  IV U5556 ( .A(n4064), .Z(n4065) );
  NOR U5557 ( .A(n4066), .B(n4065), .Z(n4559) );
  NOR U5558 ( .A(n4557), .B(n4559), .Z(n4288) );
  IV U5559 ( .A(n4067), .Z(n4071) );
  NOR U5560 ( .A(n4068), .B(n4284), .Z(n4069) );
  IV U5561 ( .A(n4069), .Z(n4070) );
  NOR U5562 ( .A(n4071), .B(n4070), .Z(n4773) );
  IV U5563 ( .A(n4072), .Z(n4073) );
  NOR U5564 ( .A(n4073), .B(n4282), .Z(n4074) );
  IV U5565 ( .A(n4074), .Z(n4566) );
  IV U5566 ( .A(n4075), .Z(n4076) );
  NOR U5567 ( .A(n4076), .B(n4282), .Z(n4570) );
  NOR U5568 ( .A(n4764), .B(n4570), .Z(n4279) );
  IV U5569 ( .A(n4077), .Z(n4078) );
  NOR U5570 ( .A(n4078), .B(n4263), .Z(n4079) );
  IV U5571 ( .A(n4079), .Z(n4270) );
  IV U5572 ( .A(n4080), .Z(n4581) );
  NOR U5573 ( .A(n4081), .B(n4581), .Z(n4268) );
  IV U5574 ( .A(n4082), .Z(n4083) );
  NOR U5575 ( .A(n4083), .B(n4259), .Z(n4740) );
  IV U5576 ( .A(n4084), .Z(n4085) );
  NOR U5577 ( .A(n4086), .B(n4085), .Z(n5169) );
  IV U5578 ( .A(n4087), .Z(n4252) );
  IV U5579 ( .A(n4088), .Z(n4089) );
  NOR U5580 ( .A(n4252), .B(n4089), .Z(n5026) );
  NOR U5581 ( .A(n5169), .B(n5026), .Z(n4584) );
  IV U5582 ( .A(n4090), .Z(n4091) );
  NOR U5583 ( .A(n4091), .B(n4252), .Z(n4591) );
  IV U5584 ( .A(n4092), .Z(n4093) );
  NOR U5585 ( .A(n4094), .B(n4093), .Z(n4598) );
  IV U5586 ( .A(n4095), .Z(n4098) );
  IV U5587 ( .A(n4096), .Z(n4097) );
  NOR U5588 ( .A(n4098), .B(n4097), .Z(n4715) );
  IV U5589 ( .A(n4099), .Z(n4100) );
  NOR U5590 ( .A(n4100), .B(n4238), .Z(n4706) );
  IV U5591 ( .A(n4101), .Z(n4103) );
  NOR U5592 ( .A(n4103), .B(n4102), .Z(n4226) );
  IV U5593 ( .A(n4104), .Z(n4221) );
  IV U5594 ( .A(n4105), .Z(n4106) );
  NOR U5595 ( .A(n4221), .B(n4106), .Z(n4223) );
  IV U5596 ( .A(n4223), .Z(n4218) );
  IV U5597 ( .A(n4107), .Z(n4109) );
  NOR U5598 ( .A(n4109), .B(n4108), .Z(n4608) );
  IV U5599 ( .A(n4110), .Z(n4111) );
  NOR U5600 ( .A(n4111), .B(n4190), .Z(n4616) );
  IV U5601 ( .A(n4112), .Z(n4113) );
  NOR U5602 ( .A(n4114), .B(n4113), .Z(n4618) );
  NOR U5603 ( .A(n4621), .B(n4618), .Z(n4183) );
  IV U5604 ( .A(n4115), .Z(n4116) );
  NOR U5605 ( .A(n4116), .B(n4122), .Z(n4623) );
  IV U5606 ( .A(n4117), .Z(n4119) );
  NOR U5607 ( .A(n4119), .B(n4118), .Z(n4628) );
  IV U5608 ( .A(n4120), .Z(n4121) );
  NOR U5609 ( .A(n4122), .B(n4121), .Z(n4626) );
  NOR U5610 ( .A(n4628), .B(n4626), .Z(n4123) );
  IV U5611 ( .A(n4123), .Z(n4182) );
  NOR U5612 ( .A(n4125), .B(n4124), .Z(n4634) );
  IV U5613 ( .A(n4126), .Z(n4128) );
  NOR U5614 ( .A(n4128), .B(n4127), .Z(n4631) );
  NOR U5615 ( .A(n4634), .B(n4631), .Z(n4181) );
  IV U5616 ( .A(n4129), .Z(n4130) );
  NOR U5617 ( .A(n4130), .B(n4172), .Z(n4637) );
  IV U5618 ( .A(n4131), .Z(n4133) );
  NOR U5619 ( .A(n4133), .B(n4132), .Z(n4137) );
  IV U5620 ( .A(n4134), .Z(n4135) );
  NOR U5621 ( .A(n4172), .B(n4135), .Z(n4136) );
  NOR U5622 ( .A(n4137), .B(n4136), .Z(n4641) );
  IV U5623 ( .A(n4641), .Z(n4169) );
  IV U5624 ( .A(n4138), .Z(n4139) );
  NOR U5625 ( .A(n4140), .B(n4139), .Z(n4145) );
  IV U5626 ( .A(n4141), .Z(n4142) );
  NOR U5627 ( .A(n4143), .B(n4142), .Z(n4144) );
  NOR U5628 ( .A(n4145), .B(n4144), .Z(n4649) );
  IV U5629 ( .A(n4146), .Z(n4147) );
  NOR U5630 ( .A(n4148), .B(n4147), .Z(n4153) );
  IV U5631 ( .A(n4149), .Z(n4150) );
  NOR U5632 ( .A(n4151), .B(n4150), .Z(n4152) );
  NOR U5633 ( .A(n4153), .B(n4152), .Z(n4654) );
  IV U5634 ( .A(n4154), .Z(n4157) );
  IV U5635 ( .A(n4155), .Z(n4156) );
  NOR U5636 ( .A(n4157), .B(n4156), .Z(n4650) );
  IV U5637 ( .A(n4158), .Z(n4160) );
  NOR U5638 ( .A(n4160), .B(n4159), .Z(n4161) );
  NOR U5639 ( .A(n4162), .B(n4161), .Z(n4659) );
  IV U5640 ( .A(n4659), .Z(n4168) );
  XOR U5641 ( .A(n4168), .B(n4658), .Z(n4651) );
  XOR U5642 ( .A(n4650), .B(n4651), .Z(n4653) );
  XOR U5643 ( .A(n4654), .B(n4653), .Z(n4647) );
  XOR U5644 ( .A(n4649), .B(n4647), .Z(n4640) );
  XOR U5645 ( .A(n4169), .B(n4640), .Z(n4662) );
  IV U5646 ( .A(n4170), .Z(n4171) );
  NOR U5647 ( .A(n4172), .B(n4171), .Z(n4660) );
  XOR U5648 ( .A(n4662), .B(n4660), .Z(n4638) );
  XOR U5649 ( .A(n4637), .B(n4638), .Z(n4642) );
  IV U5650 ( .A(n4173), .Z(n4175) );
  NOR U5651 ( .A(n4175), .B(n4174), .Z(n4180) );
  IV U5652 ( .A(n4176), .Z(n4178) );
  NOR U5653 ( .A(n4178), .B(n4177), .Z(n4179) );
  NOR U5654 ( .A(n4180), .B(n4179), .Z(n4643) );
  XOR U5655 ( .A(n4642), .B(n4643), .Z(n4632) );
  XOR U5656 ( .A(n4181), .B(n4632), .Z(n4630) );
  XOR U5657 ( .A(n4182), .B(n4630), .Z(n4624) );
  XOR U5658 ( .A(n4623), .B(n4624), .Z(n4619) );
  XOR U5659 ( .A(n4183), .B(n4619), .Z(n4615) );
  XOR U5660 ( .A(n4616), .B(n4615), .Z(n4188) );
  IV U5661 ( .A(n4184), .Z(n4186) );
  NOR U5662 ( .A(n4186), .B(n4185), .Z(n4682) );
  NOR U5663 ( .A(n4680), .B(n4682), .Z(n4187) );
  XOR U5664 ( .A(n4188), .B(n4187), .Z(n4695) );
  IV U5665 ( .A(n4695), .Z(n4196) );
  IV U5666 ( .A(n4189), .Z(n4191) );
  NOR U5667 ( .A(n4191), .B(n4190), .Z(n4688) );
  IV U5668 ( .A(n4192), .Z(n4694) );
  NOR U5669 ( .A(n4193), .B(n4694), .Z(n4194) );
  NOR U5670 ( .A(n4688), .B(n4194), .Z(n4195) );
  XOR U5671 ( .A(n4196), .B(n4195), .Z(n4692) );
  IV U5672 ( .A(n4197), .Z(n4198) );
  NOR U5673 ( .A(n4198), .B(n4694), .Z(n4690) );
  XOR U5674 ( .A(n4692), .B(n4690), .Z(n4614) );
  IV U5675 ( .A(n4199), .Z(n4200) );
  NOR U5676 ( .A(n4206), .B(n4200), .Z(n4610) );
  IV U5677 ( .A(n4201), .Z(n4203) );
  NOR U5678 ( .A(n4203), .B(n4202), .Z(n4612) );
  NOR U5679 ( .A(n4610), .B(n4612), .Z(n4204) );
  XOR U5680 ( .A(n4614), .B(n4204), .Z(n4605) );
  IV U5681 ( .A(n4605), .Z(n4210) );
  IV U5682 ( .A(n4603), .Z(n4208) );
  NOR U5683 ( .A(n4206), .B(n4205), .Z(n4207) );
  IV U5684 ( .A(n4207), .Z(n4606) );
  NOR U5685 ( .A(n4208), .B(n4606), .Z(n4211) );
  IV U5686 ( .A(n4211), .Z(n4209) );
  NOR U5687 ( .A(n4210), .B(n4209), .Z(n4215) );
  NOR U5688 ( .A(n4211), .B(n4605), .Z(n4213) );
  IV U5689 ( .A(n4604), .Z(n4602) );
  NOR U5690 ( .A(n4602), .B(n4606), .Z(n4212) );
  XOR U5691 ( .A(n4213), .B(n4212), .Z(n4214) );
  NOR U5692 ( .A(n4215), .B(n4214), .Z(n4216) );
  IV U5693 ( .A(n4216), .Z(n4609) );
  XOR U5694 ( .A(n4608), .B(n4609), .Z(n4217) );
  NOR U5695 ( .A(n4218), .B(n4217), .Z(n4601) );
  IV U5696 ( .A(n4219), .Z(n4220) );
  NOR U5697 ( .A(n4221), .B(n4220), .Z(n4607) );
  NOR U5698 ( .A(n4607), .B(n4608), .Z(n4222) );
  XOR U5699 ( .A(n4222), .B(n4609), .Z(n4227) );
  NOR U5700 ( .A(n4223), .B(n4227), .Z(n4224) );
  NOR U5701 ( .A(n4601), .B(n4224), .Z(n4225) );
  NOR U5702 ( .A(n4226), .B(n4225), .Z(n4230) );
  IV U5703 ( .A(n4226), .Z(n4229) );
  IV U5704 ( .A(n4227), .Z(n4228) );
  NOR U5705 ( .A(n4229), .B(n4228), .Z(n5053) );
  NOR U5706 ( .A(n4230), .B(n5053), .Z(n4702) );
  IV U5707 ( .A(n4231), .Z(n4232) );
  NOR U5708 ( .A(n4233), .B(n4232), .Z(n5046) );
  IV U5709 ( .A(n4234), .Z(n4235) );
  NOR U5710 ( .A(n4236), .B(n4235), .Z(n5144) );
  NOR U5711 ( .A(n5046), .B(n5144), .Z(n4703) );
  XOR U5712 ( .A(n4702), .B(n4703), .Z(n4707) );
  XOR U5713 ( .A(n4706), .B(n4707), .Z(n4713) );
  IV U5714 ( .A(n4713), .Z(n4243) );
  IV U5715 ( .A(n4237), .Z(n4239) );
  NOR U5716 ( .A(n4239), .B(n4238), .Z(n4709) );
  NOR U5717 ( .A(n4241), .B(n4240), .Z(n4712) );
  NOR U5718 ( .A(n4709), .B(n4712), .Z(n4242) );
  XOR U5719 ( .A(n4243), .B(n4242), .Z(n4717) );
  XOR U5720 ( .A(n4715), .B(n4717), .Z(n4719) );
  XOR U5721 ( .A(n4718), .B(n4719), .Z(n4599) );
  XOR U5722 ( .A(n4598), .B(n4599), .Z(n4724) );
  IV U5723 ( .A(n4244), .Z(n4246) );
  NOR U5724 ( .A(n4246), .B(n4245), .Z(n4596) );
  NOR U5725 ( .A(n4247), .B(n4725), .Z(n4248) );
  NOR U5726 ( .A(n4596), .B(n4248), .Z(n4249) );
  XOR U5727 ( .A(n4724), .B(n4249), .Z(n4250) );
  IV U5728 ( .A(n4250), .Z(n4590) );
  IV U5729 ( .A(n4251), .Z(n4253) );
  NOR U5730 ( .A(n4253), .B(n4252), .Z(n4588) );
  XOR U5731 ( .A(n4590), .B(n4588), .Z(n4592) );
  XOR U5732 ( .A(n4591), .B(n4592), .Z(n5027) );
  XOR U5733 ( .A(n4584), .B(n5027), .Z(n4586) );
  IV U5734 ( .A(n4254), .Z(n4256) );
  NOR U5735 ( .A(n4256), .B(n4255), .Z(n4585) );
  IV U5736 ( .A(n4257), .Z(n4258) );
  NOR U5737 ( .A(n4259), .B(n4258), .Z(n4737) );
  NOR U5738 ( .A(n4585), .B(n4737), .Z(n4260) );
  XOR U5739 ( .A(n4586), .B(n4260), .Z(n4741) );
  XOR U5740 ( .A(n4740), .B(n4741), .Z(n4578) );
  XOR U5741 ( .A(n4268), .B(n4578), .Z(n4261) );
  NOR U5742 ( .A(n4270), .B(n4261), .Z(n5021) );
  IV U5743 ( .A(n4262), .Z(n4264) );
  NOR U5744 ( .A(n4264), .B(n4263), .Z(n4572) );
  IV U5745 ( .A(n4265), .Z(n4267) );
  NOR U5746 ( .A(n4267), .B(n4266), .Z(n4577) );
  NOR U5747 ( .A(n4268), .B(n4577), .Z(n4269) );
  XOR U5748 ( .A(n4269), .B(n4578), .Z(n4573) );
  XOR U5749 ( .A(n4572), .B(n4573), .Z(n4272) );
  NOR U5750 ( .A(n4573), .B(n4270), .Z(n4271) );
  NOR U5751 ( .A(n4272), .B(n4271), .Z(n4273) );
  NOR U5752 ( .A(n5021), .B(n4273), .Z(n4761) );
  IV U5753 ( .A(n4274), .Z(n4277) );
  IV U5754 ( .A(n4275), .Z(n4276) );
  NOR U5755 ( .A(n4277), .B(n4276), .Z(n4278) );
  IV U5756 ( .A(n4278), .Z(n4763) );
  XOR U5757 ( .A(n4761), .B(n4763), .Z(n4765) );
  XOR U5758 ( .A(n4279), .B(n4765), .Z(n4564) );
  XOR U5759 ( .A(n4566), .B(n4564), .Z(n4569) );
  IV U5760 ( .A(n4280), .Z(n4281) );
  NOR U5761 ( .A(n4282), .B(n4281), .Z(n4567) );
  XOR U5762 ( .A(n4569), .B(n4567), .Z(n4771) );
  IV U5763 ( .A(n4283), .Z(n4285) );
  NOR U5764 ( .A(n4285), .B(n4284), .Z(n4770) );
  NOR U5765 ( .A(n4562), .B(n4770), .Z(n4286) );
  XOR U5766 ( .A(n4771), .B(n4286), .Z(n4287) );
  IV U5767 ( .A(n4287), .Z(n4774) );
  XOR U5768 ( .A(n4773), .B(n4774), .Z(n4561) );
  XOR U5769 ( .A(n4288), .B(n4561), .Z(n4539) );
  NOR U5770 ( .A(n4289), .B(n4551), .Z(n4293) );
  IV U5771 ( .A(n4290), .Z(n4540) );
  NOR U5772 ( .A(n4291), .B(n4540), .Z(n4292) );
  NOR U5773 ( .A(n4293), .B(n4292), .Z(n4294) );
  XOR U5774 ( .A(n4539), .B(n4294), .Z(n4545) );
  IV U5775 ( .A(n4295), .Z(n4296) );
  NOR U5776 ( .A(n4296), .B(n4300), .Z(n4543) );
  IV U5777 ( .A(n4308), .Z(n4298) );
  NOR U5778 ( .A(n4298), .B(n4297), .Z(n4299) );
  IV U5779 ( .A(n4299), .Z(n4301) );
  NOR U5780 ( .A(n4301), .B(n4300), .Z(n4536) );
  NOR U5781 ( .A(n4543), .B(n4536), .Z(n4302) );
  XOR U5782 ( .A(n4545), .B(n4302), .Z(n4533) );
  IV U5783 ( .A(n4303), .Z(n4304) );
  NOR U5784 ( .A(n4305), .B(n4304), .Z(n4306) );
  IV U5785 ( .A(n4306), .Z(n4307) );
  NOR U5786 ( .A(n4308), .B(n4307), .Z(n4309) );
  IV U5787 ( .A(n4309), .Z(n4534) );
  XOR U5788 ( .A(n4533), .B(n4534), .Z(n4532) );
  IV U5789 ( .A(n4310), .Z(n4312) );
  NOR U5790 ( .A(n4312), .B(n4311), .Z(n4528) );
  IV U5791 ( .A(n4313), .Z(n4314) );
  NOR U5792 ( .A(n4315), .B(n4314), .Z(n4530) );
  NOR U5793 ( .A(n4528), .B(n4530), .Z(n4316) );
  XOR U5794 ( .A(n4532), .B(n4316), .Z(n4526) );
  XOR U5795 ( .A(n4317), .B(n4526), .Z(n4523) );
  XOR U5796 ( .A(n4521), .B(n4523), .Z(n4778) );
  IV U5797 ( .A(n4318), .Z(n4319) );
  NOR U5798 ( .A(n4320), .B(n4319), .Z(n4777) );
  IV U5799 ( .A(n4321), .Z(n4323) );
  NOR U5800 ( .A(n4323), .B(n4322), .Z(n4518) );
  NOR U5801 ( .A(n4777), .B(n4518), .Z(n4324) );
  XOR U5802 ( .A(n4778), .B(n4324), .Z(n4788) );
  XOR U5803 ( .A(n4790), .B(n4788), .Z(n4791) );
  NOR U5804 ( .A(n4332), .B(n4791), .Z(n5266) );
  IV U5805 ( .A(n4325), .Z(n4327) );
  NOR U5806 ( .A(n4327), .B(n4326), .Z(n4514) );
  IV U5807 ( .A(n4328), .Z(n4329) );
  NOR U5808 ( .A(n4330), .B(n4329), .Z(n4331) );
  IV U5809 ( .A(n4331), .Z(n4792) );
  XOR U5810 ( .A(n4792), .B(n4791), .Z(n4515) );
  XOR U5811 ( .A(n4514), .B(n4515), .Z(n4334) );
  NOR U5812 ( .A(n4515), .B(n4332), .Z(n4333) );
  NOR U5813 ( .A(n4334), .B(n4333), .Z(n4335) );
  NOR U5814 ( .A(n5266), .B(n4335), .Z(n4512) );
  IV U5815 ( .A(n4336), .Z(n4338) );
  NOR U5816 ( .A(n4338), .B(n4337), .Z(n5280) );
  IV U5817 ( .A(n4339), .Z(n4340) );
  NOR U5818 ( .A(n4341), .B(n4340), .Z(n5286) );
  NOR U5819 ( .A(n5280), .B(n5286), .Z(n4513) );
  XOR U5820 ( .A(n4512), .B(n4513), .Z(n4507) );
  XOR U5821 ( .A(n4506), .B(n4507), .Z(n4510) );
  XOR U5822 ( .A(n4342), .B(n4510), .Z(n4500) );
  XOR U5823 ( .A(n4343), .B(n4500), .Z(n4496) );
  XOR U5824 ( .A(n4495), .B(n4496), .Z(n4798) );
  XOR U5825 ( .A(n4797), .B(n4798), .Z(n4491) );
  XOR U5826 ( .A(n4490), .B(n4491), .Z(n4810) );
  XOR U5827 ( .A(n4344), .B(n4810), .Z(n4813) );
  XOR U5828 ( .A(n4814), .B(n4813), .Z(n4488) );
  IV U5829 ( .A(n4345), .Z(n4346) );
  NOR U5830 ( .A(n4347), .B(n4346), .Z(n4815) );
  IV U5831 ( .A(n4348), .Z(n4350) );
  NOR U5832 ( .A(n4350), .B(n4349), .Z(n4487) );
  NOR U5833 ( .A(n4815), .B(n4487), .Z(n4351) );
  XOR U5834 ( .A(n4488), .B(n4351), .Z(n4352) );
  IV U5835 ( .A(n4352), .Z(n4486) );
  XOR U5836 ( .A(n4484), .B(n4486), .Z(n4820) );
  XOR U5837 ( .A(n4819), .B(n4820), .Z(n4823) );
  XOR U5838 ( .A(n4822), .B(n4823), .Z(n4482) );
  XOR U5839 ( .A(n4481), .B(n4482), .Z(n4952) );
  XOR U5840 ( .A(n4476), .B(n4952), .Z(n4359) );
  XOR U5841 ( .A(n4477), .B(n4359), .Z(n4355) );
  NOR U5842 ( .A(n4355), .B(n4353), .Z(n4362) );
  IV U5843 ( .A(n4354), .Z(n4357) );
  IV U5844 ( .A(n4355), .Z(n4356) );
  NOR U5845 ( .A(n4357), .B(n4356), .Z(n4938) );
  IV U5846 ( .A(n4358), .Z(n4360) );
  IV U5847 ( .A(n4359), .Z(n4478) );
  NOR U5848 ( .A(n4360), .B(n4478), .Z(n4940) );
  NOR U5849 ( .A(n4938), .B(n4940), .Z(n4827) );
  IV U5850 ( .A(n4827), .Z(n4361) );
  NOR U5851 ( .A(n4362), .B(n4361), .Z(n4363) );
  IV U5852 ( .A(n4363), .Z(n4469) );
  XOR U5853 ( .A(n4364), .B(n4469), .Z(n4376) );
  IV U5854 ( .A(n4376), .Z(n4365) );
  NOR U5855 ( .A(n4375), .B(n4365), .Z(n5310) );
  IV U5856 ( .A(n4366), .Z(n4368) );
  NOR U5857 ( .A(n4368), .B(n4367), .Z(n4373) );
  IV U5858 ( .A(n4373), .Z(n4371) );
  XOR U5859 ( .A(n4369), .B(n4469), .Z(n4370) );
  NOR U5860 ( .A(n4371), .B(n4370), .Z(n5305) );
  NOR U5861 ( .A(n5310), .B(n5305), .Z(n4372) );
  IV U5862 ( .A(n4372), .Z(n4828) );
  NOR U5863 ( .A(n4373), .B(n4376), .Z(n4374) );
  NOR U5864 ( .A(n4828), .B(n4374), .Z(n4378) );
  NOR U5865 ( .A(n4376), .B(n4375), .Z(n4377) );
  NOR U5866 ( .A(n4378), .B(n4377), .Z(n4927) );
  XOR U5867 ( .A(n4379), .B(n4927), .Z(n4461) );
  XOR U5868 ( .A(n4459), .B(n4461), .Z(n4463) );
  XOR U5869 ( .A(n4462), .B(n4463), .Z(n4455) );
  XOR U5870 ( .A(n4453), .B(n4455), .Z(n4457) );
  XOR U5871 ( .A(n4380), .B(n4457), .Z(n4444) );
  XOR U5872 ( .A(n4381), .B(n4444), .Z(n4443) );
  XOR U5873 ( .A(n4441), .B(n4443), .Z(n4834) );
  XOR U5874 ( .A(n4833), .B(n4834), .Z(n4838) );
  XOR U5875 ( .A(n4382), .B(n4838), .Z(n4433) );
  XOR U5876 ( .A(n4383), .B(n4433), .Z(n4438) );
  XOR U5877 ( .A(n4436), .B(n4438), .Z(n4426) );
  XOR U5878 ( .A(n4425), .B(n4426), .Z(n4854) );
  XOR U5879 ( .A(n4384), .B(n4854), .Z(n4416) );
  IV U5880 ( .A(n4385), .Z(n4386) );
  NOR U5881 ( .A(n4851), .B(n4386), .Z(n4387) );
  XOR U5882 ( .A(n4416), .B(n4387), .Z(n4394) );
  IV U5883 ( .A(n4394), .Z(n4389) );
  NOR U5884 ( .A(n4389), .B(n4388), .Z(n4404) );
  NOR U5885 ( .A(n4391), .B(n4390), .Z(n4392) );
  IV U5886 ( .A(n4392), .Z(n4400) );
  IV U5887 ( .A(n4393), .Z(n4395) );
  NOR U5888 ( .A(n4395), .B(n4394), .Z(n4396) );
  IV U5889 ( .A(n4396), .Z(n4397) );
  NOR U5890 ( .A(n4400), .B(n4397), .Z(n4878) );
  IV U5891 ( .A(n4398), .Z(n4399) );
  NOR U5892 ( .A(n4400), .B(n4399), .Z(n4401) );
  IV U5893 ( .A(n4401), .Z(n4402) );
  NOR U5894 ( .A(n4416), .B(n4402), .Z(n5355) );
  NOR U5895 ( .A(n4878), .B(n5355), .Z(n4403) );
  IV U5896 ( .A(n4403), .Z(n5363) );
  NOR U5897 ( .A(n4404), .B(n5363), .Z(n4405) );
  IV U5898 ( .A(n4405), .Z(n4859) );
  XOR U5899 ( .A(n4858), .B(n4859), .Z(n4864) );
  XOR U5900 ( .A(n4862), .B(n4864), .Z(n4870) );
  IV U5901 ( .A(n4870), .Z(n4414) );
  IV U5902 ( .A(n4406), .Z(n4409) );
  IV U5903 ( .A(n4407), .Z(n4408) );
  NOR U5904 ( .A(n4409), .B(n4408), .Z(n4865) );
  IV U5905 ( .A(n4410), .Z(n4411) );
  NOR U5906 ( .A(n4412), .B(n4411), .Z(n4868) );
  NOR U5907 ( .A(n4865), .B(n4868), .Z(n4413) );
  XOR U5908 ( .A(n4414), .B(n4413), .Z(n5781) );
  XOR U5909 ( .A(n4871), .B(n5781), .Z(o[3]) );
  NOR U5910 ( .A(n4416), .B(n4415), .Z(n4417) );
  IV U5911 ( .A(n4417), .Z(n4418) );
  NOR U5912 ( .A(n4851), .B(n4418), .Z(n4419) );
  IV U5913 ( .A(n4419), .Z(n4424) );
  IV U5914 ( .A(n4420), .Z(n4421) );
  NOR U5915 ( .A(n4424), .B(n4421), .Z(n4880) );
  IV U5916 ( .A(n4422), .Z(n4423) );
  NOR U5917 ( .A(n4424), .B(n4423), .Z(n4882) );
  IV U5918 ( .A(n4425), .Z(n4427) );
  NOR U5919 ( .A(n4427), .B(n4426), .Z(n4895) );
  NOR U5920 ( .A(n4854), .B(n4428), .Z(n4429) );
  IV U5921 ( .A(n4429), .Z(n4430) );
  NOR U5922 ( .A(n4431), .B(n4430), .Z(n4893) );
  NOR U5923 ( .A(n4895), .B(n4893), .Z(n4432) );
  IV U5924 ( .A(n4432), .Z(n4849) );
  IV U5925 ( .A(n4433), .Z(n4843) );
  IV U5926 ( .A(n4434), .Z(n4435) );
  NOR U5927 ( .A(n4843), .B(n4435), .Z(n4902) );
  IV U5928 ( .A(n4436), .Z(n4437) );
  NOR U5929 ( .A(n4438), .B(n4437), .Z(n4898) );
  NOR U5930 ( .A(n4902), .B(n4898), .Z(n4848) );
  IV U5931 ( .A(n4439), .Z(n4440) );
  NOR U5932 ( .A(n4440), .B(n4443), .Z(n5342) );
  IV U5933 ( .A(n4441), .Z(n4442) );
  NOR U5934 ( .A(n4443), .B(n4442), .Z(n5323) );
  IV U5935 ( .A(n4444), .Z(n4447) );
  IV U5936 ( .A(n4448), .Z(n4445) );
  NOR U5937 ( .A(n4447), .B(n4445), .Z(n5315) );
  IV U5938 ( .A(n4446), .Z(n4450) );
  XOR U5939 ( .A(n4448), .B(n4447), .Z(n4449) );
  NOR U5940 ( .A(n4450), .B(n4449), .Z(n4913) );
  NOR U5941 ( .A(n5315), .B(n4913), .Z(n5322) );
  IV U5942 ( .A(n5322), .Z(n4832) );
  IV U5943 ( .A(n4451), .Z(n4452) );
  NOR U5944 ( .A(n4452), .B(n4457), .Z(n5318) );
  IV U5945 ( .A(n4453), .Z(n4454) );
  NOR U5946 ( .A(n4455), .B(n4454), .Z(n4917) );
  IV U5947 ( .A(n4456), .Z(n4458) );
  NOR U5948 ( .A(n4458), .B(n4457), .Z(n4914) );
  NOR U5949 ( .A(n4917), .B(n4914), .Z(n4831) );
  IV U5950 ( .A(n4459), .Z(n4460) );
  NOR U5951 ( .A(n4461), .B(n4460), .Z(n4923) );
  IV U5952 ( .A(n4462), .Z(n4464) );
  NOR U5953 ( .A(n4464), .B(n4463), .Z(n4920) );
  NOR U5954 ( .A(n4923), .B(n4920), .Z(n4830) );
  NOR U5955 ( .A(n4465), .B(n4927), .Z(n4829) );
  IV U5956 ( .A(n4466), .Z(n4467) );
  NOR U5957 ( .A(n4467), .B(n4469), .Z(n5303) );
  IV U5958 ( .A(n4468), .Z(n4472) );
  NOR U5959 ( .A(n4470), .B(n4469), .Z(n4471) );
  IV U5960 ( .A(n4471), .Z(n4474) );
  NOR U5961 ( .A(n4472), .B(n4474), .Z(n4933) );
  IV U5962 ( .A(n4473), .Z(n4475) );
  NOR U5963 ( .A(n4475), .B(n4474), .Z(n4944) );
  NOR U5964 ( .A(n4476), .B(n4952), .Z(n4480) );
  IV U5965 ( .A(n4477), .Z(n4479) );
  NOR U5966 ( .A(n4479), .B(n4478), .Z(n4948) );
  NOR U5967 ( .A(n4480), .B(n4948), .Z(n4826) );
  IV U5968 ( .A(n4481), .Z(n4483) );
  NOR U5969 ( .A(n4483), .B(n4482), .Z(n4955) );
  IV U5970 ( .A(n4484), .Z(n4485) );
  NOR U5971 ( .A(n4486), .B(n4485), .Z(n4966) );
  IV U5972 ( .A(n4487), .Z(n4489) );
  NOR U5973 ( .A(n4489), .B(n4488), .Z(n4968) );
  NOR U5974 ( .A(n4966), .B(n4968), .Z(n4818) );
  IV U5975 ( .A(n4490), .Z(n4492) );
  NOR U5976 ( .A(n4492), .B(n4491), .Z(n5293) );
  IV U5977 ( .A(n4493), .Z(n4494) );
  NOR U5978 ( .A(n4494), .B(n4810), .Z(n5291) );
  NOR U5979 ( .A(n5293), .B(n5291), .Z(n4808) );
  IV U5980 ( .A(n4495), .Z(n4497) );
  NOR U5981 ( .A(n4497), .B(n4496), .Z(n4498) );
  IV U5982 ( .A(n4498), .Z(n4804) );
  IV U5983 ( .A(n4499), .Z(n4501) );
  IV U5984 ( .A(n4500), .Z(n4802) );
  NOR U5985 ( .A(n4501), .B(n4802), .Z(n4505) );
  IV U5986 ( .A(n4502), .Z(n4503) );
  NOR U5987 ( .A(n4503), .B(n4510), .Z(n4504) );
  NOR U5988 ( .A(n4505), .B(n4504), .Z(n4984) );
  IV U5989 ( .A(n4506), .Z(n4508) );
  NOR U5990 ( .A(n4508), .B(n4507), .Z(n4989) );
  IV U5991 ( .A(n4509), .Z(n4511) );
  NOR U5992 ( .A(n4511), .B(n4510), .Z(n4986) );
  NOR U5993 ( .A(n4989), .B(n4986), .Z(n4796) );
  IV U5994 ( .A(n4512), .Z(n5281) );
  NOR U5995 ( .A(n4513), .B(n5281), .Z(n4795) );
  IV U5996 ( .A(n4514), .Z(n4517) );
  IV U5997 ( .A(n4515), .Z(n4516) );
  NOR U5998 ( .A(n4517), .B(n4516), .Z(n5277) );
  IV U5999 ( .A(n4518), .Z(n4519) );
  NOR U6000 ( .A(n4519), .B(n4778), .Z(n4520) );
  IV U6001 ( .A(n4520), .Z(n5264) );
  IV U6002 ( .A(n4521), .Z(n4522) );
  NOR U6003 ( .A(n4523), .B(n4522), .Z(n4524) );
  IV U6004 ( .A(n4524), .Z(n4784) );
  IV U6005 ( .A(n4525), .Z(n4527) );
  IV U6006 ( .A(n4526), .Z(n4781) );
  NOR U6007 ( .A(n4527), .B(n4781), .Z(n5251) );
  IV U6008 ( .A(n4528), .Z(n4529) );
  NOR U6009 ( .A(n4529), .B(n4532), .Z(n5248) );
  IV U6010 ( .A(n4530), .Z(n4531) );
  NOR U6011 ( .A(n4532), .B(n4531), .Z(n5237) );
  IV U6012 ( .A(n4533), .Z(n4535) );
  NOR U6013 ( .A(n4535), .B(n4534), .Z(n5510) );
  IV U6014 ( .A(n4536), .Z(n4537) );
  NOR U6015 ( .A(n4545), .B(n4537), .Z(n5515) );
  NOR U6016 ( .A(n5510), .B(n5515), .Z(n5243) );
  IV U6017 ( .A(n4538), .Z(n4542) );
  IV U6018 ( .A(n4539), .Z(n4550) );
  NOR U6019 ( .A(n4540), .B(n4550), .Z(n4541) );
  IV U6020 ( .A(n4541), .Z(n4547) );
  NOR U6021 ( .A(n4542), .B(n4547), .Z(n5644) );
  IV U6022 ( .A(n4543), .Z(n4544) );
  NOR U6023 ( .A(n4545), .B(n4544), .Z(n5518) );
  NOR U6024 ( .A(n5644), .B(n5518), .Z(n4994) );
  IV U6025 ( .A(n4546), .Z(n4548) );
  NOR U6026 ( .A(n4548), .B(n4547), .Z(n5521) );
  IV U6027 ( .A(n4549), .Z(n4553) );
  NOR U6028 ( .A(n4551), .B(n4550), .Z(n4552) );
  IV U6029 ( .A(n4552), .Z(n4555) );
  NOR U6030 ( .A(n4553), .B(n4555), .Z(n4999) );
  IV U6031 ( .A(n4554), .Z(n4556) );
  NOR U6032 ( .A(n4556), .B(n4555), .Z(n4996) );
  IV U6033 ( .A(n4557), .Z(n4558) );
  NOR U6034 ( .A(n4558), .B(n4561), .Z(n5002) );
  IV U6035 ( .A(n4559), .Z(n4560) );
  NOR U6036 ( .A(n4561), .B(n4560), .Z(n5219) );
  IV U6037 ( .A(n4562), .Z(n4563) );
  NOR U6038 ( .A(n4563), .B(n4771), .Z(n5541) );
  IV U6039 ( .A(n4564), .Z(n4565) );
  NOR U6040 ( .A(n4566), .B(n4565), .Z(n5016) );
  IV U6041 ( .A(n4567), .Z(n4568) );
  NOR U6042 ( .A(n4569), .B(n4568), .Z(n5007) );
  NOR U6043 ( .A(n5016), .B(n5007), .Z(n4769) );
  IV U6044 ( .A(n4570), .Z(n4571) );
  NOR U6045 ( .A(n4571), .B(n4765), .Z(n5212) );
  IV U6046 ( .A(n4572), .Z(n4575) );
  IV U6047 ( .A(n4573), .Z(n4574) );
  NOR U6048 ( .A(n4575), .B(n4574), .Z(n4576) );
  IV U6049 ( .A(n4576), .Z(n5196) );
  IV U6050 ( .A(n4577), .Z(n4579) );
  NOR U6051 ( .A(n4579), .B(n4578), .Z(n5023) );
  NOR U6052 ( .A(n5023), .B(n5021), .Z(n4760) );
  IV U6053 ( .A(n4580), .Z(n4583) );
  NOR U6054 ( .A(n4581), .B(n4741), .Z(n4582) );
  IV U6055 ( .A(n4582), .Z(n4757) );
  NOR U6056 ( .A(n4583), .B(n4757), .Z(n5179) );
  NOR U6057 ( .A(n4584), .B(n5027), .Z(n4746) );
  IV U6058 ( .A(n4585), .Z(n4587) );
  IV U6059 ( .A(n4586), .Z(n4738) );
  NOR U6060 ( .A(n4587), .B(n4738), .Z(n5172) );
  NOR U6061 ( .A(n4746), .B(n5172), .Z(n4736) );
  IV U6062 ( .A(n4588), .Z(n4589) );
  NOR U6063 ( .A(n4590), .B(n4589), .Z(n4595) );
  IV U6064 ( .A(n4591), .Z(n4593) );
  NOR U6065 ( .A(n4593), .B(n4592), .Z(n4594) );
  NOR U6066 ( .A(n4595), .B(n4594), .Z(n5036) );
  IV U6067 ( .A(n4596), .Z(n4597) );
  NOR U6068 ( .A(n4597), .B(n4599), .Z(n5038) );
  IV U6069 ( .A(n4598), .Z(n4600) );
  NOR U6070 ( .A(n4600), .B(n4599), .Z(n5162) );
  IV U6071 ( .A(n4601), .Z(n5052) );
  IV U6072 ( .A(n4610), .Z(n4611) );
  NOR U6073 ( .A(n4611), .B(n4614), .Z(n5121) );
  IV U6074 ( .A(n4612), .Z(n4613) );
  NOR U6075 ( .A(n4614), .B(n4613), .Z(n5056) );
  IV U6076 ( .A(n4615), .Z(n4684) );
  IV U6077 ( .A(n4616), .Z(n4617) );
  NOR U6078 ( .A(n4684), .B(n4617), .Z(n5062) );
  IV U6079 ( .A(n4618), .Z(n4620) );
  NOR U6080 ( .A(n4620), .B(n4619), .Z(n5074) );
  IV U6081 ( .A(n4621), .Z(n4622) );
  NOR U6082 ( .A(n4622), .B(n4624), .Z(n5082) );
  IV U6083 ( .A(n4623), .Z(n4625) );
  NOR U6084 ( .A(n4625), .B(n4624), .Z(n5105) );
  IV U6085 ( .A(n4626), .Z(n4627) );
  NOR U6086 ( .A(n4630), .B(n4627), .Z(n5088) );
  IV U6087 ( .A(n4628), .Z(n4629) );
  NOR U6088 ( .A(n4630), .B(n4629), .Z(n5085) );
  IV U6089 ( .A(n4631), .Z(n4633) );
  IV U6090 ( .A(n4632), .Z(n4635) );
  NOR U6091 ( .A(n4633), .B(n4635), .Z(n5092) );
  IV U6092 ( .A(n4634), .Z(n4636) );
  NOR U6093 ( .A(n4636), .B(n4635), .Z(n4679) );
  IV U6094 ( .A(n4637), .Z(n4639) );
  NOR U6095 ( .A(n4639), .B(n4638), .Z(n4676) );
  NOR U6096 ( .A(n4641), .B(n4640), .Z(n4645) );
  NOR U6097 ( .A(n4643), .B(n4642), .Z(n4644) );
  NOR U6098 ( .A(n4645), .B(n4644), .Z(n4646) );
  IV U6099 ( .A(n4646), .Z(n4673) );
  IV U6100 ( .A(n4647), .Z(n4648) );
  NOR U6101 ( .A(n4649), .B(n4648), .Z(n4670) );
  IV U6102 ( .A(n4650), .Z(n4652) );
  NOR U6103 ( .A(n4652), .B(n4651), .Z(n4656) );
  NOR U6104 ( .A(n4654), .B(n4653), .Z(n4655) );
  NOR U6105 ( .A(n4656), .B(n4655), .Z(n4657) );
  IV U6106 ( .A(n4657), .Z(n4667) );
  NOR U6107 ( .A(n4659), .B(n4658), .Z(n4664) );
  IV U6108 ( .A(n4660), .Z(n4661) );
  NOR U6109 ( .A(n4662), .B(n4661), .Z(n4663) );
  NOR U6110 ( .A(n4664), .B(n4663), .Z(n4665) );
  IV U6111 ( .A(n4665), .Z(n4666) );
  NOR U6112 ( .A(n4667), .B(n4666), .Z(n4668) );
  IV U6113 ( .A(n4668), .Z(n4669) );
  NOR U6114 ( .A(n4670), .B(n4669), .Z(n4671) );
  IV U6115 ( .A(n4671), .Z(n4672) );
  NOR U6116 ( .A(n4673), .B(n4672), .Z(n4674) );
  IV U6117 ( .A(n4674), .Z(n4675) );
  NOR U6118 ( .A(n4676), .B(n4675), .Z(n4677) );
  IV U6119 ( .A(n4677), .Z(n4678) );
  NOR U6120 ( .A(n4679), .B(n4678), .Z(n5094) );
  XOR U6121 ( .A(n5092), .B(n5094), .Z(n5086) );
  XOR U6122 ( .A(n5085), .B(n5086), .Z(n5089) );
  XOR U6123 ( .A(n5088), .B(n5089), .Z(n5106) );
  XOR U6124 ( .A(n5105), .B(n5106), .Z(n5083) );
  XOR U6125 ( .A(n5082), .B(n5083), .Z(n5075) );
  XOR U6126 ( .A(n5074), .B(n5075), .Z(n5079) );
  IV U6127 ( .A(n4680), .Z(n4681) );
  NOR U6128 ( .A(n4684), .B(n4681), .Z(n5077) );
  XOR U6129 ( .A(n5079), .B(n5077), .Z(n5073) );
  IV U6130 ( .A(n4682), .Z(n4683) );
  NOR U6131 ( .A(n4684), .B(n4683), .Z(n5071) );
  XOR U6132 ( .A(n5073), .B(n5071), .Z(n5063) );
  XOR U6133 ( .A(n5062), .B(n5063), .Z(n5066) );
  IV U6134 ( .A(n4685), .Z(n4686) );
  NOR U6135 ( .A(n4694), .B(n4686), .Z(n4687) );
  NOR U6136 ( .A(n4688), .B(n4687), .Z(n4689) );
  NOR U6137 ( .A(n4695), .B(n4689), .Z(n5065) );
  XOR U6138 ( .A(n5066), .B(n5065), .Z(n5059) );
  IV U6139 ( .A(n4690), .Z(n4691) );
  NOR U6140 ( .A(n4692), .B(n4691), .Z(n4700) );
  IV U6141 ( .A(n4693), .Z(n4698) );
  NOR U6142 ( .A(n4695), .B(n4694), .Z(n4696) );
  IV U6143 ( .A(n4696), .Z(n4697) );
  NOR U6144 ( .A(n4698), .B(n4697), .Z(n4699) );
  NOR U6145 ( .A(n4700), .B(n4699), .Z(n5060) );
  XOR U6146 ( .A(n5059), .B(n5060), .Z(n4701) );
  IV U6147 ( .A(n4701), .Z(n5058) );
  XOR U6148 ( .A(n5056), .B(n5058), .Z(n5123) );
  XOR U6149 ( .A(n5121), .B(n5123), .Z(n5119) );
  XOR U6150 ( .A(n5120), .B(n5119), .Z(n5050) );
  XOR U6151 ( .A(n5052), .B(n5050), .Z(n5054) );
  IV U6152 ( .A(n4702), .Z(n5047) );
  NOR U6153 ( .A(n4703), .B(n5047), .Z(n4704) );
  NOR U6154 ( .A(n5053), .B(n4704), .Z(n4705) );
  XOR U6155 ( .A(n5054), .B(n4705), .Z(n5044) );
  IV U6156 ( .A(n4706), .Z(n4708) );
  NOR U6157 ( .A(n4708), .B(n4707), .Z(n5141) );
  IV U6158 ( .A(n4709), .Z(n4710) );
  NOR U6159 ( .A(n4710), .B(n4713), .Z(n5043) );
  NOR U6160 ( .A(n5141), .B(n5043), .Z(n4711) );
  XOR U6161 ( .A(n5044), .B(n4711), .Z(n5153) );
  IV U6162 ( .A(n4712), .Z(n4714) );
  NOR U6163 ( .A(n4714), .B(n4713), .Z(n5151) );
  XOR U6164 ( .A(n5153), .B(n5151), .Z(n5155) );
  IV U6165 ( .A(n4715), .Z(n4716) );
  NOR U6166 ( .A(n4717), .B(n4716), .Z(n5154) );
  IV U6167 ( .A(n4718), .Z(n4720) );
  NOR U6168 ( .A(n4720), .B(n4719), .Z(n5041) );
  NOR U6169 ( .A(n5154), .B(n5041), .Z(n4721) );
  XOR U6170 ( .A(n5155), .B(n4721), .Z(n4722) );
  IV U6171 ( .A(n4722), .Z(n5163) );
  XOR U6172 ( .A(n5162), .B(n5163), .Z(n5040) );
  XOR U6173 ( .A(n5038), .B(n5040), .Z(n4729) );
  IV U6174 ( .A(n4723), .Z(n4727) );
  NOR U6175 ( .A(n4725), .B(n4724), .Z(n4726) );
  IV U6176 ( .A(n4726), .Z(n4733) );
  NOR U6177 ( .A(n4727), .B(n4733), .Z(n4730) );
  IV U6178 ( .A(n4730), .Z(n4728) );
  NOR U6179 ( .A(n4729), .B(n4728), .Z(n5566) );
  IV U6180 ( .A(n4729), .Z(n4731) );
  NOR U6181 ( .A(n4731), .B(n4730), .Z(n5032) );
  IV U6182 ( .A(n4732), .Z(n4734) );
  NOR U6183 ( .A(n4734), .B(n4733), .Z(n5030) );
  XOR U6184 ( .A(n5032), .B(n5030), .Z(n4735) );
  NOR U6185 ( .A(n5566), .B(n4735), .Z(n5034) );
  XOR U6186 ( .A(n5036), .B(n5034), .Z(n5173) );
  XOR U6187 ( .A(n4736), .B(n5173), .Z(n4749) );
  IV U6188 ( .A(n4737), .Z(n4739) );
  NOR U6189 ( .A(n4739), .B(n4738), .Z(n4750) );
  IV U6190 ( .A(n4740), .Z(n4742) );
  NOR U6191 ( .A(n4742), .B(n4741), .Z(n4745) );
  NOR U6192 ( .A(n4750), .B(n4745), .Z(n4743) );
  IV U6193 ( .A(n4743), .Z(n4744) );
  NOR U6194 ( .A(n4749), .B(n4744), .Z(n4755) );
  IV U6195 ( .A(n4745), .Z(n4748) );
  XOR U6196 ( .A(n4746), .B(n5173), .Z(n4747) );
  NOR U6197 ( .A(n4748), .B(n4747), .Z(n4754) );
  IV U6198 ( .A(n4749), .Z(n4752) );
  IV U6199 ( .A(n4750), .Z(n4751) );
  NOR U6200 ( .A(n4752), .B(n4751), .Z(n4753) );
  NOR U6201 ( .A(n4754), .B(n4753), .Z(n5605) );
  IV U6202 ( .A(n5605), .Z(n5175) );
  NOR U6203 ( .A(n4755), .B(n5175), .Z(n5182) );
  IV U6204 ( .A(n4756), .Z(n4758) );
  NOR U6205 ( .A(n4758), .B(n4757), .Z(n4759) );
  IV U6206 ( .A(n4759), .Z(n5183) );
  XOR U6207 ( .A(n5182), .B(n5183), .Z(n5180) );
  XOR U6208 ( .A(n5179), .B(n5180), .Z(n5024) );
  XOR U6209 ( .A(n4760), .B(n5024), .Z(n5194) );
  XOR U6210 ( .A(n5196), .B(n5194), .Z(n5210) );
  IV U6211 ( .A(n4761), .Z(n4762) );
  NOR U6212 ( .A(n4763), .B(n4762), .Z(n5019) );
  IV U6213 ( .A(n4764), .Z(n4766) );
  NOR U6214 ( .A(n4766), .B(n4765), .Z(n5209) );
  NOR U6215 ( .A(n5019), .B(n5209), .Z(n4767) );
  XOR U6216 ( .A(n5210), .B(n4767), .Z(n4768) );
  IV U6217 ( .A(n4768), .Z(n5213) );
  XOR U6218 ( .A(n5212), .B(n5213), .Z(n5017) );
  IV U6219 ( .A(n5017), .Z(n5010) );
  XOR U6220 ( .A(n4769), .B(n5010), .Z(n5542) );
  XOR U6221 ( .A(n5541), .B(n5542), .Z(n5529) );
  IV U6222 ( .A(n4770), .Z(n4772) );
  NOR U6223 ( .A(n4772), .B(n4771), .Z(n5008) );
  IV U6224 ( .A(n4773), .Z(n4775) );
  NOR U6225 ( .A(n4775), .B(n4774), .Z(n5005) );
  NOR U6226 ( .A(n5008), .B(n5005), .Z(n5530) );
  XOR U6227 ( .A(n5529), .B(n5530), .Z(n4776) );
  IV U6228 ( .A(n4776), .Z(n5220) );
  XOR U6229 ( .A(n5219), .B(n5220), .Z(n5003) );
  XOR U6230 ( .A(n5002), .B(n5003), .Z(n4998) );
  XOR U6231 ( .A(n4996), .B(n4998), .Z(n5001) );
  XOR U6232 ( .A(n4999), .B(n5001), .Z(n5519) );
  XOR U6233 ( .A(n5521), .B(n5519), .Z(n4993) );
  XOR U6234 ( .A(n4994), .B(n4993), .Z(n5242) );
  XOR U6235 ( .A(n5243), .B(n5242), .Z(n5238) );
  XOR U6236 ( .A(n5237), .B(n5238), .Z(n5249) );
  XOR U6237 ( .A(n5248), .B(n5249), .Z(n5253) );
  XOR U6238 ( .A(n5251), .B(n5253), .Z(n5255) );
  NOR U6239 ( .A(n4784), .B(n5255), .Z(n5493) );
  IV U6240 ( .A(n4777), .Z(n4779) );
  NOR U6241 ( .A(n4779), .B(n4778), .Z(n5258) );
  IV U6242 ( .A(n4780), .Z(n4782) );
  NOR U6243 ( .A(n4782), .B(n4781), .Z(n4783) );
  IV U6244 ( .A(n4783), .Z(n5256) );
  XOR U6245 ( .A(n5256), .B(n5255), .Z(n5259) );
  XOR U6246 ( .A(n5258), .B(n5259), .Z(n4786) );
  NOR U6247 ( .A(n5259), .B(n4784), .Z(n4785) );
  NOR U6248 ( .A(n4786), .B(n4785), .Z(n4787) );
  NOR U6249 ( .A(n5493), .B(n4787), .Z(n5262) );
  XOR U6250 ( .A(n5264), .B(n5262), .Z(n5273) );
  IV U6251 ( .A(n4788), .Z(n4789) );
  NOR U6252 ( .A(n4790), .B(n4789), .Z(n5272) );
  NOR U6253 ( .A(n4792), .B(n4791), .Z(n5269) );
  NOR U6254 ( .A(n5272), .B(n5269), .Z(n4793) );
  XOR U6255 ( .A(n5273), .B(n4793), .Z(n4794) );
  IV U6256 ( .A(n4794), .Z(n5282) );
  XOR U6257 ( .A(n5266), .B(n5282), .Z(n5278) );
  XOR U6258 ( .A(n5277), .B(n5278), .Z(n4990) );
  XOR U6259 ( .A(n4795), .B(n4990), .Z(n4987) );
  XOR U6260 ( .A(n4796), .B(n4987), .Z(n4983) );
  XOR U6261 ( .A(n4984), .B(n4983), .Z(n4981) );
  NOR U6262 ( .A(n4804), .B(n4981), .Z(n5675) );
  IV U6263 ( .A(n4797), .Z(n4799) );
  NOR U6264 ( .A(n4799), .B(n4798), .Z(n4976) );
  IV U6265 ( .A(n4800), .Z(n4801) );
  NOR U6266 ( .A(n4802), .B(n4801), .Z(n4803) );
  IV U6267 ( .A(n4803), .Z(n4982) );
  XOR U6268 ( .A(n4982), .B(n4981), .Z(n4977) );
  XOR U6269 ( .A(n4976), .B(n4977), .Z(n4806) );
  NOR U6270 ( .A(n4977), .B(n4804), .Z(n4805) );
  NOR U6271 ( .A(n4806), .B(n4805), .Z(n4807) );
  NOR U6272 ( .A(n5675), .B(n4807), .Z(n5290) );
  XOR U6273 ( .A(n4808), .B(n5290), .Z(n4972) );
  IV U6274 ( .A(n4809), .Z(n4811) );
  NOR U6275 ( .A(n4811), .B(n4810), .Z(n4812) );
  IV U6276 ( .A(n4812), .Z(n4971) );
  XOR U6277 ( .A(n4972), .B(n4971), .Z(n4973) );
  IV U6278 ( .A(n4813), .Z(n4817) );
  NOR U6279 ( .A(n4817), .B(n4814), .Z(n5461) );
  IV U6280 ( .A(n4815), .Z(n4816) );
  NOR U6281 ( .A(n4817), .B(n4816), .Z(n5456) );
  NOR U6282 ( .A(n5461), .B(n5456), .Z(n4974) );
  XOR U6283 ( .A(n4973), .B(n4974), .Z(n4970) );
  XOR U6284 ( .A(n4818), .B(n4970), .Z(n4964) );
  IV U6285 ( .A(n4819), .Z(n4821) );
  NOR U6286 ( .A(n4821), .B(n4820), .Z(n4963) );
  IV U6287 ( .A(n4822), .Z(n4824) );
  NOR U6288 ( .A(n4824), .B(n4823), .Z(n5298) );
  NOR U6289 ( .A(n4963), .B(n5298), .Z(n4825) );
  XOR U6290 ( .A(n4964), .B(n4825), .Z(n4957) );
  XOR U6291 ( .A(n4955), .B(n4957), .Z(n4949) );
  XOR U6292 ( .A(n4826), .B(n4949), .Z(n4937) );
  XOR U6293 ( .A(n4827), .B(n4937), .Z(n4946) );
  XOR U6294 ( .A(n4944), .B(n4946), .Z(n4935) );
  XOR U6295 ( .A(n4933), .B(n4935), .Z(n5311) );
  XOR U6296 ( .A(n5303), .B(n5311), .Z(n5306) );
  XOR U6297 ( .A(n4828), .B(n5306), .Z(n4926) );
  XOR U6298 ( .A(n4829), .B(n4926), .Z(n4922) );
  XOR U6299 ( .A(n4830), .B(n4922), .Z(n4915) );
  XOR U6300 ( .A(n4831), .B(n4915), .Z(n5320) );
  XOR U6301 ( .A(n5318), .B(n5320), .Z(n5321) );
  XOR U6302 ( .A(n4832), .B(n5321), .Z(n5324) );
  XOR U6303 ( .A(n5323), .B(n5324), .Z(n5347) );
  IV U6304 ( .A(n5347), .Z(n4840) );
  IV U6305 ( .A(n4833), .Z(n4835) );
  NOR U6306 ( .A(n4835), .B(n4834), .Z(n4911) );
  IV U6307 ( .A(n4836), .Z(n4837) );
  NOR U6308 ( .A(n4838), .B(n4837), .Z(n5345) );
  NOR U6309 ( .A(n4911), .B(n5345), .Z(n4839) );
  XOR U6310 ( .A(n4840), .B(n4839), .Z(n5344) );
  XOR U6311 ( .A(n5342), .B(n5344), .Z(n4908) );
  IV U6312 ( .A(n4842), .Z(n4841) );
  NOR U6313 ( .A(n4843), .B(n4841), .Z(n4907) );
  XOR U6314 ( .A(n4843), .B(n4842), .Z(n4846) );
  IV U6315 ( .A(n4844), .Z(n4845) );
  NOR U6316 ( .A(n4846), .B(n4845), .Z(n4905) );
  NOR U6317 ( .A(n4907), .B(n4905), .Z(n4847) );
  XOR U6318 ( .A(n4908), .B(n4847), .Z(n4899) );
  XOR U6319 ( .A(n4848), .B(n4899), .Z(n4897) );
  XOR U6320 ( .A(n4849), .B(n4897), .Z(n4886) );
  NOR U6321 ( .A(n4851), .B(n4850), .Z(n4852) );
  IV U6322 ( .A(n4852), .Z(n4853) );
  NOR U6323 ( .A(n4854), .B(n4853), .Z(n4855) );
  IV U6324 ( .A(n4855), .Z(n4887) );
  NOR U6325 ( .A(n4856), .B(n4887), .Z(n4857) );
  XOR U6326 ( .A(n4886), .B(n4857), .Z(n4884) );
  XOR U6327 ( .A(n4882), .B(n4884), .Z(n5357) );
  XOR U6328 ( .A(n4880), .B(n5357), .Z(n5364) );
  IV U6329 ( .A(n4858), .Z(n4860) );
  NOR U6330 ( .A(n4860), .B(n4859), .Z(n5361) );
  NOR U6331 ( .A(n5361), .B(n5363), .Z(n4861) );
  XOR U6332 ( .A(n5364), .B(n4861), .Z(n5369) );
  IV U6333 ( .A(n4862), .Z(n4863) );
  NOR U6334 ( .A(n4864), .B(n4863), .Z(n5365) );
  IV U6335 ( .A(n4865), .Z(n4866) );
  NOR U6336 ( .A(n4866), .B(n4870), .Z(n5370) );
  NOR U6337 ( .A(n5365), .B(n5370), .Z(n4867) );
  XOR U6338 ( .A(n5369), .B(n4867), .Z(n4875) );
  IV U6339 ( .A(n4868), .Z(n4869) );
  NOR U6340 ( .A(n4870), .B(n4869), .Z(n4873) );
  XOR U6341 ( .A(n4875), .B(n4873), .Z(n5782) );
  NOR U6342 ( .A(n4871), .B(n5781), .Z(n4872) );
  IV U6343 ( .A(n4872), .Z(n4876) );
  XOR U6344 ( .A(n5782), .B(n4876), .Z(o[4]) );
  IV U6345 ( .A(n4873), .Z(n4874) );
  NOR U6346 ( .A(n4875), .B(n4874), .Z(n5790) );
  NOR U6347 ( .A(n5782), .B(n4876), .Z(n4877) );
  NOR U6348 ( .A(n5790), .B(n4877), .Z(n5373) );
  IV U6349 ( .A(n4878), .Z(n4879) );
  NOR U6350 ( .A(n5364), .B(n4879), .Z(n5359) );
  IV U6351 ( .A(n5359), .Z(n5354) );
  IV U6352 ( .A(n4880), .Z(n4881) );
  NOR U6353 ( .A(n5357), .B(n4881), .Z(n5767) );
  IV U6354 ( .A(n4882), .Z(n4883) );
  NOR U6355 ( .A(n4884), .B(n4883), .Z(n5385) );
  IV U6356 ( .A(n4885), .Z(n4889) );
  NOR U6357 ( .A(n4887), .B(n4886), .Z(n4888) );
  IV U6358 ( .A(n4888), .Z(n4891) );
  NOR U6359 ( .A(n4889), .B(n4891), .Z(n5387) );
  NOR U6360 ( .A(n5385), .B(n5387), .Z(n5352) );
  IV U6361 ( .A(n4890), .Z(n4892) );
  NOR U6362 ( .A(n4892), .B(n4891), .Z(n5390) );
  IV U6363 ( .A(n4893), .Z(n4894) );
  NOR U6364 ( .A(n4897), .B(n4894), .Z(n5763) );
  NOR U6365 ( .A(n5390), .B(n5763), .Z(n5351) );
  IV U6366 ( .A(n4895), .Z(n4896) );
  NOR U6367 ( .A(n4897), .B(n4896), .Z(n5757) );
  IV U6368 ( .A(n4898), .Z(n4901) );
  IV U6369 ( .A(n4899), .Z(n4900) );
  NOR U6370 ( .A(n4901), .B(n4900), .Z(n5755) );
  IV U6371 ( .A(n4902), .Z(n4904) );
  XOR U6372 ( .A(n4907), .B(n4908), .Z(n4903) );
  NOR U6373 ( .A(n4904), .B(n4903), .Z(n5393) );
  IV U6374 ( .A(n4905), .Z(n4906) );
  NOR U6375 ( .A(n4906), .B(n4908), .Z(n5396) );
  IV U6376 ( .A(n4907), .Z(n4909) );
  NOR U6377 ( .A(n4909), .B(n4908), .Z(n5398) );
  XOR U6378 ( .A(n5396), .B(n5398), .Z(n4910) );
  NOR U6379 ( .A(n5393), .B(n4910), .Z(n5349) );
  IV U6380 ( .A(n4911), .Z(n4912) );
  NOR U6381 ( .A(n4912), .B(n5324), .Z(n5336) );
  IV U6382 ( .A(n4913), .Z(n5314) );
  IV U6383 ( .A(n4914), .Z(n4916) );
  IV U6384 ( .A(n4915), .Z(n4918) );
  NOR U6385 ( .A(n4916), .B(n4918), .Z(n5717) );
  IV U6386 ( .A(n4917), .Z(n4919) );
  NOR U6387 ( .A(n4919), .B(n4918), .Z(n5720) );
  IV U6388 ( .A(n4920), .Z(n4921) );
  NOR U6389 ( .A(n4922), .B(n4921), .Z(n5412) );
  IV U6390 ( .A(n4923), .Z(n4924) );
  NOR U6391 ( .A(n4926), .B(n4924), .Z(n5708) );
  IV U6392 ( .A(n4925), .Z(n4929) );
  NOR U6393 ( .A(n4927), .B(n4926), .Z(n4928) );
  IV U6394 ( .A(n4928), .Z(n4931) );
  NOR U6395 ( .A(n4929), .B(n4931), .Z(n5415) );
  IV U6396 ( .A(n4930), .Z(n4932) );
  NOR U6397 ( .A(n4932), .B(n4931), .Z(n5421) );
  IV U6398 ( .A(n4933), .Z(n4934) );
  NOR U6399 ( .A(n4935), .B(n4934), .Z(n4936) );
  IV U6400 ( .A(n4936), .Z(n5699) );
  IV U6401 ( .A(n4937), .Z(n4942) );
  IV U6402 ( .A(n4938), .Z(n4939) );
  NOR U6403 ( .A(n4942), .B(n4939), .Z(n5436) );
  IV U6404 ( .A(n4940), .Z(n4941) );
  NOR U6405 ( .A(n4942), .B(n4941), .Z(n5433) );
  NOR U6406 ( .A(n5436), .B(n5433), .Z(n4943) );
  IV U6407 ( .A(n4943), .Z(n4947) );
  IV U6408 ( .A(n4944), .Z(n4945) );
  NOR U6409 ( .A(n4946), .B(n4945), .Z(n5431) );
  NOR U6410 ( .A(n4947), .B(n5431), .Z(n5302) );
  IV U6411 ( .A(n4948), .Z(n4950) );
  NOR U6412 ( .A(n4950), .B(n4949), .Z(n5441) );
  IV U6413 ( .A(n4951), .Z(n4954) );
  NOR U6414 ( .A(n4957), .B(n4952), .Z(n4953) );
  IV U6415 ( .A(n4953), .Z(n4959) );
  NOR U6416 ( .A(n4954), .B(n4959), .Z(n5438) );
  IV U6417 ( .A(n4955), .Z(n4956) );
  NOR U6418 ( .A(n4957), .B(n4956), .Z(n4962) );
  IV U6419 ( .A(n4958), .Z(n4960) );
  NOR U6420 ( .A(n4960), .B(n4959), .Z(n4961) );
  NOR U6421 ( .A(n4962), .B(n4961), .Z(n5450) );
  IV U6422 ( .A(n5450), .Z(n5301) );
  IV U6423 ( .A(n4963), .Z(n4965) );
  IV U6424 ( .A(n4964), .Z(n5299) );
  NOR U6425 ( .A(n4965), .B(n5299), .Z(n5453) );
  IV U6426 ( .A(n4966), .Z(n4967) );
  NOR U6427 ( .A(n4967), .B(n4970), .Z(n5692) );
  IV U6428 ( .A(n4968), .Z(n4969) );
  NOR U6429 ( .A(n4970), .B(n4969), .Z(n5689) );
  NOR U6430 ( .A(n4972), .B(n4971), .Z(n5469) );
  IV U6431 ( .A(n4973), .Z(n5463) );
  NOR U6432 ( .A(n4974), .B(n5463), .Z(n4975) );
  NOR U6433 ( .A(n5469), .B(n4975), .Z(n5297) );
  IV U6434 ( .A(n4976), .Z(n4979) );
  IV U6435 ( .A(n4977), .Z(n4978) );
  NOR U6436 ( .A(n4979), .B(n4978), .Z(n4980) );
  IV U6437 ( .A(n4980), .Z(n5473) );
  NOR U6438 ( .A(n4982), .B(n4981), .Z(n5480) );
  NOR U6439 ( .A(n5480), .B(n5675), .Z(n5289) );
  IV U6440 ( .A(n4983), .Z(n4985) );
  NOR U6441 ( .A(n4985), .B(n4984), .Z(n5678) );
  IV U6442 ( .A(n4986), .Z(n4988) );
  NOR U6443 ( .A(n4988), .B(n4987), .Z(n5485) );
  IV U6444 ( .A(n4989), .Z(n4991) );
  NOR U6445 ( .A(n4991), .B(n4990), .Z(n5482) );
  IV U6446 ( .A(n5521), .Z(n4992) );
  NOR U6447 ( .A(n4992), .B(n5519), .Z(n5645) );
  NOR U6448 ( .A(n4994), .B(n4993), .Z(n4995) );
  NOR U6449 ( .A(n5645), .B(n4995), .Z(n5236) );
  IV U6450 ( .A(n4996), .Z(n4997) );
  NOR U6451 ( .A(n4998), .B(n4997), .Z(n5636) );
  IV U6452 ( .A(n4999), .Z(n5000) );
  NOR U6453 ( .A(n5001), .B(n5000), .Z(n5527) );
  NOR U6454 ( .A(n5636), .B(n5527), .Z(n5235) );
  IV U6455 ( .A(n5002), .Z(n5004) );
  NOR U6456 ( .A(n5004), .B(n5003), .Z(n5224) );
  IV U6457 ( .A(n5005), .Z(n5006) );
  NOR U6458 ( .A(n5006), .B(n5529), .Z(n5218) );
  IV U6459 ( .A(n5007), .Z(n5009) );
  NOR U6460 ( .A(n5009), .B(n5017), .Z(n5534) );
  NOR U6461 ( .A(n5541), .B(n5008), .Z(n5014) );
  XOR U6462 ( .A(n5016), .B(n5010), .Z(n5012) );
  NOR U6463 ( .A(n5010), .B(n5009), .Z(n5011) );
  NOR U6464 ( .A(n5012), .B(n5011), .Z(n5013) );
  NOR U6465 ( .A(n5014), .B(n5013), .Z(n5015) );
  NOR U6466 ( .A(n5534), .B(n5015), .Z(n5217) );
  IV U6467 ( .A(n5016), .Z(n5018) );
  NOR U6468 ( .A(n5018), .B(n5017), .Z(n5545) );
  IV U6469 ( .A(n5019), .Z(n5020) );
  NOR U6470 ( .A(n5020), .B(n5210), .Z(n5537) );
  IV U6471 ( .A(n5021), .Z(n5022) );
  NOR U6472 ( .A(n5022), .B(n5024), .Z(n5202) );
  IV U6473 ( .A(n5023), .Z(n5025) );
  NOR U6474 ( .A(n5025), .B(n5024), .Z(n5191) );
  IV U6475 ( .A(n5191), .Z(n5178) );
  IV U6476 ( .A(n5026), .Z(n5029) );
  NOR U6477 ( .A(n5027), .B(n5173), .Z(n5028) );
  IV U6478 ( .A(n5028), .Z(n5170) );
  NOR U6479 ( .A(n5029), .B(n5170), .Z(n5569) );
  IV U6480 ( .A(n5030), .Z(n5031) );
  NOR U6481 ( .A(n5032), .B(n5031), .Z(n5573) );
  NOR U6482 ( .A(n5566), .B(n5573), .Z(n5033) );
  IV U6483 ( .A(n5033), .Z(n5037) );
  IV U6484 ( .A(n5034), .Z(n5035) );
  NOR U6485 ( .A(n5036), .B(n5035), .Z(n5572) );
  NOR U6486 ( .A(n5037), .B(n5572), .Z(n5168) );
  IV U6487 ( .A(n5038), .Z(n5039) );
  NOR U6488 ( .A(n5040), .B(n5039), .Z(n5166) );
  IV U6489 ( .A(n5166), .Z(n5161) );
  IV U6490 ( .A(n5041), .Z(n5042) );
  NOR U6491 ( .A(n5042), .B(n5155), .Z(n5580) );
  IV U6492 ( .A(n5043), .Z(n5045) );
  IV U6493 ( .A(n5044), .Z(n5142) );
  NOR U6494 ( .A(n5045), .B(n5142), .Z(n5150) );
  IV U6495 ( .A(n5046), .Z(n5049) );
  NOR U6496 ( .A(n5047), .B(n5054), .Z(n5048) );
  IV U6497 ( .A(n5048), .Z(n5145) );
  NOR U6498 ( .A(n5049), .B(n5145), .Z(n5140) );
  IV U6499 ( .A(n5050), .Z(n5051) );
  NOR U6500 ( .A(n5052), .B(n5051), .Z(n5137) );
  IV U6501 ( .A(n5053), .Z(n5055) );
  NOR U6502 ( .A(n5055), .B(n5054), .Z(n5134) );
  IV U6503 ( .A(n5056), .Z(n5057) );
  NOR U6504 ( .A(n5058), .B(n5057), .Z(n5131) );
  NOR U6505 ( .A(n5060), .B(n5059), .Z(n5061) );
  IV U6506 ( .A(n5061), .Z(n5118) );
  IV U6507 ( .A(n5062), .Z(n5064) );
  NOR U6508 ( .A(n5064), .B(n5063), .Z(n5069) );
  IV U6509 ( .A(n5065), .Z(n5067) );
  NOR U6510 ( .A(n5067), .B(n5066), .Z(n5068) );
  NOR U6511 ( .A(n5069), .B(n5068), .Z(n5070) );
  IV U6512 ( .A(n5070), .Z(n5116) );
  IV U6513 ( .A(n5071), .Z(n5072) );
  NOR U6514 ( .A(n5073), .B(n5072), .Z(n5113) );
  IV U6515 ( .A(n5074), .Z(n5076) );
  NOR U6516 ( .A(n5076), .B(n5075), .Z(n5081) );
  IV U6517 ( .A(n5077), .Z(n5078) );
  NOR U6518 ( .A(n5079), .B(n5078), .Z(n5080) );
  NOR U6519 ( .A(n5081), .B(n5080), .Z(n5111) );
  IV U6520 ( .A(n5082), .Z(n5084) );
  NOR U6521 ( .A(n5084), .B(n5083), .Z(n5103) );
  IV U6522 ( .A(n5085), .Z(n5087) );
  NOR U6523 ( .A(n5087), .B(n5086), .Z(n5091) );
  IV U6524 ( .A(n5088), .Z(n5090) );
  NOR U6525 ( .A(n5090), .B(n5089), .Z(n5098) );
  NOR U6526 ( .A(n5091), .B(n5098), .Z(n5095) );
  IV U6527 ( .A(n5092), .Z(n5093) );
  NOR U6528 ( .A(n5094), .B(n5093), .Z(n5096) );
  NOR U6529 ( .A(n5095), .B(n5096), .Z(n5100) );
  IV U6530 ( .A(n5096), .Z(n5097) );
  NOR U6531 ( .A(n5098), .B(n5097), .Z(n5099) );
  NOR U6532 ( .A(n5100), .B(n5099), .Z(n5101) );
  IV U6533 ( .A(n5101), .Z(n5102) );
  NOR U6534 ( .A(n5103), .B(n5102), .Z(n5104) );
  IV U6535 ( .A(n5104), .Z(n5109) );
  IV U6536 ( .A(n5105), .Z(n5107) );
  NOR U6537 ( .A(n5107), .B(n5106), .Z(n5108) );
  NOR U6538 ( .A(n5109), .B(n5108), .Z(n5110) );
  XOR U6539 ( .A(n5111), .B(n5110), .Z(n5112) );
  NOR U6540 ( .A(n5113), .B(n5112), .Z(n5114) );
  IV U6541 ( .A(n5114), .Z(n5115) );
  NOR U6542 ( .A(n5116), .B(n5115), .Z(n5117) );
  XOR U6543 ( .A(n5118), .B(n5117), .Z(n5128) );
  NOR U6544 ( .A(n5120), .B(n5119), .Z(n5125) );
  IV U6545 ( .A(n5121), .Z(n5122) );
  NOR U6546 ( .A(n5123), .B(n5122), .Z(n5124) );
  NOR U6547 ( .A(n5125), .B(n5124), .Z(n5126) );
  IV U6548 ( .A(n5126), .Z(n5127) );
  NOR U6549 ( .A(n5128), .B(n5127), .Z(n5129) );
  IV U6550 ( .A(n5129), .Z(n5130) );
  NOR U6551 ( .A(n5131), .B(n5130), .Z(n5132) );
  IV U6552 ( .A(n5132), .Z(n5133) );
  NOR U6553 ( .A(n5134), .B(n5133), .Z(n5135) );
  IV U6554 ( .A(n5135), .Z(n5136) );
  NOR U6555 ( .A(n5137), .B(n5136), .Z(n5138) );
  IV U6556 ( .A(n5138), .Z(n5139) );
  NOR U6557 ( .A(n5140), .B(n5139), .Z(n5587) );
  IV U6558 ( .A(n5141), .Z(n5143) );
  NOR U6559 ( .A(n5143), .B(n5142), .Z(n5148) );
  IV U6560 ( .A(n5144), .Z(n5146) );
  NOR U6561 ( .A(n5146), .B(n5145), .Z(n5147) );
  NOR U6562 ( .A(n5148), .B(n5147), .Z(n5588) );
  XOR U6563 ( .A(n5587), .B(n5588), .Z(n5149) );
  NOR U6564 ( .A(n5150), .B(n5149), .Z(n5583) );
  IV U6565 ( .A(n5583), .Z(n5159) );
  IV U6566 ( .A(n5151), .Z(n5152) );
  NOR U6567 ( .A(n5153), .B(n5152), .Z(n5158) );
  IV U6568 ( .A(n5154), .Z(n5156) );
  NOR U6569 ( .A(n5156), .B(n5155), .Z(n5157) );
  NOR U6570 ( .A(n5158), .B(n5157), .Z(n5582) );
  XOR U6571 ( .A(n5159), .B(n5582), .Z(n5590) );
  XOR U6572 ( .A(n5580), .B(n5590), .Z(n5160) );
  NOR U6573 ( .A(n5161), .B(n5160), .Z(n5584) );
  IV U6574 ( .A(n5162), .Z(n5164) );
  NOR U6575 ( .A(n5164), .B(n5163), .Z(n5589) );
  NOR U6576 ( .A(n5580), .B(n5589), .Z(n5165) );
  XOR U6577 ( .A(n5165), .B(n5590), .Z(n5565) );
  NOR U6578 ( .A(n5166), .B(n5565), .Z(n5167) );
  NOR U6579 ( .A(n5584), .B(n5167), .Z(n5574) );
  XOR U6580 ( .A(n5168), .B(n5574), .Z(n5571) );
  XOR U6581 ( .A(n5569), .B(n5571), .Z(n5561) );
  IV U6582 ( .A(n5169), .Z(n5171) );
  NOR U6583 ( .A(n5171), .B(n5170), .Z(n5559) );
  XOR U6584 ( .A(n5561), .B(n5559), .Z(n5604) );
  IV U6585 ( .A(n5172), .Z(n5174) );
  NOR U6586 ( .A(n5174), .B(n5173), .Z(n5557) );
  NOR U6587 ( .A(n5557), .B(n5175), .Z(n5176) );
  XOR U6588 ( .A(n5604), .B(n5176), .Z(n5187) );
  IV U6589 ( .A(n5187), .Z(n5177) );
  NOR U6590 ( .A(n5178), .B(n5177), .Z(n5623) );
  IV U6591 ( .A(n5179), .Z(n5181) );
  NOR U6592 ( .A(n5181), .B(n5180), .Z(n5612) );
  IV U6593 ( .A(n5182), .Z(n5184) );
  NOR U6594 ( .A(n5184), .B(n5183), .Z(n5188) );
  IV U6595 ( .A(n5188), .Z(n5186) );
  XOR U6596 ( .A(n5557), .B(n5604), .Z(n5185) );
  NOR U6597 ( .A(n5186), .B(n5185), .Z(n5555) );
  NOR U6598 ( .A(n5188), .B(n5187), .Z(n5189) );
  NOR U6599 ( .A(n5555), .B(n5189), .Z(n5613) );
  XOR U6600 ( .A(n5612), .B(n5613), .Z(n5190) );
  NOR U6601 ( .A(n5191), .B(n5190), .Z(n5192) );
  NOR U6602 ( .A(n5623), .B(n5192), .Z(n5199) );
  NOR U6603 ( .A(n5202), .B(n5199), .Z(n5193) );
  IV U6604 ( .A(n5193), .Z(n5197) );
  IV U6605 ( .A(n5194), .Z(n5195) );
  NOR U6606 ( .A(n5196), .B(n5195), .Z(n5198) );
  NOR U6607 ( .A(n5197), .B(n5198), .Z(n5208) );
  IV U6608 ( .A(n5198), .Z(n5203) );
  XOR U6609 ( .A(n5202), .B(n5203), .Z(n5201) );
  IV U6610 ( .A(n5199), .Z(n5200) );
  NOR U6611 ( .A(n5201), .B(n5200), .Z(n5206) );
  IV U6612 ( .A(n5202), .Z(n5204) );
  NOR U6613 ( .A(n5204), .B(n5203), .Z(n5205) );
  NOR U6614 ( .A(n5206), .B(n5205), .Z(n5207) );
  IV U6615 ( .A(n5207), .Z(n5628) );
  NOR U6616 ( .A(n5208), .B(n5628), .Z(n5538) );
  XOR U6617 ( .A(n5537), .B(n5538), .Z(n5551) );
  IV U6618 ( .A(n5209), .Z(n5211) );
  NOR U6619 ( .A(n5211), .B(n5210), .Z(n5216) );
  IV U6620 ( .A(n5212), .Z(n5214) );
  NOR U6621 ( .A(n5214), .B(n5213), .Z(n5215) );
  NOR U6622 ( .A(n5216), .B(n5215), .Z(n5553) );
  XOR U6623 ( .A(n5551), .B(n5553), .Z(n5546) );
  XOR U6624 ( .A(n5545), .B(n5546), .Z(n5535) );
  XOR U6625 ( .A(n5217), .B(n5535), .Z(n5228) );
  XOR U6626 ( .A(n5218), .B(n5228), .Z(n5532) );
  IV U6627 ( .A(n5219), .Z(n5221) );
  NOR U6628 ( .A(n5221), .B(n5220), .Z(n5227) );
  NOR U6629 ( .A(n5532), .B(n5227), .Z(n5222) );
  IV U6630 ( .A(n5222), .Z(n5223) );
  NOR U6631 ( .A(n5224), .B(n5223), .Z(n5234) );
  IV U6632 ( .A(n5224), .Z(n5226) );
  IV U6633 ( .A(n5532), .Z(n5225) );
  NOR U6634 ( .A(n5226), .B(n5225), .Z(n5232) );
  IV U6635 ( .A(n5227), .Z(n5230) );
  IV U6636 ( .A(n5228), .Z(n5229) );
  NOR U6637 ( .A(n5230), .B(n5229), .Z(n5231) );
  NOR U6638 ( .A(n5232), .B(n5231), .Z(n5233) );
  IV U6639 ( .A(n5233), .Z(n5927) );
  NOR U6640 ( .A(n5234), .B(n5927), .Z(n5526) );
  XOR U6641 ( .A(n5235), .B(n5526), .Z(n5522) );
  XOR U6642 ( .A(n5236), .B(n5522), .Z(n5244) );
  IV U6643 ( .A(n5244), .Z(n5241) );
  IV U6644 ( .A(n5237), .Z(n5239) );
  NOR U6645 ( .A(n5239), .B(n5238), .Z(n5246) );
  IV U6646 ( .A(n5246), .Z(n5240) );
  NOR U6647 ( .A(n5241), .B(n5240), .Z(n5946) );
  IV U6648 ( .A(n5242), .Z(n5511) );
  NOR U6649 ( .A(n5243), .B(n5511), .Z(n5245) );
  XOR U6650 ( .A(n5245), .B(n5244), .Z(n5506) );
  NOR U6651 ( .A(n5246), .B(n5506), .Z(n5247) );
  NOR U6652 ( .A(n5946), .B(n5247), .Z(n5503) );
  IV U6653 ( .A(n5248), .Z(n5250) );
  NOR U6654 ( .A(n5250), .B(n5249), .Z(n5507) );
  IV U6655 ( .A(n5251), .Z(n5252) );
  NOR U6656 ( .A(n5253), .B(n5252), .Z(n5502) );
  NOR U6657 ( .A(n5507), .B(n5502), .Z(n5254) );
  XOR U6658 ( .A(n5503), .B(n5254), .Z(n5501) );
  NOR U6659 ( .A(n5256), .B(n5255), .Z(n5499) );
  NOR U6660 ( .A(n5499), .B(n5493), .Z(n5257) );
  XOR U6661 ( .A(n5501), .B(n5257), .Z(n5491) );
  IV U6662 ( .A(n5258), .Z(n5261) );
  IV U6663 ( .A(n5259), .Z(n5260) );
  NOR U6664 ( .A(n5261), .B(n5260), .Z(n5495) );
  IV U6665 ( .A(n5262), .Z(n5263) );
  NOR U6666 ( .A(n5264), .B(n5263), .Z(n5490) );
  NOR U6667 ( .A(n5495), .B(n5490), .Z(n5265) );
  XOR U6668 ( .A(n5491), .B(n5265), .Z(n5651) );
  IV U6669 ( .A(n5266), .Z(n5267) );
  NOR U6670 ( .A(n5282), .B(n5267), .Z(n5275) );
  IV U6671 ( .A(n5275), .Z(n5268) );
  NOR U6672 ( .A(n5651), .B(n5268), .Z(n5667) );
  IV U6673 ( .A(n5269), .Z(n5270) );
  NOR U6674 ( .A(n5270), .B(n5273), .Z(n5271) );
  IV U6675 ( .A(n5271), .Z(n5653) );
  IV U6676 ( .A(n5272), .Z(n5274) );
  NOR U6677 ( .A(n5274), .B(n5273), .Z(n5649) );
  XOR U6678 ( .A(n5649), .B(n5651), .Z(n5652) );
  XOR U6679 ( .A(n5653), .B(n5652), .Z(n5656) );
  NOR U6680 ( .A(n5275), .B(n5656), .Z(n5276) );
  NOR U6681 ( .A(n5667), .B(n5276), .Z(n5663) );
  IV U6682 ( .A(n5277), .Z(n5279) );
  NOR U6683 ( .A(n5279), .B(n5278), .Z(n5662) );
  IV U6684 ( .A(n5280), .Z(n5284) );
  NOR U6685 ( .A(n5282), .B(n5281), .Z(n5283) );
  IV U6686 ( .A(n5283), .Z(n5287) );
  NOR U6687 ( .A(n5284), .B(n5287), .Z(n5657) );
  NOR U6688 ( .A(n5662), .B(n5657), .Z(n5285) );
  XOR U6689 ( .A(n5663), .B(n5285), .Z(n5673) );
  IV U6690 ( .A(n5286), .Z(n5288) );
  NOR U6691 ( .A(n5288), .B(n5287), .Z(n5671) );
  XOR U6692 ( .A(n5673), .B(n5671), .Z(n5483) );
  XOR U6693 ( .A(n5482), .B(n5483), .Z(n5487) );
  XOR U6694 ( .A(n5485), .B(n5487), .Z(n5679) );
  XOR U6695 ( .A(n5678), .B(n5679), .Z(n5676) );
  XOR U6696 ( .A(n5289), .B(n5676), .Z(n5472) );
  XOR U6697 ( .A(n5473), .B(n5472), .Z(n5476) );
  IV U6698 ( .A(n5290), .Z(n5294) );
  IV U6699 ( .A(n5291), .Z(n5292) );
  NOR U6700 ( .A(n5294), .B(n5292), .Z(n5467) );
  IV U6701 ( .A(n5293), .Z(n5295) );
  NOR U6702 ( .A(n5295), .B(n5294), .Z(n5475) );
  NOR U6703 ( .A(n5467), .B(n5475), .Z(n5296) );
  XOR U6704 ( .A(n5476), .B(n5296), .Z(n5457) );
  XOR U6705 ( .A(n5297), .B(n5457), .Z(n5691) );
  XOR U6706 ( .A(n5689), .B(n5691), .Z(n5693) );
  XOR U6707 ( .A(n5692), .B(n5693), .Z(n5454) );
  XOR U6708 ( .A(n5453), .B(n5454), .Z(n5448) );
  IV U6709 ( .A(n5298), .Z(n5300) );
  NOR U6710 ( .A(n5300), .B(n5299), .Z(n5446) );
  XOR U6711 ( .A(n5448), .B(n5446), .Z(n5449) );
  XOR U6712 ( .A(n5301), .B(n5449), .Z(n5440) );
  XOR U6713 ( .A(n5438), .B(n5440), .Z(n5443) );
  XOR U6714 ( .A(n5441), .B(n5443), .Z(n5434) );
  XOR U6715 ( .A(n5302), .B(n5434), .Z(n5427) );
  XOR U6716 ( .A(n5699), .B(n5427), .Z(n5426) );
  IV U6717 ( .A(n5303), .Z(n5304) );
  NOR U6718 ( .A(n5304), .B(n5311), .Z(n5428) );
  IV U6719 ( .A(n5305), .Z(n5307) );
  NOR U6720 ( .A(n5307), .B(n5306), .Z(n5424) );
  NOR U6721 ( .A(n5428), .B(n5424), .Z(n5308) );
  XOR U6722 ( .A(n5426), .B(n5308), .Z(n5309) );
  IV U6723 ( .A(n5309), .Z(n5420) );
  IV U6724 ( .A(n5310), .Z(n5312) );
  NOR U6725 ( .A(n5312), .B(n5311), .Z(n5418) );
  XOR U6726 ( .A(n5420), .B(n5418), .Z(n5423) );
  XOR U6727 ( .A(n5421), .B(n5423), .Z(n5417) );
  XOR U6728 ( .A(n5415), .B(n5417), .Z(n5710) );
  XOR U6729 ( .A(n5708), .B(n5710), .Z(n5414) );
  XOR U6730 ( .A(n5412), .B(n5414), .Z(n5722) );
  XOR U6731 ( .A(n5720), .B(n5722), .Z(n5719) );
  XOR U6732 ( .A(n5717), .B(n5719), .Z(n5410) );
  NOR U6733 ( .A(n5321), .B(n5410), .Z(n5313) );
  IV U6734 ( .A(n5313), .Z(n5316) );
  NOR U6735 ( .A(n5314), .B(n5316), .Z(n5737) );
  IV U6736 ( .A(n5315), .Z(n5317) );
  NOR U6737 ( .A(n5317), .B(n5316), .Z(n5743) );
  IV U6738 ( .A(n5318), .Z(n5319) );
  NOR U6739 ( .A(n5320), .B(n5319), .Z(n5409) );
  XOR U6740 ( .A(n5409), .B(n5410), .Z(n5338) );
  IV U6741 ( .A(n5338), .Z(n5329) );
  NOR U6742 ( .A(n5322), .B(n5321), .Z(n5326) );
  IV U6743 ( .A(n5323), .Z(n5325) );
  NOR U6744 ( .A(n5325), .B(n5324), .Z(n5334) );
  NOR U6745 ( .A(n5326), .B(n5334), .Z(n5327) );
  IV U6746 ( .A(n5327), .Z(n5328) );
  NOR U6747 ( .A(n5329), .B(n5328), .Z(n5330) );
  NOR U6748 ( .A(n5743), .B(n5330), .Z(n5331) );
  IV U6749 ( .A(n5331), .Z(n5332) );
  NOR U6750 ( .A(n5737), .B(n5332), .Z(n5333) );
  NOR U6751 ( .A(n5336), .B(n5333), .Z(n5341) );
  IV U6752 ( .A(n5334), .Z(n5335) );
  NOR U6753 ( .A(n5335), .B(n5338), .Z(n5874) );
  IV U6754 ( .A(n5336), .Z(n5337) );
  NOR U6755 ( .A(n5338), .B(n5337), .Z(n5871) );
  NOR U6756 ( .A(n5874), .B(n5871), .Z(n5339) );
  IV U6757 ( .A(n5339), .Z(n5340) );
  NOR U6758 ( .A(n5341), .B(n5340), .Z(n5404) );
  IV U6759 ( .A(n5342), .Z(n5343) );
  NOR U6760 ( .A(n5344), .B(n5343), .Z(n5403) );
  IV U6761 ( .A(n5345), .Z(n5346) );
  NOR U6762 ( .A(n5347), .B(n5346), .Z(n5406) );
  NOR U6763 ( .A(n5403), .B(n5406), .Z(n5348) );
  XOR U6764 ( .A(n5404), .B(n5348), .Z(n5397) );
  XOR U6765 ( .A(n5349), .B(n5397), .Z(n5350) );
  IV U6766 ( .A(n5350), .Z(n5764) );
  XOR U6767 ( .A(n5755), .B(n5764), .Z(n5758) );
  XOR U6768 ( .A(n5757), .B(n5758), .Z(n5391) );
  XOR U6769 ( .A(n5351), .B(n5391), .Z(n5384) );
  XOR U6770 ( .A(n5352), .B(n5384), .Z(n5768) );
  XOR U6771 ( .A(n5767), .B(n5768), .Z(n5353) );
  NOR U6772 ( .A(n5354), .B(n5353), .Z(n5779) );
  IV U6773 ( .A(n5355), .Z(n5356) );
  NOR U6774 ( .A(n5357), .B(n5356), .Z(n5381) );
  NOR U6775 ( .A(n5767), .B(n5381), .Z(n5358) );
  XOR U6776 ( .A(n5358), .B(n5768), .Z(n5774) );
  NOR U6777 ( .A(n5359), .B(n5774), .Z(n5360) );
  NOR U6778 ( .A(n5779), .B(n5360), .Z(n5377) );
  IV U6779 ( .A(n5361), .Z(n5362) );
  NOR U6780 ( .A(n5364), .B(n5362), .Z(n5775) );
  XOR U6781 ( .A(n5364), .B(n5363), .Z(n5367) );
  IV U6782 ( .A(n5365), .Z(n5366) );
  NOR U6783 ( .A(n5367), .B(n5366), .Z(n5378) );
  NOR U6784 ( .A(n5775), .B(n5378), .Z(n5368) );
  XOR U6785 ( .A(n5377), .B(n5368), .Z(n5376) );
  IV U6786 ( .A(n5369), .Z(n5372) );
  IV U6787 ( .A(n5370), .Z(n5371) );
  NOR U6788 ( .A(n5372), .B(n5371), .Z(n5374) );
  XOR U6789 ( .A(n5376), .B(n5374), .Z(n5792) );
  XOR U6790 ( .A(n5373), .B(n5792), .Z(o[5]) );
  IV U6791 ( .A(n5374), .Z(n5375) );
  NOR U6792 ( .A(n5376), .B(n5375), .Z(n5794) );
  IV U6793 ( .A(n5377), .Z(n5380) );
  IV U6794 ( .A(n5378), .Z(n5379) );
  NOR U6795 ( .A(n5380), .B(n5379), .Z(n5805) );
  IV U6796 ( .A(n5381), .Z(n5382) );
  NOR U6797 ( .A(n5768), .B(n5382), .Z(n5383) );
  IV U6798 ( .A(n5383), .Z(n5817) );
  IV U6799 ( .A(n5384), .Z(n5389) );
  IV U6800 ( .A(n5385), .Z(n5386) );
  NOR U6801 ( .A(n5389), .B(n5386), .Z(n5772) );
  IV U6802 ( .A(n5772), .Z(n5766) );
  IV U6803 ( .A(n5387), .Z(n5388) );
  NOR U6804 ( .A(n5389), .B(n5388), .Z(n5834) );
  IV U6805 ( .A(n5390), .Z(n5392) );
  NOR U6806 ( .A(n5392), .B(n5391), .Z(n5828) );
  IV U6807 ( .A(n5393), .Z(n5394) );
  NOR U6808 ( .A(n5397), .B(n5394), .Z(n5850) );
  IV U6809 ( .A(n5398), .Z(n5395) );
  NOR U6810 ( .A(n5395), .B(n5397), .Z(n5402) );
  IV U6811 ( .A(n5396), .Z(n5400) );
  XOR U6812 ( .A(n5398), .B(n5397), .Z(n5399) );
  NOR U6813 ( .A(n5400), .B(n5399), .Z(n5401) );
  NOR U6814 ( .A(n5402), .B(n5401), .Z(n5842) );
  IV U6815 ( .A(n5403), .Z(n5405) );
  IV U6816 ( .A(n5404), .Z(n5408) );
  NOR U6817 ( .A(n5405), .B(n5408), .Z(n5844) );
  IV U6818 ( .A(n5406), .Z(n5407) );
  NOR U6819 ( .A(n5408), .B(n5407), .Z(n5839) );
  NOR U6820 ( .A(n5871), .B(n5839), .Z(n5754) );
  IV U6821 ( .A(n5409), .Z(n5411) );
  NOR U6822 ( .A(n5411), .B(n5410), .Z(n5740) );
  IV U6823 ( .A(n5412), .Z(n5413) );
  NOR U6824 ( .A(n5414), .B(n5413), .Z(n5715) );
  IV U6825 ( .A(n5715), .Z(n5707) );
  IV U6826 ( .A(n5415), .Z(n5416) );
  NOR U6827 ( .A(n5417), .B(n5416), .Z(n5712) );
  IV U6828 ( .A(n5418), .Z(n5419) );
  NOR U6829 ( .A(n5420), .B(n5419), .Z(n6052) );
  IV U6830 ( .A(n5421), .Z(n5422) );
  NOR U6831 ( .A(n5423), .B(n5422), .Z(n6048) );
  NOR U6832 ( .A(n6052), .B(n6048), .Z(n5705) );
  IV U6833 ( .A(n5424), .Z(n5425) );
  NOR U6834 ( .A(n5426), .B(n5425), .Z(n6051) );
  IV U6835 ( .A(n5427), .Z(n5700) );
  IV U6836 ( .A(n5428), .Z(n5429) );
  NOR U6837 ( .A(n5700), .B(n5429), .Z(n5430) );
  IV U6838 ( .A(n5430), .Z(n6039) );
  IV U6839 ( .A(n5431), .Z(n5432) );
  NOR U6840 ( .A(n5432), .B(n5434), .Z(n6035) );
  IV U6841 ( .A(n6035), .Z(n6042) );
  IV U6842 ( .A(n5433), .Z(n5435) );
  NOR U6843 ( .A(n5435), .B(n5434), .Z(n5975) );
  IV U6844 ( .A(n5436), .Z(n5437) );
  NOR U6845 ( .A(n5437), .B(n5443), .Z(n5978) );
  IV U6846 ( .A(n5438), .Z(n5439) );
  NOR U6847 ( .A(n5440), .B(n5439), .Z(n5445) );
  IV U6848 ( .A(n5441), .Z(n5442) );
  NOR U6849 ( .A(n5443), .B(n5442), .Z(n5444) );
  NOR U6850 ( .A(n5445), .B(n5444), .Z(n5984) );
  IV U6851 ( .A(n5446), .Z(n5447) );
  NOR U6852 ( .A(n5448), .B(n5447), .Z(n5452) );
  NOR U6853 ( .A(n5450), .B(n5449), .Z(n5451) );
  NOR U6854 ( .A(n5452), .B(n5451), .Z(n5986) );
  IV U6855 ( .A(n5453), .Z(n5455) );
  NOR U6856 ( .A(n5455), .B(n5454), .Z(n5990) );
  IV U6857 ( .A(n5456), .Z(n5458) );
  IV U6858 ( .A(n5457), .Z(n5470) );
  NOR U6859 ( .A(n5458), .B(n5470), .Z(n5459) );
  IV U6860 ( .A(n5459), .Z(n5460) );
  NOR U6861 ( .A(n5463), .B(n5460), .Z(n6014) );
  IV U6862 ( .A(n5461), .Z(n5466) );
  XOR U6863 ( .A(n5475), .B(n5476), .Z(n5462) );
  NOR U6864 ( .A(n5463), .B(n5462), .Z(n5464) );
  IV U6865 ( .A(n5464), .Z(n5465) );
  NOR U6866 ( .A(n5466), .B(n5465), .Z(n5993) );
  IV U6867 ( .A(n5467), .Z(n5468) );
  NOR U6868 ( .A(n5468), .B(n5476), .Z(n6004) );
  IV U6869 ( .A(n5469), .Z(n5471) );
  NOR U6870 ( .A(n5471), .B(n5470), .Z(n5997) );
  NOR U6871 ( .A(n6004), .B(n5997), .Z(n5688) );
  IV U6872 ( .A(n5472), .Z(n5474) );
  NOR U6873 ( .A(n5474), .B(n5473), .Z(n5479) );
  IV U6874 ( .A(n5475), .Z(n5477) );
  NOR U6875 ( .A(n5477), .B(n5476), .Z(n5478) );
  NOR U6876 ( .A(n5479), .B(n5478), .Z(n6007) );
  IV U6877 ( .A(n5480), .Z(n5481) );
  NOR U6878 ( .A(n5481), .B(n5676), .Z(n5888) );
  IV U6879 ( .A(n5482), .Z(n5484) );
  NOR U6880 ( .A(n5484), .B(n5483), .Z(n5489) );
  IV U6881 ( .A(n5485), .Z(n5486) );
  NOR U6882 ( .A(n5487), .B(n5486), .Z(n5488) );
  NOR U6883 ( .A(n5489), .B(n5488), .Z(n5899) );
  IV U6884 ( .A(n5490), .Z(n5492) );
  IV U6885 ( .A(n5491), .Z(n5496) );
  NOR U6886 ( .A(n5492), .B(n5496), .Z(n5913) );
  IV U6887 ( .A(n5493), .Z(n5494) );
  NOR U6888 ( .A(n5501), .B(n5494), .Z(n5912) );
  IV U6889 ( .A(n5495), .Z(n5497) );
  NOR U6890 ( .A(n5497), .B(n5496), .Z(n5909) );
  XOR U6891 ( .A(n5912), .B(n5909), .Z(n5498) );
  NOR U6892 ( .A(n5913), .B(n5498), .Z(n5648) );
  IV U6893 ( .A(n5499), .Z(n5500) );
  NOR U6894 ( .A(n5501), .B(n5500), .Z(n5919) );
  IV U6895 ( .A(n5502), .Z(n5505) );
  IV U6896 ( .A(n5503), .Z(n5504) );
  NOR U6897 ( .A(n5505), .B(n5504), .Z(n5916) );
  IV U6898 ( .A(n5506), .Z(n5509) );
  IV U6899 ( .A(n5507), .Z(n5508) );
  NOR U6900 ( .A(n5509), .B(n5508), .Z(n5943) );
  IV U6901 ( .A(n5510), .Z(n5514) );
  XOR U6902 ( .A(n5645), .B(n5522), .Z(n5512) );
  NOR U6903 ( .A(n5512), .B(n5511), .Z(n5513) );
  IV U6904 ( .A(n5513), .Z(n5516) );
  NOR U6905 ( .A(n5514), .B(n5516), .Z(n5935) );
  IV U6906 ( .A(n5515), .Z(n5517) );
  NOR U6907 ( .A(n5517), .B(n5516), .Z(n5955) );
  IV U6908 ( .A(n5518), .Z(n5525) );
  IV U6909 ( .A(n5519), .Z(n5520) );
  NOR U6910 ( .A(n5521), .B(n5520), .Z(n5523) );
  NOR U6911 ( .A(n5523), .B(n5522), .Z(n5524) );
  IV U6912 ( .A(n5524), .Z(n5646) );
  NOR U6913 ( .A(n5525), .B(n5646), .Z(n5938) );
  IV U6914 ( .A(n5526), .Z(n5637) );
  IV U6915 ( .A(n5527), .Z(n5528) );
  NOR U6916 ( .A(n5637), .B(n5528), .Z(n5643) );
  NOR U6917 ( .A(n5530), .B(n5529), .Z(n5531) );
  IV U6918 ( .A(n5531), .Z(n5533) );
  NOR U6919 ( .A(n5533), .B(n5532), .Z(n5928) );
  IV U6920 ( .A(n5534), .Z(n5536) );
  NOR U6921 ( .A(n5536), .B(n5535), .Z(n5635) );
  IV U6922 ( .A(n5537), .Z(n5540) );
  IV U6923 ( .A(n5538), .Z(n5539) );
  NOR U6924 ( .A(n5540), .B(n5539), .Z(n5549) );
  IV U6925 ( .A(n5541), .Z(n5543) );
  NOR U6926 ( .A(n5543), .B(n5542), .Z(n5544) );
  NOR U6927 ( .A(n5545), .B(n5544), .Z(n5547) );
  NOR U6928 ( .A(n5547), .B(n5546), .Z(n5548) );
  NOR U6929 ( .A(n5549), .B(n5548), .Z(n5550) );
  IV U6930 ( .A(n5550), .Z(n5632) );
  IV U6931 ( .A(n5551), .Z(n5552) );
  NOR U6932 ( .A(n5553), .B(n5552), .Z(n5554) );
  NOR U6933 ( .A(n5555), .B(n5554), .Z(n5556) );
  IV U6934 ( .A(n5556), .Z(n5626) );
  IV U6935 ( .A(n5557), .Z(n5558) );
  NOR U6936 ( .A(n5558), .B(n5604), .Z(n5563) );
  IV U6937 ( .A(n5559), .Z(n5560) );
  NOR U6938 ( .A(n5561), .B(n5560), .Z(n5562) );
  NOR U6939 ( .A(n5563), .B(n5562), .Z(n5564) );
  IV U6940 ( .A(n5564), .Z(n5620) );
  IV U6941 ( .A(n5565), .Z(n5568) );
  IV U6942 ( .A(n5566), .Z(n5567) );
  NOR U6943 ( .A(n5568), .B(n5567), .Z(n5610) );
  IV U6944 ( .A(n5569), .Z(n5570) );
  NOR U6945 ( .A(n5571), .B(n5570), .Z(n5578) );
  NOR U6946 ( .A(n5573), .B(n5572), .Z(n5576) );
  IV U6947 ( .A(n5574), .Z(n5575) );
  NOR U6948 ( .A(n5576), .B(n5575), .Z(n5577) );
  NOR U6949 ( .A(n5578), .B(n5577), .Z(n5579) );
  IV U6950 ( .A(n5579), .Z(n5602) );
  IV U6951 ( .A(n5580), .Z(n5581) );
  NOR U6952 ( .A(n5581), .B(n5590), .Z(n5599) );
  NOR U6953 ( .A(n5583), .B(n5582), .Z(n5585) );
  NOR U6954 ( .A(n5585), .B(n5584), .Z(n5586) );
  IV U6955 ( .A(n5586), .Z(n5596) );
  NOR U6956 ( .A(n5588), .B(n5587), .Z(n5593) );
  IV U6957 ( .A(n5589), .Z(n5591) );
  NOR U6958 ( .A(n5591), .B(n5590), .Z(n5592) );
  NOR U6959 ( .A(n5593), .B(n5592), .Z(n5594) );
  IV U6960 ( .A(n5594), .Z(n5595) );
  NOR U6961 ( .A(n5596), .B(n5595), .Z(n5597) );
  IV U6962 ( .A(n5597), .Z(n5598) );
  NOR U6963 ( .A(n5599), .B(n5598), .Z(n5600) );
  IV U6964 ( .A(n5600), .Z(n5601) );
  NOR U6965 ( .A(n5602), .B(n5601), .Z(n5603) );
  IV U6966 ( .A(n5603), .Z(n5607) );
  NOR U6967 ( .A(n5605), .B(n5604), .Z(n5606) );
  NOR U6968 ( .A(n5607), .B(n5606), .Z(n5608) );
  IV U6969 ( .A(n5608), .Z(n5609) );
  NOR U6970 ( .A(n5610), .B(n5609), .Z(n5611) );
  IV U6971 ( .A(n5611), .Z(n5617) );
  IV U6972 ( .A(n5612), .Z(n5615) );
  IV U6973 ( .A(n5613), .Z(n5614) );
  NOR U6974 ( .A(n5615), .B(n5614), .Z(n5616) );
  NOR U6975 ( .A(n5617), .B(n5616), .Z(n5618) );
  IV U6976 ( .A(n5618), .Z(n5619) );
  NOR U6977 ( .A(n5620), .B(n5619), .Z(n5621) );
  IV U6978 ( .A(n5621), .Z(n5622) );
  NOR U6979 ( .A(n5623), .B(n5622), .Z(n5624) );
  IV U6980 ( .A(n5624), .Z(n5625) );
  NOR U6981 ( .A(n5626), .B(n5625), .Z(n5627) );
  IV U6982 ( .A(n5627), .Z(n5629) );
  NOR U6983 ( .A(n5629), .B(n5628), .Z(n5630) );
  IV U6984 ( .A(n5630), .Z(n5631) );
  NOR U6985 ( .A(n5632), .B(n5631), .Z(n5633) );
  IV U6986 ( .A(n5633), .Z(n5634) );
  NOR U6987 ( .A(n5635), .B(n5634), .Z(n5930) );
  XOR U6988 ( .A(n5928), .B(n5930), .Z(n5641) );
  IV U6989 ( .A(n5636), .Z(n5638) );
  NOR U6990 ( .A(n5638), .B(n5637), .Z(n5639) );
  NOR U6991 ( .A(n5639), .B(n5927), .Z(n5640) );
  XOR U6992 ( .A(n5641), .B(n5640), .Z(n5642) );
  NOR U6993 ( .A(n5643), .B(n5642), .Z(n5925) );
  NOR U6994 ( .A(n5645), .B(n5644), .Z(n5647) );
  NOR U6995 ( .A(n5647), .B(n5646), .Z(n5924) );
  XOR U6996 ( .A(n5925), .B(n5924), .Z(n5939) );
  XOR U6997 ( .A(n5938), .B(n5939), .Z(n5956) );
  XOR U6998 ( .A(n5955), .B(n5956), .Z(n5937) );
  XOR U6999 ( .A(n5935), .B(n5937), .Z(n5947) );
  XOR U7000 ( .A(n5946), .B(n5947), .Z(n5945) );
  XOR U7001 ( .A(n5943), .B(n5945), .Z(n5917) );
  XOR U7002 ( .A(n5916), .B(n5917), .Z(n5920) );
  XOR U7003 ( .A(n5919), .B(n5920), .Z(n5915) );
  XOR U7004 ( .A(n5648), .B(n5915), .Z(n5906) );
  IV U7005 ( .A(n5649), .Z(n5650) );
  NOR U7006 ( .A(n5651), .B(n5650), .Z(n5655) );
  NOR U7007 ( .A(n5653), .B(n5652), .Z(n5654) );
  NOR U7008 ( .A(n5655), .B(n5654), .Z(n5907) );
  XOR U7009 ( .A(n5906), .B(n5907), .Z(n5896) );
  XOR U7010 ( .A(n5667), .B(n5896), .Z(n5661) );
  IV U7011 ( .A(n5656), .Z(n5659) );
  IV U7012 ( .A(n5657), .Z(n5658) );
  NOR U7013 ( .A(n5659), .B(n5658), .Z(n5669) );
  IV U7014 ( .A(n5669), .Z(n5660) );
  NOR U7015 ( .A(n5661), .B(n5660), .Z(n5898) );
  IV U7016 ( .A(n5662), .Z(n5665) );
  IV U7017 ( .A(n5663), .Z(n5664) );
  NOR U7018 ( .A(n5665), .B(n5664), .Z(n5666) );
  NOR U7019 ( .A(n5667), .B(n5666), .Z(n5895) );
  XOR U7020 ( .A(n5896), .B(n5895), .Z(n5668) );
  NOR U7021 ( .A(n5669), .B(n5668), .Z(n5670) );
  NOR U7022 ( .A(n5898), .B(n5670), .Z(n5901) );
  IV U7023 ( .A(n5671), .Z(n5672) );
  NOR U7024 ( .A(n5673), .B(n5672), .Z(n5674) );
  IV U7025 ( .A(n5674), .Z(n5903) );
  XOR U7026 ( .A(n5901), .B(n5903), .Z(n5900) );
  XOR U7027 ( .A(n5899), .B(n5900), .Z(n5885) );
  IV U7028 ( .A(n5675), .Z(n5677) );
  NOR U7029 ( .A(n5677), .B(n5676), .Z(n5683) );
  IV U7030 ( .A(n5683), .Z(n5887) );
  XOR U7031 ( .A(n5885), .B(n5887), .Z(n5681) );
  IV U7032 ( .A(n5678), .Z(n5680) );
  NOR U7033 ( .A(n5680), .B(n5679), .Z(n5889) );
  XOR U7034 ( .A(n5681), .B(n5889), .Z(n5682) );
  NOR U7035 ( .A(n5888), .B(n5682), .Z(n5687) );
  IV U7036 ( .A(n5888), .Z(n5685) );
  NOR U7037 ( .A(n5683), .B(n5885), .Z(n5894) );
  IV U7038 ( .A(n5894), .Z(n5684) );
  NOR U7039 ( .A(n5685), .B(n5684), .Z(n5686) );
  NOR U7040 ( .A(n5687), .B(n5686), .Z(n6008) );
  IV U7041 ( .A(n6008), .Z(n6002) );
  XOR U7042 ( .A(n6007), .B(n6002), .Z(n5999) );
  XOR U7043 ( .A(n5688), .B(n5999), .Z(n5994) );
  XOR U7044 ( .A(n5993), .B(n5994), .Z(n6013) );
  XOR U7045 ( .A(n6014), .B(n6013), .Z(n5697) );
  IV U7046 ( .A(n5689), .Z(n5690) );
  NOR U7047 ( .A(n5691), .B(n5690), .Z(n5696) );
  IV U7048 ( .A(n5692), .Z(n5694) );
  NOR U7049 ( .A(n5694), .B(n5693), .Z(n5695) );
  NOR U7050 ( .A(n5696), .B(n5695), .Z(n6017) );
  XOR U7051 ( .A(n5697), .B(n6017), .Z(n5991) );
  XOR U7052 ( .A(n5990), .B(n5991), .Z(n5987) );
  XOR U7053 ( .A(n5986), .B(n5987), .Z(n5983) );
  XOR U7054 ( .A(n5984), .B(n5983), .Z(n5980) );
  XOR U7055 ( .A(n5978), .B(n5980), .Z(n5977) );
  XOR U7056 ( .A(n5975), .B(n5977), .Z(n6037) );
  NOR U7057 ( .A(n6042), .B(n6037), .Z(n5703) );
  IV U7058 ( .A(n6037), .Z(n5698) );
  NOR U7059 ( .A(n6035), .B(n5698), .Z(n5701) );
  NOR U7060 ( .A(n5700), .B(n5699), .Z(n6038) );
  XOR U7061 ( .A(n5701), .B(n6038), .Z(n5702) );
  NOR U7062 ( .A(n5703), .B(n5702), .Z(n5704) );
  XOR U7063 ( .A(n6039), .B(n5704), .Z(n6053) );
  XOR U7064 ( .A(n6051), .B(n6053), .Z(n6049) );
  XOR U7065 ( .A(n5705), .B(n6049), .Z(n5713) );
  IV U7066 ( .A(n5713), .Z(n6056) );
  XOR U7067 ( .A(n5712), .B(n6056), .Z(n5706) );
  NOR U7068 ( .A(n5707), .B(n5706), .Z(n5878) );
  IV U7069 ( .A(n5708), .Z(n5709) );
  NOR U7070 ( .A(n5710), .B(n5709), .Z(n5711) );
  NOR U7071 ( .A(n5712), .B(n5711), .Z(n6055) );
  XOR U7072 ( .A(n6055), .B(n5713), .Z(n5723) );
  IV U7073 ( .A(n5723), .Z(n5714) );
  NOR U7074 ( .A(n5715), .B(n5714), .Z(n5716) );
  NOR U7075 ( .A(n5878), .B(n5716), .Z(n5866) );
  IV U7076 ( .A(n5717), .Z(n5718) );
  NOR U7077 ( .A(n5719), .B(n5718), .Z(n5729) );
  IV U7078 ( .A(n5729), .Z(n5868) );
  NOR U7079 ( .A(n5866), .B(n5868), .Z(n5731) );
  IV U7080 ( .A(n5720), .Z(n5721) );
  NOR U7081 ( .A(n5722), .B(n5721), .Z(n5725) );
  IV U7082 ( .A(n5725), .Z(n5724) );
  NOR U7083 ( .A(n5724), .B(n5723), .Z(n5883) );
  NOR U7084 ( .A(n5866), .B(n5725), .Z(n5726) );
  NOR U7085 ( .A(n5883), .B(n5726), .Z(n5727) );
  IV U7086 ( .A(n5727), .Z(n5728) );
  NOR U7087 ( .A(n5729), .B(n5728), .Z(n5730) );
  NOR U7088 ( .A(n5731), .B(n5730), .Z(n5739) );
  IV U7089 ( .A(n5739), .Z(n5732) );
  NOR U7090 ( .A(n5740), .B(n5732), .Z(n5733) );
  IV U7091 ( .A(n5733), .Z(n5734) );
  NOR U7092 ( .A(n5743), .B(n5734), .Z(n5735) );
  IV U7093 ( .A(n5735), .Z(n5736) );
  NOR U7094 ( .A(n5736), .B(n5737), .Z(n5752) );
  IV U7095 ( .A(n5737), .Z(n5741) );
  XOR U7096 ( .A(n5740), .B(n5741), .Z(n5744) );
  XOR U7097 ( .A(n5743), .B(n5744), .Z(n5738) );
  NOR U7098 ( .A(n5739), .B(n5738), .Z(n5750) );
  IV U7099 ( .A(n5740), .Z(n5742) );
  NOR U7100 ( .A(n5742), .B(n5741), .Z(n5747) );
  IV U7101 ( .A(n5743), .Z(n5745) );
  NOR U7102 ( .A(n5745), .B(n5744), .Z(n5746) );
  NOR U7103 ( .A(n5747), .B(n5746), .Z(n5748) );
  IV U7104 ( .A(n5748), .Z(n5749) );
  NOR U7105 ( .A(n5750), .B(n5749), .Z(n5751) );
  IV U7106 ( .A(n5751), .Z(n5860) );
  NOR U7107 ( .A(n5752), .B(n5860), .Z(n5840) );
  XOR U7108 ( .A(n5874), .B(n5840), .Z(n5753) );
  XOR U7109 ( .A(n5754), .B(n5753), .Z(n5845) );
  XOR U7110 ( .A(n5844), .B(n5845), .Z(n5843) );
  XOR U7111 ( .A(n5842), .B(n5843), .Z(n5853) );
  XOR U7112 ( .A(n5850), .B(n5853), .Z(n5762) );
  IV U7113 ( .A(n5755), .Z(n5756) );
  NOR U7114 ( .A(n5764), .B(n5756), .Z(n5761) );
  IV U7115 ( .A(n5757), .Z(n5759) );
  NOR U7116 ( .A(n5759), .B(n5758), .Z(n5760) );
  NOR U7117 ( .A(n5761), .B(n5760), .Z(n5854) );
  XOR U7118 ( .A(n5762), .B(n5854), .Z(n5826) );
  IV U7119 ( .A(n5763), .Z(n5765) );
  NOR U7120 ( .A(n5765), .B(n5764), .Z(n5825) );
  XOR U7121 ( .A(n5826), .B(n5825), .Z(n5829) );
  XOR U7122 ( .A(n5828), .B(n5829), .Z(n5835) );
  XOR U7123 ( .A(n5834), .B(n5835), .Z(n5770) );
  NOR U7124 ( .A(n5766), .B(n5770), .Z(n5823) );
  IV U7125 ( .A(n5767), .Z(n5769) );
  NOR U7126 ( .A(n5769), .B(n5768), .Z(n5820) );
  IV U7127 ( .A(n5770), .Z(n5771) );
  NOR U7128 ( .A(n5772), .B(n5771), .Z(n5822) );
  XOR U7129 ( .A(n5820), .B(n5822), .Z(n5773) );
  NOR U7130 ( .A(n5823), .B(n5773), .Z(n5815) );
  XOR U7131 ( .A(n5817), .B(n5815), .Z(n5814) );
  IV U7132 ( .A(n5774), .Z(n5777) );
  IV U7133 ( .A(n5775), .Z(n5776) );
  NOR U7134 ( .A(n5777), .B(n5776), .Z(n5778) );
  NOR U7135 ( .A(n5779), .B(n5778), .Z(n5813) );
  XOR U7136 ( .A(n5814), .B(n5813), .Z(n5780) );
  IV U7137 ( .A(n5780), .Z(n5807) );
  XOR U7138 ( .A(n5805), .B(n5807), .Z(n6072) );
  XOR U7139 ( .A(n5794), .B(n6072), .Z(n5789) );
  NOR U7140 ( .A(n5782), .B(n5781), .Z(n5783) );
  IV U7141 ( .A(n5783), .Z(n5784) );
  NOR U7142 ( .A(n5792), .B(n5784), .Z(n5785) );
  IV U7143 ( .A(n5785), .Z(n5797) );
  IV U7144 ( .A(n5786), .Z(n5787) );
  NOR U7145 ( .A(n5797), .B(n5787), .Z(n5799) );
  IV U7146 ( .A(n5799), .Z(n5788) );
  NOR U7147 ( .A(n5789), .B(n5788), .Z(n5812) );
  IV U7148 ( .A(n5790), .Z(n5791) );
  NOR U7149 ( .A(n5792), .B(n5791), .Z(n5793) );
  NOR U7150 ( .A(n5794), .B(n5793), .Z(n6073) );
  XOR U7151 ( .A(n6073), .B(n6072), .Z(n5801) );
  IV U7152 ( .A(n5795), .Z(n5796) );
  NOR U7153 ( .A(n5797), .B(n5796), .Z(n5802) );
  XOR U7154 ( .A(n5801), .B(n5802), .Z(n5798) );
  NOR U7155 ( .A(n5799), .B(n5798), .Z(n5800) );
  NOR U7156 ( .A(n5812), .B(n5800), .Z(o[6]) );
  IV U7157 ( .A(n5801), .Z(n5804) );
  IV U7158 ( .A(n5802), .Z(n5803) );
  NOR U7159 ( .A(n5804), .B(n5803), .Z(n5809) );
  IV U7160 ( .A(n5805), .Z(n5806) );
  NOR U7161 ( .A(n5807), .B(n5806), .Z(n5808) );
  NOR U7162 ( .A(n5809), .B(n5808), .Z(n5810) );
  IV U7163 ( .A(n5810), .Z(n5811) );
  NOR U7164 ( .A(n5812), .B(n5811), .Z(n6079) );
  NOR U7165 ( .A(n5814), .B(n5813), .Z(n5819) );
  IV U7166 ( .A(n5815), .Z(n5816) );
  NOR U7167 ( .A(n5817), .B(n5816), .Z(n5818) );
  NOR U7168 ( .A(n5819), .B(n5818), .Z(n6077) );
  IV U7169 ( .A(n5820), .Z(n5821) );
  NOR U7170 ( .A(n5822), .B(n5821), .Z(n5824) );
  NOR U7171 ( .A(n5824), .B(n5823), .Z(n6071) );
  IV U7172 ( .A(n5825), .Z(n5827) );
  NOR U7173 ( .A(n5827), .B(n5826), .Z(n5832) );
  IV U7174 ( .A(n5828), .Z(n5830) );
  NOR U7175 ( .A(n5830), .B(n5829), .Z(n5831) );
  NOR U7176 ( .A(n5832), .B(n5831), .Z(n5833) );
  IV U7177 ( .A(n5833), .Z(n5838) );
  IV U7178 ( .A(n5834), .Z(n5836) );
  NOR U7179 ( .A(n5836), .B(n5835), .Z(n5837) );
  NOR U7180 ( .A(n5838), .B(n5837), .Z(n6069) );
  IV U7181 ( .A(n5839), .Z(n5841) );
  IV U7182 ( .A(n5840), .Z(n5872) );
  NOR U7183 ( .A(n5841), .B(n5872), .Z(n5864) );
  NOR U7184 ( .A(n5843), .B(n5842), .Z(n5848) );
  IV U7185 ( .A(n5844), .Z(n5846) );
  NOR U7186 ( .A(n5846), .B(n5845), .Z(n5847) );
  NOR U7187 ( .A(n5848), .B(n5847), .Z(n5859) );
  IV U7188 ( .A(n5854), .Z(n5849) );
  NOR U7189 ( .A(n5849), .B(n5853), .Z(n5852) );
  IV U7190 ( .A(n5850), .Z(n5851) );
  NOR U7191 ( .A(n5852), .B(n5851), .Z(n5857) );
  IV U7192 ( .A(n5853), .Z(n5855) );
  NOR U7193 ( .A(n5855), .B(n5854), .Z(n5856) );
  NOR U7194 ( .A(n5857), .B(n5856), .Z(n5858) );
  XOR U7195 ( .A(n5859), .B(n5858), .Z(n5861) );
  NOR U7196 ( .A(n5861), .B(n5860), .Z(n5862) );
  IV U7197 ( .A(n5862), .Z(n5863) );
  NOR U7198 ( .A(n5864), .B(n5863), .Z(n5865) );
  IV U7199 ( .A(n5865), .Z(n5870) );
  IV U7200 ( .A(n5866), .Z(n5867) );
  NOR U7201 ( .A(n5868), .B(n5867), .Z(n5869) );
  NOR U7202 ( .A(n5870), .B(n5869), .Z(n6067) );
  IV U7203 ( .A(n5871), .Z(n5875) );
  XOR U7204 ( .A(n5874), .B(n5875), .Z(n5873) );
  NOR U7205 ( .A(n5873), .B(n5872), .Z(n5881) );
  IV U7206 ( .A(n5874), .Z(n5876) );
  NOR U7207 ( .A(n5876), .B(n5875), .Z(n5877) );
  NOR U7208 ( .A(n5878), .B(n5877), .Z(n5879) );
  IV U7209 ( .A(n5879), .Z(n5880) );
  NOR U7210 ( .A(n5881), .B(n5880), .Z(n5882) );
  IV U7211 ( .A(n5882), .Z(n5884) );
  NOR U7212 ( .A(n5884), .B(n5883), .Z(n6034) );
  IV U7213 ( .A(n5885), .Z(n5886) );
  NOR U7214 ( .A(n5887), .B(n5886), .Z(n5892) );
  NOR U7215 ( .A(n5889), .B(n5888), .Z(n5890) );
  IV U7216 ( .A(n5890), .Z(n5891) );
  NOR U7217 ( .A(n5892), .B(n5891), .Z(n5893) );
  NOR U7218 ( .A(n5894), .B(n5893), .Z(n5974) );
  NOR U7219 ( .A(n5896), .B(n5895), .Z(n5897) );
  NOR U7220 ( .A(n5898), .B(n5897), .Z(n5972) );
  NOR U7221 ( .A(n5900), .B(n5899), .Z(n5905) );
  IV U7222 ( .A(n5901), .Z(n5902) );
  NOR U7223 ( .A(n5903), .B(n5902), .Z(n5904) );
  NOR U7224 ( .A(n5905), .B(n5904), .Z(n5970) );
  IV U7225 ( .A(n5906), .Z(n5908) );
  NOR U7226 ( .A(n5908), .B(n5907), .Z(n5968) );
  IV U7227 ( .A(n5909), .Z(n5911) );
  XOR U7228 ( .A(n5915), .B(n5912), .Z(n5910) );
  NOR U7229 ( .A(n5911), .B(n5910), .Z(n5965) );
  NOR U7230 ( .A(n5913), .B(n5912), .Z(n5914) );
  NOR U7231 ( .A(n5915), .B(n5914), .Z(n5962) );
  IV U7232 ( .A(n5916), .Z(n5918) );
  NOR U7233 ( .A(n5918), .B(n5917), .Z(n5923) );
  IV U7234 ( .A(n5919), .Z(n5921) );
  NOR U7235 ( .A(n5921), .B(n5920), .Z(n5922) );
  NOR U7236 ( .A(n5923), .B(n5922), .Z(n5934) );
  IV U7237 ( .A(n5924), .Z(n5926) );
  NOR U7238 ( .A(n5926), .B(n5925), .Z(n5932) );
  NOR U7239 ( .A(n5928), .B(n5927), .Z(n5929) );
  NOR U7240 ( .A(n5930), .B(n5929), .Z(n5931) );
  NOR U7241 ( .A(n5932), .B(n5931), .Z(n5933) );
  XOR U7242 ( .A(n5934), .B(n5933), .Z(n5954) );
  IV U7243 ( .A(n5935), .Z(n5936) );
  NOR U7244 ( .A(n5937), .B(n5936), .Z(n5942) );
  IV U7245 ( .A(n5938), .Z(n5940) );
  NOR U7246 ( .A(n5940), .B(n5939), .Z(n5941) );
  NOR U7247 ( .A(n5942), .B(n5941), .Z(n5952) );
  IV U7248 ( .A(n5943), .Z(n5944) );
  NOR U7249 ( .A(n5945), .B(n5944), .Z(n5950) );
  IV U7250 ( .A(n5946), .Z(n5948) );
  NOR U7251 ( .A(n5948), .B(n5947), .Z(n5949) );
  NOR U7252 ( .A(n5950), .B(n5949), .Z(n5951) );
  XOR U7253 ( .A(n5952), .B(n5951), .Z(n5953) );
  XOR U7254 ( .A(n5954), .B(n5953), .Z(n5959) );
  IV U7255 ( .A(n5955), .Z(n5957) );
  NOR U7256 ( .A(n5957), .B(n5956), .Z(n5958) );
  NOR U7257 ( .A(n5959), .B(n5958), .Z(n5960) );
  IV U7258 ( .A(n5960), .Z(n5961) );
  NOR U7259 ( .A(n5962), .B(n5961), .Z(n5963) );
  IV U7260 ( .A(n5963), .Z(n5964) );
  NOR U7261 ( .A(n5965), .B(n5964), .Z(n5966) );
  IV U7262 ( .A(n5966), .Z(n5967) );
  NOR U7263 ( .A(n5968), .B(n5967), .Z(n5969) );
  XOR U7264 ( .A(n5970), .B(n5969), .Z(n5971) );
  XOR U7265 ( .A(n5972), .B(n5971), .Z(n5973) );
  XOR U7266 ( .A(n5974), .B(n5973), .Z(n6032) );
  IV U7267 ( .A(n5975), .Z(n5976) );
  NOR U7268 ( .A(n5977), .B(n5976), .Z(n5982) );
  IV U7269 ( .A(n5978), .Z(n5979) );
  NOR U7270 ( .A(n5980), .B(n5979), .Z(n5981) );
  NOR U7271 ( .A(n5982), .B(n5981), .Z(n6030) );
  IV U7272 ( .A(n5983), .Z(n5985) );
  NOR U7273 ( .A(n5985), .B(n5984), .Z(n5989) );
  NOR U7274 ( .A(n5987), .B(n5986), .Z(n5988) );
  NOR U7275 ( .A(n5989), .B(n5988), .Z(n6028) );
  IV U7276 ( .A(n5990), .Z(n5992) );
  NOR U7277 ( .A(n5992), .B(n5991), .Z(n6026) );
  IV U7278 ( .A(n5993), .Z(n5996) );
  IV U7279 ( .A(n5994), .Z(n5995) );
  NOR U7280 ( .A(n5996), .B(n5995), .Z(n6001) );
  IV U7281 ( .A(n5997), .Z(n5998) );
  NOR U7282 ( .A(n5999), .B(n5998), .Z(n6000) );
  NOR U7283 ( .A(n6001), .B(n6000), .Z(n6012) );
  IV U7284 ( .A(n6007), .Z(n6003) );
  NOR U7285 ( .A(n6003), .B(n6002), .Z(n6006) );
  IV U7286 ( .A(n6004), .Z(n6005) );
  NOR U7287 ( .A(n6006), .B(n6005), .Z(n6010) );
  NOR U7288 ( .A(n6008), .B(n6007), .Z(n6009) );
  NOR U7289 ( .A(n6010), .B(n6009), .Z(n6011) );
  XOR U7290 ( .A(n6012), .B(n6011), .Z(n6023) );
  NOR U7291 ( .A(n6013), .B(n6014), .Z(n6021) );
  IV U7292 ( .A(n6013), .Z(n6016) );
  IV U7293 ( .A(n6014), .Z(n6015) );
  NOR U7294 ( .A(n6016), .B(n6015), .Z(n6019) );
  IV U7295 ( .A(n6017), .Z(n6018) );
  NOR U7296 ( .A(n6019), .B(n6018), .Z(n6020) );
  NOR U7297 ( .A(n6021), .B(n6020), .Z(n6022) );
  NOR U7298 ( .A(n6023), .B(n6022), .Z(n6024) );
  IV U7299 ( .A(n6024), .Z(n6025) );
  NOR U7300 ( .A(n6026), .B(n6025), .Z(n6027) );
  XOR U7301 ( .A(n6028), .B(n6027), .Z(n6029) );
  XOR U7302 ( .A(n6030), .B(n6029), .Z(n6031) );
  XOR U7303 ( .A(n6032), .B(n6031), .Z(n6033) );
  XOR U7304 ( .A(n6034), .B(n6033), .Z(n6065) );
  XOR U7305 ( .A(n6038), .B(n6039), .Z(n6041) );
  XOR U7306 ( .A(n6035), .B(n6041), .Z(n6036) );
  NOR U7307 ( .A(n6037), .B(n6036), .Z(n6047) );
  IV U7308 ( .A(n6038), .Z(n6040) );
  NOR U7309 ( .A(n6040), .B(n6039), .Z(n6044) );
  NOR U7310 ( .A(n6042), .B(n6041), .Z(n6043) );
  NOR U7311 ( .A(n6044), .B(n6043), .Z(n6045) );
  IV U7312 ( .A(n6045), .Z(n6046) );
  NOR U7313 ( .A(n6047), .B(n6046), .Z(n6063) );
  IV U7314 ( .A(n6048), .Z(n6050) );
  NOR U7315 ( .A(n6050), .B(n6049), .Z(n6061) );
  NOR U7316 ( .A(n6052), .B(n6051), .Z(n6054) );
  NOR U7317 ( .A(n6054), .B(n6053), .Z(n6058) );
  NOR U7318 ( .A(n6056), .B(n6055), .Z(n6057) );
  NOR U7319 ( .A(n6058), .B(n6057), .Z(n6059) );
  IV U7320 ( .A(n6059), .Z(n6060) );
  NOR U7321 ( .A(n6061), .B(n6060), .Z(n6062) );
  XOR U7322 ( .A(n6063), .B(n6062), .Z(n6064) );
  XOR U7323 ( .A(n6065), .B(n6064), .Z(n6066) );
  XOR U7324 ( .A(n6067), .B(n6066), .Z(n6068) );
  XOR U7325 ( .A(n6069), .B(n6068), .Z(n6070) );
  XOR U7326 ( .A(n6071), .B(n6070), .Z(n6075) );
  NOR U7327 ( .A(n6073), .B(n6072), .Z(n6074) );
  XOR U7328 ( .A(n6075), .B(n6074), .Z(n6076) );
  XOR U7329 ( .A(n6077), .B(n6076), .Z(n6078) );
  XOR U7330 ( .A(n6079), .B(n6078), .Z(o[7]) );
endmodule

