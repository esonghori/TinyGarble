
module sum_N1024_CC1 ( clk, rst, a, b, c );
  input [1023:0] a;
  input [1023:0] b;
  output [1023:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090;

  XNOR U2 ( .A(a[2]), .B(n4086), .Z(n778) );
  XNOR U3 ( .A(a[5]), .B(n4077), .Z(n445) );
  XNOR U4 ( .A(a[8]), .B(n4068), .Z(n112) );
  XNOR U5 ( .A(a[11]), .B(n4059), .Z(n978) );
  XNOR U6 ( .A(a[14]), .B(n4050), .Z(n945) );
  XNOR U7 ( .A(a[17]), .B(n4041), .Z(n912) );
  XNOR U8 ( .A(a[20]), .B(n4032), .Z(n878) );
  XNOR U9 ( .A(a[23]), .B(n4023), .Z(n845) );
  XNOR U10 ( .A(a[26]), .B(n4014), .Z(n812) );
  XNOR U11 ( .A(a[29]), .B(n4005), .Z(n779) );
  XNOR U12 ( .A(a[32]), .B(n3996), .Z(n745) );
  XNOR U13 ( .A(a[35]), .B(n3987), .Z(n712) );
  XNOR U14 ( .A(a[38]), .B(n3978), .Z(n679) );
  XNOR U15 ( .A(a[41]), .B(n3969), .Z(n645) );
  XNOR U16 ( .A(a[44]), .B(n3960), .Z(n612) );
  XNOR U17 ( .A(a[47]), .B(n3951), .Z(n579) );
  XNOR U18 ( .A(a[50]), .B(n3942), .Z(n545) );
  XNOR U19 ( .A(a[53]), .B(n3933), .Z(n512) );
  XNOR U20 ( .A(a[56]), .B(n3924), .Z(n479) );
  XNOR U21 ( .A(a[59]), .B(n3915), .Z(n446) );
  XNOR U22 ( .A(a[62]), .B(n3906), .Z(n412) );
  XNOR U23 ( .A(a[65]), .B(n3897), .Z(n379) );
  XNOR U24 ( .A(a[68]), .B(n3888), .Z(n346) );
  XNOR U25 ( .A(a[71]), .B(n3879), .Z(n312) );
  XNOR U26 ( .A(a[74]), .B(n3870), .Z(n279) );
  XNOR U27 ( .A(a[77]), .B(n3861), .Z(n246) );
  XNOR U28 ( .A(a[80]), .B(n3852), .Z(n212) );
  XNOR U29 ( .A(a[83]), .B(n3843), .Z(n179) );
  XNOR U30 ( .A(a[86]), .B(n3834), .Z(n146) );
  XNOR U31 ( .A(a[89]), .B(n3825), .Z(n113) );
  XNOR U32 ( .A(a[92]), .B(n3816), .Z(n79) );
  XNOR U33 ( .A(a[95]), .B(n3807), .Z(n46) );
  XNOR U34 ( .A(a[98]), .B(n3798), .Z(n13) );
  XNOR U35 ( .A(a[101]), .B(n3789), .Z(n1016) );
  XNOR U36 ( .A(a[104]), .B(n3780), .Z(n995) );
  XNOR U37 ( .A(a[107]), .B(n3771), .Z(n992) );
  XNOR U38 ( .A(a[110]), .B(n3762), .Z(n988) );
  XNOR U39 ( .A(a[113]), .B(n3753), .Z(n985) );
  XNOR U40 ( .A(a[116]), .B(n3744), .Z(n982) );
  XNOR U41 ( .A(a[119]), .B(n3735), .Z(n979) );
  XNOR U42 ( .A(a[122]), .B(n3726), .Z(n975) );
  XNOR U43 ( .A(a[125]), .B(n3717), .Z(n972) );
  XNOR U44 ( .A(a[128]), .B(n3708), .Z(n969) );
  XNOR U45 ( .A(a[131]), .B(n3699), .Z(n965) );
  XNOR U46 ( .A(a[134]), .B(n3690), .Z(n962) );
  XNOR U47 ( .A(a[137]), .B(n3681), .Z(n959) );
  XNOR U48 ( .A(a[140]), .B(n3672), .Z(n955) );
  XNOR U49 ( .A(a[143]), .B(n3663), .Z(n952) );
  XNOR U50 ( .A(a[146]), .B(n3654), .Z(n949) );
  XNOR U51 ( .A(a[149]), .B(n3645), .Z(n946) );
  XNOR U52 ( .A(a[152]), .B(n3636), .Z(n942) );
  XNOR U53 ( .A(a[155]), .B(n3627), .Z(n939) );
  XNOR U54 ( .A(a[158]), .B(n3618), .Z(n936) );
  XNOR U55 ( .A(a[161]), .B(n3609), .Z(n932) );
  XNOR U56 ( .A(a[164]), .B(n3600), .Z(n929) );
  XNOR U57 ( .A(a[167]), .B(n3591), .Z(n926) );
  XNOR U58 ( .A(a[170]), .B(n3582), .Z(n922) );
  XNOR U59 ( .A(a[173]), .B(n3573), .Z(n919) );
  XNOR U60 ( .A(a[176]), .B(n3564), .Z(n916) );
  XNOR U61 ( .A(a[179]), .B(n3555), .Z(n913) );
  XNOR U62 ( .A(a[182]), .B(n3546), .Z(n909) );
  XNOR U63 ( .A(a[185]), .B(n3537), .Z(n906) );
  XNOR U64 ( .A(a[188]), .B(n3528), .Z(n903) );
  XNOR U65 ( .A(a[191]), .B(n3519), .Z(n899) );
  XNOR U66 ( .A(a[194]), .B(n3510), .Z(n896) );
  XNOR U67 ( .A(a[197]), .B(n3501), .Z(n893) );
  XNOR U68 ( .A(a[200]), .B(n3492), .Z(n888) );
  XNOR U69 ( .A(a[203]), .B(n3483), .Z(n885) );
  XNOR U70 ( .A(a[206]), .B(n3474), .Z(n882) );
  XNOR U71 ( .A(a[209]), .B(n3465), .Z(n879) );
  XNOR U72 ( .A(a[212]), .B(n3456), .Z(n875) );
  XNOR U73 ( .A(a[215]), .B(n3447), .Z(n872) );
  XNOR U74 ( .A(a[218]), .B(n3438), .Z(n869) );
  XNOR U75 ( .A(a[221]), .B(n3429), .Z(n865) );
  XNOR U76 ( .A(a[224]), .B(n3420), .Z(n862) );
  XNOR U77 ( .A(a[227]), .B(n3411), .Z(n859) );
  XNOR U78 ( .A(a[230]), .B(n3402), .Z(n855) );
  XNOR U79 ( .A(a[233]), .B(n3393), .Z(n852) );
  XNOR U80 ( .A(a[236]), .B(n3384), .Z(n849) );
  XNOR U81 ( .A(a[239]), .B(n3375), .Z(n846) );
  XNOR U82 ( .A(a[242]), .B(n3366), .Z(n842) );
  XNOR U83 ( .A(a[245]), .B(n3357), .Z(n839) );
  XNOR U84 ( .A(a[248]), .B(n3348), .Z(n836) );
  XNOR U85 ( .A(a[251]), .B(n3339), .Z(n832) );
  XNOR U86 ( .A(a[254]), .B(n3330), .Z(n829) );
  XNOR U87 ( .A(a[257]), .B(n3321), .Z(n826) );
  XNOR U88 ( .A(a[260]), .B(n3312), .Z(n822) );
  XNOR U89 ( .A(a[263]), .B(n3303), .Z(n819) );
  XNOR U90 ( .A(a[266]), .B(n3294), .Z(n816) );
  XNOR U91 ( .A(a[269]), .B(n3285), .Z(n813) );
  XNOR U92 ( .A(a[272]), .B(n3276), .Z(n809) );
  XNOR U93 ( .A(a[275]), .B(n3267), .Z(n806) );
  XNOR U94 ( .A(a[278]), .B(n3258), .Z(n803) );
  XNOR U95 ( .A(a[281]), .B(n3249), .Z(n799) );
  XNOR U96 ( .A(a[284]), .B(n3240), .Z(n796) );
  XNOR U97 ( .A(a[287]), .B(n3231), .Z(n793) );
  XNOR U98 ( .A(a[290]), .B(n3222), .Z(n789) );
  XNOR U99 ( .A(a[293]), .B(n3213), .Z(n786) );
  XNOR U100 ( .A(a[296]), .B(n3204), .Z(n783) );
  XNOR U101 ( .A(a[299]), .B(n3195), .Z(n780) );
  XNOR U102 ( .A(a[302]), .B(n3186), .Z(n775) );
  XNOR U103 ( .A(a[305]), .B(n3177), .Z(n772) );
  XNOR U104 ( .A(a[308]), .B(n3168), .Z(n769) );
  XNOR U105 ( .A(a[311]), .B(n3159), .Z(n765) );
  XNOR U106 ( .A(a[314]), .B(n3150), .Z(n762) );
  XNOR U107 ( .A(a[317]), .B(n3141), .Z(n759) );
  XNOR U108 ( .A(a[320]), .B(n3132), .Z(n755) );
  XNOR U109 ( .A(a[323]), .B(n3123), .Z(n752) );
  XNOR U110 ( .A(a[326]), .B(n3114), .Z(n749) );
  XNOR U111 ( .A(a[329]), .B(n3105), .Z(n746) );
  XNOR U112 ( .A(a[332]), .B(n3096), .Z(n742) );
  XNOR U113 ( .A(a[335]), .B(n3087), .Z(n739) );
  XNOR U114 ( .A(a[338]), .B(n3078), .Z(n736) );
  XNOR U115 ( .A(a[341]), .B(n3069), .Z(n732) );
  XNOR U116 ( .A(a[344]), .B(n3060), .Z(n729) );
  XNOR U117 ( .A(a[347]), .B(n3051), .Z(n726) );
  XNOR U118 ( .A(a[350]), .B(n3042), .Z(n722) );
  XNOR U119 ( .A(a[353]), .B(n3033), .Z(n719) );
  XNOR U120 ( .A(a[356]), .B(n3024), .Z(n716) );
  XNOR U121 ( .A(a[359]), .B(n3015), .Z(n713) );
  XNOR U122 ( .A(a[362]), .B(n3006), .Z(n709) );
  XNOR U123 ( .A(a[365]), .B(n2997), .Z(n706) );
  XNOR U124 ( .A(a[368]), .B(n2988), .Z(n703) );
  XNOR U125 ( .A(a[371]), .B(n2979), .Z(n699) );
  XNOR U126 ( .A(a[374]), .B(n2970), .Z(n696) );
  XNOR U127 ( .A(a[377]), .B(n2961), .Z(n693) );
  XNOR U128 ( .A(a[380]), .B(n2952), .Z(n689) );
  XNOR U129 ( .A(a[383]), .B(n2943), .Z(n686) );
  XNOR U130 ( .A(a[386]), .B(n2934), .Z(n683) );
  XNOR U131 ( .A(a[389]), .B(n2925), .Z(n680) );
  XNOR U132 ( .A(a[392]), .B(n2916), .Z(n676) );
  XNOR U133 ( .A(a[395]), .B(n2907), .Z(n673) );
  XNOR U134 ( .A(a[398]), .B(n2898), .Z(n670) );
  XNOR U135 ( .A(a[401]), .B(n2889), .Z(n665) );
  XNOR U136 ( .A(a[404]), .B(n2880), .Z(n662) );
  XNOR U137 ( .A(a[407]), .B(n2871), .Z(n659) );
  XNOR U138 ( .A(a[410]), .B(n2862), .Z(n655) );
  XNOR U139 ( .A(a[413]), .B(n2853), .Z(n652) );
  XNOR U140 ( .A(a[416]), .B(n2844), .Z(n649) );
  XNOR U141 ( .A(a[419]), .B(n2835), .Z(n646) );
  XNOR U142 ( .A(a[422]), .B(n2826), .Z(n642) );
  XNOR U143 ( .A(a[425]), .B(n2817), .Z(n639) );
  XNOR U144 ( .A(a[428]), .B(n2808), .Z(n636) );
  XNOR U145 ( .A(a[431]), .B(n2799), .Z(n632) );
  XNOR U146 ( .A(a[434]), .B(n2790), .Z(n629) );
  XNOR U147 ( .A(a[437]), .B(n2781), .Z(n626) );
  XNOR U148 ( .A(a[440]), .B(n2772), .Z(n622) );
  XNOR U149 ( .A(a[443]), .B(n2763), .Z(n619) );
  XNOR U150 ( .A(a[446]), .B(n2754), .Z(n616) );
  XNOR U151 ( .A(a[449]), .B(n2745), .Z(n613) );
  XNOR U152 ( .A(a[452]), .B(n2736), .Z(n609) );
  XNOR U153 ( .A(a[455]), .B(n2727), .Z(n606) );
  XNOR U154 ( .A(a[458]), .B(n2718), .Z(n603) );
  XNOR U155 ( .A(a[461]), .B(n2709), .Z(n599) );
  XNOR U156 ( .A(a[464]), .B(n2700), .Z(n596) );
  XNOR U157 ( .A(a[467]), .B(n2691), .Z(n593) );
  XNOR U158 ( .A(a[470]), .B(n2682), .Z(n589) );
  XNOR U159 ( .A(a[473]), .B(n2673), .Z(n586) );
  XNOR U160 ( .A(a[476]), .B(n2664), .Z(n583) );
  XNOR U161 ( .A(a[479]), .B(n2655), .Z(n580) );
  XNOR U162 ( .A(a[482]), .B(n2646), .Z(n576) );
  XNOR U163 ( .A(a[485]), .B(n2637), .Z(n573) );
  XNOR U164 ( .A(a[488]), .B(n2628), .Z(n570) );
  XNOR U165 ( .A(a[491]), .B(n2619), .Z(n566) );
  XNOR U166 ( .A(a[494]), .B(n2610), .Z(n563) );
  XNOR U167 ( .A(a[497]), .B(n2601), .Z(n560) );
  XNOR U168 ( .A(a[500]), .B(n2592), .Z(n555) );
  XNOR U169 ( .A(a[503]), .B(n2583), .Z(n552) );
  XNOR U170 ( .A(a[506]), .B(n2574), .Z(n549) );
  XNOR U171 ( .A(a[509]), .B(n2565), .Z(n546) );
  XNOR U172 ( .A(a[512]), .B(n2556), .Z(n542) );
  XNOR U173 ( .A(a[515]), .B(n2547), .Z(n539) );
  XNOR U174 ( .A(a[518]), .B(n2538), .Z(n536) );
  XNOR U175 ( .A(a[521]), .B(n2529), .Z(n532) );
  XNOR U176 ( .A(a[524]), .B(n2520), .Z(n529) );
  XNOR U177 ( .A(a[527]), .B(n2511), .Z(n526) );
  XNOR U178 ( .A(a[530]), .B(n2502), .Z(n522) );
  XNOR U179 ( .A(a[533]), .B(n2493), .Z(n519) );
  XNOR U180 ( .A(a[536]), .B(n2484), .Z(n516) );
  XNOR U181 ( .A(a[539]), .B(n2475), .Z(n513) );
  XNOR U182 ( .A(a[542]), .B(n2466), .Z(n509) );
  XNOR U183 ( .A(a[545]), .B(n2457), .Z(n506) );
  XNOR U184 ( .A(a[548]), .B(n2448), .Z(n503) );
  XNOR U185 ( .A(a[551]), .B(n2439), .Z(n499) );
  XNOR U186 ( .A(a[554]), .B(n2430), .Z(n496) );
  XNOR U187 ( .A(a[557]), .B(n2421), .Z(n493) );
  XNOR U188 ( .A(a[560]), .B(n2412), .Z(n489) );
  XNOR U189 ( .A(a[563]), .B(n2403), .Z(n486) );
  XNOR U190 ( .A(a[566]), .B(n2394), .Z(n483) );
  XNOR U191 ( .A(a[569]), .B(n2385), .Z(n480) );
  XNOR U192 ( .A(a[572]), .B(n2376), .Z(n476) );
  XNOR U193 ( .A(a[575]), .B(n2367), .Z(n473) );
  XNOR U194 ( .A(a[578]), .B(n2358), .Z(n470) );
  XNOR U195 ( .A(a[581]), .B(n2349), .Z(n466) );
  XNOR U196 ( .A(a[584]), .B(n2340), .Z(n463) );
  XNOR U197 ( .A(a[587]), .B(n2331), .Z(n460) );
  XNOR U198 ( .A(a[590]), .B(n2322), .Z(n456) );
  XNOR U199 ( .A(a[593]), .B(n2313), .Z(n453) );
  XNOR U200 ( .A(a[596]), .B(n2304), .Z(n450) );
  XNOR U201 ( .A(a[599]), .B(n2295), .Z(n447) );
  XNOR U202 ( .A(a[602]), .B(n2286), .Z(n442) );
  XNOR U203 ( .A(a[605]), .B(n2277), .Z(n439) );
  XNOR U204 ( .A(a[608]), .B(n2268), .Z(n436) );
  XNOR U205 ( .A(a[611]), .B(n2259), .Z(n432) );
  XNOR U206 ( .A(a[614]), .B(n2250), .Z(n429) );
  XNOR U207 ( .A(a[617]), .B(n2241), .Z(n426) );
  XNOR U208 ( .A(a[620]), .B(n2232), .Z(n422) );
  XNOR U209 ( .A(a[623]), .B(n2223), .Z(n419) );
  XNOR U210 ( .A(a[626]), .B(n2214), .Z(n416) );
  XNOR U211 ( .A(a[629]), .B(n2205), .Z(n413) );
  XNOR U212 ( .A(a[632]), .B(n2196), .Z(n409) );
  XNOR U213 ( .A(a[635]), .B(n2187), .Z(n406) );
  XNOR U214 ( .A(a[638]), .B(n2178), .Z(n403) );
  XNOR U215 ( .A(a[641]), .B(n2169), .Z(n399) );
  XNOR U216 ( .A(a[644]), .B(n2160), .Z(n396) );
  XNOR U217 ( .A(a[647]), .B(n2151), .Z(n393) );
  XNOR U218 ( .A(a[650]), .B(n2142), .Z(n389) );
  XNOR U219 ( .A(a[653]), .B(n2133), .Z(n386) );
  XNOR U220 ( .A(a[656]), .B(n2124), .Z(n383) );
  XNOR U221 ( .A(a[659]), .B(n2115), .Z(n380) );
  XNOR U222 ( .A(a[662]), .B(n2106), .Z(n376) );
  XNOR U223 ( .A(a[665]), .B(n2097), .Z(n373) );
  XNOR U224 ( .A(a[668]), .B(n2088), .Z(n370) );
  XNOR U225 ( .A(a[671]), .B(n2079), .Z(n366) );
  XNOR U226 ( .A(a[674]), .B(n2070), .Z(n363) );
  XNOR U227 ( .A(a[677]), .B(n2061), .Z(n360) );
  XNOR U228 ( .A(a[680]), .B(n2052), .Z(n356) );
  XNOR U229 ( .A(a[683]), .B(n2043), .Z(n353) );
  XNOR U230 ( .A(a[686]), .B(n2034), .Z(n350) );
  XNOR U231 ( .A(a[689]), .B(n2025), .Z(n347) );
  XNOR U232 ( .A(a[692]), .B(n2016), .Z(n343) );
  XNOR U233 ( .A(a[695]), .B(n2007), .Z(n340) );
  XNOR U234 ( .A(a[698]), .B(n1998), .Z(n337) );
  XNOR U235 ( .A(a[701]), .B(n1989), .Z(n332) );
  XNOR U236 ( .A(a[704]), .B(n1980), .Z(n329) );
  XNOR U237 ( .A(a[707]), .B(n1971), .Z(n326) );
  XNOR U238 ( .A(a[710]), .B(n1962), .Z(n322) );
  XNOR U239 ( .A(a[713]), .B(n1953), .Z(n319) );
  XNOR U240 ( .A(a[716]), .B(n1944), .Z(n316) );
  XNOR U241 ( .A(a[719]), .B(n1935), .Z(n313) );
  XNOR U242 ( .A(a[722]), .B(n1926), .Z(n309) );
  XNOR U243 ( .A(a[725]), .B(n1917), .Z(n306) );
  XNOR U244 ( .A(a[728]), .B(n1908), .Z(n303) );
  XNOR U245 ( .A(a[731]), .B(n1899), .Z(n299) );
  XNOR U246 ( .A(a[734]), .B(n1890), .Z(n296) );
  XNOR U247 ( .A(a[737]), .B(n1881), .Z(n293) );
  XNOR U248 ( .A(a[740]), .B(n1872), .Z(n289) );
  XNOR U249 ( .A(a[743]), .B(n1863), .Z(n286) );
  XNOR U250 ( .A(a[746]), .B(n1854), .Z(n283) );
  XNOR U251 ( .A(a[749]), .B(n1845), .Z(n280) );
  XNOR U252 ( .A(a[752]), .B(n1836), .Z(n276) );
  XNOR U253 ( .A(a[755]), .B(n1827), .Z(n273) );
  XNOR U254 ( .A(a[758]), .B(n1818), .Z(n270) );
  XNOR U255 ( .A(a[761]), .B(n1809), .Z(n266) );
  XNOR U256 ( .A(a[764]), .B(n1800), .Z(n263) );
  XNOR U257 ( .A(a[767]), .B(n1791), .Z(n260) );
  XNOR U258 ( .A(a[770]), .B(n1782), .Z(n256) );
  XNOR U259 ( .A(a[773]), .B(n1773), .Z(n253) );
  XNOR U260 ( .A(a[776]), .B(n1764), .Z(n250) );
  XNOR U261 ( .A(a[779]), .B(n1755), .Z(n247) );
  XNOR U262 ( .A(a[782]), .B(n1746), .Z(n243) );
  XNOR U263 ( .A(a[785]), .B(n1737), .Z(n240) );
  XNOR U264 ( .A(a[788]), .B(n1728), .Z(n237) );
  XNOR U265 ( .A(a[791]), .B(n1719), .Z(n233) );
  XNOR U266 ( .A(a[794]), .B(n1710), .Z(n230) );
  XNOR U267 ( .A(a[797]), .B(n1701), .Z(n227) );
  XNOR U268 ( .A(a[800]), .B(n1692), .Z(n222) );
  XNOR U269 ( .A(a[803]), .B(n1683), .Z(n219) );
  XNOR U270 ( .A(a[806]), .B(n1674), .Z(n216) );
  XNOR U271 ( .A(a[809]), .B(n1665), .Z(n213) );
  XNOR U272 ( .A(a[812]), .B(n1656), .Z(n209) );
  XNOR U273 ( .A(a[815]), .B(n1647), .Z(n206) );
  XNOR U274 ( .A(a[818]), .B(n1638), .Z(n203) );
  XNOR U275 ( .A(a[821]), .B(n1629), .Z(n199) );
  XNOR U276 ( .A(a[824]), .B(n1620), .Z(n196) );
  XNOR U277 ( .A(a[827]), .B(n1611), .Z(n193) );
  XNOR U278 ( .A(a[830]), .B(n1602), .Z(n189) );
  XNOR U279 ( .A(a[833]), .B(n1593), .Z(n186) );
  XNOR U280 ( .A(a[836]), .B(n1584), .Z(n183) );
  XNOR U281 ( .A(a[839]), .B(n1575), .Z(n180) );
  XNOR U282 ( .A(a[842]), .B(n1566), .Z(n176) );
  XNOR U283 ( .A(a[845]), .B(n1557), .Z(n173) );
  XNOR U284 ( .A(a[848]), .B(n1548), .Z(n170) );
  XNOR U285 ( .A(a[851]), .B(n1539), .Z(n166) );
  XNOR U286 ( .A(a[854]), .B(n1530), .Z(n163) );
  XNOR U287 ( .A(a[857]), .B(n1521), .Z(n160) );
  XNOR U288 ( .A(a[860]), .B(n1512), .Z(n156) );
  XNOR U289 ( .A(a[863]), .B(n1503), .Z(n153) );
  XNOR U290 ( .A(a[866]), .B(n1494), .Z(n150) );
  XNOR U291 ( .A(a[869]), .B(n1485), .Z(n147) );
  XNOR U292 ( .A(a[872]), .B(n1476), .Z(n143) );
  XNOR U293 ( .A(a[875]), .B(n1467), .Z(n140) );
  XNOR U294 ( .A(a[878]), .B(n1458), .Z(n137) );
  XNOR U295 ( .A(a[881]), .B(n1449), .Z(n133) );
  XNOR U296 ( .A(a[884]), .B(n1440), .Z(n130) );
  XNOR U297 ( .A(a[887]), .B(n1431), .Z(n127) );
  XNOR U298 ( .A(a[890]), .B(n1422), .Z(n123) );
  XNOR U299 ( .A(a[893]), .B(n1413), .Z(n120) );
  XNOR U300 ( .A(a[896]), .B(n1404), .Z(n117) );
  XNOR U301 ( .A(a[899]), .B(n1395), .Z(n114) );
  XNOR U302 ( .A(a[902]), .B(n1386), .Z(n109) );
  XNOR U303 ( .A(a[905]), .B(n1377), .Z(n106) );
  XNOR U304 ( .A(a[908]), .B(n1368), .Z(n103) );
  XNOR U305 ( .A(a[911]), .B(n1359), .Z(n99) );
  XNOR U306 ( .A(a[914]), .B(n1350), .Z(n96) );
  XNOR U307 ( .A(a[917]), .B(n1341), .Z(n93) );
  XNOR U308 ( .A(a[920]), .B(n1332), .Z(n89) );
  XNOR U309 ( .A(a[923]), .B(n1323), .Z(n86) );
  XNOR U310 ( .A(a[926]), .B(n1314), .Z(n83) );
  XNOR U311 ( .A(a[929]), .B(n1305), .Z(n80) );
  XNOR U312 ( .A(a[932]), .B(n1296), .Z(n76) );
  XNOR U313 ( .A(a[935]), .B(n1287), .Z(n73) );
  XNOR U314 ( .A(a[938]), .B(n1278), .Z(n70) );
  XNOR U315 ( .A(a[941]), .B(n1269), .Z(n66) );
  XNOR U316 ( .A(a[944]), .B(n1260), .Z(n63) );
  XNOR U317 ( .A(a[947]), .B(n1251), .Z(n60) );
  XNOR U318 ( .A(a[950]), .B(n1242), .Z(n56) );
  XNOR U319 ( .A(a[953]), .B(n1233), .Z(n53) );
  XNOR U320 ( .A(a[956]), .B(n1224), .Z(n50) );
  XNOR U321 ( .A(a[959]), .B(n1215), .Z(n47) );
  XNOR U322 ( .A(a[962]), .B(n1206), .Z(n43) );
  XNOR U323 ( .A(a[965]), .B(n1197), .Z(n40) );
  XNOR U324 ( .A(a[968]), .B(n1188), .Z(n37) );
  XNOR U325 ( .A(a[971]), .B(n1179), .Z(n33) );
  XNOR U326 ( .A(a[974]), .B(n1170), .Z(n30) );
  XNOR U327 ( .A(a[977]), .B(n1161), .Z(n27) );
  XNOR U328 ( .A(a[980]), .B(n1152), .Z(n23) );
  XNOR U329 ( .A(a[983]), .B(n1143), .Z(n20) );
  XNOR U330 ( .A(a[986]), .B(n1134), .Z(n17) );
  XNOR U331 ( .A(a[989]), .B(n1125), .Z(n14) );
  XNOR U332 ( .A(a[992]), .B(n1116), .Z(n10) );
  XNOR U333 ( .A(a[995]), .B(n1107), .Z(n7) );
  XNOR U334 ( .A(a[998]), .B(n1098), .Z(n4) );
  XNOR U335 ( .A(a[1001]), .B(n1087), .Z(n1089) );
  XNOR U336 ( .A(a[1004]), .B(n1075), .Z(n1077) );
  XNOR U337 ( .A(a[1007]), .B(n1063), .Z(n1065) );
  XNOR U338 ( .A(a[1010]), .B(n1050), .Z(n1052) );
  XNOR U339 ( .A(a[1013]), .B(n1038), .Z(n1040) );
  XNOR U340 ( .A(a[1016]), .B(n1026), .Z(n1028) );
  XNOR U341 ( .A(a[1019]), .B(n1013), .Z(n1015) );
  XNOR U342 ( .A(a[3]), .B(n4083), .Z(n667) );
  XNOR U343 ( .A(a[6]), .B(n4074), .Z(n334) );
  XNOR U344 ( .A(a[9]), .B(n4065), .Z(n1) );
  XNOR U345 ( .A(a[12]), .B(n4056), .Z(n967) );
  XNOR U346 ( .A(a[15]), .B(n4047), .Z(n934) );
  XNOR U347 ( .A(a[18]), .B(n4038), .Z(n901) );
  XNOR U348 ( .A(a[21]), .B(n4029), .Z(n867) );
  XNOR U349 ( .A(a[24]), .B(n4020), .Z(n834) );
  XNOR U350 ( .A(a[27]), .B(n4011), .Z(n801) );
  XNOR U351 ( .A(a[30]), .B(n4002), .Z(n767) );
  XNOR U352 ( .A(a[33]), .B(n3993), .Z(n734) );
  XNOR U353 ( .A(a[36]), .B(n3984), .Z(n701) );
  XNOR U354 ( .A(a[39]), .B(n3975), .Z(n668) );
  XNOR U355 ( .A(a[42]), .B(n3966), .Z(n634) );
  XNOR U356 ( .A(a[45]), .B(n3957), .Z(n601) );
  XNOR U357 ( .A(a[48]), .B(n3948), .Z(n568) );
  XNOR U358 ( .A(a[51]), .B(n3939), .Z(n534) );
  XNOR U359 ( .A(a[54]), .B(n3930), .Z(n501) );
  XNOR U360 ( .A(a[57]), .B(n3921), .Z(n468) );
  XNOR U361 ( .A(a[60]), .B(n3912), .Z(n434) );
  XNOR U362 ( .A(a[63]), .B(n3903), .Z(n401) );
  XNOR U363 ( .A(a[66]), .B(n3894), .Z(n368) );
  XNOR U364 ( .A(a[69]), .B(n3885), .Z(n335) );
  XNOR U365 ( .A(a[72]), .B(n3876), .Z(n301) );
  XNOR U366 ( .A(a[75]), .B(n3867), .Z(n268) );
  XNOR U367 ( .A(a[78]), .B(n3858), .Z(n235) );
  XNOR U368 ( .A(a[81]), .B(n3849), .Z(n201) );
  XNOR U369 ( .A(a[84]), .B(n3840), .Z(n168) );
  XNOR U370 ( .A(a[87]), .B(n3831), .Z(n135) );
  XNOR U371 ( .A(a[90]), .B(n3822), .Z(n101) );
  XNOR U372 ( .A(a[93]), .B(n3813), .Z(n68) );
  XNOR U373 ( .A(a[96]), .B(n3804), .Z(n35) );
  XNOR U374 ( .A(a[99]), .B(n3795), .Z(n2) );
  XNOR U375 ( .A(a[102]), .B(n3786), .Z(n997) );
  XNOR U376 ( .A(a[105]), .B(n3777), .Z(n994) );
  XNOR U377 ( .A(a[108]), .B(n3768), .Z(n991) );
  XNOR U378 ( .A(a[111]), .B(n3759), .Z(n987) );
  XNOR U379 ( .A(a[114]), .B(n3750), .Z(n984) );
  XNOR U380 ( .A(a[117]), .B(n3741), .Z(n981) );
  XNOR U381 ( .A(a[120]), .B(n3732), .Z(n977) );
  XNOR U382 ( .A(a[123]), .B(n3723), .Z(n974) );
  XNOR U383 ( .A(a[126]), .B(n3714), .Z(n971) );
  XNOR U384 ( .A(a[129]), .B(n3705), .Z(n968) );
  XNOR U385 ( .A(a[132]), .B(n3696), .Z(n964) );
  XNOR U386 ( .A(a[135]), .B(n3687), .Z(n961) );
  XNOR U387 ( .A(a[138]), .B(n3678), .Z(n958) );
  XNOR U388 ( .A(a[141]), .B(n3669), .Z(n954) );
  XNOR U389 ( .A(a[144]), .B(n3660), .Z(n951) );
  XNOR U390 ( .A(a[147]), .B(n3651), .Z(n948) );
  XNOR U391 ( .A(a[150]), .B(n3642), .Z(n944) );
  XNOR U392 ( .A(a[153]), .B(n3633), .Z(n941) );
  XNOR U393 ( .A(a[156]), .B(n3624), .Z(n938) );
  XNOR U394 ( .A(a[159]), .B(n3615), .Z(n935) );
  XNOR U395 ( .A(a[162]), .B(n3606), .Z(n931) );
  XNOR U396 ( .A(a[165]), .B(n3597), .Z(n928) );
  XNOR U397 ( .A(a[168]), .B(n3588), .Z(n925) );
  XNOR U398 ( .A(a[171]), .B(n3579), .Z(n921) );
  XNOR U399 ( .A(a[174]), .B(n3570), .Z(n918) );
  XNOR U400 ( .A(a[177]), .B(n3561), .Z(n915) );
  XNOR U401 ( .A(a[180]), .B(n3552), .Z(n911) );
  XNOR U402 ( .A(a[183]), .B(n3543), .Z(n908) );
  XNOR U403 ( .A(a[186]), .B(n3534), .Z(n905) );
  XNOR U404 ( .A(a[189]), .B(n3525), .Z(n902) );
  XNOR U405 ( .A(a[192]), .B(n3516), .Z(n898) );
  XNOR U406 ( .A(a[195]), .B(n3507), .Z(n895) );
  XNOR U407 ( .A(a[198]), .B(n3498), .Z(n892) );
  XNOR U408 ( .A(a[201]), .B(n3489), .Z(n887) );
  XNOR U409 ( .A(a[204]), .B(n3480), .Z(n884) );
  XNOR U410 ( .A(a[207]), .B(n3471), .Z(n881) );
  XNOR U411 ( .A(a[210]), .B(n3462), .Z(n877) );
  XNOR U412 ( .A(a[213]), .B(n3453), .Z(n874) );
  XNOR U413 ( .A(a[216]), .B(n3444), .Z(n871) );
  XNOR U414 ( .A(a[219]), .B(n3435), .Z(n868) );
  XNOR U415 ( .A(a[222]), .B(n3426), .Z(n864) );
  XNOR U416 ( .A(a[225]), .B(n3417), .Z(n861) );
  XNOR U417 ( .A(a[228]), .B(n3408), .Z(n858) );
  XNOR U418 ( .A(a[231]), .B(n3399), .Z(n854) );
  XNOR U419 ( .A(a[234]), .B(n3390), .Z(n851) );
  XNOR U420 ( .A(a[237]), .B(n3381), .Z(n848) );
  XNOR U421 ( .A(a[240]), .B(n3372), .Z(n844) );
  XNOR U422 ( .A(a[243]), .B(n3363), .Z(n841) );
  XNOR U423 ( .A(a[246]), .B(n3354), .Z(n838) );
  XNOR U424 ( .A(a[249]), .B(n3345), .Z(n835) );
  XNOR U425 ( .A(a[252]), .B(n3336), .Z(n831) );
  XNOR U426 ( .A(a[255]), .B(n3327), .Z(n828) );
  XNOR U427 ( .A(a[258]), .B(n3318), .Z(n825) );
  XNOR U428 ( .A(a[261]), .B(n3309), .Z(n821) );
  XNOR U429 ( .A(a[264]), .B(n3300), .Z(n818) );
  XNOR U430 ( .A(a[267]), .B(n3291), .Z(n815) );
  XNOR U431 ( .A(a[270]), .B(n3282), .Z(n811) );
  XNOR U432 ( .A(a[273]), .B(n3273), .Z(n808) );
  XNOR U433 ( .A(a[276]), .B(n3264), .Z(n805) );
  XNOR U434 ( .A(a[279]), .B(n3255), .Z(n802) );
  XNOR U435 ( .A(a[282]), .B(n3246), .Z(n798) );
  XNOR U436 ( .A(a[285]), .B(n3237), .Z(n795) );
  XNOR U437 ( .A(a[288]), .B(n3228), .Z(n792) );
  XNOR U438 ( .A(a[291]), .B(n3219), .Z(n788) );
  XNOR U439 ( .A(a[294]), .B(n3210), .Z(n785) );
  XNOR U440 ( .A(a[297]), .B(n3201), .Z(n782) );
  XNOR U441 ( .A(a[300]), .B(n3192), .Z(n777) );
  XNOR U442 ( .A(a[303]), .B(n3183), .Z(n774) );
  XNOR U443 ( .A(a[306]), .B(n3174), .Z(n771) );
  XNOR U444 ( .A(a[309]), .B(n3165), .Z(n768) );
  XNOR U445 ( .A(a[312]), .B(n3156), .Z(n764) );
  XNOR U446 ( .A(a[315]), .B(n3147), .Z(n761) );
  XNOR U447 ( .A(a[318]), .B(n3138), .Z(n758) );
  XNOR U448 ( .A(a[321]), .B(n3129), .Z(n754) );
  XNOR U449 ( .A(a[324]), .B(n3120), .Z(n751) );
  XNOR U450 ( .A(a[327]), .B(n3111), .Z(n748) );
  XNOR U451 ( .A(a[330]), .B(n3102), .Z(n744) );
  XNOR U452 ( .A(a[333]), .B(n3093), .Z(n741) );
  XNOR U453 ( .A(a[336]), .B(n3084), .Z(n738) );
  XNOR U454 ( .A(a[339]), .B(n3075), .Z(n735) );
  XNOR U455 ( .A(a[342]), .B(n3066), .Z(n731) );
  XNOR U456 ( .A(a[345]), .B(n3057), .Z(n728) );
  XNOR U457 ( .A(a[348]), .B(n3048), .Z(n725) );
  XNOR U458 ( .A(a[351]), .B(n3039), .Z(n721) );
  XNOR U459 ( .A(a[354]), .B(n3030), .Z(n718) );
  XNOR U460 ( .A(a[357]), .B(n3021), .Z(n715) );
  XNOR U461 ( .A(a[360]), .B(n3012), .Z(n711) );
  XNOR U462 ( .A(a[363]), .B(n3003), .Z(n708) );
  XNOR U463 ( .A(a[366]), .B(n2994), .Z(n705) );
  XNOR U464 ( .A(a[369]), .B(n2985), .Z(n702) );
  XNOR U465 ( .A(a[372]), .B(n2976), .Z(n698) );
  XNOR U466 ( .A(a[375]), .B(n2967), .Z(n695) );
  XNOR U467 ( .A(a[378]), .B(n2958), .Z(n692) );
  XNOR U468 ( .A(a[381]), .B(n2949), .Z(n688) );
  XNOR U469 ( .A(a[384]), .B(n2940), .Z(n685) );
  XNOR U470 ( .A(a[387]), .B(n2931), .Z(n682) );
  XNOR U471 ( .A(a[390]), .B(n2922), .Z(n678) );
  XNOR U472 ( .A(a[393]), .B(n2913), .Z(n675) );
  XNOR U473 ( .A(a[396]), .B(n2904), .Z(n672) );
  XNOR U474 ( .A(a[399]), .B(n2895), .Z(n669) );
  XNOR U475 ( .A(a[402]), .B(n2886), .Z(n664) );
  XNOR U476 ( .A(a[405]), .B(n2877), .Z(n661) );
  XNOR U477 ( .A(a[408]), .B(n2868), .Z(n658) );
  XNOR U478 ( .A(a[411]), .B(n2859), .Z(n654) );
  XNOR U479 ( .A(a[414]), .B(n2850), .Z(n651) );
  XNOR U480 ( .A(a[417]), .B(n2841), .Z(n648) );
  XNOR U481 ( .A(a[420]), .B(n2832), .Z(n644) );
  XNOR U482 ( .A(a[423]), .B(n2823), .Z(n641) );
  XNOR U483 ( .A(a[426]), .B(n2814), .Z(n638) );
  XNOR U484 ( .A(a[429]), .B(n2805), .Z(n635) );
  XNOR U485 ( .A(a[432]), .B(n2796), .Z(n631) );
  XNOR U486 ( .A(a[435]), .B(n2787), .Z(n628) );
  XNOR U487 ( .A(a[438]), .B(n2778), .Z(n625) );
  XNOR U488 ( .A(a[441]), .B(n2769), .Z(n621) );
  XNOR U489 ( .A(a[444]), .B(n2760), .Z(n618) );
  XNOR U490 ( .A(a[447]), .B(n2751), .Z(n615) );
  XNOR U491 ( .A(a[450]), .B(n2742), .Z(n611) );
  XNOR U492 ( .A(a[453]), .B(n2733), .Z(n608) );
  XNOR U493 ( .A(a[456]), .B(n2724), .Z(n605) );
  XNOR U494 ( .A(a[459]), .B(n2715), .Z(n602) );
  XNOR U495 ( .A(a[462]), .B(n2706), .Z(n598) );
  XNOR U496 ( .A(a[465]), .B(n2697), .Z(n595) );
  XNOR U497 ( .A(a[468]), .B(n2688), .Z(n592) );
  XNOR U498 ( .A(a[471]), .B(n2679), .Z(n588) );
  XNOR U499 ( .A(a[474]), .B(n2670), .Z(n585) );
  XNOR U500 ( .A(a[477]), .B(n2661), .Z(n582) );
  XNOR U501 ( .A(a[480]), .B(n2652), .Z(n578) );
  XNOR U502 ( .A(a[483]), .B(n2643), .Z(n575) );
  XNOR U503 ( .A(a[486]), .B(n2634), .Z(n572) );
  XNOR U504 ( .A(a[489]), .B(n2625), .Z(n569) );
  XNOR U505 ( .A(a[492]), .B(n2616), .Z(n565) );
  XNOR U506 ( .A(a[495]), .B(n2607), .Z(n562) );
  XNOR U507 ( .A(a[498]), .B(n2598), .Z(n559) );
  XNOR U508 ( .A(a[501]), .B(n2589), .Z(n554) );
  XNOR U509 ( .A(a[504]), .B(n2580), .Z(n551) );
  XNOR U510 ( .A(a[507]), .B(n2571), .Z(n548) );
  XNOR U511 ( .A(a[510]), .B(n2562), .Z(n544) );
  XNOR U512 ( .A(a[513]), .B(n2553), .Z(n541) );
  XNOR U513 ( .A(a[516]), .B(n2544), .Z(n538) );
  XNOR U514 ( .A(a[519]), .B(n2535), .Z(n535) );
  XNOR U515 ( .A(a[522]), .B(n2526), .Z(n531) );
  XNOR U516 ( .A(a[525]), .B(n2517), .Z(n528) );
  XNOR U517 ( .A(a[528]), .B(n2508), .Z(n525) );
  XNOR U518 ( .A(a[531]), .B(n2499), .Z(n521) );
  XNOR U519 ( .A(a[534]), .B(n2490), .Z(n518) );
  XNOR U520 ( .A(a[537]), .B(n2481), .Z(n515) );
  XNOR U521 ( .A(a[540]), .B(n2472), .Z(n511) );
  XNOR U522 ( .A(a[543]), .B(n2463), .Z(n508) );
  XNOR U523 ( .A(a[546]), .B(n2454), .Z(n505) );
  XNOR U524 ( .A(a[549]), .B(n2445), .Z(n502) );
  XNOR U525 ( .A(a[552]), .B(n2436), .Z(n498) );
  XNOR U526 ( .A(a[555]), .B(n2427), .Z(n495) );
  XNOR U527 ( .A(a[558]), .B(n2418), .Z(n492) );
  XNOR U528 ( .A(a[561]), .B(n2409), .Z(n488) );
  XNOR U529 ( .A(a[564]), .B(n2400), .Z(n485) );
  XNOR U530 ( .A(a[567]), .B(n2391), .Z(n482) );
  XNOR U531 ( .A(a[570]), .B(n2382), .Z(n478) );
  XNOR U532 ( .A(a[573]), .B(n2373), .Z(n475) );
  XNOR U533 ( .A(a[576]), .B(n2364), .Z(n472) );
  XNOR U534 ( .A(a[579]), .B(n2355), .Z(n469) );
  XNOR U535 ( .A(a[582]), .B(n2346), .Z(n465) );
  XNOR U536 ( .A(a[585]), .B(n2337), .Z(n462) );
  XNOR U537 ( .A(a[588]), .B(n2328), .Z(n459) );
  XNOR U538 ( .A(a[591]), .B(n2319), .Z(n455) );
  XNOR U539 ( .A(a[594]), .B(n2310), .Z(n452) );
  XNOR U540 ( .A(a[597]), .B(n2301), .Z(n449) );
  XNOR U541 ( .A(a[600]), .B(n2292), .Z(n444) );
  XNOR U542 ( .A(a[603]), .B(n2283), .Z(n441) );
  XNOR U543 ( .A(a[606]), .B(n2274), .Z(n438) );
  XNOR U544 ( .A(a[609]), .B(n2265), .Z(n435) );
  XNOR U545 ( .A(a[612]), .B(n2256), .Z(n431) );
  XNOR U546 ( .A(a[615]), .B(n2247), .Z(n428) );
  XNOR U547 ( .A(a[618]), .B(n2238), .Z(n425) );
  XNOR U548 ( .A(a[621]), .B(n2229), .Z(n421) );
  XNOR U549 ( .A(a[624]), .B(n2220), .Z(n418) );
  XNOR U550 ( .A(a[627]), .B(n2211), .Z(n415) );
  XNOR U551 ( .A(a[630]), .B(n2202), .Z(n411) );
  XNOR U552 ( .A(a[633]), .B(n2193), .Z(n408) );
  XNOR U553 ( .A(a[636]), .B(n2184), .Z(n405) );
  XNOR U554 ( .A(a[639]), .B(n2175), .Z(n402) );
  XNOR U555 ( .A(a[642]), .B(n2166), .Z(n398) );
  XNOR U556 ( .A(a[645]), .B(n2157), .Z(n395) );
  XNOR U557 ( .A(a[648]), .B(n2148), .Z(n392) );
  XNOR U558 ( .A(a[651]), .B(n2139), .Z(n388) );
  XNOR U559 ( .A(a[654]), .B(n2130), .Z(n385) );
  XNOR U560 ( .A(a[657]), .B(n2121), .Z(n382) );
  XNOR U561 ( .A(a[660]), .B(n2112), .Z(n378) );
  XNOR U562 ( .A(a[663]), .B(n2103), .Z(n375) );
  XNOR U563 ( .A(a[666]), .B(n2094), .Z(n372) );
  XNOR U564 ( .A(a[669]), .B(n2085), .Z(n369) );
  XNOR U565 ( .A(a[672]), .B(n2076), .Z(n365) );
  XNOR U566 ( .A(a[675]), .B(n2067), .Z(n362) );
  XNOR U567 ( .A(a[678]), .B(n2058), .Z(n359) );
  XNOR U568 ( .A(a[681]), .B(n2049), .Z(n355) );
  XNOR U569 ( .A(a[684]), .B(n2040), .Z(n352) );
  XNOR U570 ( .A(a[687]), .B(n2031), .Z(n349) );
  XNOR U571 ( .A(a[690]), .B(n2022), .Z(n345) );
  XNOR U572 ( .A(a[693]), .B(n2013), .Z(n342) );
  XNOR U573 ( .A(a[696]), .B(n2004), .Z(n339) );
  XNOR U574 ( .A(a[699]), .B(n1995), .Z(n336) );
  XNOR U575 ( .A(a[702]), .B(n1986), .Z(n331) );
  XNOR U576 ( .A(a[705]), .B(n1977), .Z(n328) );
  XNOR U577 ( .A(a[708]), .B(n1968), .Z(n325) );
  XNOR U578 ( .A(a[711]), .B(n1959), .Z(n321) );
  XNOR U579 ( .A(a[714]), .B(n1950), .Z(n318) );
  XNOR U580 ( .A(a[717]), .B(n1941), .Z(n315) );
  XNOR U581 ( .A(a[720]), .B(n1932), .Z(n311) );
  XNOR U582 ( .A(a[723]), .B(n1923), .Z(n308) );
  XNOR U583 ( .A(a[726]), .B(n1914), .Z(n305) );
  XNOR U584 ( .A(a[729]), .B(n1905), .Z(n302) );
  XNOR U585 ( .A(a[732]), .B(n1896), .Z(n298) );
  XNOR U586 ( .A(a[735]), .B(n1887), .Z(n295) );
  XNOR U587 ( .A(a[738]), .B(n1878), .Z(n292) );
  XNOR U588 ( .A(a[741]), .B(n1869), .Z(n288) );
  XNOR U589 ( .A(a[744]), .B(n1860), .Z(n285) );
  XNOR U590 ( .A(a[747]), .B(n1851), .Z(n282) );
  XNOR U591 ( .A(a[750]), .B(n1842), .Z(n278) );
  XNOR U592 ( .A(a[753]), .B(n1833), .Z(n275) );
  XNOR U593 ( .A(a[756]), .B(n1824), .Z(n272) );
  XNOR U594 ( .A(a[759]), .B(n1815), .Z(n269) );
  XNOR U595 ( .A(a[762]), .B(n1806), .Z(n265) );
  XNOR U596 ( .A(a[765]), .B(n1797), .Z(n262) );
  XNOR U597 ( .A(a[768]), .B(n1788), .Z(n259) );
  XNOR U598 ( .A(a[771]), .B(n1779), .Z(n255) );
  XNOR U599 ( .A(a[774]), .B(n1770), .Z(n252) );
  XNOR U600 ( .A(a[777]), .B(n1761), .Z(n249) );
  XNOR U601 ( .A(a[780]), .B(n1752), .Z(n245) );
  XNOR U602 ( .A(a[783]), .B(n1743), .Z(n242) );
  XNOR U603 ( .A(a[786]), .B(n1734), .Z(n239) );
  XNOR U604 ( .A(a[789]), .B(n1725), .Z(n236) );
  XNOR U605 ( .A(a[792]), .B(n1716), .Z(n232) );
  XNOR U606 ( .A(a[795]), .B(n1707), .Z(n229) );
  XNOR U607 ( .A(a[798]), .B(n1698), .Z(n226) );
  XNOR U608 ( .A(a[801]), .B(n1689), .Z(n221) );
  XNOR U609 ( .A(a[804]), .B(n1680), .Z(n218) );
  XNOR U610 ( .A(a[807]), .B(n1671), .Z(n215) );
  XNOR U611 ( .A(a[810]), .B(n1662), .Z(n211) );
  XNOR U612 ( .A(a[813]), .B(n1653), .Z(n208) );
  XNOR U613 ( .A(a[816]), .B(n1644), .Z(n205) );
  XNOR U614 ( .A(a[819]), .B(n1635), .Z(n202) );
  XNOR U615 ( .A(a[822]), .B(n1626), .Z(n198) );
  XNOR U616 ( .A(a[825]), .B(n1617), .Z(n195) );
  XNOR U617 ( .A(a[828]), .B(n1608), .Z(n192) );
  XNOR U618 ( .A(a[831]), .B(n1599), .Z(n188) );
  XNOR U619 ( .A(a[834]), .B(n1590), .Z(n185) );
  XNOR U620 ( .A(a[837]), .B(n1581), .Z(n182) );
  XNOR U621 ( .A(a[840]), .B(n1572), .Z(n178) );
  XNOR U622 ( .A(a[843]), .B(n1563), .Z(n175) );
  XNOR U623 ( .A(a[846]), .B(n1554), .Z(n172) );
  XNOR U624 ( .A(a[849]), .B(n1545), .Z(n169) );
  XNOR U625 ( .A(a[852]), .B(n1536), .Z(n165) );
  XNOR U626 ( .A(a[855]), .B(n1527), .Z(n162) );
  XNOR U627 ( .A(a[858]), .B(n1518), .Z(n159) );
  XNOR U628 ( .A(a[861]), .B(n1509), .Z(n155) );
  XNOR U629 ( .A(a[864]), .B(n1500), .Z(n152) );
  XNOR U630 ( .A(a[867]), .B(n1491), .Z(n149) );
  XNOR U631 ( .A(a[870]), .B(n1482), .Z(n145) );
  XNOR U632 ( .A(a[873]), .B(n1473), .Z(n142) );
  XNOR U633 ( .A(a[876]), .B(n1464), .Z(n139) );
  XNOR U634 ( .A(a[879]), .B(n1455), .Z(n136) );
  XNOR U635 ( .A(a[882]), .B(n1446), .Z(n132) );
  XNOR U636 ( .A(a[885]), .B(n1437), .Z(n129) );
  XNOR U637 ( .A(a[888]), .B(n1428), .Z(n126) );
  XNOR U638 ( .A(a[891]), .B(n1419), .Z(n122) );
  XNOR U639 ( .A(a[894]), .B(n1410), .Z(n119) );
  XNOR U640 ( .A(a[897]), .B(n1401), .Z(n116) );
  XNOR U641 ( .A(a[900]), .B(n1392), .Z(n111) );
  XNOR U642 ( .A(a[903]), .B(n1383), .Z(n108) );
  XNOR U643 ( .A(a[906]), .B(n1374), .Z(n105) );
  XNOR U644 ( .A(a[909]), .B(n1365), .Z(n102) );
  XNOR U645 ( .A(a[912]), .B(n1356), .Z(n98) );
  XNOR U646 ( .A(a[915]), .B(n1347), .Z(n95) );
  XNOR U647 ( .A(a[918]), .B(n1338), .Z(n92) );
  XNOR U648 ( .A(a[921]), .B(n1329), .Z(n88) );
  XNOR U649 ( .A(a[924]), .B(n1320), .Z(n85) );
  XNOR U650 ( .A(a[927]), .B(n1311), .Z(n82) );
  XNOR U651 ( .A(a[930]), .B(n1302), .Z(n78) );
  XNOR U652 ( .A(a[933]), .B(n1293), .Z(n75) );
  XNOR U653 ( .A(a[936]), .B(n1284), .Z(n72) );
  XNOR U654 ( .A(a[939]), .B(n1275), .Z(n69) );
  XNOR U655 ( .A(a[942]), .B(n1266), .Z(n65) );
  XNOR U656 ( .A(a[945]), .B(n1257), .Z(n62) );
  XNOR U657 ( .A(a[948]), .B(n1248), .Z(n59) );
  XNOR U658 ( .A(a[951]), .B(n1239), .Z(n55) );
  XNOR U659 ( .A(a[954]), .B(n1230), .Z(n52) );
  XNOR U660 ( .A(a[957]), .B(n1221), .Z(n49) );
  XNOR U661 ( .A(a[960]), .B(n1212), .Z(n45) );
  XNOR U662 ( .A(a[963]), .B(n1203), .Z(n42) );
  XNOR U663 ( .A(a[966]), .B(n1194), .Z(n39) );
  XNOR U664 ( .A(a[969]), .B(n1185), .Z(n36) );
  XNOR U665 ( .A(a[972]), .B(n1176), .Z(n32) );
  XNOR U666 ( .A(a[975]), .B(n1167), .Z(n29) );
  XNOR U667 ( .A(a[978]), .B(n1158), .Z(n26) );
  XNOR U668 ( .A(a[981]), .B(n1149), .Z(n22) );
  XNOR U669 ( .A(a[984]), .B(n1140), .Z(n19) );
  XNOR U670 ( .A(a[987]), .B(n1131), .Z(n16) );
  XNOR U671 ( .A(a[990]), .B(n1122), .Z(n12) );
  XNOR U672 ( .A(a[993]), .B(n1113), .Z(n9) );
  XNOR U673 ( .A(a[996]), .B(n1104), .Z(n6) );
  XNOR U674 ( .A(a[999]), .B(n1095), .Z(n3) );
  XNOR U675 ( .A(a[1002]), .B(n1083), .Z(n1085) );
  XNOR U676 ( .A(a[1005]), .B(n1071), .Z(n1073) );
  XNOR U677 ( .A(a[1008]), .B(n1059), .Z(n1061) );
  XNOR U678 ( .A(a[1011]), .B(n1046), .Z(n1048) );
  XNOR U679 ( .A(a[1014]), .B(n1034), .Z(n1036) );
  XNOR U680 ( .A(a[1017]), .B(n1022), .Z(n1024) );
  XNOR U681 ( .A(a[1020]), .B(n1009), .Z(n1011) );
  XNOR U682 ( .A(a[4]), .B(n4080), .Z(n556) );
  XNOR U683 ( .A(a[7]), .B(n4071), .Z(n223) );
  XNOR U684 ( .A(a[10]), .B(n4062), .Z(n989) );
  XNOR U685 ( .A(a[13]), .B(n4053), .Z(n956) );
  XNOR U686 ( .A(a[16]), .B(n4044), .Z(n923) );
  XNOR U687 ( .A(a[19]), .B(n4035), .Z(n890) );
  XNOR U688 ( .A(a[22]), .B(n4026), .Z(n856) );
  XNOR U689 ( .A(a[25]), .B(n4017), .Z(n823) );
  XNOR U690 ( .A(a[28]), .B(n4008), .Z(n790) );
  XNOR U691 ( .A(a[31]), .B(n3999), .Z(n756) );
  XNOR U692 ( .A(a[34]), .B(n3990), .Z(n723) );
  XNOR U693 ( .A(a[37]), .B(n3981), .Z(n690) );
  XNOR U694 ( .A(a[40]), .B(n3972), .Z(n656) );
  XNOR U695 ( .A(a[43]), .B(n3963), .Z(n623) );
  XNOR U696 ( .A(a[46]), .B(n3954), .Z(n590) );
  XNOR U697 ( .A(a[49]), .B(n3945), .Z(n557) );
  XNOR U698 ( .A(a[52]), .B(n3936), .Z(n523) );
  XNOR U699 ( .A(a[55]), .B(n3927), .Z(n490) );
  XNOR U700 ( .A(a[58]), .B(n3918), .Z(n457) );
  XNOR U701 ( .A(a[61]), .B(n3909), .Z(n423) );
  XNOR U702 ( .A(a[64]), .B(n3900), .Z(n390) );
  XNOR U703 ( .A(a[67]), .B(n3891), .Z(n357) );
  XNOR U704 ( .A(a[70]), .B(n3882), .Z(n323) );
  XNOR U705 ( .A(a[73]), .B(n3873), .Z(n290) );
  XNOR U706 ( .A(a[76]), .B(n3864), .Z(n257) );
  XNOR U707 ( .A(a[79]), .B(n3855), .Z(n224) );
  XNOR U708 ( .A(a[82]), .B(n3846), .Z(n190) );
  XNOR U709 ( .A(a[85]), .B(n3837), .Z(n157) );
  XNOR U710 ( .A(a[88]), .B(n3828), .Z(n124) );
  XNOR U711 ( .A(a[91]), .B(n3819), .Z(n90) );
  XNOR U712 ( .A(a[94]), .B(n3810), .Z(n57) );
  XNOR U713 ( .A(a[97]), .B(n3801), .Z(n24) );
  XNOR U714 ( .A(a[100]), .B(n3792), .Z(n1057) );
  XNOR U715 ( .A(a[103]), .B(n3783), .Z(n996) );
  XNOR U716 ( .A(a[106]), .B(n3774), .Z(n993) );
  XNOR U717 ( .A(a[109]), .B(n3765), .Z(n990) );
  XNOR U718 ( .A(a[112]), .B(n3756), .Z(n986) );
  XNOR U719 ( .A(a[115]), .B(n3747), .Z(n983) );
  XNOR U720 ( .A(a[118]), .B(n3738), .Z(n980) );
  XNOR U721 ( .A(a[121]), .B(n3729), .Z(n976) );
  XNOR U722 ( .A(a[124]), .B(n3720), .Z(n973) );
  XNOR U723 ( .A(a[127]), .B(n3711), .Z(n970) );
  XNOR U724 ( .A(a[130]), .B(n3702), .Z(n966) );
  XNOR U725 ( .A(a[133]), .B(n3693), .Z(n963) );
  XNOR U726 ( .A(a[136]), .B(n3684), .Z(n960) );
  XNOR U727 ( .A(a[139]), .B(n3675), .Z(n957) );
  XNOR U728 ( .A(a[142]), .B(n3666), .Z(n953) );
  XNOR U729 ( .A(a[145]), .B(n3657), .Z(n950) );
  XNOR U730 ( .A(a[148]), .B(n3648), .Z(n947) );
  XNOR U731 ( .A(a[151]), .B(n3639), .Z(n943) );
  XNOR U732 ( .A(a[154]), .B(n3630), .Z(n940) );
  XNOR U733 ( .A(a[157]), .B(n3621), .Z(n937) );
  XNOR U734 ( .A(a[160]), .B(n3612), .Z(n933) );
  XNOR U735 ( .A(a[163]), .B(n3603), .Z(n930) );
  XNOR U736 ( .A(a[166]), .B(n3594), .Z(n927) );
  XNOR U737 ( .A(a[169]), .B(n3585), .Z(n924) );
  XNOR U738 ( .A(a[172]), .B(n3576), .Z(n920) );
  XNOR U739 ( .A(a[175]), .B(n3567), .Z(n917) );
  XNOR U740 ( .A(a[178]), .B(n3558), .Z(n914) );
  XNOR U741 ( .A(a[181]), .B(n3549), .Z(n910) );
  XNOR U742 ( .A(a[184]), .B(n3540), .Z(n907) );
  XNOR U743 ( .A(a[187]), .B(n3531), .Z(n904) );
  XNOR U744 ( .A(a[190]), .B(n3522), .Z(n900) );
  XNOR U745 ( .A(a[193]), .B(n3513), .Z(n897) );
  XNOR U746 ( .A(a[196]), .B(n3504), .Z(n894) );
  XNOR U747 ( .A(a[199]), .B(n3495), .Z(n891) );
  XNOR U748 ( .A(a[202]), .B(n3486), .Z(n886) );
  XNOR U749 ( .A(a[205]), .B(n3477), .Z(n883) );
  XNOR U750 ( .A(a[208]), .B(n3468), .Z(n880) );
  XNOR U751 ( .A(a[211]), .B(n3459), .Z(n876) );
  XNOR U752 ( .A(a[214]), .B(n3450), .Z(n873) );
  XNOR U753 ( .A(a[217]), .B(n3441), .Z(n870) );
  XNOR U754 ( .A(a[220]), .B(n3432), .Z(n866) );
  XNOR U755 ( .A(a[223]), .B(n3423), .Z(n863) );
  XNOR U756 ( .A(a[226]), .B(n3414), .Z(n860) );
  XNOR U757 ( .A(a[229]), .B(n3405), .Z(n857) );
  XNOR U758 ( .A(a[232]), .B(n3396), .Z(n853) );
  XNOR U759 ( .A(a[235]), .B(n3387), .Z(n850) );
  XNOR U760 ( .A(a[238]), .B(n3378), .Z(n847) );
  XNOR U761 ( .A(a[241]), .B(n3369), .Z(n843) );
  XNOR U762 ( .A(a[244]), .B(n3360), .Z(n840) );
  XNOR U763 ( .A(a[247]), .B(n3351), .Z(n837) );
  XNOR U764 ( .A(a[250]), .B(n3342), .Z(n833) );
  XNOR U765 ( .A(a[253]), .B(n3333), .Z(n830) );
  XNOR U766 ( .A(a[256]), .B(n3324), .Z(n827) );
  XNOR U767 ( .A(a[259]), .B(n3315), .Z(n824) );
  XNOR U768 ( .A(a[262]), .B(n3306), .Z(n820) );
  XNOR U769 ( .A(a[265]), .B(n3297), .Z(n817) );
  XNOR U770 ( .A(a[268]), .B(n3288), .Z(n814) );
  XNOR U771 ( .A(a[271]), .B(n3279), .Z(n810) );
  XNOR U772 ( .A(a[274]), .B(n3270), .Z(n807) );
  XNOR U773 ( .A(a[277]), .B(n3261), .Z(n804) );
  XNOR U774 ( .A(a[280]), .B(n3252), .Z(n800) );
  XNOR U775 ( .A(a[283]), .B(n3243), .Z(n797) );
  XNOR U776 ( .A(a[286]), .B(n3234), .Z(n794) );
  XNOR U777 ( .A(a[289]), .B(n3225), .Z(n791) );
  XNOR U778 ( .A(a[292]), .B(n3216), .Z(n787) );
  XNOR U779 ( .A(a[295]), .B(n3207), .Z(n784) );
  XNOR U780 ( .A(a[298]), .B(n3198), .Z(n781) );
  XNOR U781 ( .A(a[301]), .B(n3189), .Z(n776) );
  XNOR U782 ( .A(a[304]), .B(n3180), .Z(n773) );
  XNOR U783 ( .A(a[307]), .B(n3171), .Z(n770) );
  XNOR U784 ( .A(a[310]), .B(n3162), .Z(n766) );
  XNOR U785 ( .A(a[313]), .B(n3153), .Z(n763) );
  XNOR U786 ( .A(a[316]), .B(n3144), .Z(n760) );
  XNOR U787 ( .A(a[319]), .B(n3135), .Z(n757) );
  XNOR U788 ( .A(a[322]), .B(n3126), .Z(n753) );
  XNOR U789 ( .A(a[325]), .B(n3117), .Z(n750) );
  XNOR U790 ( .A(a[328]), .B(n3108), .Z(n747) );
  XNOR U791 ( .A(a[331]), .B(n3099), .Z(n743) );
  XNOR U792 ( .A(a[334]), .B(n3090), .Z(n740) );
  XNOR U793 ( .A(a[337]), .B(n3081), .Z(n737) );
  XNOR U794 ( .A(a[340]), .B(n3072), .Z(n733) );
  XNOR U795 ( .A(a[343]), .B(n3063), .Z(n730) );
  XNOR U796 ( .A(a[346]), .B(n3054), .Z(n727) );
  XNOR U797 ( .A(a[349]), .B(n3045), .Z(n724) );
  XNOR U798 ( .A(a[352]), .B(n3036), .Z(n720) );
  XNOR U799 ( .A(a[355]), .B(n3027), .Z(n717) );
  XNOR U800 ( .A(a[358]), .B(n3018), .Z(n714) );
  XNOR U801 ( .A(a[361]), .B(n3009), .Z(n710) );
  XNOR U802 ( .A(a[364]), .B(n3000), .Z(n707) );
  XNOR U803 ( .A(a[367]), .B(n2991), .Z(n704) );
  XNOR U804 ( .A(a[370]), .B(n2982), .Z(n700) );
  XNOR U805 ( .A(a[373]), .B(n2973), .Z(n697) );
  XNOR U806 ( .A(a[376]), .B(n2964), .Z(n694) );
  XNOR U807 ( .A(a[379]), .B(n2955), .Z(n691) );
  XNOR U808 ( .A(a[382]), .B(n2946), .Z(n687) );
  XNOR U809 ( .A(a[385]), .B(n2937), .Z(n684) );
  XNOR U810 ( .A(a[388]), .B(n2928), .Z(n681) );
  XNOR U811 ( .A(a[391]), .B(n2919), .Z(n677) );
  XNOR U812 ( .A(a[394]), .B(n2910), .Z(n674) );
  XNOR U813 ( .A(a[397]), .B(n2901), .Z(n671) );
  XNOR U814 ( .A(a[400]), .B(n2892), .Z(n666) );
  XNOR U815 ( .A(a[403]), .B(n2883), .Z(n663) );
  XNOR U816 ( .A(a[406]), .B(n2874), .Z(n660) );
  XNOR U817 ( .A(a[409]), .B(n2865), .Z(n657) );
  XNOR U818 ( .A(a[412]), .B(n2856), .Z(n653) );
  XNOR U819 ( .A(a[415]), .B(n2847), .Z(n650) );
  XNOR U820 ( .A(a[418]), .B(n2838), .Z(n647) );
  XNOR U821 ( .A(a[421]), .B(n2829), .Z(n643) );
  XNOR U822 ( .A(a[424]), .B(n2820), .Z(n640) );
  XNOR U823 ( .A(a[427]), .B(n2811), .Z(n637) );
  XNOR U824 ( .A(a[430]), .B(n2802), .Z(n633) );
  XNOR U825 ( .A(a[433]), .B(n2793), .Z(n630) );
  XNOR U826 ( .A(a[436]), .B(n2784), .Z(n627) );
  XNOR U827 ( .A(a[439]), .B(n2775), .Z(n624) );
  XNOR U828 ( .A(a[442]), .B(n2766), .Z(n620) );
  XNOR U829 ( .A(a[445]), .B(n2757), .Z(n617) );
  XNOR U830 ( .A(a[448]), .B(n2748), .Z(n614) );
  XNOR U831 ( .A(a[451]), .B(n2739), .Z(n610) );
  XNOR U832 ( .A(a[454]), .B(n2730), .Z(n607) );
  XNOR U833 ( .A(a[457]), .B(n2721), .Z(n604) );
  XNOR U834 ( .A(a[460]), .B(n2712), .Z(n600) );
  XNOR U835 ( .A(a[463]), .B(n2703), .Z(n597) );
  XNOR U836 ( .A(a[466]), .B(n2694), .Z(n594) );
  XNOR U837 ( .A(a[469]), .B(n2685), .Z(n591) );
  XNOR U838 ( .A(a[472]), .B(n2676), .Z(n587) );
  XNOR U839 ( .A(a[475]), .B(n2667), .Z(n584) );
  XNOR U840 ( .A(a[478]), .B(n2658), .Z(n581) );
  XNOR U841 ( .A(a[481]), .B(n2649), .Z(n577) );
  XNOR U842 ( .A(a[484]), .B(n2640), .Z(n574) );
  XNOR U843 ( .A(a[487]), .B(n2631), .Z(n571) );
  XNOR U844 ( .A(a[490]), .B(n2622), .Z(n567) );
  XNOR U845 ( .A(a[493]), .B(n2613), .Z(n564) );
  XNOR U846 ( .A(a[496]), .B(n2604), .Z(n561) );
  XNOR U847 ( .A(a[499]), .B(n2595), .Z(n558) );
  XNOR U848 ( .A(a[502]), .B(n2586), .Z(n553) );
  XNOR U849 ( .A(a[505]), .B(n2577), .Z(n550) );
  XNOR U850 ( .A(a[508]), .B(n2568), .Z(n547) );
  XNOR U851 ( .A(a[511]), .B(n2559), .Z(n543) );
  XNOR U852 ( .A(a[514]), .B(n2550), .Z(n540) );
  XNOR U853 ( .A(a[517]), .B(n2541), .Z(n537) );
  XNOR U854 ( .A(a[520]), .B(n2532), .Z(n533) );
  XNOR U855 ( .A(a[523]), .B(n2523), .Z(n530) );
  XNOR U856 ( .A(a[526]), .B(n2514), .Z(n527) );
  XNOR U857 ( .A(a[529]), .B(n2505), .Z(n524) );
  XNOR U858 ( .A(a[532]), .B(n2496), .Z(n520) );
  XNOR U859 ( .A(a[535]), .B(n2487), .Z(n517) );
  XNOR U860 ( .A(a[538]), .B(n2478), .Z(n514) );
  XNOR U861 ( .A(a[541]), .B(n2469), .Z(n510) );
  XNOR U862 ( .A(a[544]), .B(n2460), .Z(n507) );
  XNOR U863 ( .A(a[547]), .B(n2451), .Z(n504) );
  XNOR U864 ( .A(a[550]), .B(n2442), .Z(n500) );
  XNOR U865 ( .A(a[553]), .B(n2433), .Z(n497) );
  XNOR U866 ( .A(a[556]), .B(n2424), .Z(n494) );
  XNOR U867 ( .A(a[559]), .B(n2415), .Z(n491) );
  XNOR U868 ( .A(a[562]), .B(n2406), .Z(n487) );
  XNOR U869 ( .A(a[565]), .B(n2397), .Z(n484) );
  XNOR U870 ( .A(a[568]), .B(n2388), .Z(n481) );
  XNOR U871 ( .A(a[571]), .B(n2379), .Z(n477) );
  XNOR U872 ( .A(a[574]), .B(n2370), .Z(n474) );
  XNOR U873 ( .A(a[577]), .B(n2361), .Z(n471) );
  XNOR U874 ( .A(a[580]), .B(n2352), .Z(n467) );
  XNOR U875 ( .A(a[583]), .B(n2343), .Z(n464) );
  XNOR U876 ( .A(a[586]), .B(n2334), .Z(n461) );
  XNOR U877 ( .A(a[589]), .B(n2325), .Z(n458) );
  XNOR U878 ( .A(a[592]), .B(n2316), .Z(n454) );
  XNOR U879 ( .A(a[595]), .B(n2307), .Z(n451) );
  XNOR U880 ( .A(a[598]), .B(n2298), .Z(n448) );
  XNOR U881 ( .A(a[601]), .B(n2289), .Z(n443) );
  XNOR U882 ( .A(a[604]), .B(n2280), .Z(n440) );
  XNOR U883 ( .A(a[607]), .B(n2271), .Z(n437) );
  XNOR U884 ( .A(a[610]), .B(n2262), .Z(n433) );
  XNOR U885 ( .A(a[613]), .B(n2253), .Z(n430) );
  XNOR U886 ( .A(a[616]), .B(n2244), .Z(n427) );
  XNOR U887 ( .A(a[619]), .B(n2235), .Z(n424) );
  XNOR U888 ( .A(a[622]), .B(n2226), .Z(n420) );
  XNOR U889 ( .A(a[625]), .B(n2217), .Z(n417) );
  XNOR U890 ( .A(a[628]), .B(n2208), .Z(n414) );
  XNOR U891 ( .A(a[631]), .B(n2199), .Z(n410) );
  XNOR U892 ( .A(a[634]), .B(n2190), .Z(n407) );
  XNOR U893 ( .A(a[637]), .B(n2181), .Z(n404) );
  XNOR U894 ( .A(a[640]), .B(n2172), .Z(n400) );
  XNOR U895 ( .A(a[643]), .B(n2163), .Z(n397) );
  XNOR U896 ( .A(a[646]), .B(n2154), .Z(n394) );
  XNOR U897 ( .A(a[649]), .B(n2145), .Z(n391) );
  XNOR U898 ( .A(a[652]), .B(n2136), .Z(n387) );
  XNOR U899 ( .A(a[655]), .B(n2127), .Z(n384) );
  XNOR U900 ( .A(a[658]), .B(n2118), .Z(n381) );
  XNOR U901 ( .A(a[661]), .B(n2109), .Z(n377) );
  XNOR U902 ( .A(a[664]), .B(n2100), .Z(n374) );
  XNOR U903 ( .A(a[667]), .B(n2091), .Z(n371) );
  XNOR U904 ( .A(a[670]), .B(n2082), .Z(n367) );
  XNOR U905 ( .A(a[673]), .B(n2073), .Z(n364) );
  XNOR U906 ( .A(a[676]), .B(n2064), .Z(n361) );
  XNOR U907 ( .A(a[679]), .B(n2055), .Z(n358) );
  XNOR U908 ( .A(a[682]), .B(n2046), .Z(n354) );
  XNOR U909 ( .A(a[685]), .B(n2037), .Z(n351) );
  XNOR U910 ( .A(a[688]), .B(n2028), .Z(n348) );
  XNOR U911 ( .A(a[691]), .B(n2019), .Z(n344) );
  XNOR U912 ( .A(a[694]), .B(n2010), .Z(n341) );
  XNOR U913 ( .A(a[697]), .B(n2001), .Z(n338) );
  XNOR U914 ( .A(a[700]), .B(n1992), .Z(n333) );
  XNOR U915 ( .A(a[703]), .B(n1983), .Z(n330) );
  XNOR U916 ( .A(a[706]), .B(n1974), .Z(n327) );
  XNOR U917 ( .A(a[709]), .B(n1965), .Z(n324) );
  XNOR U918 ( .A(a[712]), .B(n1956), .Z(n320) );
  XNOR U919 ( .A(a[715]), .B(n1947), .Z(n317) );
  XNOR U920 ( .A(a[718]), .B(n1938), .Z(n314) );
  XNOR U921 ( .A(a[721]), .B(n1929), .Z(n310) );
  XNOR U922 ( .A(a[724]), .B(n1920), .Z(n307) );
  XNOR U923 ( .A(a[727]), .B(n1911), .Z(n304) );
  XNOR U924 ( .A(a[730]), .B(n1902), .Z(n300) );
  XNOR U925 ( .A(a[733]), .B(n1893), .Z(n297) );
  XNOR U926 ( .A(a[736]), .B(n1884), .Z(n294) );
  XNOR U927 ( .A(a[739]), .B(n1875), .Z(n291) );
  XNOR U928 ( .A(a[742]), .B(n1866), .Z(n287) );
  XNOR U929 ( .A(a[745]), .B(n1857), .Z(n284) );
  XNOR U930 ( .A(a[748]), .B(n1848), .Z(n281) );
  XNOR U931 ( .A(a[751]), .B(n1839), .Z(n277) );
  XNOR U932 ( .A(a[754]), .B(n1830), .Z(n274) );
  XNOR U933 ( .A(a[757]), .B(n1821), .Z(n271) );
  XNOR U934 ( .A(a[760]), .B(n1812), .Z(n267) );
  XNOR U935 ( .A(a[763]), .B(n1803), .Z(n264) );
  XNOR U936 ( .A(a[766]), .B(n1794), .Z(n261) );
  XNOR U937 ( .A(a[769]), .B(n1785), .Z(n258) );
  XNOR U938 ( .A(a[772]), .B(n1776), .Z(n254) );
  XNOR U939 ( .A(a[775]), .B(n1767), .Z(n251) );
  XNOR U940 ( .A(a[778]), .B(n1758), .Z(n248) );
  XNOR U941 ( .A(a[781]), .B(n1749), .Z(n244) );
  XNOR U942 ( .A(a[784]), .B(n1740), .Z(n241) );
  XNOR U943 ( .A(a[787]), .B(n1731), .Z(n238) );
  XNOR U944 ( .A(a[790]), .B(n1722), .Z(n234) );
  XNOR U945 ( .A(a[793]), .B(n1713), .Z(n231) );
  XNOR U946 ( .A(a[796]), .B(n1704), .Z(n228) );
  XNOR U947 ( .A(a[799]), .B(n1695), .Z(n225) );
  XNOR U948 ( .A(a[802]), .B(n1686), .Z(n220) );
  XNOR U949 ( .A(a[805]), .B(n1677), .Z(n217) );
  XNOR U950 ( .A(a[808]), .B(n1668), .Z(n214) );
  XNOR U951 ( .A(a[811]), .B(n1659), .Z(n210) );
  XNOR U952 ( .A(a[814]), .B(n1650), .Z(n207) );
  XNOR U953 ( .A(a[817]), .B(n1641), .Z(n204) );
  XNOR U954 ( .A(a[820]), .B(n1632), .Z(n200) );
  XNOR U955 ( .A(a[823]), .B(n1623), .Z(n197) );
  XNOR U956 ( .A(a[826]), .B(n1614), .Z(n194) );
  XNOR U957 ( .A(a[829]), .B(n1605), .Z(n191) );
  XNOR U958 ( .A(a[832]), .B(n1596), .Z(n187) );
  XNOR U959 ( .A(a[835]), .B(n1587), .Z(n184) );
  XNOR U960 ( .A(a[838]), .B(n1578), .Z(n181) );
  XNOR U961 ( .A(a[841]), .B(n1569), .Z(n177) );
  XNOR U962 ( .A(a[844]), .B(n1560), .Z(n174) );
  XNOR U963 ( .A(a[847]), .B(n1551), .Z(n171) );
  XNOR U964 ( .A(a[850]), .B(n1542), .Z(n167) );
  XNOR U965 ( .A(a[853]), .B(n1533), .Z(n164) );
  XNOR U966 ( .A(a[856]), .B(n1524), .Z(n161) );
  XNOR U967 ( .A(a[859]), .B(n1515), .Z(n158) );
  XNOR U968 ( .A(a[862]), .B(n1506), .Z(n154) );
  XNOR U969 ( .A(a[865]), .B(n1497), .Z(n151) );
  XNOR U970 ( .A(a[868]), .B(n1488), .Z(n148) );
  XNOR U971 ( .A(a[871]), .B(n1479), .Z(n144) );
  XNOR U972 ( .A(a[874]), .B(n1470), .Z(n141) );
  XNOR U973 ( .A(a[877]), .B(n1461), .Z(n138) );
  XNOR U974 ( .A(a[880]), .B(n1452), .Z(n134) );
  XNOR U975 ( .A(a[883]), .B(n1443), .Z(n131) );
  XNOR U976 ( .A(a[886]), .B(n1434), .Z(n128) );
  XNOR U977 ( .A(a[889]), .B(n1425), .Z(n125) );
  XNOR U978 ( .A(a[892]), .B(n1416), .Z(n121) );
  XNOR U979 ( .A(a[895]), .B(n1407), .Z(n118) );
  XNOR U980 ( .A(a[898]), .B(n1398), .Z(n115) );
  XNOR U981 ( .A(a[901]), .B(n1389), .Z(n110) );
  XNOR U982 ( .A(a[904]), .B(n1380), .Z(n107) );
  XNOR U983 ( .A(a[907]), .B(n1371), .Z(n104) );
  XNOR U984 ( .A(a[910]), .B(n1362), .Z(n100) );
  XNOR U985 ( .A(a[913]), .B(n1353), .Z(n97) );
  XNOR U986 ( .A(a[916]), .B(n1344), .Z(n94) );
  XNOR U987 ( .A(a[919]), .B(n1335), .Z(n91) );
  XNOR U988 ( .A(a[922]), .B(n1326), .Z(n87) );
  XNOR U989 ( .A(a[925]), .B(n1317), .Z(n84) );
  XNOR U990 ( .A(a[928]), .B(n1308), .Z(n81) );
  XNOR U991 ( .A(a[931]), .B(n1299), .Z(n77) );
  XNOR U992 ( .A(a[934]), .B(n1290), .Z(n74) );
  XNOR U993 ( .A(a[937]), .B(n1281), .Z(n71) );
  XNOR U994 ( .A(a[940]), .B(n1272), .Z(n67) );
  XNOR U995 ( .A(a[943]), .B(n1263), .Z(n64) );
  XNOR U996 ( .A(a[946]), .B(n1254), .Z(n61) );
  XNOR U997 ( .A(a[949]), .B(n1245), .Z(n58) );
  XNOR U998 ( .A(a[952]), .B(n1236), .Z(n54) );
  XNOR U999 ( .A(a[955]), .B(n1227), .Z(n51) );
  XNOR U1000 ( .A(a[958]), .B(n1218), .Z(n48) );
  XNOR U1001 ( .A(a[961]), .B(n1209), .Z(n44) );
  XNOR U1002 ( .A(a[964]), .B(n1200), .Z(n41) );
  XNOR U1003 ( .A(a[967]), .B(n1191), .Z(n38) );
  XNOR U1004 ( .A(a[970]), .B(n1182), .Z(n34) );
  XNOR U1005 ( .A(a[973]), .B(n1173), .Z(n31) );
  XNOR U1006 ( .A(a[976]), .B(n1164), .Z(n28) );
  XNOR U1007 ( .A(a[979]), .B(n1155), .Z(n25) );
  XNOR U1008 ( .A(a[982]), .B(n1146), .Z(n21) );
  XNOR U1009 ( .A(a[985]), .B(n1137), .Z(n18) );
  XNOR U1010 ( .A(a[988]), .B(n1128), .Z(n15) );
  XNOR U1011 ( .A(a[991]), .B(n1119), .Z(n11) );
  XNOR U1012 ( .A(a[994]), .B(n1110), .Z(n8) );
  XNOR U1013 ( .A(a[997]), .B(n1101), .Z(n5) );
  XNOR U1014 ( .A(a[1000]), .B(n1091), .Z(n1093) );
  XNOR U1015 ( .A(a[1003]), .B(n1079), .Z(n1081) );
  XNOR U1016 ( .A(a[1006]), .B(n1067), .Z(n1069) );
  XNOR U1017 ( .A(a[1009]), .B(n1054), .Z(n1056) );
  XNOR U1018 ( .A(a[1012]), .B(n1042), .Z(n1044) );
  XNOR U1019 ( .A(a[1015]), .B(n1030), .Z(n1032) );
  XNOR U1020 ( .A(a[1018]), .B(n1018), .Z(n1020) );
  XNOR U1021 ( .A(a[1021]), .B(n1005), .Z(n1007) );
  XNOR U1022 ( .A(b[9]), .B(n1), .Z(c[9]) );
  XNOR U1023 ( .A(b[99]), .B(n2), .Z(c[99]) );
  XNOR U1024 ( .A(b[999]), .B(n3), .Z(c[999]) );
  XNOR U1025 ( .A(b[998]), .B(n4), .Z(c[998]) );
  XNOR U1026 ( .A(b[997]), .B(n5), .Z(c[997]) );
  XNOR U1027 ( .A(b[996]), .B(n6), .Z(c[996]) );
  XNOR U1028 ( .A(b[995]), .B(n7), .Z(c[995]) );
  XNOR U1029 ( .A(b[994]), .B(n8), .Z(c[994]) );
  XNOR U1030 ( .A(b[993]), .B(n9), .Z(c[993]) );
  XNOR U1031 ( .A(b[992]), .B(n10), .Z(c[992]) );
  XNOR U1032 ( .A(b[991]), .B(n11), .Z(c[991]) );
  XNOR U1033 ( .A(b[990]), .B(n12), .Z(c[990]) );
  XNOR U1034 ( .A(b[98]), .B(n13), .Z(c[98]) );
  XNOR U1035 ( .A(b[989]), .B(n14), .Z(c[989]) );
  XNOR U1036 ( .A(b[988]), .B(n15), .Z(c[988]) );
  XNOR U1037 ( .A(b[987]), .B(n16), .Z(c[987]) );
  XNOR U1038 ( .A(b[986]), .B(n17), .Z(c[986]) );
  XNOR U1039 ( .A(b[985]), .B(n18), .Z(c[985]) );
  XNOR U1040 ( .A(b[984]), .B(n19), .Z(c[984]) );
  XNOR U1041 ( .A(b[983]), .B(n20), .Z(c[983]) );
  XNOR U1042 ( .A(b[982]), .B(n21), .Z(c[982]) );
  XNOR U1043 ( .A(b[981]), .B(n22), .Z(c[981]) );
  XNOR U1044 ( .A(b[980]), .B(n23), .Z(c[980]) );
  XNOR U1045 ( .A(b[97]), .B(n24), .Z(c[97]) );
  XNOR U1046 ( .A(b[979]), .B(n25), .Z(c[979]) );
  XNOR U1047 ( .A(b[978]), .B(n26), .Z(c[978]) );
  XNOR U1048 ( .A(b[977]), .B(n27), .Z(c[977]) );
  XNOR U1049 ( .A(b[976]), .B(n28), .Z(c[976]) );
  XNOR U1050 ( .A(b[975]), .B(n29), .Z(c[975]) );
  XNOR U1051 ( .A(b[974]), .B(n30), .Z(c[974]) );
  XNOR U1052 ( .A(b[973]), .B(n31), .Z(c[973]) );
  XNOR U1053 ( .A(b[972]), .B(n32), .Z(c[972]) );
  XNOR U1054 ( .A(b[971]), .B(n33), .Z(c[971]) );
  XNOR U1055 ( .A(b[970]), .B(n34), .Z(c[970]) );
  XNOR U1056 ( .A(b[96]), .B(n35), .Z(c[96]) );
  XNOR U1057 ( .A(b[969]), .B(n36), .Z(c[969]) );
  XNOR U1058 ( .A(b[968]), .B(n37), .Z(c[968]) );
  XNOR U1059 ( .A(b[967]), .B(n38), .Z(c[967]) );
  XNOR U1060 ( .A(b[966]), .B(n39), .Z(c[966]) );
  XNOR U1061 ( .A(b[965]), .B(n40), .Z(c[965]) );
  XNOR U1062 ( .A(b[964]), .B(n41), .Z(c[964]) );
  XNOR U1063 ( .A(b[963]), .B(n42), .Z(c[963]) );
  XNOR U1064 ( .A(b[962]), .B(n43), .Z(c[962]) );
  XNOR U1065 ( .A(b[961]), .B(n44), .Z(c[961]) );
  XNOR U1066 ( .A(b[960]), .B(n45), .Z(c[960]) );
  XNOR U1067 ( .A(b[95]), .B(n46), .Z(c[95]) );
  XNOR U1068 ( .A(b[959]), .B(n47), .Z(c[959]) );
  XNOR U1069 ( .A(b[958]), .B(n48), .Z(c[958]) );
  XNOR U1070 ( .A(b[957]), .B(n49), .Z(c[957]) );
  XNOR U1071 ( .A(b[956]), .B(n50), .Z(c[956]) );
  XNOR U1072 ( .A(b[955]), .B(n51), .Z(c[955]) );
  XNOR U1073 ( .A(b[954]), .B(n52), .Z(c[954]) );
  XNOR U1074 ( .A(b[953]), .B(n53), .Z(c[953]) );
  XNOR U1075 ( .A(b[952]), .B(n54), .Z(c[952]) );
  XNOR U1076 ( .A(b[951]), .B(n55), .Z(c[951]) );
  XNOR U1077 ( .A(b[950]), .B(n56), .Z(c[950]) );
  XNOR U1078 ( .A(b[94]), .B(n57), .Z(c[94]) );
  XNOR U1079 ( .A(b[949]), .B(n58), .Z(c[949]) );
  XNOR U1080 ( .A(b[948]), .B(n59), .Z(c[948]) );
  XNOR U1081 ( .A(b[947]), .B(n60), .Z(c[947]) );
  XNOR U1082 ( .A(b[946]), .B(n61), .Z(c[946]) );
  XNOR U1083 ( .A(b[945]), .B(n62), .Z(c[945]) );
  XNOR U1084 ( .A(b[944]), .B(n63), .Z(c[944]) );
  XNOR U1085 ( .A(b[943]), .B(n64), .Z(c[943]) );
  XNOR U1086 ( .A(b[942]), .B(n65), .Z(c[942]) );
  XNOR U1087 ( .A(b[941]), .B(n66), .Z(c[941]) );
  XNOR U1088 ( .A(b[940]), .B(n67), .Z(c[940]) );
  XNOR U1089 ( .A(b[93]), .B(n68), .Z(c[93]) );
  XNOR U1090 ( .A(b[939]), .B(n69), .Z(c[939]) );
  XNOR U1091 ( .A(b[938]), .B(n70), .Z(c[938]) );
  XNOR U1092 ( .A(b[937]), .B(n71), .Z(c[937]) );
  XNOR U1093 ( .A(b[936]), .B(n72), .Z(c[936]) );
  XNOR U1094 ( .A(b[935]), .B(n73), .Z(c[935]) );
  XNOR U1095 ( .A(b[934]), .B(n74), .Z(c[934]) );
  XNOR U1096 ( .A(b[933]), .B(n75), .Z(c[933]) );
  XNOR U1097 ( .A(b[932]), .B(n76), .Z(c[932]) );
  XNOR U1098 ( .A(b[931]), .B(n77), .Z(c[931]) );
  XNOR U1099 ( .A(b[930]), .B(n78), .Z(c[930]) );
  XNOR U1100 ( .A(b[92]), .B(n79), .Z(c[92]) );
  XNOR U1101 ( .A(b[929]), .B(n80), .Z(c[929]) );
  XNOR U1102 ( .A(b[928]), .B(n81), .Z(c[928]) );
  XNOR U1103 ( .A(b[927]), .B(n82), .Z(c[927]) );
  XNOR U1104 ( .A(b[926]), .B(n83), .Z(c[926]) );
  XNOR U1105 ( .A(b[925]), .B(n84), .Z(c[925]) );
  XNOR U1106 ( .A(b[924]), .B(n85), .Z(c[924]) );
  XNOR U1107 ( .A(b[923]), .B(n86), .Z(c[923]) );
  XNOR U1108 ( .A(b[922]), .B(n87), .Z(c[922]) );
  XNOR U1109 ( .A(b[921]), .B(n88), .Z(c[921]) );
  XNOR U1110 ( .A(b[920]), .B(n89), .Z(c[920]) );
  XNOR U1111 ( .A(b[91]), .B(n90), .Z(c[91]) );
  XNOR U1112 ( .A(b[919]), .B(n91), .Z(c[919]) );
  XNOR U1113 ( .A(b[918]), .B(n92), .Z(c[918]) );
  XNOR U1114 ( .A(b[917]), .B(n93), .Z(c[917]) );
  XNOR U1115 ( .A(b[916]), .B(n94), .Z(c[916]) );
  XNOR U1116 ( .A(b[915]), .B(n95), .Z(c[915]) );
  XNOR U1117 ( .A(b[914]), .B(n96), .Z(c[914]) );
  XNOR U1118 ( .A(b[913]), .B(n97), .Z(c[913]) );
  XNOR U1119 ( .A(b[912]), .B(n98), .Z(c[912]) );
  XNOR U1120 ( .A(b[911]), .B(n99), .Z(c[911]) );
  XNOR U1121 ( .A(b[910]), .B(n100), .Z(c[910]) );
  XNOR U1122 ( .A(b[90]), .B(n101), .Z(c[90]) );
  XNOR U1123 ( .A(b[909]), .B(n102), .Z(c[909]) );
  XNOR U1124 ( .A(b[908]), .B(n103), .Z(c[908]) );
  XNOR U1125 ( .A(b[907]), .B(n104), .Z(c[907]) );
  XNOR U1126 ( .A(b[906]), .B(n105), .Z(c[906]) );
  XNOR U1127 ( .A(b[905]), .B(n106), .Z(c[905]) );
  XNOR U1128 ( .A(b[904]), .B(n107), .Z(c[904]) );
  XNOR U1129 ( .A(b[903]), .B(n108), .Z(c[903]) );
  XNOR U1130 ( .A(b[902]), .B(n109), .Z(c[902]) );
  XNOR U1131 ( .A(b[901]), .B(n110), .Z(c[901]) );
  XNOR U1132 ( .A(b[900]), .B(n111), .Z(c[900]) );
  XNOR U1133 ( .A(b[8]), .B(n112), .Z(c[8]) );
  XNOR U1134 ( .A(b[89]), .B(n113), .Z(c[89]) );
  XNOR U1135 ( .A(b[899]), .B(n114), .Z(c[899]) );
  XNOR U1136 ( .A(b[898]), .B(n115), .Z(c[898]) );
  XNOR U1137 ( .A(b[897]), .B(n116), .Z(c[897]) );
  XNOR U1138 ( .A(b[896]), .B(n117), .Z(c[896]) );
  XNOR U1139 ( .A(b[895]), .B(n118), .Z(c[895]) );
  XNOR U1140 ( .A(b[894]), .B(n119), .Z(c[894]) );
  XNOR U1141 ( .A(b[893]), .B(n120), .Z(c[893]) );
  XNOR U1142 ( .A(b[892]), .B(n121), .Z(c[892]) );
  XNOR U1143 ( .A(b[891]), .B(n122), .Z(c[891]) );
  XNOR U1144 ( .A(b[890]), .B(n123), .Z(c[890]) );
  XNOR U1145 ( .A(b[88]), .B(n124), .Z(c[88]) );
  XNOR U1146 ( .A(b[889]), .B(n125), .Z(c[889]) );
  XNOR U1147 ( .A(b[888]), .B(n126), .Z(c[888]) );
  XNOR U1148 ( .A(b[887]), .B(n127), .Z(c[887]) );
  XNOR U1149 ( .A(b[886]), .B(n128), .Z(c[886]) );
  XNOR U1150 ( .A(b[885]), .B(n129), .Z(c[885]) );
  XNOR U1151 ( .A(b[884]), .B(n130), .Z(c[884]) );
  XNOR U1152 ( .A(b[883]), .B(n131), .Z(c[883]) );
  XNOR U1153 ( .A(b[882]), .B(n132), .Z(c[882]) );
  XNOR U1154 ( .A(b[881]), .B(n133), .Z(c[881]) );
  XNOR U1155 ( .A(b[880]), .B(n134), .Z(c[880]) );
  XNOR U1156 ( .A(b[87]), .B(n135), .Z(c[87]) );
  XNOR U1157 ( .A(b[879]), .B(n136), .Z(c[879]) );
  XNOR U1158 ( .A(b[878]), .B(n137), .Z(c[878]) );
  XNOR U1159 ( .A(b[877]), .B(n138), .Z(c[877]) );
  XNOR U1160 ( .A(b[876]), .B(n139), .Z(c[876]) );
  XNOR U1161 ( .A(b[875]), .B(n140), .Z(c[875]) );
  XNOR U1162 ( .A(b[874]), .B(n141), .Z(c[874]) );
  XNOR U1163 ( .A(b[873]), .B(n142), .Z(c[873]) );
  XNOR U1164 ( .A(b[872]), .B(n143), .Z(c[872]) );
  XNOR U1165 ( .A(b[871]), .B(n144), .Z(c[871]) );
  XNOR U1166 ( .A(b[870]), .B(n145), .Z(c[870]) );
  XNOR U1167 ( .A(b[86]), .B(n146), .Z(c[86]) );
  XNOR U1168 ( .A(b[869]), .B(n147), .Z(c[869]) );
  XNOR U1169 ( .A(b[868]), .B(n148), .Z(c[868]) );
  XNOR U1170 ( .A(b[867]), .B(n149), .Z(c[867]) );
  XNOR U1171 ( .A(b[866]), .B(n150), .Z(c[866]) );
  XNOR U1172 ( .A(b[865]), .B(n151), .Z(c[865]) );
  XNOR U1173 ( .A(b[864]), .B(n152), .Z(c[864]) );
  XNOR U1174 ( .A(b[863]), .B(n153), .Z(c[863]) );
  XNOR U1175 ( .A(b[862]), .B(n154), .Z(c[862]) );
  XNOR U1176 ( .A(b[861]), .B(n155), .Z(c[861]) );
  XNOR U1177 ( .A(b[860]), .B(n156), .Z(c[860]) );
  XNOR U1178 ( .A(b[85]), .B(n157), .Z(c[85]) );
  XNOR U1179 ( .A(b[859]), .B(n158), .Z(c[859]) );
  XNOR U1180 ( .A(b[858]), .B(n159), .Z(c[858]) );
  XNOR U1181 ( .A(b[857]), .B(n160), .Z(c[857]) );
  XNOR U1182 ( .A(b[856]), .B(n161), .Z(c[856]) );
  XNOR U1183 ( .A(b[855]), .B(n162), .Z(c[855]) );
  XNOR U1184 ( .A(b[854]), .B(n163), .Z(c[854]) );
  XNOR U1185 ( .A(b[853]), .B(n164), .Z(c[853]) );
  XNOR U1186 ( .A(b[852]), .B(n165), .Z(c[852]) );
  XNOR U1187 ( .A(b[851]), .B(n166), .Z(c[851]) );
  XNOR U1188 ( .A(b[850]), .B(n167), .Z(c[850]) );
  XNOR U1189 ( .A(b[84]), .B(n168), .Z(c[84]) );
  XNOR U1190 ( .A(b[849]), .B(n169), .Z(c[849]) );
  XNOR U1191 ( .A(b[848]), .B(n170), .Z(c[848]) );
  XNOR U1192 ( .A(b[847]), .B(n171), .Z(c[847]) );
  XNOR U1193 ( .A(b[846]), .B(n172), .Z(c[846]) );
  XNOR U1194 ( .A(b[845]), .B(n173), .Z(c[845]) );
  XNOR U1195 ( .A(b[844]), .B(n174), .Z(c[844]) );
  XNOR U1196 ( .A(b[843]), .B(n175), .Z(c[843]) );
  XNOR U1197 ( .A(b[842]), .B(n176), .Z(c[842]) );
  XNOR U1198 ( .A(b[841]), .B(n177), .Z(c[841]) );
  XNOR U1199 ( .A(b[840]), .B(n178), .Z(c[840]) );
  XNOR U1200 ( .A(b[83]), .B(n179), .Z(c[83]) );
  XNOR U1201 ( .A(b[839]), .B(n180), .Z(c[839]) );
  XNOR U1202 ( .A(b[838]), .B(n181), .Z(c[838]) );
  XNOR U1203 ( .A(b[837]), .B(n182), .Z(c[837]) );
  XNOR U1204 ( .A(b[836]), .B(n183), .Z(c[836]) );
  XNOR U1205 ( .A(b[835]), .B(n184), .Z(c[835]) );
  XNOR U1206 ( .A(b[834]), .B(n185), .Z(c[834]) );
  XNOR U1207 ( .A(b[833]), .B(n186), .Z(c[833]) );
  XNOR U1208 ( .A(b[832]), .B(n187), .Z(c[832]) );
  XNOR U1209 ( .A(b[831]), .B(n188), .Z(c[831]) );
  XNOR U1210 ( .A(b[830]), .B(n189), .Z(c[830]) );
  XNOR U1211 ( .A(b[82]), .B(n190), .Z(c[82]) );
  XNOR U1212 ( .A(b[829]), .B(n191), .Z(c[829]) );
  XNOR U1213 ( .A(b[828]), .B(n192), .Z(c[828]) );
  XNOR U1214 ( .A(b[827]), .B(n193), .Z(c[827]) );
  XNOR U1215 ( .A(b[826]), .B(n194), .Z(c[826]) );
  XNOR U1216 ( .A(b[825]), .B(n195), .Z(c[825]) );
  XNOR U1217 ( .A(b[824]), .B(n196), .Z(c[824]) );
  XNOR U1218 ( .A(b[823]), .B(n197), .Z(c[823]) );
  XNOR U1219 ( .A(b[822]), .B(n198), .Z(c[822]) );
  XNOR U1220 ( .A(b[821]), .B(n199), .Z(c[821]) );
  XNOR U1221 ( .A(b[820]), .B(n200), .Z(c[820]) );
  XNOR U1222 ( .A(b[81]), .B(n201), .Z(c[81]) );
  XNOR U1223 ( .A(b[819]), .B(n202), .Z(c[819]) );
  XNOR U1224 ( .A(b[818]), .B(n203), .Z(c[818]) );
  XNOR U1225 ( .A(b[817]), .B(n204), .Z(c[817]) );
  XNOR U1226 ( .A(b[816]), .B(n205), .Z(c[816]) );
  XNOR U1227 ( .A(b[815]), .B(n206), .Z(c[815]) );
  XNOR U1228 ( .A(b[814]), .B(n207), .Z(c[814]) );
  XNOR U1229 ( .A(b[813]), .B(n208), .Z(c[813]) );
  XNOR U1230 ( .A(b[812]), .B(n209), .Z(c[812]) );
  XNOR U1231 ( .A(b[811]), .B(n210), .Z(c[811]) );
  XNOR U1232 ( .A(b[810]), .B(n211), .Z(c[810]) );
  XNOR U1233 ( .A(b[80]), .B(n212), .Z(c[80]) );
  XNOR U1234 ( .A(b[809]), .B(n213), .Z(c[809]) );
  XNOR U1235 ( .A(b[808]), .B(n214), .Z(c[808]) );
  XNOR U1236 ( .A(b[807]), .B(n215), .Z(c[807]) );
  XNOR U1237 ( .A(b[806]), .B(n216), .Z(c[806]) );
  XNOR U1238 ( .A(b[805]), .B(n217), .Z(c[805]) );
  XNOR U1239 ( .A(b[804]), .B(n218), .Z(c[804]) );
  XNOR U1240 ( .A(b[803]), .B(n219), .Z(c[803]) );
  XNOR U1241 ( .A(b[802]), .B(n220), .Z(c[802]) );
  XNOR U1242 ( .A(b[801]), .B(n221), .Z(c[801]) );
  XNOR U1243 ( .A(b[800]), .B(n222), .Z(c[800]) );
  XNOR U1244 ( .A(b[7]), .B(n223), .Z(c[7]) );
  XNOR U1245 ( .A(b[79]), .B(n224), .Z(c[79]) );
  XNOR U1246 ( .A(b[799]), .B(n225), .Z(c[799]) );
  XNOR U1247 ( .A(b[798]), .B(n226), .Z(c[798]) );
  XNOR U1248 ( .A(b[797]), .B(n227), .Z(c[797]) );
  XNOR U1249 ( .A(b[796]), .B(n228), .Z(c[796]) );
  XNOR U1250 ( .A(b[795]), .B(n229), .Z(c[795]) );
  XNOR U1251 ( .A(b[794]), .B(n230), .Z(c[794]) );
  XNOR U1252 ( .A(b[793]), .B(n231), .Z(c[793]) );
  XNOR U1253 ( .A(b[792]), .B(n232), .Z(c[792]) );
  XNOR U1254 ( .A(b[791]), .B(n233), .Z(c[791]) );
  XNOR U1255 ( .A(b[790]), .B(n234), .Z(c[790]) );
  XNOR U1256 ( .A(b[78]), .B(n235), .Z(c[78]) );
  XNOR U1257 ( .A(b[789]), .B(n236), .Z(c[789]) );
  XNOR U1258 ( .A(b[788]), .B(n237), .Z(c[788]) );
  XNOR U1259 ( .A(b[787]), .B(n238), .Z(c[787]) );
  XNOR U1260 ( .A(b[786]), .B(n239), .Z(c[786]) );
  XNOR U1261 ( .A(b[785]), .B(n240), .Z(c[785]) );
  XNOR U1262 ( .A(b[784]), .B(n241), .Z(c[784]) );
  XNOR U1263 ( .A(b[783]), .B(n242), .Z(c[783]) );
  XNOR U1264 ( .A(b[782]), .B(n243), .Z(c[782]) );
  XNOR U1265 ( .A(b[781]), .B(n244), .Z(c[781]) );
  XNOR U1266 ( .A(b[780]), .B(n245), .Z(c[780]) );
  XNOR U1267 ( .A(b[77]), .B(n246), .Z(c[77]) );
  XNOR U1268 ( .A(b[779]), .B(n247), .Z(c[779]) );
  XNOR U1269 ( .A(b[778]), .B(n248), .Z(c[778]) );
  XNOR U1270 ( .A(b[777]), .B(n249), .Z(c[777]) );
  XNOR U1271 ( .A(b[776]), .B(n250), .Z(c[776]) );
  XNOR U1272 ( .A(b[775]), .B(n251), .Z(c[775]) );
  XNOR U1273 ( .A(b[774]), .B(n252), .Z(c[774]) );
  XNOR U1274 ( .A(b[773]), .B(n253), .Z(c[773]) );
  XNOR U1275 ( .A(b[772]), .B(n254), .Z(c[772]) );
  XNOR U1276 ( .A(b[771]), .B(n255), .Z(c[771]) );
  XNOR U1277 ( .A(b[770]), .B(n256), .Z(c[770]) );
  XNOR U1278 ( .A(b[76]), .B(n257), .Z(c[76]) );
  XNOR U1279 ( .A(b[769]), .B(n258), .Z(c[769]) );
  XNOR U1280 ( .A(b[768]), .B(n259), .Z(c[768]) );
  XNOR U1281 ( .A(b[767]), .B(n260), .Z(c[767]) );
  XNOR U1282 ( .A(b[766]), .B(n261), .Z(c[766]) );
  XNOR U1283 ( .A(b[765]), .B(n262), .Z(c[765]) );
  XNOR U1284 ( .A(b[764]), .B(n263), .Z(c[764]) );
  XNOR U1285 ( .A(b[763]), .B(n264), .Z(c[763]) );
  XNOR U1286 ( .A(b[762]), .B(n265), .Z(c[762]) );
  XNOR U1287 ( .A(b[761]), .B(n266), .Z(c[761]) );
  XNOR U1288 ( .A(b[760]), .B(n267), .Z(c[760]) );
  XNOR U1289 ( .A(b[75]), .B(n268), .Z(c[75]) );
  XNOR U1290 ( .A(b[759]), .B(n269), .Z(c[759]) );
  XNOR U1291 ( .A(b[758]), .B(n270), .Z(c[758]) );
  XNOR U1292 ( .A(b[757]), .B(n271), .Z(c[757]) );
  XNOR U1293 ( .A(b[756]), .B(n272), .Z(c[756]) );
  XNOR U1294 ( .A(b[755]), .B(n273), .Z(c[755]) );
  XNOR U1295 ( .A(b[754]), .B(n274), .Z(c[754]) );
  XNOR U1296 ( .A(b[753]), .B(n275), .Z(c[753]) );
  XNOR U1297 ( .A(b[752]), .B(n276), .Z(c[752]) );
  XNOR U1298 ( .A(b[751]), .B(n277), .Z(c[751]) );
  XNOR U1299 ( .A(b[750]), .B(n278), .Z(c[750]) );
  XNOR U1300 ( .A(b[74]), .B(n279), .Z(c[74]) );
  XNOR U1301 ( .A(b[749]), .B(n280), .Z(c[749]) );
  XNOR U1302 ( .A(b[748]), .B(n281), .Z(c[748]) );
  XNOR U1303 ( .A(b[747]), .B(n282), .Z(c[747]) );
  XNOR U1304 ( .A(b[746]), .B(n283), .Z(c[746]) );
  XNOR U1305 ( .A(b[745]), .B(n284), .Z(c[745]) );
  XNOR U1306 ( .A(b[744]), .B(n285), .Z(c[744]) );
  XNOR U1307 ( .A(b[743]), .B(n286), .Z(c[743]) );
  XNOR U1308 ( .A(b[742]), .B(n287), .Z(c[742]) );
  XNOR U1309 ( .A(b[741]), .B(n288), .Z(c[741]) );
  XNOR U1310 ( .A(b[740]), .B(n289), .Z(c[740]) );
  XNOR U1311 ( .A(b[73]), .B(n290), .Z(c[73]) );
  XNOR U1312 ( .A(b[739]), .B(n291), .Z(c[739]) );
  XNOR U1313 ( .A(b[738]), .B(n292), .Z(c[738]) );
  XNOR U1314 ( .A(b[737]), .B(n293), .Z(c[737]) );
  XNOR U1315 ( .A(b[736]), .B(n294), .Z(c[736]) );
  XNOR U1316 ( .A(b[735]), .B(n295), .Z(c[735]) );
  XNOR U1317 ( .A(b[734]), .B(n296), .Z(c[734]) );
  XNOR U1318 ( .A(b[733]), .B(n297), .Z(c[733]) );
  XNOR U1319 ( .A(b[732]), .B(n298), .Z(c[732]) );
  XNOR U1320 ( .A(b[731]), .B(n299), .Z(c[731]) );
  XNOR U1321 ( .A(b[730]), .B(n300), .Z(c[730]) );
  XNOR U1322 ( .A(b[72]), .B(n301), .Z(c[72]) );
  XNOR U1323 ( .A(b[729]), .B(n302), .Z(c[729]) );
  XNOR U1324 ( .A(b[728]), .B(n303), .Z(c[728]) );
  XNOR U1325 ( .A(b[727]), .B(n304), .Z(c[727]) );
  XNOR U1326 ( .A(b[726]), .B(n305), .Z(c[726]) );
  XNOR U1327 ( .A(b[725]), .B(n306), .Z(c[725]) );
  XNOR U1328 ( .A(b[724]), .B(n307), .Z(c[724]) );
  XNOR U1329 ( .A(b[723]), .B(n308), .Z(c[723]) );
  XNOR U1330 ( .A(b[722]), .B(n309), .Z(c[722]) );
  XNOR U1331 ( .A(b[721]), .B(n310), .Z(c[721]) );
  XNOR U1332 ( .A(b[720]), .B(n311), .Z(c[720]) );
  XNOR U1333 ( .A(b[71]), .B(n312), .Z(c[71]) );
  XNOR U1334 ( .A(b[719]), .B(n313), .Z(c[719]) );
  XNOR U1335 ( .A(b[718]), .B(n314), .Z(c[718]) );
  XNOR U1336 ( .A(b[717]), .B(n315), .Z(c[717]) );
  XNOR U1337 ( .A(b[716]), .B(n316), .Z(c[716]) );
  XNOR U1338 ( .A(b[715]), .B(n317), .Z(c[715]) );
  XNOR U1339 ( .A(b[714]), .B(n318), .Z(c[714]) );
  XNOR U1340 ( .A(b[713]), .B(n319), .Z(c[713]) );
  XNOR U1341 ( .A(b[712]), .B(n320), .Z(c[712]) );
  XNOR U1342 ( .A(b[711]), .B(n321), .Z(c[711]) );
  XNOR U1343 ( .A(b[710]), .B(n322), .Z(c[710]) );
  XNOR U1344 ( .A(b[70]), .B(n323), .Z(c[70]) );
  XNOR U1345 ( .A(b[709]), .B(n324), .Z(c[709]) );
  XNOR U1346 ( .A(b[708]), .B(n325), .Z(c[708]) );
  XNOR U1347 ( .A(b[707]), .B(n326), .Z(c[707]) );
  XNOR U1348 ( .A(b[706]), .B(n327), .Z(c[706]) );
  XNOR U1349 ( .A(b[705]), .B(n328), .Z(c[705]) );
  XNOR U1350 ( .A(b[704]), .B(n329), .Z(c[704]) );
  XNOR U1351 ( .A(b[703]), .B(n330), .Z(c[703]) );
  XNOR U1352 ( .A(b[702]), .B(n331), .Z(c[702]) );
  XNOR U1353 ( .A(b[701]), .B(n332), .Z(c[701]) );
  XNOR U1354 ( .A(b[700]), .B(n333), .Z(c[700]) );
  XNOR U1355 ( .A(b[6]), .B(n334), .Z(c[6]) );
  XNOR U1356 ( .A(b[69]), .B(n335), .Z(c[69]) );
  XNOR U1357 ( .A(b[699]), .B(n336), .Z(c[699]) );
  XNOR U1358 ( .A(b[698]), .B(n337), .Z(c[698]) );
  XNOR U1359 ( .A(b[697]), .B(n338), .Z(c[697]) );
  XNOR U1360 ( .A(b[696]), .B(n339), .Z(c[696]) );
  XNOR U1361 ( .A(b[695]), .B(n340), .Z(c[695]) );
  XNOR U1362 ( .A(b[694]), .B(n341), .Z(c[694]) );
  XNOR U1363 ( .A(b[693]), .B(n342), .Z(c[693]) );
  XNOR U1364 ( .A(b[692]), .B(n343), .Z(c[692]) );
  XNOR U1365 ( .A(b[691]), .B(n344), .Z(c[691]) );
  XNOR U1366 ( .A(b[690]), .B(n345), .Z(c[690]) );
  XNOR U1367 ( .A(b[68]), .B(n346), .Z(c[68]) );
  XNOR U1368 ( .A(b[689]), .B(n347), .Z(c[689]) );
  XNOR U1369 ( .A(b[688]), .B(n348), .Z(c[688]) );
  XNOR U1370 ( .A(b[687]), .B(n349), .Z(c[687]) );
  XNOR U1371 ( .A(b[686]), .B(n350), .Z(c[686]) );
  XNOR U1372 ( .A(b[685]), .B(n351), .Z(c[685]) );
  XNOR U1373 ( .A(b[684]), .B(n352), .Z(c[684]) );
  XNOR U1374 ( .A(b[683]), .B(n353), .Z(c[683]) );
  XNOR U1375 ( .A(b[682]), .B(n354), .Z(c[682]) );
  XNOR U1376 ( .A(b[681]), .B(n355), .Z(c[681]) );
  XNOR U1377 ( .A(b[680]), .B(n356), .Z(c[680]) );
  XNOR U1378 ( .A(b[67]), .B(n357), .Z(c[67]) );
  XNOR U1379 ( .A(b[679]), .B(n358), .Z(c[679]) );
  XNOR U1380 ( .A(b[678]), .B(n359), .Z(c[678]) );
  XNOR U1381 ( .A(b[677]), .B(n360), .Z(c[677]) );
  XNOR U1382 ( .A(b[676]), .B(n361), .Z(c[676]) );
  XNOR U1383 ( .A(b[675]), .B(n362), .Z(c[675]) );
  XNOR U1384 ( .A(b[674]), .B(n363), .Z(c[674]) );
  XNOR U1385 ( .A(b[673]), .B(n364), .Z(c[673]) );
  XNOR U1386 ( .A(b[672]), .B(n365), .Z(c[672]) );
  XNOR U1387 ( .A(b[671]), .B(n366), .Z(c[671]) );
  XNOR U1388 ( .A(b[670]), .B(n367), .Z(c[670]) );
  XNOR U1389 ( .A(b[66]), .B(n368), .Z(c[66]) );
  XNOR U1390 ( .A(b[669]), .B(n369), .Z(c[669]) );
  XNOR U1391 ( .A(b[668]), .B(n370), .Z(c[668]) );
  XNOR U1392 ( .A(b[667]), .B(n371), .Z(c[667]) );
  XNOR U1393 ( .A(b[666]), .B(n372), .Z(c[666]) );
  XNOR U1394 ( .A(b[665]), .B(n373), .Z(c[665]) );
  XNOR U1395 ( .A(b[664]), .B(n374), .Z(c[664]) );
  XNOR U1396 ( .A(b[663]), .B(n375), .Z(c[663]) );
  XNOR U1397 ( .A(b[662]), .B(n376), .Z(c[662]) );
  XNOR U1398 ( .A(b[661]), .B(n377), .Z(c[661]) );
  XNOR U1399 ( .A(b[660]), .B(n378), .Z(c[660]) );
  XNOR U1400 ( .A(b[65]), .B(n379), .Z(c[65]) );
  XNOR U1401 ( .A(b[659]), .B(n380), .Z(c[659]) );
  XNOR U1402 ( .A(b[658]), .B(n381), .Z(c[658]) );
  XNOR U1403 ( .A(b[657]), .B(n382), .Z(c[657]) );
  XNOR U1404 ( .A(b[656]), .B(n383), .Z(c[656]) );
  XNOR U1405 ( .A(b[655]), .B(n384), .Z(c[655]) );
  XNOR U1406 ( .A(b[654]), .B(n385), .Z(c[654]) );
  XNOR U1407 ( .A(b[653]), .B(n386), .Z(c[653]) );
  XNOR U1408 ( .A(b[652]), .B(n387), .Z(c[652]) );
  XNOR U1409 ( .A(b[651]), .B(n388), .Z(c[651]) );
  XNOR U1410 ( .A(b[650]), .B(n389), .Z(c[650]) );
  XNOR U1411 ( .A(b[64]), .B(n390), .Z(c[64]) );
  XNOR U1412 ( .A(b[649]), .B(n391), .Z(c[649]) );
  XNOR U1413 ( .A(b[648]), .B(n392), .Z(c[648]) );
  XNOR U1414 ( .A(b[647]), .B(n393), .Z(c[647]) );
  XNOR U1415 ( .A(b[646]), .B(n394), .Z(c[646]) );
  XNOR U1416 ( .A(b[645]), .B(n395), .Z(c[645]) );
  XNOR U1417 ( .A(b[644]), .B(n396), .Z(c[644]) );
  XNOR U1418 ( .A(b[643]), .B(n397), .Z(c[643]) );
  XNOR U1419 ( .A(b[642]), .B(n398), .Z(c[642]) );
  XNOR U1420 ( .A(b[641]), .B(n399), .Z(c[641]) );
  XNOR U1421 ( .A(b[640]), .B(n400), .Z(c[640]) );
  XNOR U1422 ( .A(b[63]), .B(n401), .Z(c[63]) );
  XNOR U1423 ( .A(b[639]), .B(n402), .Z(c[639]) );
  XNOR U1424 ( .A(b[638]), .B(n403), .Z(c[638]) );
  XNOR U1425 ( .A(b[637]), .B(n404), .Z(c[637]) );
  XNOR U1426 ( .A(b[636]), .B(n405), .Z(c[636]) );
  XNOR U1427 ( .A(b[635]), .B(n406), .Z(c[635]) );
  XNOR U1428 ( .A(b[634]), .B(n407), .Z(c[634]) );
  XNOR U1429 ( .A(b[633]), .B(n408), .Z(c[633]) );
  XNOR U1430 ( .A(b[632]), .B(n409), .Z(c[632]) );
  XNOR U1431 ( .A(b[631]), .B(n410), .Z(c[631]) );
  XNOR U1432 ( .A(b[630]), .B(n411), .Z(c[630]) );
  XNOR U1433 ( .A(b[62]), .B(n412), .Z(c[62]) );
  XNOR U1434 ( .A(b[629]), .B(n413), .Z(c[629]) );
  XNOR U1435 ( .A(b[628]), .B(n414), .Z(c[628]) );
  XNOR U1436 ( .A(b[627]), .B(n415), .Z(c[627]) );
  XNOR U1437 ( .A(b[626]), .B(n416), .Z(c[626]) );
  XNOR U1438 ( .A(b[625]), .B(n417), .Z(c[625]) );
  XNOR U1439 ( .A(b[624]), .B(n418), .Z(c[624]) );
  XNOR U1440 ( .A(b[623]), .B(n419), .Z(c[623]) );
  XNOR U1441 ( .A(b[622]), .B(n420), .Z(c[622]) );
  XNOR U1442 ( .A(b[621]), .B(n421), .Z(c[621]) );
  XNOR U1443 ( .A(b[620]), .B(n422), .Z(c[620]) );
  XNOR U1444 ( .A(b[61]), .B(n423), .Z(c[61]) );
  XNOR U1445 ( .A(b[619]), .B(n424), .Z(c[619]) );
  XNOR U1446 ( .A(b[618]), .B(n425), .Z(c[618]) );
  XNOR U1447 ( .A(b[617]), .B(n426), .Z(c[617]) );
  XNOR U1448 ( .A(b[616]), .B(n427), .Z(c[616]) );
  XNOR U1449 ( .A(b[615]), .B(n428), .Z(c[615]) );
  XNOR U1450 ( .A(b[614]), .B(n429), .Z(c[614]) );
  XNOR U1451 ( .A(b[613]), .B(n430), .Z(c[613]) );
  XNOR U1452 ( .A(b[612]), .B(n431), .Z(c[612]) );
  XNOR U1453 ( .A(b[611]), .B(n432), .Z(c[611]) );
  XNOR U1454 ( .A(b[610]), .B(n433), .Z(c[610]) );
  XNOR U1455 ( .A(b[60]), .B(n434), .Z(c[60]) );
  XNOR U1456 ( .A(b[609]), .B(n435), .Z(c[609]) );
  XNOR U1457 ( .A(b[608]), .B(n436), .Z(c[608]) );
  XNOR U1458 ( .A(b[607]), .B(n437), .Z(c[607]) );
  XNOR U1459 ( .A(b[606]), .B(n438), .Z(c[606]) );
  XNOR U1460 ( .A(b[605]), .B(n439), .Z(c[605]) );
  XNOR U1461 ( .A(b[604]), .B(n440), .Z(c[604]) );
  XNOR U1462 ( .A(b[603]), .B(n441), .Z(c[603]) );
  XNOR U1463 ( .A(b[602]), .B(n442), .Z(c[602]) );
  XNOR U1464 ( .A(b[601]), .B(n443), .Z(c[601]) );
  XNOR U1465 ( .A(b[600]), .B(n444), .Z(c[600]) );
  XNOR U1466 ( .A(b[5]), .B(n445), .Z(c[5]) );
  XNOR U1467 ( .A(b[59]), .B(n446), .Z(c[59]) );
  XNOR U1468 ( .A(b[599]), .B(n447), .Z(c[599]) );
  XNOR U1469 ( .A(b[598]), .B(n448), .Z(c[598]) );
  XNOR U1470 ( .A(b[597]), .B(n449), .Z(c[597]) );
  XNOR U1471 ( .A(b[596]), .B(n450), .Z(c[596]) );
  XNOR U1472 ( .A(b[595]), .B(n451), .Z(c[595]) );
  XNOR U1473 ( .A(b[594]), .B(n452), .Z(c[594]) );
  XNOR U1474 ( .A(b[593]), .B(n453), .Z(c[593]) );
  XNOR U1475 ( .A(b[592]), .B(n454), .Z(c[592]) );
  XNOR U1476 ( .A(b[591]), .B(n455), .Z(c[591]) );
  XNOR U1477 ( .A(b[590]), .B(n456), .Z(c[590]) );
  XNOR U1478 ( .A(b[58]), .B(n457), .Z(c[58]) );
  XNOR U1479 ( .A(b[589]), .B(n458), .Z(c[589]) );
  XNOR U1480 ( .A(b[588]), .B(n459), .Z(c[588]) );
  XNOR U1481 ( .A(b[587]), .B(n460), .Z(c[587]) );
  XNOR U1482 ( .A(b[586]), .B(n461), .Z(c[586]) );
  XNOR U1483 ( .A(b[585]), .B(n462), .Z(c[585]) );
  XNOR U1484 ( .A(b[584]), .B(n463), .Z(c[584]) );
  XNOR U1485 ( .A(b[583]), .B(n464), .Z(c[583]) );
  XNOR U1486 ( .A(b[582]), .B(n465), .Z(c[582]) );
  XNOR U1487 ( .A(b[581]), .B(n466), .Z(c[581]) );
  XNOR U1488 ( .A(b[580]), .B(n467), .Z(c[580]) );
  XNOR U1489 ( .A(b[57]), .B(n468), .Z(c[57]) );
  XNOR U1490 ( .A(b[579]), .B(n469), .Z(c[579]) );
  XNOR U1491 ( .A(b[578]), .B(n470), .Z(c[578]) );
  XNOR U1492 ( .A(b[577]), .B(n471), .Z(c[577]) );
  XNOR U1493 ( .A(b[576]), .B(n472), .Z(c[576]) );
  XNOR U1494 ( .A(b[575]), .B(n473), .Z(c[575]) );
  XNOR U1495 ( .A(b[574]), .B(n474), .Z(c[574]) );
  XNOR U1496 ( .A(b[573]), .B(n475), .Z(c[573]) );
  XNOR U1497 ( .A(b[572]), .B(n476), .Z(c[572]) );
  XNOR U1498 ( .A(b[571]), .B(n477), .Z(c[571]) );
  XNOR U1499 ( .A(b[570]), .B(n478), .Z(c[570]) );
  XNOR U1500 ( .A(b[56]), .B(n479), .Z(c[56]) );
  XNOR U1501 ( .A(b[569]), .B(n480), .Z(c[569]) );
  XNOR U1502 ( .A(b[568]), .B(n481), .Z(c[568]) );
  XNOR U1503 ( .A(b[567]), .B(n482), .Z(c[567]) );
  XNOR U1504 ( .A(b[566]), .B(n483), .Z(c[566]) );
  XNOR U1505 ( .A(b[565]), .B(n484), .Z(c[565]) );
  XNOR U1506 ( .A(b[564]), .B(n485), .Z(c[564]) );
  XNOR U1507 ( .A(b[563]), .B(n486), .Z(c[563]) );
  XNOR U1508 ( .A(b[562]), .B(n487), .Z(c[562]) );
  XNOR U1509 ( .A(b[561]), .B(n488), .Z(c[561]) );
  XNOR U1510 ( .A(b[560]), .B(n489), .Z(c[560]) );
  XNOR U1511 ( .A(b[55]), .B(n490), .Z(c[55]) );
  XNOR U1512 ( .A(b[559]), .B(n491), .Z(c[559]) );
  XNOR U1513 ( .A(b[558]), .B(n492), .Z(c[558]) );
  XNOR U1514 ( .A(b[557]), .B(n493), .Z(c[557]) );
  XNOR U1515 ( .A(b[556]), .B(n494), .Z(c[556]) );
  XNOR U1516 ( .A(b[555]), .B(n495), .Z(c[555]) );
  XNOR U1517 ( .A(b[554]), .B(n496), .Z(c[554]) );
  XNOR U1518 ( .A(b[553]), .B(n497), .Z(c[553]) );
  XNOR U1519 ( .A(b[552]), .B(n498), .Z(c[552]) );
  XNOR U1520 ( .A(b[551]), .B(n499), .Z(c[551]) );
  XNOR U1521 ( .A(b[550]), .B(n500), .Z(c[550]) );
  XNOR U1522 ( .A(b[54]), .B(n501), .Z(c[54]) );
  XNOR U1523 ( .A(b[549]), .B(n502), .Z(c[549]) );
  XNOR U1524 ( .A(b[548]), .B(n503), .Z(c[548]) );
  XNOR U1525 ( .A(b[547]), .B(n504), .Z(c[547]) );
  XNOR U1526 ( .A(b[546]), .B(n505), .Z(c[546]) );
  XNOR U1527 ( .A(b[545]), .B(n506), .Z(c[545]) );
  XNOR U1528 ( .A(b[544]), .B(n507), .Z(c[544]) );
  XNOR U1529 ( .A(b[543]), .B(n508), .Z(c[543]) );
  XNOR U1530 ( .A(b[542]), .B(n509), .Z(c[542]) );
  XNOR U1531 ( .A(b[541]), .B(n510), .Z(c[541]) );
  XNOR U1532 ( .A(b[540]), .B(n511), .Z(c[540]) );
  XNOR U1533 ( .A(b[53]), .B(n512), .Z(c[53]) );
  XNOR U1534 ( .A(b[539]), .B(n513), .Z(c[539]) );
  XNOR U1535 ( .A(b[538]), .B(n514), .Z(c[538]) );
  XNOR U1536 ( .A(b[537]), .B(n515), .Z(c[537]) );
  XNOR U1537 ( .A(b[536]), .B(n516), .Z(c[536]) );
  XNOR U1538 ( .A(b[535]), .B(n517), .Z(c[535]) );
  XNOR U1539 ( .A(b[534]), .B(n518), .Z(c[534]) );
  XNOR U1540 ( .A(b[533]), .B(n519), .Z(c[533]) );
  XNOR U1541 ( .A(b[532]), .B(n520), .Z(c[532]) );
  XNOR U1542 ( .A(b[531]), .B(n521), .Z(c[531]) );
  XNOR U1543 ( .A(b[530]), .B(n522), .Z(c[530]) );
  XNOR U1544 ( .A(b[52]), .B(n523), .Z(c[52]) );
  XNOR U1545 ( .A(b[529]), .B(n524), .Z(c[529]) );
  XNOR U1546 ( .A(b[528]), .B(n525), .Z(c[528]) );
  XNOR U1547 ( .A(b[527]), .B(n526), .Z(c[527]) );
  XNOR U1548 ( .A(b[526]), .B(n527), .Z(c[526]) );
  XNOR U1549 ( .A(b[525]), .B(n528), .Z(c[525]) );
  XNOR U1550 ( .A(b[524]), .B(n529), .Z(c[524]) );
  XNOR U1551 ( .A(b[523]), .B(n530), .Z(c[523]) );
  XNOR U1552 ( .A(b[522]), .B(n531), .Z(c[522]) );
  XNOR U1553 ( .A(b[521]), .B(n532), .Z(c[521]) );
  XNOR U1554 ( .A(b[520]), .B(n533), .Z(c[520]) );
  XNOR U1555 ( .A(b[51]), .B(n534), .Z(c[51]) );
  XNOR U1556 ( .A(b[519]), .B(n535), .Z(c[519]) );
  XNOR U1557 ( .A(b[518]), .B(n536), .Z(c[518]) );
  XNOR U1558 ( .A(b[517]), .B(n537), .Z(c[517]) );
  XNOR U1559 ( .A(b[516]), .B(n538), .Z(c[516]) );
  XNOR U1560 ( .A(b[515]), .B(n539), .Z(c[515]) );
  XNOR U1561 ( .A(b[514]), .B(n540), .Z(c[514]) );
  XNOR U1562 ( .A(b[513]), .B(n541), .Z(c[513]) );
  XNOR U1563 ( .A(b[512]), .B(n542), .Z(c[512]) );
  XNOR U1564 ( .A(b[511]), .B(n543), .Z(c[511]) );
  XNOR U1565 ( .A(b[510]), .B(n544), .Z(c[510]) );
  XNOR U1566 ( .A(b[50]), .B(n545), .Z(c[50]) );
  XNOR U1567 ( .A(b[509]), .B(n546), .Z(c[509]) );
  XNOR U1568 ( .A(b[508]), .B(n547), .Z(c[508]) );
  XNOR U1569 ( .A(b[507]), .B(n548), .Z(c[507]) );
  XNOR U1570 ( .A(b[506]), .B(n549), .Z(c[506]) );
  XNOR U1571 ( .A(b[505]), .B(n550), .Z(c[505]) );
  XNOR U1572 ( .A(b[504]), .B(n551), .Z(c[504]) );
  XNOR U1573 ( .A(b[503]), .B(n552), .Z(c[503]) );
  XNOR U1574 ( .A(b[502]), .B(n553), .Z(c[502]) );
  XNOR U1575 ( .A(b[501]), .B(n554), .Z(c[501]) );
  XNOR U1576 ( .A(b[500]), .B(n555), .Z(c[500]) );
  XNOR U1577 ( .A(b[4]), .B(n556), .Z(c[4]) );
  XNOR U1578 ( .A(b[49]), .B(n557), .Z(c[49]) );
  XNOR U1579 ( .A(b[499]), .B(n558), .Z(c[499]) );
  XNOR U1580 ( .A(b[498]), .B(n559), .Z(c[498]) );
  XNOR U1581 ( .A(b[497]), .B(n560), .Z(c[497]) );
  XNOR U1582 ( .A(b[496]), .B(n561), .Z(c[496]) );
  XNOR U1583 ( .A(b[495]), .B(n562), .Z(c[495]) );
  XNOR U1584 ( .A(b[494]), .B(n563), .Z(c[494]) );
  XNOR U1585 ( .A(b[493]), .B(n564), .Z(c[493]) );
  XNOR U1586 ( .A(b[492]), .B(n565), .Z(c[492]) );
  XNOR U1587 ( .A(b[491]), .B(n566), .Z(c[491]) );
  XNOR U1588 ( .A(b[490]), .B(n567), .Z(c[490]) );
  XNOR U1589 ( .A(b[48]), .B(n568), .Z(c[48]) );
  XNOR U1590 ( .A(b[489]), .B(n569), .Z(c[489]) );
  XNOR U1591 ( .A(b[488]), .B(n570), .Z(c[488]) );
  XNOR U1592 ( .A(b[487]), .B(n571), .Z(c[487]) );
  XNOR U1593 ( .A(b[486]), .B(n572), .Z(c[486]) );
  XNOR U1594 ( .A(b[485]), .B(n573), .Z(c[485]) );
  XNOR U1595 ( .A(b[484]), .B(n574), .Z(c[484]) );
  XNOR U1596 ( .A(b[483]), .B(n575), .Z(c[483]) );
  XNOR U1597 ( .A(b[482]), .B(n576), .Z(c[482]) );
  XNOR U1598 ( .A(b[481]), .B(n577), .Z(c[481]) );
  XNOR U1599 ( .A(b[480]), .B(n578), .Z(c[480]) );
  XNOR U1600 ( .A(b[47]), .B(n579), .Z(c[47]) );
  XNOR U1601 ( .A(b[479]), .B(n580), .Z(c[479]) );
  XNOR U1602 ( .A(b[478]), .B(n581), .Z(c[478]) );
  XNOR U1603 ( .A(b[477]), .B(n582), .Z(c[477]) );
  XNOR U1604 ( .A(b[476]), .B(n583), .Z(c[476]) );
  XNOR U1605 ( .A(b[475]), .B(n584), .Z(c[475]) );
  XNOR U1606 ( .A(b[474]), .B(n585), .Z(c[474]) );
  XNOR U1607 ( .A(b[473]), .B(n586), .Z(c[473]) );
  XNOR U1608 ( .A(b[472]), .B(n587), .Z(c[472]) );
  XNOR U1609 ( .A(b[471]), .B(n588), .Z(c[471]) );
  XNOR U1610 ( .A(b[470]), .B(n589), .Z(c[470]) );
  XNOR U1611 ( .A(b[46]), .B(n590), .Z(c[46]) );
  XNOR U1612 ( .A(b[469]), .B(n591), .Z(c[469]) );
  XNOR U1613 ( .A(b[468]), .B(n592), .Z(c[468]) );
  XNOR U1614 ( .A(b[467]), .B(n593), .Z(c[467]) );
  XNOR U1615 ( .A(b[466]), .B(n594), .Z(c[466]) );
  XNOR U1616 ( .A(b[465]), .B(n595), .Z(c[465]) );
  XNOR U1617 ( .A(b[464]), .B(n596), .Z(c[464]) );
  XNOR U1618 ( .A(b[463]), .B(n597), .Z(c[463]) );
  XNOR U1619 ( .A(b[462]), .B(n598), .Z(c[462]) );
  XNOR U1620 ( .A(b[461]), .B(n599), .Z(c[461]) );
  XNOR U1621 ( .A(b[460]), .B(n600), .Z(c[460]) );
  XNOR U1622 ( .A(b[45]), .B(n601), .Z(c[45]) );
  XNOR U1623 ( .A(b[459]), .B(n602), .Z(c[459]) );
  XNOR U1624 ( .A(b[458]), .B(n603), .Z(c[458]) );
  XNOR U1625 ( .A(b[457]), .B(n604), .Z(c[457]) );
  XNOR U1626 ( .A(b[456]), .B(n605), .Z(c[456]) );
  XNOR U1627 ( .A(b[455]), .B(n606), .Z(c[455]) );
  XNOR U1628 ( .A(b[454]), .B(n607), .Z(c[454]) );
  XNOR U1629 ( .A(b[453]), .B(n608), .Z(c[453]) );
  XNOR U1630 ( .A(b[452]), .B(n609), .Z(c[452]) );
  XNOR U1631 ( .A(b[451]), .B(n610), .Z(c[451]) );
  XNOR U1632 ( .A(b[450]), .B(n611), .Z(c[450]) );
  XNOR U1633 ( .A(b[44]), .B(n612), .Z(c[44]) );
  XNOR U1634 ( .A(b[449]), .B(n613), .Z(c[449]) );
  XNOR U1635 ( .A(b[448]), .B(n614), .Z(c[448]) );
  XNOR U1636 ( .A(b[447]), .B(n615), .Z(c[447]) );
  XNOR U1637 ( .A(b[446]), .B(n616), .Z(c[446]) );
  XNOR U1638 ( .A(b[445]), .B(n617), .Z(c[445]) );
  XNOR U1639 ( .A(b[444]), .B(n618), .Z(c[444]) );
  XNOR U1640 ( .A(b[443]), .B(n619), .Z(c[443]) );
  XNOR U1641 ( .A(b[442]), .B(n620), .Z(c[442]) );
  XNOR U1642 ( .A(b[441]), .B(n621), .Z(c[441]) );
  XNOR U1643 ( .A(b[440]), .B(n622), .Z(c[440]) );
  XNOR U1644 ( .A(b[43]), .B(n623), .Z(c[43]) );
  XNOR U1645 ( .A(b[439]), .B(n624), .Z(c[439]) );
  XNOR U1646 ( .A(b[438]), .B(n625), .Z(c[438]) );
  XNOR U1647 ( .A(b[437]), .B(n626), .Z(c[437]) );
  XNOR U1648 ( .A(b[436]), .B(n627), .Z(c[436]) );
  XNOR U1649 ( .A(b[435]), .B(n628), .Z(c[435]) );
  XNOR U1650 ( .A(b[434]), .B(n629), .Z(c[434]) );
  XNOR U1651 ( .A(b[433]), .B(n630), .Z(c[433]) );
  XNOR U1652 ( .A(b[432]), .B(n631), .Z(c[432]) );
  XNOR U1653 ( .A(b[431]), .B(n632), .Z(c[431]) );
  XNOR U1654 ( .A(b[430]), .B(n633), .Z(c[430]) );
  XNOR U1655 ( .A(b[42]), .B(n634), .Z(c[42]) );
  XNOR U1656 ( .A(b[429]), .B(n635), .Z(c[429]) );
  XNOR U1657 ( .A(b[428]), .B(n636), .Z(c[428]) );
  XNOR U1658 ( .A(b[427]), .B(n637), .Z(c[427]) );
  XNOR U1659 ( .A(b[426]), .B(n638), .Z(c[426]) );
  XNOR U1660 ( .A(b[425]), .B(n639), .Z(c[425]) );
  XNOR U1661 ( .A(b[424]), .B(n640), .Z(c[424]) );
  XNOR U1662 ( .A(b[423]), .B(n641), .Z(c[423]) );
  XNOR U1663 ( .A(b[422]), .B(n642), .Z(c[422]) );
  XNOR U1664 ( .A(b[421]), .B(n643), .Z(c[421]) );
  XNOR U1665 ( .A(b[420]), .B(n644), .Z(c[420]) );
  XNOR U1666 ( .A(b[41]), .B(n645), .Z(c[41]) );
  XNOR U1667 ( .A(b[419]), .B(n646), .Z(c[419]) );
  XNOR U1668 ( .A(b[418]), .B(n647), .Z(c[418]) );
  XNOR U1669 ( .A(b[417]), .B(n648), .Z(c[417]) );
  XNOR U1670 ( .A(b[416]), .B(n649), .Z(c[416]) );
  XNOR U1671 ( .A(b[415]), .B(n650), .Z(c[415]) );
  XNOR U1672 ( .A(b[414]), .B(n651), .Z(c[414]) );
  XNOR U1673 ( .A(b[413]), .B(n652), .Z(c[413]) );
  XNOR U1674 ( .A(b[412]), .B(n653), .Z(c[412]) );
  XNOR U1675 ( .A(b[411]), .B(n654), .Z(c[411]) );
  XNOR U1676 ( .A(b[410]), .B(n655), .Z(c[410]) );
  XNOR U1677 ( .A(b[40]), .B(n656), .Z(c[40]) );
  XNOR U1678 ( .A(b[409]), .B(n657), .Z(c[409]) );
  XNOR U1679 ( .A(b[408]), .B(n658), .Z(c[408]) );
  XNOR U1680 ( .A(b[407]), .B(n659), .Z(c[407]) );
  XNOR U1681 ( .A(b[406]), .B(n660), .Z(c[406]) );
  XNOR U1682 ( .A(b[405]), .B(n661), .Z(c[405]) );
  XNOR U1683 ( .A(b[404]), .B(n662), .Z(c[404]) );
  XNOR U1684 ( .A(b[403]), .B(n663), .Z(c[403]) );
  XNOR U1685 ( .A(b[402]), .B(n664), .Z(c[402]) );
  XNOR U1686 ( .A(b[401]), .B(n665), .Z(c[401]) );
  XNOR U1687 ( .A(b[400]), .B(n666), .Z(c[400]) );
  XNOR U1688 ( .A(b[3]), .B(n667), .Z(c[3]) );
  XNOR U1689 ( .A(b[39]), .B(n668), .Z(c[39]) );
  XNOR U1690 ( .A(b[399]), .B(n669), .Z(c[399]) );
  XNOR U1691 ( .A(b[398]), .B(n670), .Z(c[398]) );
  XNOR U1692 ( .A(b[397]), .B(n671), .Z(c[397]) );
  XNOR U1693 ( .A(b[396]), .B(n672), .Z(c[396]) );
  XNOR U1694 ( .A(b[395]), .B(n673), .Z(c[395]) );
  XNOR U1695 ( .A(b[394]), .B(n674), .Z(c[394]) );
  XNOR U1696 ( .A(b[393]), .B(n675), .Z(c[393]) );
  XNOR U1697 ( .A(b[392]), .B(n676), .Z(c[392]) );
  XNOR U1698 ( .A(b[391]), .B(n677), .Z(c[391]) );
  XNOR U1699 ( .A(b[390]), .B(n678), .Z(c[390]) );
  XNOR U1700 ( .A(b[38]), .B(n679), .Z(c[38]) );
  XNOR U1701 ( .A(b[389]), .B(n680), .Z(c[389]) );
  XNOR U1702 ( .A(b[388]), .B(n681), .Z(c[388]) );
  XNOR U1703 ( .A(b[387]), .B(n682), .Z(c[387]) );
  XNOR U1704 ( .A(b[386]), .B(n683), .Z(c[386]) );
  XNOR U1705 ( .A(b[385]), .B(n684), .Z(c[385]) );
  XNOR U1706 ( .A(b[384]), .B(n685), .Z(c[384]) );
  XNOR U1707 ( .A(b[383]), .B(n686), .Z(c[383]) );
  XNOR U1708 ( .A(b[382]), .B(n687), .Z(c[382]) );
  XNOR U1709 ( .A(b[381]), .B(n688), .Z(c[381]) );
  XNOR U1710 ( .A(b[380]), .B(n689), .Z(c[380]) );
  XNOR U1711 ( .A(b[37]), .B(n690), .Z(c[37]) );
  XNOR U1712 ( .A(b[379]), .B(n691), .Z(c[379]) );
  XNOR U1713 ( .A(b[378]), .B(n692), .Z(c[378]) );
  XNOR U1714 ( .A(b[377]), .B(n693), .Z(c[377]) );
  XNOR U1715 ( .A(b[376]), .B(n694), .Z(c[376]) );
  XNOR U1716 ( .A(b[375]), .B(n695), .Z(c[375]) );
  XNOR U1717 ( .A(b[374]), .B(n696), .Z(c[374]) );
  XNOR U1718 ( .A(b[373]), .B(n697), .Z(c[373]) );
  XNOR U1719 ( .A(b[372]), .B(n698), .Z(c[372]) );
  XNOR U1720 ( .A(b[371]), .B(n699), .Z(c[371]) );
  XNOR U1721 ( .A(b[370]), .B(n700), .Z(c[370]) );
  XNOR U1722 ( .A(b[36]), .B(n701), .Z(c[36]) );
  XNOR U1723 ( .A(b[369]), .B(n702), .Z(c[369]) );
  XNOR U1724 ( .A(b[368]), .B(n703), .Z(c[368]) );
  XNOR U1725 ( .A(b[367]), .B(n704), .Z(c[367]) );
  XNOR U1726 ( .A(b[366]), .B(n705), .Z(c[366]) );
  XNOR U1727 ( .A(b[365]), .B(n706), .Z(c[365]) );
  XNOR U1728 ( .A(b[364]), .B(n707), .Z(c[364]) );
  XNOR U1729 ( .A(b[363]), .B(n708), .Z(c[363]) );
  XNOR U1730 ( .A(b[362]), .B(n709), .Z(c[362]) );
  XNOR U1731 ( .A(b[361]), .B(n710), .Z(c[361]) );
  XNOR U1732 ( .A(b[360]), .B(n711), .Z(c[360]) );
  XNOR U1733 ( .A(b[35]), .B(n712), .Z(c[35]) );
  XNOR U1734 ( .A(b[359]), .B(n713), .Z(c[359]) );
  XNOR U1735 ( .A(b[358]), .B(n714), .Z(c[358]) );
  XNOR U1736 ( .A(b[357]), .B(n715), .Z(c[357]) );
  XNOR U1737 ( .A(b[356]), .B(n716), .Z(c[356]) );
  XNOR U1738 ( .A(b[355]), .B(n717), .Z(c[355]) );
  XNOR U1739 ( .A(b[354]), .B(n718), .Z(c[354]) );
  XNOR U1740 ( .A(b[353]), .B(n719), .Z(c[353]) );
  XNOR U1741 ( .A(b[352]), .B(n720), .Z(c[352]) );
  XNOR U1742 ( .A(b[351]), .B(n721), .Z(c[351]) );
  XNOR U1743 ( .A(b[350]), .B(n722), .Z(c[350]) );
  XNOR U1744 ( .A(b[34]), .B(n723), .Z(c[34]) );
  XNOR U1745 ( .A(b[349]), .B(n724), .Z(c[349]) );
  XNOR U1746 ( .A(b[348]), .B(n725), .Z(c[348]) );
  XNOR U1747 ( .A(b[347]), .B(n726), .Z(c[347]) );
  XNOR U1748 ( .A(b[346]), .B(n727), .Z(c[346]) );
  XNOR U1749 ( .A(b[345]), .B(n728), .Z(c[345]) );
  XNOR U1750 ( .A(b[344]), .B(n729), .Z(c[344]) );
  XNOR U1751 ( .A(b[343]), .B(n730), .Z(c[343]) );
  XNOR U1752 ( .A(b[342]), .B(n731), .Z(c[342]) );
  XNOR U1753 ( .A(b[341]), .B(n732), .Z(c[341]) );
  XNOR U1754 ( .A(b[340]), .B(n733), .Z(c[340]) );
  XNOR U1755 ( .A(b[33]), .B(n734), .Z(c[33]) );
  XNOR U1756 ( .A(b[339]), .B(n735), .Z(c[339]) );
  XNOR U1757 ( .A(b[338]), .B(n736), .Z(c[338]) );
  XNOR U1758 ( .A(b[337]), .B(n737), .Z(c[337]) );
  XNOR U1759 ( .A(b[336]), .B(n738), .Z(c[336]) );
  XNOR U1760 ( .A(b[335]), .B(n739), .Z(c[335]) );
  XNOR U1761 ( .A(b[334]), .B(n740), .Z(c[334]) );
  XNOR U1762 ( .A(b[333]), .B(n741), .Z(c[333]) );
  XNOR U1763 ( .A(b[332]), .B(n742), .Z(c[332]) );
  XNOR U1764 ( .A(b[331]), .B(n743), .Z(c[331]) );
  XNOR U1765 ( .A(b[330]), .B(n744), .Z(c[330]) );
  XNOR U1766 ( .A(b[32]), .B(n745), .Z(c[32]) );
  XNOR U1767 ( .A(b[329]), .B(n746), .Z(c[329]) );
  XNOR U1768 ( .A(b[328]), .B(n747), .Z(c[328]) );
  XNOR U1769 ( .A(b[327]), .B(n748), .Z(c[327]) );
  XNOR U1770 ( .A(b[326]), .B(n749), .Z(c[326]) );
  XNOR U1771 ( .A(b[325]), .B(n750), .Z(c[325]) );
  XNOR U1772 ( .A(b[324]), .B(n751), .Z(c[324]) );
  XNOR U1773 ( .A(b[323]), .B(n752), .Z(c[323]) );
  XNOR U1774 ( .A(b[322]), .B(n753), .Z(c[322]) );
  XNOR U1775 ( .A(b[321]), .B(n754), .Z(c[321]) );
  XNOR U1776 ( .A(b[320]), .B(n755), .Z(c[320]) );
  XNOR U1777 ( .A(b[31]), .B(n756), .Z(c[31]) );
  XNOR U1778 ( .A(b[319]), .B(n757), .Z(c[319]) );
  XNOR U1779 ( .A(b[318]), .B(n758), .Z(c[318]) );
  XNOR U1780 ( .A(b[317]), .B(n759), .Z(c[317]) );
  XNOR U1781 ( .A(b[316]), .B(n760), .Z(c[316]) );
  XNOR U1782 ( .A(b[315]), .B(n761), .Z(c[315]) );
  XNOR U1783 ( .A(b[314]), .B(n762), .Z(c[314]) );
  XNOR U1784 ( .A(b[313]), .B(n763), .Z(c[313]) );
  XNOR U1785 ( .A(b[312]), .B(n764), .Z(c[312]) );
  XNOR U1786 ( .A(b[311]), .B(n765), .Z(c[311]) );
  XNOR U1787 ( .A(b[310]), .B(n766), .Z(c[310]) );
  XNOR U1788 ( .A(b[30]), .B(n767), .Z(c[30]) );
  XNOR U1789 ( .A(b[309]), .B(n768), .Z(c[309]) );
  XNOR U1790 ( .A(b[308]), .B(n769), .Z(c[308]) );
  XNOR U1791 ( .A(b[307]), .B(n770), .Z(c[307]) );
  XNOR U1792 ( .A(b[306]), .B(n771), .Z(c[306]) );
  XNOR U1793 ( .A(b[305]), .B(n772), .Z(c[305]) );
  XNOR U1794 ( .A(b[304]), .B(n773), .Z(c[304]) );
  XNOR U1795 ( .A(b[303]), .B(n774), .Z(c[303]) );
  XNOR U1796 ( .A(b[302]), .B(n775), .Z(c[302]) );
  XNOR U1797 ( .A(b[301]), .B(n776), .Z(c[301]) );
  XNOR U1798 ( .A(b[300]), .B(n777), .Z(c[300]) );
  XNOR U1799 ( .A(b[2]), .B(n778), .Z(c[2]) );
  XNOR U1800 ( .A(b[29]), .B(n779), .Z(c[29]) );
  XNOR U1801 ( .A(b[299]), .B(n780), .Z(c[299]) );
  XNOR U1802 ( .A(b[298]), .B(n781), .Z(c[298]) );
  XNOR U1803 ( .A(b[297]), .B(n782), .Z(c[297]) );
  XNOR U1804 ( .A(b[296]), .B(n783), .Z(c[296]) );
  XNOR U1805 ( .A(b[295]), .B(n784), .Z(c[295]) );
  XNOR U1806 ( .A(b[294]), .B(n785), .Z(c[294]) );
  XNOR U1807 ( .A(b[293]), .B(n786), .Z(c[293]) );
  XNOR U1808 ( .A(b[292]), .B(n787), .Z(c[292]) );
  XNOR U1809 ( .A(b[291]), .B(n788), .Z(c[291]) );
  XNOR U1810 ( .A(b[290]), .B(n789), .Z(c[290]) );
  XNOR U1811 ( .A(b[28]), .B(n790), .Z(c[28]) );
  XNOR U1812 ( .A(b[289]), .B(n791), .Z(c[289]) );
  XNOR U1813 ( .A(b[288]), .B(n792), .Z(c[288]) );
  XNOR U1814 ( .A(b[287]), .B(n793), .Z(c[287]) );
  XNOR U1815 ( .A(b[286]), .B(n794), .Z(c[286]) );
  XNOR U1816 ( .A(b[285]), .B(n795), .Z(c[285]) );
  XNOR U1817 ( .A(b[284]), .B(n796), .Z(c[284]) );
  XNOR U1818 ( .A(b[283]), .B(n797), .Z(c[283]) );
  XNOR U1819 ( .A(b[282]), .B(n798), .Z(c[282]) );
  XNOR U1820 ( .A(b[281]), .B(n799), .Z(c[281]) );
  XNOR U1821 ( .A(b[280]), .B(n800), .Z(c[280]) );
  XNOR U1822 ( .A(b[27]), .B(n801), .Z(c[27]) );
  XNOR U1823 ( .A(b[279]), .B(n802), .Z(c[279]) );
  XNOR U1824 ( .A(b[278]), .B(n803), .Z(c[278]) );
  XNOR U1825 ( .A(b[277]), .B(n804), .Z(c[277]) );
  XNOR U1826 ( .A(b[276]), .B(n805), .Z(c[276]) );
  XNOR U1827 ( .A(b[275]), .B(n806), .Z(c[275]) );
  XNOR U1828 ( .A(b[274]), .B(n807), .Z(c[274]) );
  XNOR U1829 ( .A(b[273]), .B(n808), .Z(c[273]) );
  XNOR U1830 ( .A(b[272]), .B(n809), .Z(c[272]) );
  XNOR U1831 ( .A(b[271]), .B(n810), .Z(c[271]) );
  XNOR U1832 ( .A(b[270]), .B(n811), .Z(c[270]) );
  XNOR U1833 ( .A(b[26]), .B(n812), .Z(c[26]) );
  XNOR U1834 ( .A(b[269]), .B(n813), .Z(c[269]) );
  XNOR U1835 ( .A(b[268]), .B(n814), .Z(c[268]) );
  XNOR U1836 ( .A(b[267]), .B(n815), .Z(c[267]) );
  XNOR U1837 ( .A(b[266]), .B(n816), .Z(c[266]) );
  XNOR U1838 ( .A(b[265]), .B(n817), .Z(c[265]) );
  XNOR U1839 ( .A(b[264]), .B(n818), .Z(c[264]) );
  XNOR U1840 ( .A(b[263]), .B(n819), .Z(c[263]) );
  XNOR U1841 ( .A(b[262]), .B(n820), .Z(c[262]) );
  XNOR U1842 ( .A(b[261]), .B(n821), .Z(c[261]) );
  XNOR U1843 ( .A(b[260]), .B(n822), .Z(c[260]) );
  XNOR U1844 ( .A(b[25]), .B(n823), .Z(c[25]) );
  XNOR U1845 ( .A(b[259]), .B(n824), .Z(c[259]) );
  XNOR U1846 ( .A(b[258]), .B(n825), .Z(c[258]) );
  XNOR U1847 ( .A(b[257]), .B(n826), .Z(c[257]) );
  XNOR U1848 ( .A(b[256]), .B(n827), .Z(c[256]) );
  XNOR U1849 ( .A(b[255]), .B(n828), .Z(c[255]) );
  XNOR U1850 ( .A(b[254]), .B(n829), .Z(c[254]) );
  XNOR U1851 ( .A(b[253]), .B(n830), .Z(c[253]) );
  XNOR U1852 ( .A(b[252]), .B(n831), .Z(c[252]) );
  XNOR U1853 ( .A(b[251]), .B(n832), .Z(c[251]) );
  XNOR U1854 ( .A(b[250]), .B(n833), .Z(c[250]) );
  XNOR U1855 ( .A(b[24]), .B(n834), .Z(c[24]) );
  XNOR U1856 ( .A(b[249]), .B(n835), .Z(c[249]) );
  XNOR U1857 ( .A(b[248]), .B(n836), .Z(c[248]) );
  XNOR U1858 ( .A(b[247]), .B(n837), .Z(c[247]) );
  XNOR U1859 ( .A(b[246]), .B(n838), .Z(c[246]) );
  XNOR U1860 ( .A(b[245]), .B(n839), .Z(c[245]) );
  XNOR U1861 ( .A(b[244]), .B(n840), .Z(c[244]) );
  XNOR U1862 ( .A(b[243]), .B(n841), .Z(c[243]) );
  XNOR U1863 ( .A(b[242]), .B(n842), .Z(c[242]) );
  XNOR U1864 ( .A(b[241]), .B(n843), .Z(c[241]) );
  XNOR U1865 ( .A(b[240]), .B(n844), .Z(c[240]) );
  XNOR U1866 ( .A(b[23]), .B(n845), .Z(c[23]) );
  XNOR U1867 ( .A(b[239]), .B(n846), .Z(c[239]) );
  XNOR U1868 ( .A(b[238]), .B(n847), .Z(c[238]) );
  XNOR U1869 ( .A(b[237]), .B(n848), .Z(c[237]) );
  XNOR U1870 ( .A(b[236]), .B(n849), .Z(c[236]) );
  XNOR U1871 ( .A(b[235]), .B(n850), .Z(c[235]) );
  XNOR U1872 ( .A(b[234]), .B(n851), .Z(c[234]) );
  XNOR U1873 ( .A(b[233]), .B(n852), .Z(c[233]) );
  XNOR U1874 ( .A(b[232]), .B(n853), .Z(c[232]) );
  XNOR U1875 ( .A(b[231]), .B(n854), .Z(c[231]) );
  XNOR U1876 ( .A(b[230]), .B(n855), .Z(c[230]) );
  XNOR U1877 ( .A(b[22]), .B(n856), .Z(c[22]) );
  XNOR U1878 ( .A(b[229]), .B(n857), .Z(c[229]) );
  XNOR U1879 ( .A(b[228]), .B(n858), .Z(c[228]) );
  XNOR U1880 ( .A(b[227]), .B(n859), .Z(c[227]) );
  XNOR U1881 ( .A(b[226]), .B(n860), .Z(c[226]) );
  XNOR U1882 ( .A(b[225]), .B(n861), .Z(c[225]) );
  XNOR U1883 ( .A(b[224]), .B(n862), .Z(c[224]) );
  XNOR U1884 ( .A(b[223]), .B(n863), .Z(c[223]) );
  XNOR U1885 ( .A(b[222]), .B(n864), .Z(c[222]) );
  XNOR U1886 ( .A(b[221]), .B(n865), .Z(c[221]) );
  XNOR U1887 ( .A(b[220]), .B(n866), .Z(c[220]) );
  XNOR U1888 ( .A(b[21]), .B(n867), .Z(c[21]) );
  XNOR U1889 ( .A(b[219]), .B(n868), .Z(c[219]) );
  XNOR U1890 ( .A(b[218]), .B(n869), .Z(c[218]) );
  XNOR U1891 ( .A(b[217]), .B(n870), .Z(c[217]) );
  XNOR U1892 ( .A(b[216]), .B(n871), .Z(c[216]) );
  XNOR U1893 ( .A(b[215]), .B(n872), .Z(c[215]) );
  XNOR U1894 ( .A(b[214]), .B(n873), .Z(c[214]) );
  XNOR U1895 ( .A(b[213]), .B(n874), .Z(c[213]) );
  XNOR U1896 ( .A(b[212]), .B(n875), .Z(c[212]) );
  XNOR U1897 ( .A(b[211]), .B(n876), .Z(c[211]) );
  XNOR U1898 ( .A(b[210]), .B(n877), .Z(c[210]) );
  XNOR U1899 ( .A(b[20]), .B(n878), .Z(c[20]) );
  XNOR U1900 ( .A(b[209]), .B(n879), .Z(c[209]) );
  XNOR U1901 ( .A(b[208]), .B(n880), .Z(c[208]) );
  XNOR U1902 ( .A(b[207]), .B(n881), .Z(c[207]) );
  XNOR U1903 ( .A(b[206]), .B(n882), .Z(c[206]) );
  XNOR U1904 ( .A(b[205]), .B(n883), .Z(c[205]) );
  XNOR U1905 ( .A(b[204]), .B(n884), .Z(c[204]) );
  XNOR U1906 ( .A(b[203]), .B(n885), .Z(c[203]) );
  XNOR U1907 ( .A(b[202]), .B(n886), .Z(c[202]) );
  XNOR U1908 ( .A(b[201]), .B(n887), .Z(c[201]) );
  XNOR U1909 ( .A(b[200]), .B(n888), .Z(c[200]) );
  XNOR U1910 ( .A(b[1]), .B(n889), .Z(c[1]) );
  XNOR U1911 ( .A(b[19]), .B(n890), .Z(c[19]) );
  XNOR U1912 ( .A(b[199]), .B(n891), .Z(c[199]) );
  XNOR U1913 ( .A(b[198]), .B(n892), .Z(c[198]) );
  XNOR U1914 ( .A(b[197]), .B(n893), .Z(c[197]) );
  XNOR U1915 ( .A(b[196]), .B(n894), .Z(c[196]) );
  XNOR U1916 ( .A(b[195]), .B(n895), .Z(c[195]) );
  XNOR U1917 ( .A(b[194]), .B(n896), .Z(c[194]) );
  XNOR U1918 ( .A(b[193]), .B(n897), .Z(c[193]) );
  XNOR U1919 ( .A(b[192]), .B(n898), .Z(c[192]) );
  XNOR U1920 ( .A(b[191]), .B(n899), .Z(c[191]) );
  XNOR U1921 ( .A(b[190]), .B(n900), .Z(c[190]) );
  XNOR U1922 ( .A(b[18]), .B(n901), .Z(c[18]) );
  XNOR U1923 ( .A(b[189]), .B(n902), .Z(c[189]) );
  XNOR U1924 ( .A(b[188]), .B(n903), .Z(c[188]) );
  XNOR U1925 ( .A(b[187]), .B(n904), .Z(c[187]) );
  XNOR U1926 ( .A(b[186]), .B(n905), .Z(c[186]) );
  XNOR U1927 ( .A(b[185]), .B(n906), .Z(c[185]) );
  XNOR U1928 ( .A(b[184]), .B(n907), .Z(c[184]) );
  XNOR U1929 ( .A(b[183]), .B(n908), .Z(c[183]) );
  XNOR U1930 ( .A(b[182]), .B(n909), .Z(c[182]) );
  XNOR U1931 ( .A(b[181]), .B(n910), .Z(c[181]) );
  XNOR U1932 ( .A(b[180]), .B(n911), .Z(c[180]) );
  XNOR U1933 ( .A(b[17]), .B(n912), .Z(c[17]) );
  XNOR U1934 ( .A(b[179]), .B(n913), .Z(c[179]) );
  XNOR U1935 ( .A(b[178]), .B(n914), .Z(c[178]) );
  XNOR U1936 ( .A(b[177]), .B(n915), .Z(c[177]) );
  XNOR U1937 ( .A(b[176]), .B(n916), .Z(c[176]) );
  XNOR U1938 ( .A(b[175]), .B(n917), .Z(c[175]) );
  XNOR U1939 ( .A(b[174]), .B(n918), .Z(c[174]) );
  XNOR U1940 ( .A(b[173]), .B(n919), .Z(c[173]) );
  XNOR U1941 ( .A(b[172]), .B(n920), .Z(c[172]) );
  XNOR U1942 ( .A(b[171]), .B(n921), .Z(c[171]) );
  XNOR U1943 ( .A(b[170]), .B(n922), .Z(c[170]) );
  XNOR U1944 ( .A(b[16]), .B(n923), .Z(c[16]) );
  XNOR U1945 ( .A(b[169]), .B(n924), .Z(c[169]) );
  XNOR U1946 ( .A(b[168]), .B(n925), .Z(c[168]) );
  XNOR U1947 ( .A(b[167]), .B(n926), .Z(c[167]) );
  XNOR U1948 ( .A(b[166]), .B(n927), .Z(c[166]) );
  XNOR U1949 ( .A(b[165]), .B(n928), .Z(c[165]) );
  XNOR U1950 ( .A(b[164]), .B(n929), .Z(c[164]) );
  XNOR U1951 ( .A(b[163]), .B(n930), .Z(c[163]) );
  XNOR U1952 ( .A(b[162]), .B(n931), .Z(c[162]) );
  XNOR U1953 ( .A(b[161]), .B(n932), .Z(c[161]) );
  XNOR U1954 ( .A(b[160]), .B(n933), .Z(c[160]) );
  XNOR U1955 ( .A(b[15]), .B(n934), .Z(c[15]) );
  XNOR U1956 ( .A(b[159]), .B(n935), .Z(c[159]) );
  XNOR U1957 ( .A(b[158]), .B(n936), .Z(c[158]) );
  XNOR U1958 ( .A(b[157]), .B(n937), .Z(c[157]) );
  XNOR U1959 ( .A(b[156]), .B(n938), .Z(c[156]) );
  XNOR U1960 ( .A(b[155]), .B(n939), .Z(c[155]) );
  XNOR U1961 ( .A(b[154]), .B(n940), .Z(c[154]) );
  XNOR U1962 ( .A(b[153]), .B(n941), .Z(c[153]) );
  XNOR U1963 ( .A(b[152]), .B(n942), .Z(c[152]) );
  XNOR U1964 ( .A(b[151]), .B(n943), .Z(c[151]) );
  XNOR U1965 ( .A(b[150]), .B(n944), .Z(c[150]) );
  XNOR U1966 ( .A(b[14]), .B(n945), .Z(c[14]) );
  XNOR U1967 ( .A(b[149]), .B(n946), .Z(c[149]) );
  XNOR U1968 ( .A(b[148]), .B(n947), .Z(c[148]) );
  XNOR U1969 ( .A(b[147]), .B(n948), .Z(c[147]) );
  XNOR U1970 ( .A(b[146]), .B(n949), .Z(c[146]) );
  XNOR U1971 ( .A(b[145]), .B(n950), .Z(c[145]) );
  XNOR U1972 ( .A(b[144]), .B(n951), .Z(c[144]) );
  XNOR U1973 ( .A(b[143]), .B(n952), .Z(c[143]) );
  XNOR U1974 ( .A(b[142]), .B(n953), .Z(c[142]) );
  XNOR U1975 ( .A(b[141]), .B(n954), .Z(c[141]) );
  XNOR U1976 ( .A(b[140]), .B(n955), .Z(c[140]) );
  XNOR U1977 ( .A(b[13]), .B(n956), .Z(c[13]) );
  XNOR U1978 ( .A(b[139]), .B(n957), .Z(c[139]) );
  XNOR U1979 ( .A(b[138]), .B(n958), .Z(c[138]) );
  XNOR U1980 ( .A(b[137]), .B(n959), .Z(c[137]) );
  XNOR U1981 ( .A(b[136]), .B(n960), .Z(c[136]) );
  XNOR U1982 ( .A(b[135]), .B(n961), .Z(c[135]) );
  XNOR U1983 ( .A(b[134]), .B(n962), .Z(c[134]) );
  XNOR U1984 ( .A(b[133]), .B(n963), .Z(c[133]) );
  XNOR U1985 ( .A(b[132]), .B(n964), .Z(c[132]) );
  XNOR U1986 ( .A(b[131]), .B(n965), .Z(c[131]) );
  XNOR U1987 ( .A(b[130]), .B(n966), .Z(c[130]) );
  XNOR U1988 ( .A(b[12]), .B(n967), .Z(c[12]) );
  XNOR U1989 ( .A(b[129]), .B(n968), .Z(c[129]) );
  XNOR U1990 ( .A(b[128]), .B(n969), .Z(c[128]) );
  XNOR U1991 ( .A(b[127]), .B(n970), .Z(c[127]) );
  XNOR U1992 ( .A(b[126]), .B(n971), .Z(c[126]) );
  XNOR U1993 ( .A(b[125]), .B(n972), .Z(c[125]) );
  XNOR U1994 ( .A(b[124]), .B(n973), .Z(c[124]) );
  XNOR U1995 ( .A(b[123]), .B(n974), .Z(c[123]) );
  XNOR U1996 ( .A(b[122]), .B(n975), .Z(c[122]) );
  XNOR U1997 ( .A(b[121]), .B(n976), .Z(c[121]) );
  XNOR U1998 ( .A(b[120]), .B(n977), .Z(c[120]) );
  XNOR U1999 ( .A(b[11]), .B(n978), .Z(c[11]) );
  XNOR U2000 ( .A(b[119]), .B(n979), .Z(c[119]) );
  XNOR U2001 ( .A(b[118]), .B(n980), .Z(c[118]) );
  XNOR U2002 ( .A(b[117]), .B(n981), .Z(c[117]) );
  XNOR U2003 ( .A(b[116]), .B(n982), .Z(c[116]) );
  XNOR U2004 ( .A(b[115]), .B(n983), .Z(c[115]) );
  XNOR U2005 ( .A(b[114]), .B(n984), .Z(c[114]) );
  XNOR U2006 ( .A(b[113]), .B(n985), .Z(c[113]) );
  XNOR U2007 ( .A(b[112]), .B(n986), .Z(c[112]) );
  XNOR U2008 ( .A(b[111]), .B(n987), .Z(c[111]) );
  XNOR U2009 ( .A(b[110]), .B(n988), .Z(c[110]) );
  XNOR U2010 ( .A(b[10]), .B(n989), .Z(c[10]) );
  XNOR U2011 ( .A(b[109]), .B(n990), .Z(c[109]) );
  XNOR U2012 ( .A(b[108]), .B(n991), .Z(c[108]) );
  XNOR U2013 ( .A(b[107]), .B(n992), .Z(c[107]) );
  XNOR U2014 ( .A(b[106]), .B(n993), .Z(c[106]) );
  XNOR U2015 ( .A(b[105]), .B(n994), .Z(c[105]) );
  XNOR U2016 ( .A(b[104]), .B(n995), .Z(c[104]) );
  XNOR U2017 ( .A(b[103]), .B(n996), .Z(c[103]) );
  XNOR U2018 ( .A(b[102]), .B(n997), .Z(c[102]) );
  XOR U2019 ( .A(n998), .B(n999), .Z(c[1023]) );
  XOR U2020 ( .A(n1000), .B(n1001), .Z(n999) );
  ANDN U2021 ( .B(n1002), .A(n1003), .Z(n1000) );
  XOR U2022 ( .A(b[1022]), .B(n1001), .Z(n1002) );
  XOR U2023 ( .A(b[1023]), .B(a[1023]), .Z(n998) );
  XNOR U2024 ( .A(b[1022]), .B(n1003), .Z(c[1022]) );
  XNOR U2025 ( .A(a[1022]), .B(n1001), .Z(n1003) );
  XOR U2026 ( .A(n1004), .B(n1005), .Z(n1001) );
  ANDN U2027 ( .B(n1006), .A(n1007), .Z(n1004) );
  XOR U2028 ( .A(b[1021]), .B(n1005), .Z(n1006) );
  XNOR U2029 ( .A(b[1021]), .B(n1007), .Z(c[1021]) );
  XOR U2030 ( .A(n1008), .B(n1009), .Z(n1005) );
  ANDN U2031 ( .B(n1010), .A(n1011), .Z(n1008) );
  XOR U2032 ( .A(b[1020]), .B(n1009), .Z(n1010) );
  XNOR U2033 ( .A(b[1020]), .B(n1011), .Z(c[1020]) );
  XOR U2034 ( .A(n1012), .B(n1013), .Z(n1009) );
  ANDN U2035 ( .B(n1014), .A(n1015), .Z(n1012) );
  XOR U2036 ( .A(b[1019]), .B(n1013), .Z(n1014) );
  XNOR U2037 ( .A(b[101]), .B(n1016), .Z(c[101]) );
  XNOR U2038 ( .A(b[1019]), .B(n1015), .Z(c[1019]) );
  XOR U2039 ( .A(n1017), .B(n1018), .Z(n1013) );
  ANDN U2040 ( .B(n1019), .A(n1020), .Z(n1017) );
  XOR U2041 ( .A(b[1018]), .B(n1018), .Z(n1019) );
  XNOR U2042 ( .A(b[1018]), .B(n1020), .Z(c[1018]) );
  XOR U2043 ( .A(n1021), .B(n1022), .Z(n1018) );
  ANDN U2044 ( .B(n1023), .A(n1024), .Z(n1021) );
  XOR U2045 ( .A(b[1017]), .B(n1022), .Z(n1023) );
  XNOR U2046 ( .A(b[1017]), .B(n1024), .Z(c[1017]) );
  XOR U2047 ( .A(n1025), .B(n1026), .Z(n1022) );
  ANDN U2048 ( .B(n1027), .A(n1028), .Z(n1025) );
  XOR U2049 ( .A(b[1016]), .B(n1026), .Z(n1027) );
  XNOR U2050 ( .A(b[1016]), .B(n1028), .Z(c[1016]) );
  XOR U2051 ( .A(n1029), .B(n1030), .Z(n1026) );
  ANDN U2052 ( .B(n1031), .A(n1032), .Z(n1029) );
  XOR U2053 ( .A(b[1015]), .B(n1030), .Z(n1031) );
  XNOR U2054 ( .A(b[1015]), .B(n1032), .Z(c[1015]) );
  XOR U2055 ( .A(n1033), .B(n1034), .Z(n1030) );
  ANDN U2056 ( .B(n1035), .A(n1036), .Z(n1033) );
  XOR U2057 ( .A(b[1014]), .B(n1034), .Z(n1035) );
  XNOR U2058 ( .A(b[1014]), .B(n1036), .Z(c[1014]) );
  XOR U2059 ( .A(n1037), .B(n1038), .Z(n1034) );
  ANDN U2060 ( .B(n1039), .A(n1040), .Z(n1037) );
  XOR U2061 ( .A(b[1013]), .B(n1038), .Z(n1039) );
  XNOR U2062 ( .A(b[1013]), .B(n1040), .Z(c[1013]) );
  XOR U2063 ( .A(n1041), .B(n1042), .Z(n1038) );
  ANDN U2064 ( .B(n1043), .A(n1044), .Z(n1041) );
  XOR U2065 ( .A(b[1012]), .B(n1042), .Z(n1043) );
  XNOR U2066 ( .A(b[1012]), .B(n1044), .Z(c[1012]) );
  XOR U2067 ( .A(n1045), .B(n1046), .Z(n1042) );
  ANDN U2068 ( .B(n1047), .A(n1048), .Z(n1045) );
  XOR U2069 ( .A(b[1011]), .B(n1046), .Z(n1047) );
  XNOR U2070 ( .A(b[1011]), .B(n1048), .Z(c[1011]) );
  XOR U2071 ( .A(n1049), .B(n1050), .Z(n1046) );
  ANDN U2072 ( .B(n1051), .A(n1052), .Z(n1049) );
  XOR U2073 ( .A(b[1010]), .B(n1050), .Z(n1051) );
  XNOR U2074 ( .A(b[1010]), .B(n1052), .Z(c[1010]) );
  XOR U2075 ( .A(n1053), .B(n1054), .Z(n1050) );
  ANDN U2076 ( .B(n1055), .A(n1056), .Z(n1053) );
  XOR U2077 ( .A(b[1009]), .B(n1054), .Z(n1055) );
  XNOR U2078 ( .A(b[100]), .B(n1057), .Z(c[100]) );
  XNOR U2079 ( .A(b[1009]), .B(n1056), .Z(c[1009]) );
  XOR U2080 ( .A(n1058), .B(n1059), .Z(n1054) );
  ANDN U2081 ( .B(n1060), .A(n1061), .Z(n1058) );
  XOR U2082 ( .A(b[1008]), .B(n1059), .Z(n1060) );
  XNOR U2083 ( .A(b[1008]), .B(n1061), .Z(c[1008]) );
  XOR U2084 ( .A(n1062), .B(n1063), .Z(n1059) );
  ANDN U2085 ( .B(n1064), .A(n1065), .Z(n1062) );
  XOR U2086 ( .A(b[1007]), .B(n1063), .Z(n1064) );
  XNOR U2087 ( .A(b[1007]), .B(n1065), .Z(c[1007]) );
  XOR U2088 ( .A(n1066), .B(n1067), .Z(n1063) );
  ANDN U2089 ( .B(n1068), .A(n1069), .Z(n1066) );
  XOR U2090 ( .A(b[1006]), .B(n1067), .Z(n1068) );
  XNOR U2091 ( .A(b[1006]), .B(n1069), .Z(c[1006]) );
  XOR U2092 ( .A(n1070), .B(n1071), .Z(n1067) );
  ANDN U2093 ( .B(n1072), .A(n1073), .Z(n1070) );
  XOR U2094 ( .A(b[1005]), .B(n1071), .Z(n1072) );
  XNOR U2095 ( .A(b[1005]), .B(n1073), .Z(c[1005]) );
  XOR U2096 ( .A(n1074), .B(n1075), .Z(n1071) );
  ANDN U2097 ( .B(n1076), .A(n1077), .Z(n1074) );
  XOR U2098 ( .A(b[1004]), .B(n1075), .Z(n1076) );
  XNOR U2099 ( .A(b[1004]), .B(n1077), .Z(c[1004]) );
  XOR U2100 ( .A(n1078), .B(n1079), .Z(n1075) );
  ANDN U2101 ( .B(n1080), .A(n1081), .Z(n1078) );
  XOR U2102 ( .A(b[1003]), .B(n1079), .Z(n1080) );
  XNOR U2103 ( .A(b[1003]), .B(n1081), .Z(c[1003]) );
  XOR U2104 ( .A(n1082), .B(n1083), .Z(n1079) );
  ANDN U2105 ( .B(n1084), .A(n1085), .Z(n1082) );
  XOR U2106 ( .A(b[1002]), .B(n1083), .Z(n1084) );
  XNOR U2107 ( .A(b[1002]), .B(n1085), .Z(c[1002]) );
  XOR U2108 ( .A(n1086), .B(n1087), .Z(n1083) );
  ANDN U2109 ( .B(n1088), .A(n1089), .Z(n1086) );
  XOR U2110 ( .A(b[1001]), .B(n1087), .Z(n1088) );
  XNOR U2111 ( .A(b[1001]), .B(n1089), .Z(c[1001]) );
  XOR U2112 ( .A(n1090), .B(n1091), .Z(n1087) );
  ANDN U2113 ( .B(n1092), .A(n1093), .Z(n1090) );
  XOR U2114 ( .A(b[1000]), .B(n1091), .Z(n1092) );
  XNOR U2115 ( .A(b[1000]), .B(n1093), .Z(c[1000]) );
  XOR U2116 ( .A(n1094), .B(n1095), .Z(n1091) );
  ANDN U2117 ( .B(n1096), .A(n3), .Z(n1094) );
  XOR U2118 ( .A(b[999]), .B(n1095), .Z(n1096) );
  XOR U2119 ( .A(n1097), .B(n1098), .Z(n1095) );
  ANDN U2120 ( .B(n1099), .A(n4), .Z(n1097) );
  XOR U2121 ( .A(b[998]), .B(n1098), .Z(n1099) );
  XOR U2122 ( .A(n1100), .B(n1101), .Z(n1098) );
  ANDN U2123 ( .B(n1102), .A(n5), .Z(n1100) );
  XOR U2124 ( .A(b[997]), .B(n1101), .Z(n1102) );
  XOR U2125 ( .A(n1103), .B(n1104), .Z(n1101) );
  ANDN U2126 ( .B(n1105), .A(n6), .Z(n1103) );
  XOR U2127 ( .A(b[996]), .B(n1104), .Z(n1105) );
  XOR U2128 ( .A(n1106), .B(n1107), .Z(n1104) );
  ANDN U2129 ( .B(n1108), .A(n7), .Z(n1106) );
  XOR U2130 ( .A(b[995]), .B(n1107), .Z(n1108) );
  XOR U2131 ( .A(n1109), .B(n1110), .Z(n1107) );
  ANDN U2132 ( .B(n1111), .A(n8), .Z(n1109) );
  XOR U2133 ( .A(b[994]), .B(n1110), .Z(n1111) );
  XOR U2134 ( .A(n1112), .B(n1113), .Z(n1110) );
  ANDN U2135 ( .B(n1114), .A(n9), .Z(n1112) );
  XOR U2136 ( .A(b[993]), .B(n1113), .Z(n1114) );
  XOR U2137 ( .A(n1115), .B(n1116), .Z(n1113) );
  ANDN U2138 ( .B(n1117), .A(n10), .Z(n1115) );
  XOR U2139 ( .A(b[992]), .B(n1116), .Z(n1117) );
  XOR U2140 ( .A(n1118), .B(n1119), .Z(n1116) );
  ANDN U2141 ( .B(n1120), .A(n11), .Z(n1118) );
  XOR U2142 ( .A(b[991]), .B(n1119), .Z(n1120) );
  XOR U2143 ( .A(n1121), .B(n1122), .Z(n1119) );
  ANDN U2144 ( .B(n1123), .A(n12), .Z(n1121) );
  XOR U2145 ( .A(b[990]), .B(n1122), .Z(n1123) );
  XOR U2146 ( .A(n1124), .B(n1125), .Z(n1122) );
  ANDN U2147 ( .B(n1126), .A(n14), .Z(n1124) );
  XOR U2148 ( .A(b[989]), .B(n1125), .Z(n1126) );
  XOR U2149 ( .A(n1127), .B(n1128), .Z(n1125) );
  ANDN U2150 ( .B(n1129), .A(n15), .Z(n1127) );
  XOR U2151 ( .A(b[988]), .B(n1128), .Z(n1129) );
  XOR U2152 ( .A(n1130), .B(n1131), .Z(n1128) );
  ANDN U2153 ( .B(n1132), .A(n16), .Z(n1130) );
  XOR U2154 ( .A(b[987]), .B(n1131), .Z(n1132) );
  XOR U2155 ( .A(n1133), .B(n1134), .Z(n1131) );
  ANDN U2156 ( .B(n1135), .A(n17), .Z(n1133) );
  XOR U2157 ( .A(b[986]), .B(n1134), .Z(n1135) );
  XOR U2158 ( .A(n1136), .B(n1137), .Z(n1134) );
  ANDN U2159 ( .B(n1138), .A(n18), .Z(n1136) );
  XOR U2160 ( .A(b[985]), .B(n1137), .Z(n1138) );
  XOR U2161 ( .A(n1139), .B(n1140), .Z(n1137) );
  ANDN U2162 ( .B(n1141), .A(n19), .Z(n1139) );
  XOR U2163 ( .A(b[984]), .B(n1140), .Z(n1141) );
  XOR U2164 ( .A(n1142), .B(n1143), .Z(n1140) );
  ANDN U2165 ( .B(n1144), .A(n20), .Z(n1142) );
  XOR U2166 ( .A(b[983]), .B(n1143), .Z(n1144) );
  XOR U2167 ( .A(n1145), .B(n1146), .Z(n1143) );
  ANDN U2168 ( .B(n1147), .A(n21), .Z(n1145) );
  XOR U2169 ( .A(b[982]), .B(n1146), .Z(n1147) );
  XOR U2170 ( .A(n1148), .B(n1149), .Z(n1146) );
  ANDN U2171 ( .B(n1150), .A(n22), .Z(n1148) );
  XOR U2172 ( .A(b[981]), .B(n1149), .Z(n1150) );
  XOR U2173 ( .A(n1151), .B(n1152), .Z(n1149) );
  ANDN U2174 ( .B(n1153), .A(n23), .Z(n1151) );
  XOR U2175 ( .A(b[980]), .B(n1152), .Z(n1153) );
  XOR U2176 ( .A(n1154), .B(n1155), .Z(n1152) );
  ANDN U2177 ( .B(n1156), .A(n25), .Z(n1154) );
  XOR U2178 ( .A(b[979]), .B(n1155), .Z(n1156) );
  XOR U2179 ( .A(n1157), .B(n1158), .Z(n1155) );
  ANDN U2180 ( .B(n1159), .A(n26), .Z(n1157) );
  XOR U2181 ( .A(b[978]), .B(n1158), .Z(n1159) );
  XOR U2182 ( .A(n1160), .B(n1161), .Z(n1158) );
  ANDN U2183 ( .B(n1162), .A(n27), .Z(n1160) );
  XOR U2184 ( .A(b[977]), .B(n1161), .Z(n1162) );
  XOR U2185 ( .A(n1163), .B(n1164), .Z(n1161) );
  ANDN U2186 ( .B(n1165), .A(n28), .Z(n1163) );
  XOR U2187 ( .A(b[976]), .B(n1164), .Z(n1165) );
  XOR U2188 ( .A(n1166), .B(n1167), .Z(n1164) );
  ANDN U2189 ( .B(n1168), .A(n29), .Z(n1166) );
  XOR U2190 ( .A(b[975]), .B(n1167), .Z(n1168) );
  XOR U2191 ( .A(n1169), .B(n1170), .Z(n1167) );
  ANDN U2192 ( .B(n1171), .A(n30), .Z(n1169) );
  XOR U2193 ( .A(b[974]), .B(n1170), .Z(n1171) );
  XOR U2194 ( .A(n1172), .B(n1173), .Z(n1170) );
  ANDN U2195 ( .B(n1174), .A(n31), .Z(n1172) );
  XOR U2196 ( .A(b[973]), .B(n1173), .Z(n1174) );
  XOR U2197 ( .A(n1175), .B(n1176), .Z(n1173) );
  ANDN U2198 ( .B(n1177), .A(n32), .Z(n1175) );
  XOR U2199 ( .A(b[972]), .B(n1176), .Z(n1177) );
  XOR U2200 ( .A(n1178), .B(n1179), .Z(n1176) );
  ANDN U2201 ( .B(n1180), .A(n33), .Z(n1178) );
  XOR U2202 ( .A(b[971]), .B(n1179), .Z(n1180) );
  XOR U2203 ( .A(n1181), .B(n1182), .Z(n1179) );
  ANDN U2204 ( .B(n1183), .A(n34), .Z(n1181) );
  XOR U2205 ( .A(b[970]), .B(n1182), .Z(n1183) );
  XOR U2206 ( .A(n1184), .B(n1185), .Z(n1182) );
  ANDN U2207 ( .B(n1186), .A(n36), .Z(n1184) );
  XOR U2208 ( .A(b[969]), .B(n1185), .Z(n1186) );
  XOR U2209 ( .A(n1187), .B(n1188), .Z(n1185) );
  ANDN U2210 ( .B(n1189), .A(n37), .Z(n1187) );
  XOR U2211 ( .A(b[968]), .B(n1188), .Z(n1189) );
  XOR U2212 ( .A(n1190), .B(n1191), .Z(n1188) );
  ANDN U2213 ( .B(n1192), .A(n38), .Z(n1190) );
  XOR U2214 ( .A(b[967]), .B(n1191), .Z(n1192) );
  XOR U2215 ( .A(n1193), .B(n1194), .Z(n1191) );
  ANDN U2216 ( .B(n1195), .A(n39), .Z(n1193) );
  XOR U2217 ( .A(b[966]), .B(n1194), .Z(n1195) );
  XOR U2218 ( .A(n1196), .B(n1197), .Z(n1194) );
  ANDN U2219 ( .B(n1198), .A(n40), .Z(n1196) );
  XOR U2220 ( .A(b[965]), .B(n1197), .Z(n1198) );
  XOR U2221 ( .A(n1199), .B(n1200), .Z(n1197) );
  ANDN U2222 ( .B(n1201), .A(n41), .Z(n1199) );
  XOR U2223 ( .A(b[964]), .B(n1200), .Z(n1201) );
  XOR U2224 ( .A(n1202), .B(n1203), .Z(n1200) );
  ANDN U2225 ( .B(n1204), .A(n42), .Z(n1202) );
  XOR U2226 ( .A(b[963]), .B(n1203), .Z(n1204) );
  XOR U2227 ( .A(n1205), .B(n1206), .Z(n1203) );
  ANDN U2228 ( .B(n1207), .A(n43), .Z(n1205) );
  XOR U2229 ( .A(b[962]), .B(n1206), .Z(n1207) );
  XOR U2230 ( .A(n1208), .B(n1209), .Z(n1206) );
  ANDN U2231 ( .B(n1210), .A(n44), .Z(n1208) );
  XOR U2232 ( .A(b[961]), .B(n1209), .Z(n1210) );
  XOR U2233 ( .A(n1211), .B(n1212), .Z(n1209) );
  ANDN U2234 ( .B(n1213), .A(n45), .Z(n1211) );
  XOR U2235 ( .A(b[960]), .B(n1212), .Z(n1213) );
  XOR U2236 ( .A(n1214), .B(n1215), .Z(n1212) );
  ANDN U2237 ( .B(n1216), .A(n47), .Z(n1214) );
  XOR U2238 ( .A(b[959]), .B(n1215), .Z(n1216) );
  XOR U2239 ( .A(n1217), .B(n1218), .Z(n1215) );
  ANDN U2240 ( .B(n1219), .A(n48), .Z(n1217) );
  XOR U2241 ( .A(b[958]), .B(n1218), .Z(n1219) );
  XOR U2242 ( .A(n1220), .B(n1221), .Z(n1218) );
  ANDN U2243 ( .B(n1222), .A(n49), .Z(n1220) );
  XOR U2244 ( .A(b[957]), .B(n1221), .Z(n1222) );
  XOR U2245 ( .A(n1223), .B(n1224), .Z(n1221) );
  ANDN U2246 ( .B(n1225), .A(n50), .Z(n1223) );
  XOR U2247 ( .A(b[956]), .B(n1224), .Z(n1225) );
  XOR U2248 ( .A(n1226), .B(n1227), .Z(n1224) );
  ANDN U2249 ( .B(n1228), .A(n51), .Z(n1226) );
  XOR U2250 ( .A(b[955]), .B(n1227), .Z(n1228) );
  XOR U2251 ( .A(n1229), .B(n1230), .Z(n1227) );
  ANDN U2252 ( .B(n1231), .A(n52), .Z(n1229) );
  XOR U2253 ( .A(b[954]), .B(n1230), .Z(n1231) );
  XOR U2254 ( .A(n1232), .B(n1233), .Z(n1230) );
  ANDN U2255 ( .B(n1234), .A(n53), .Z(n1232) );
  XOR U2256 ( .A(b[953]), .B(n1233), .Z(n1234) );
  XOR U2257 ( .A(n1235), .B(n1236), .Z(n1233) );
  ANDN U2258 ( .B(n1237), .A(n54), .Z(n1235) );
  XOR U2259 ( .A(b[952]), .B(n1236), .Z(n1237) );
  XOR U2260 ( .A(n1238), .B(n1239), .Z(n1236) );
  ANDN U2261 ( .B(n1240), .A(n55), .Z(n1238) );
  XOR U2262 ( .A(b[951]), .B(n1239), .Z(n1240) );
  XOR U2263 ( .A(n1241), .B(n1242), .Z(n1239) );
  ANDN U2264 ( .B(n1243), .A(n56), .Z(n1241) );
  XOR U2265 ( .A(b[950]), .B(n1242), .Z(n1243) );
  XOR U2266 ( .A(n1244), .B(n1245), .Z(n1242) );
  ANDN U2267 ( .B(n1246), .A(n58), .Z(n1244) );
  XOR U2268 ( .A(b[949]), .B(n1245), .Z(n1246) );
  XOR U2269 ( .A(n1247), .B(n1248), .Z(n1245) );
  ANDN U2270 ( .B(n1249), .A(n59), .Z(n1247) );
  XOR U2271 ( .A(b[948]), .B(n1248), .Z(n1249) );
  XOR U2272 ( .A(n1250), .B(n1251), .Z(n1248) );
  ANDN U2273 ( .B(n1252), .A(n60), .Z(n1250) );
  XOR U2274 ( .A(b[947]), .B(n1251), .Z(n1252) );
  XOR U2275 ( .A(n1253), .B(n1254), .Z(n1251) );
  ANDN U2276 ( .B(n1255), .A(n61), .Z(n1253) );
  XOR U2277 ( .A(b[946]), .B(n1254), .Z(n1255) );
  XOR U2278 ( .A(n1256), .B(n1257), .Z(n1254) );
  ANDN U2279 ( .B(n1258), .A(n62), .Z(n1256) );
  XOR U2280 ( .A(b[945]), .B(n1257), .Z(n1258) );
  XOR U2281 ( .A(n1259), .B(n1260), .Z(n1257) );
  ANDN U2282 ( .B(n1261), .A(n63), .Z(n1259) );
  XOR U2283 ( .A(b[944]), .B(n1260), .Z(n1261) );
  XOR U2284 ( .A(n1262), .B(n1263), .Z(n1260) );
  ANDN U2285 ( .B(n1264), .A(n64), .Z(n1262) );
  XOR U2286 ( .A(b[943]), .B(n1263), .Z(n1264) );
  XOR U2287 ( .A(n1265), .B(n1266), .Z(n1263) );
  ANDN U2288 ( .B(n1267), .A(n65), .Z(n1265) );
  XOR U2289 ( .A(b[942]), .B(n1266), .Z(n1267) );
  XOR U2290 ( .A(n1268), .B(n1269), .Z(n1266) );
  ANDN U2291 ( .B(n1270), .A(n66), .Z(n1268) );
  XOR U2292 ( .A(b[941]), .B(n1269), .Z(n1270) );
  XOR U2293 ( .A(n1271), .B(n1272), .Z(n1269) );
  ANDN U2294 ( .B(n1273), .A(n67), .Z(n1271) );
  XOR U2295 ( .A(b[940]), .B(n1272), .Z(n1273) );
  XOR U2296 ( .A(n1274), .B(n1275), .Z(n1272) );
  ANDN U2297 ( .B(n1276), .A(n69), .Z(n1274) );
  XOR U2298 ( .A(b[939]), .B(n1275), .Z(n1276) );
  XOR U2299 ( .A(n1277), .B(n1278), .Z(n1275) );
  ANDN U2300 ( .B(n1279), .A(n70), .Z(n1277) );
  XOR U2301 ( .A(b[938]), .B(n1278), .Z(n1279) );
  XOR U2302 ( .A(n1280), .B(n1281), .Z(n1278) );
  ANDN U2303 ( .B(n1282), .A(n71), .Z(n1280) );
  XOR U2304 ( .A(b[937]), .B(n1281), .Z(n1282) );
  XOR U2305 ( .A(n1283), .B(n1284), .Z(n1281) );
  ANDN U2306 ( .B(n1285), .A(n72), .Z(n1283) );
  XOR U2307 ( .A(b[936]), .B(n1284), .Z(n1285) );
  XOR U2308 ( .A(n1286), .B(n1287), .Z(n1284) );
  ANDN U2309 ( .B(n1288), .A(n73), .Z(n1286) );
  XOR U2310 ( .A(b[935]), .B(n1287), .Z(n1288) );
  XOR U2311 ( .A(n1289), .B(n1290), .Z(n1287) );
  ANDN U2312 ( .B(n1291), .A(n74), .Z(n1289) );
  XOR U2313 ( .A(b[934]), .B(n1290), .Z(n1291) );
  XOR U2314 ( .A(n1292), .B(n1293), .Z(n1290) );
  ANDN U2315 ( .B(n1294), .A(n75), .Z(n1292) );
  XOR U2316 ( .A(b[933]), .B(n1293), .Z(n1294) );
  XOR U2317 ( .A(n1295), .B(n1296), .Z(n1293) );
  ANDN U2318 ( .B(n1297), .A(n76), .Z(n1295) );
  XOR U2319 ( .A(b[932]), .B(n1296), .Z(n1297) );
  XOR U2320 ( .A(n1298), .B(n1299), .Z(n1296) );
  ANDN U2321 ( .B(n1300), .A(n77), .Z(n1298) );
  XOR U2322 ( .A(b[931]), .B(n1299), .Z(n1300) );
  XOR U2323 ( .A(n1301), .B(n1302), .Z(n1299) );
  ANDN U2324 ( .B(n1303), .A(n78), .Z(n1301) );
  XOR U2325 ( .A(b[930]), .B(n1302), .Z(n1303) );
  XOR U2326 ( .A(n1304), .B(n1305), .Z(n1302) );
  ANDN U2327 ( .B(n1306), .A(n80), .Z(n1304) );
  XOR U2328 ( .A(b[929]), .B(n1305), .Z(n1306) );
  XOR U2329 ( .A(n1307), .B(n1308), .Z(n1305) );
  ANDN U2330 ( .B(n1309), .A(n81), .Z(n1307) );
  XOR U2331 ( .A(b[928]), .B(n1308), .Z(n1309) );
  XOR U2332 ( .A(n1310), .B(n1311), .Z(n1308) );
  ANDN U2333 ( .B(n1312), .A(n82), .Z(n1310) );
  XOR U2334 ( .A(b[927]), .B(n1311), .Z(n1312) );
  XOR U2335 ( .A(n1313), .B(n1314), .Z(n1311) );
  ANDN U2336 ( .B(n1315), .A(n83), .Z(n1313) );
  XOR U2337 ( .A(b[926]), .B(n1314), .Z(n1315) );
  XOR U2338 ( .A(n1316), .B(n1317), .Z(n1314) );
  ANDN U2339 ( .B(n1318), .A(n84), .Z(n1316) );
  XOR U2340 ( .A(b[925]), .B(n1317), .Z(n1318) );
  XOR U2341 ( .A(n1319), .B(n1320), .Z(n1317) );
  ANDN U2342 ( .B(n1321), .A(n85), .Z(n1319) );
  XOR U2343 ( .A(b[924]), .B(n1320), .Z(n1321) );
  XOR U2344 ( .A(n1322), .B(n1323), .Z(n1320) );
  ANDN U2345 ( .B(n1324), .A(n86), .Z(n1322) );
  XOR U2346 ( .A(b[923]), .B(n1323), .Z(n1324) );
  XOR U2347 ( .A(n1325), .B(n1326), .Z(n1323) );
  ANDN U2348 ( .B(n1327), .A(n87), .Z(n1325) );
  XOR U2349 ( .A(b[922]), .B(n1326), .Z(n1327) );
  XOR U2350 ( .A(n1328), .B(n1329), .Z(n1326) );
  ANDN U2351 ( .B(n1330), .A(n88), .Z(n1328) );
  XOR U2352 ( .A(b[921]), .B(n1329), .Z(n1330) );
  XOR U2353 ( .A(n1331), .B(n1332), .Z(n1329) );
  ANDN U2354 ( .B(n1333), .A(n89), .Z(n1331) );
  XOR U2355 ( .A(b[920]), .B(n1332), .Z(n1333) );
  XOR U2356 ( .A(n1334), .B(n1335), .Z(n1332) );
  ANDN U2357 ( .B(n1336), .A(n91), .Z(n1334) );
  XOR U2358 ( .A(b[919]), .B(n1335), .Z(n1336) );
  XOR U2359 ( .A(n1337), .B(n1338), .Z(n1335) );
  ANDN U2360 ( .B(n1339), .A(n92), .Z(n1337) );
  XOR U2361 ( .A(b[918]), .B(n1338), .Z(n1339) );
  XOR U2362 ( .A(n1340), .B(n1341), .Z(n1338) );
  ANDN U2363 ( .B(n1342), .A(n93), .Z(n1340) );
  XOR U2364 ( .A(b[917]), .B(n1341), .Z(n1342) );
  XOR U2365 ( .A(n1343), .B(n1344), .Z(n1341) );
  ANDN U2366 ( .B(n1345), .A(n94), .Z(n1343) );
  XOR U2367 ( .A(b[916]), .B(n1344), .Z(n1345) );
  XOR U2368 ( .A(n1346), .B(n1347), .Z(n1344) );
  ANDN U2369 ( .B(n1348), .A(n95), .Z(n1346) );
  XOR U2370 ( .A(b[915]), .B(n1347), .Z(n1348) );
  XOR U2371 ( .A(n1349), .B(n1350), .Z(n1347) );
  ANDN U2372 ( .B(n1351), .A(n96), .Z(n1349) );
  XOR U2373 ( .A(b[914]), .B(n1350), .Z(n1351) );
  XOR U2374 ( .A(n1352), .B(n1353), .Z(n1350) );
  ANDN U2375 ( .B(n1354), .A(n97), .Z(n1352) );
  XOR U2376 ( .A(b[913]), .B(n1353), .Z(n1354) );
  XOR U2377 ( .A(n1355), .B(n1356), .Z(n1353) );
  ANDN U2378 ( .B(n1357), .A(n98), .Z(n1355) );
  XOR U2379 ( .A(b[912]), .B(n1356), .Z(n1357) );
  XOR U2380 ( .A(n1358), .B(n1359), .Z(n1356) );
  ANDN U2381 ( .B(n1360), .A(n99), .Z(n1358) );
  XOR U2382 ( .A(b[911]), .B(n1359), .Z(n1360) );
  XOR U2383 ( .A(n1361), .B(n1362), .Z(n1359) );
  ANDN U2384 ( .B(n1363), .A(n100), .Z(n1361) );
  XOR U2385 ( .A(b[910]), .B(n1362), .Z(n1363) );
  XOR U2386 ( .A(n1364), .B(n1365), .Z(n1362) );
  ANDN U2387 ( .B(n1366), .A(n102), .Z(n1364) );
  XOR U2388 ( .A(b[909]), .B(n1365), .Z(n1366) );
  XOR U2389 ( .A(n1367), .B(n1368), .Z(n1365) );
  ANDN U2390 ( .B(n1369), .A(n103), .Z(n1367) );
  XOR U2391 ( .A(b[908]), .B(n1368), .Z(n1369) );
  XOR U2392 ( .A(n1370), .B(n1371), .Z(n1368) );
  ANDN U2393 ( .B(n1372), .A(n104), .Z(n1370) );
  XOR U2394 ( .A(b[907]), .B(n1371), .Z(n1372) );
  XOR U2395 ( .A(n1373), .B(n1374), .Z(n1371) );
  ANDN U2396 ( .B(n1375), .A(n105), .Z(n1373) );
  XOR U2397 ( .A(b[906]), .B(n1374), .Z(n1375) );
  XOR U2398 ( .A(n1376), .B(n1377), .Z(n1374) );
  ANDN U2399 ( .B(n1378), .A(n106), .Z(n1376) );
  XOR U2400 ( .A(b[905]), .B(n1377), .Z(n1378) );
  XOR U2401 ( .A(n1379), .B(n1380), .Z(n1377) );
  ANDN U2402 ( .B(n1381), .A(n107), .Z(n1379) );
  XOR U2403 ( .A(b[904]), .B(n1380), .Z(n1381) );
  XOR U2404 ( .A(n1382), .B(n1383), .Z(n1380) );
  ANDN U2405 ( .B(n1384), .A(n108), .Z(n1382) );
  XOR U2406 ( .A(b[903]), .B(n1383), .Z(n1384) );
  XOR U2407 ( .A(n1385), .B(n1386), .Z(n1383) );
  ANDN U2408 ( .B(n1387), .A(n109), .Z(n1385) );
  XOR U2409 ( .A(b[902]), .B(n1386), .Z(n1387) );
  XOR U2410 ( .A(n1388), .B(n1389), .Z(n1386) );
  ANDN U2411 ( .B(n1390), .A(n110), .Z(n1388) );
  XOR U2412 ( .A(b[901]), .B(n1389), .Z(n1390) );
  XOR U2413 ( .A(n1391), .B(n1392), .Z(n1389) );
  ANDN U2414 ( .B(n1393), .A(n111), .Z(n1391) );
  XOR U2415 ( .A(b[900]), .B(n1392), .Z(n1393) );
  XOR U2416 ( .A(n1394), .B(n1395), .Z(n1392) );
  ANDN U2417 ( .B(n1396), .A(n114), .Z(n1394) );
  XOR U2418 ( .A(b[899]), .B(n1395), .Z(n1396) );
  XOR U2419 ( .A(n1397), .B(n1398), .Z(n1395) );
  ANDN U2420 ( .B(n1399), .A(n115), .Z(n1397) );
  XOR U2421 ( .A(b[898]), .B(n1398), .Z(n1399) );
  XOR U2422 ( .A(n1400), .B(n1401), .Z(n1398) );
  ANDN U2423 ( .B(n1402), .A(n116), .Z(n1400) );
  XOR U2424 ( .A(b[897]), .B(n1401), .Z(n1402) );
  XOR U2425 ( .A(n1403), .B(n1404), .Z(n1401) );
  ANDN U2426 ( .B(n1405), .A(n117), .Z(n1403) );
  XOR U2427 ( .A(b[896]), .B(n1404), .Z(n1405) );
  XOR U2428 ( .A(n1406), .B(n1407), .Z(n1404) );
  ANDN U2429 ( .B(n1408), .A(n118), .Z(n1406) );
  XOR U2430 ( .A(b[895]), .B(n1407), .Z(n1408) );
  XOR U2431 ( .A(n1409), .B(n1410), .Z(n1407) );
  ANDN U2432 ( .B(n1411), .A(n119), .Z(n1409) );
  XOR U2433 ( .A(b[894]), .B(n1410), .Z(n1411) );
  XOR U2434 ( .A(n1412), .B(n1413), .Z(n1410) );
  ANDN U2435 ( .B(n1414), .A(n120), .Z(n1412) );
  XOR U2436 ( .A(b[893]), .B(n1413), .Z(n1414) );
  XOR U2437 ( .A(n1415), .B(n1416), .Z(n1413) );
  ANDN U2438 ( .B(n1417), .A(n121), .Z(n1415) );
  XOR U2439 ( .A(b[892]), .B(n1416), .Z(n1417) );
  XOR U2440 ( .A(n1418), .B(n1419), .Z(n1416) );
  ANDN U2441 ( .B(n1420), .A(n122), .Z(n1418) );
  XOR U2442 ( .A(b[891]), .B(n1419), .Z(n1420) );
  XOR U2443 ( .A(n1421), .B(n1422), .Z(n1419) );
  ANDN U2444 ( .B(n1423), .A(n123), .Z(n1421) );
  XOR U2445 ( .A(b[890]), .B(n1422), .Z(n1423) );
  XOR U2446 ( .A(n1424), .B(n1425), .Z(n1422) );
  ANDN U2447 ( .B(n1426), .A(n125), .Z(n1424) );
  XOR U2448 ( .A(b[889]), .B(n1425), .Z(n1426) );
  XOR U2449 ( .A(n1427), .B(n1428), .Z(n1425) );
  ANDN U2450 ( .B(n1429), .A(n126), .Z(n1427) );
  XOR U2451 ( .A(b[888]), .B(n1428), .Z(n1429) );
  XOR U2452 ( .A(n1430), .B(n1431), .Z(n1428) );
  ANDN U2453 ( .B(n1432), .A(n127), .Z(n1430) );
  XOR U2454 ( .A(b[887]), .B(n1431), .Z(n1432) );
  XOR U2455 ( .A(n1433), .B(n1434), .Z(n1431) );
  ANDN U2456 ( .B(n1435), .A(n128), .Z(n1433) );
  XOR U2457 ( .A(b[886]), .B(n1434), .Z(n1435) );
  XOR U2458 ( .A(n1436), .B(n1437), .Z(n1434) );
  ANDN U2459 ( .B(n1438), .A(n129), .Z(n1436) );
  XOR U2460 ( .A(b[885]), .B(n1437), .Z(n1438) );
  XOR U2461 ( .A(n1439), .B(n1440), .Z(n1437) );
  ANDN U2462 ( .B(n1441), .A(n130), .Z(n1439) );
  XOR U2463 ( .A(b[884]), .B(n1440), .Z(n1441) );
  XOR U2464 ( .A(n1442), .B(n1443), .Z(n1440) );
  ANDN U2465 ( .B(n1444), .A(n131), .Z(n1442) );
  XOR U2466 ( .A(b[883]), .B(n1443), .Z(n1444) );
  XOR U2467 ( .A(n1445), .B(n1446), .Z(n1443) );
  ANDN U2468 ( .B(n1447), .A(n132), .Z(n1445) );
  XOR U2469 ( .A(b[882]), .B(n1446), .Z(n1447) );
  XOR U2470 ( .A(n1448), .B(n1449), .Z(n1446) );
  ANDN U2471 ( .B(n1450), .A(n133), .Z(n1448) );
  XOR U2472 ( .A(b[881]), .B(n1449), .Z(n1450) );
  XOR U2473 ( .A(n1451), .B(n1452), .Z(n1449) );
  ANDN U2474 ( .B(n1453), .A(n134), .Z(n1451) );
  XOR U2475 ( .A(b[880]), .B(n1452), .Z(n1453) );
  XOR U2476 ( .A(n1454), .B(n1455), .Z(n1452) );
  ANDN U2477 ( .B(n1456), .A(n136), .Z(n1454) );
  XOR U2478 ( .A(b[879]), .B(n1455), .Z(n1456) );
  XOR U2479 ( .A(n1457), .B(n1458), .Z(n1455) );
  ANDN U2480 ( .B(n1459), .A(n137), .Z(n1457) );
  XOR U2481 ( .A(b[878]), .B(n1458), .Z(n1459) );
  XOR U2482 ( .A(n1460), .B(n1461), .Z(n1458) );
  ANDN U2483 ( .B(n1462), .A(n138), .Z(n1460) );
  XOR U2484 ( .A(b[877]), .B(n1461), .Z(n1462) );
  XOR U2485 ( .A(n1463), .B(n1464), .Z(n1461) );
  ANDN U2486 ( .B(n1465), .A(n139), .Z(n1463) );
  XOR U2487 ( .A(b[876]), .B(n1464), .Z(n1465) );
  XOR U2488 ( .A(n1466), .B(n1467), .Z(n1464) );
  ANDN U2489 ( .B(n1468), .A(n140), .Z(n1466) );
  XOR U2490 ( .A(b[875]), .B(n1467), .Z(n1468) );
  XOR U2491 ( .A(n1469), .B(n1470), .Z(n1467) );
  ANDN U2492 ( .B(n1471), .A(n141), .Z(n1469) );
  XOR U2493 ( .A(b[874]), .B(n1470), .Z(n1471) );
  XOR U2494 ( .A(n1472), .B(n1473), .Z(n1470) );
  ANDN U2495 ( .B(n1474), .A(n142), .Z(n1472) );
  XOR U2496 ( .A(b[873]), .B(n1473), .Z(n1474) );
  XOR U2497 ( .A(n1475), .B(n1476), .Z(n1473) );
  ANDN U2498 ( .B(n1477), .A(n143), .Z(n1475) );
  XOR U2499 ( .A(b[872]), .B(n1476), .Z(n1477) );
  XOR U2500 ( .A(n1478), .B(n1479), .Z(n1476) );
  ANDN U2501 ( .B(n1480), .A(n144), .Z(n1478) );
  XOR U2502 ( .A(b[871]), .B(n1479), .Z(n1480) );
  XOR U2503 ( .A(n1481), .B(n1482), .Z(n1479) );
  ANDN U2504 ( .B(n1483), .A(n145), .Z(n1481) );
  XOR U2505 ( .A(b[870]), .B(n1482), .Z(n1483) );
  XOR U2506 ( .A(n1484), .B(n1485), .Z(n1482) );
  ANDN U2507 ( .B(n1486), .A(n147), .Z(n1484) );
  XOR U2508 ( .A(b[869]), .B(n1485), .Z(n1486) );
  XOR U2509 ( .A(n1487), .B(n1488), .Z(n1485) );
  ANDN U2510 ( .B(n1489), .A(n148), .Z(n1487) );
  XOR U2511 ( .A(b[868]), .B(n1488), .Z(n1489) );
  XOR U2512 ( .A(n1490), .B(n1491), .Z(n1488) );
  ANDN U2513 ( .B(n1492), .A(n149), .Z(n1490) );
  XOR U2514 ( .A(b[867]), .B(n1491), .Z(n1492) );
  XOR U2515 ( .A(n1493), .B(n1494), .Z(n1491) );
  ANDN U2516 ( .B(n1495), .A(n150), .Z(n1493) );
  XOR U2517 ( .A(b[866]), .B(n1494), .Z(n1495) );
  XOR U2518 ( .A(n1496), .B(n1497), .Z(n1494) );
  ANDN U2519 ( .B(n1498), .A(n151), .Z(n1496) );
  XOR U2520 ( .A(b[865]), .B(n1497), .Z(n1498) );
  XOR U2521 ( .A(n1499), .B(n1500), .Z(n1497) );
  ANDN U2522 ( .B(n1501), .A(n152), .Z(n1499) );
  XOR U2523 ( .A(b[864]), .B(n1500), .Z(n1501) );
  XOR U2524 ( .A(n1502), .B(n1503), .Z(n1500) );
  ANDN U2525 ( .B(n1504), .A(n153), .Z(n1502) );
  XOR U2526 ( .A(b[863]), .B(n1503), .Z(n1504) );
  XOR U2527 ( .A(n1505), .B(n1506), .Z(n1503) );
  ANDN U2528 ( .B(n1507), .A(n154), .Z(n1505) );
  XOR U2529 ( .A(b[862]), .B(n1506), .Z(n1507) );
  XOR U2530 ( .A(n1508), .B(n1509), .Z(n1506) );
  ANDN U2531 ( .B(n1510), .A(n155), .Z(n1508) );
  XOR U2532 ( .A(b[861]), .B(n1509), .Z(n1510) );
  XOR U2533 ( .A(n1511), .B(n1512), .Z(n1509) );
  ANDN U2534 ( .B(n1513), .A(n156), .Z(n1511) );
  XOR U2535 ( .A(b[860]), .B(n1512), .Z(n1513) );
  XOR U2536 ( .A(n1514), .B(n1515), .Z(n1512) );
  ANDN U2537 ( .B(n1516), .A(n158), .Z(n1514) );
  XOR U2538 ( .A(b[859]), .B(n1515), .Z(n1516) );
  XOR U2539 ( .A(n1517), .B(n1518), .Z(n1515) );
  ANDN U2540 ( .B(n1519), .A(n159), .Z(n1517) );
  XOR U2541 ( .A(b[858]), .B(n1518), .Z(n1519) );
  XOR U2542 ( .A(n1520), .B(n1521), .Z(n1518) );
  ANDN U2543 ( .B(n1522), .A(n160), .Z(n1520) );
  XOR U2544 ( .A(b[857]), .B(n1521), .Z(n1522) );
  XOR U2545 ( .A(n1523), .B(n1524), .Z(n1521) );
  ANDN U2546 ( .B(n1525), .A(n161), .Z(n1523) );
  XOR U2547 ( .A(b[856]), .B(n1524), .Z(n1525) );
  XOR U2548 ( .A(n1526), .B(n1527), .Z(n1524) );
  ANDN U2549 ( .B(n1528), .A(n162), .Z(n1526) );
  XOR U2550 ( .A(b[855]), .B(n1527), .Z(n1528) );
  XOR U2551 ( .A(n1529), .B(n1530), .Z(n1527) );
  ANDN U2552 ( .B(n1531), .A(n163), .Z(n1529) );
  XOR U2553 ( .A(b[854]), .B(n1530), .Z(n1531) );
  XOR U2554 ( .A(n1532), .B(n1533), .Z(n1530) );
  ANDN U2555 ( .B(n1534), .A(n164), .Z(n1532) );
  XOR U2556 ( .A(b[853]), .B(n1533), .Z(n1534) );
  XOR U2557 ( .A(n1535), .B(n1536), .Z(n1533) );
  ANDN U2558 ( .B(n1537), .A(n165), .Z(n1535) );
  XOR U2559 ( .A(b[852]), .B(n1536), .Z(n1537) );
  XOR U2560 ( .A(n1538), .B(n1539), .Z(n1536) );
  ANDN U2561 ( .B(n1540), .A(n166), .Z(n1538) );
  XOR U2562 ( .A(b[851]), .B(n1539), .Z(n1540) );
  XOR U2563 ( .A(n1541), .B(n1542), .Z(n1539) );
  ANDN U2564 ( .B(n1543), .A(n167), .Z(n1541) );
  XOR U2565 ( .A(b[850]), .B(n1542), .Z(n1543) );
  XOR U2566 ( .A(n1544), .B(n1545), .Z(n1542) );
  ANDN U2567 ( .B(n1546), .A(n169), .Z(n1544) );
  XOR U2568 ( .A(b[849]), .B(n1545), .Z(n1546) );
  XOR U2569 ( .A(n1547), .B(n1548), .Z(n1545) );
  ANDN U2570 ( .B(n1549), .A(n170), .Z(n1547) );
  XOR U2571 ( .A(b[848]), .B(n1548), .Z(n1549) );
  XOR U2572 ( .A(n1550), .B(n1551), .Z(n1548) );
  ANDN U2573 ( .B(n1552), .A(n171), .Z(n1550) );
  XOR U2574 ( .A(b[847]), .B(n1551), .Z(n1552) );
  XOR U2575 ( .A(n1553), .B(n1554), .Z(n1551) );
  ANDN U2576 ( .B(n1555), .A(n172), .Z(n1553) );
  XOR U2577 ( .A(b[846]), .B(n1554), .Z(n1555) );
  XOR U2578 ( .A(n1556), .B(n1557), .Z(n1554) );
  ANDN U2579 ( .B(n1558), .A(n173), .Z(n1556) );
  XOR U2580 ( .A(b[845]), .B(n1557), .Z(n1558) );
  XOR U2581 ( .A(n1559), .B(n1560), .Z(n1557) );
  ANDN U2582 ( .B(n1561), .A(n174), .Z(n1559) );
  XOR U2583 ( .A(b[844]), .B(n1560), .Z(n1561) );
  XOR U2584 ( .A(n1562), .B(n1563), .Z(n1560) );
  ANDN U2585 ( .B(n1564), .A(n175), .Z(n1562) );
  XOR U2586 ( .A(b[843]), .B(n1563), .Z(n1564) );
  XOR U2587 ( .A(n1565), .B(n1566), .Z(n1563) );
  ANDN U2588 ( .B(n1567), .A(n176), .Z(n1565) );
  XOR U2589 ( .A(b[842]), .B(n1566), .Z(n1567) );
  XOR U2590 ( .A(n1568), .B(n1569), .Z(n1566) );
  ANDN U2591 ( .B(n1570), .A(n177), .Z(n1568) );
  XOR U2592 ( .A(b[841]), .B(n1569), .Z(n1570) );
  XOR U2593 ( .A(n1571), .B(n1572), .Z(n1569) );
  ANDN U2594 ( .B(n1573), .A(n178), .Z(n1571) );
  XOR U2595 ( .A(b[840]), .B(n1572), .Z(n1573) );
  XOR U2596 ( .A(n1574), .B(n1575), .Z(n1572) );
  ANDN U2597 ( .B(n1576), .A(n180), .Z(n1574) );
  XOR U2598 ( .A(b[839]), .B(n1575), .Z(n1576) );
  XOR U2599 ( .A(n1577), .B(n1578), .Z(n1575) );
  ANDN U2600 ( .B(n1579), .A(n181), .Z(n1577) );
  XOR U2601 ( .A(b[838]), .B(n1578), .Z(n1579) );
  XOR U2602 ( .A(n1580), .B(n1581), .Z(n1578) );
  ANDN U2603 ( .B(n1582), .A(n182), .Z(n1580) );
  XOR U2604 ( .A(b[837]), .B(n1581), .Z(n1582) );
  XOR U2605 ( .A(n1583), .B(n1584), .Z(n1581) );
  ANDN U2606 ( .B(n1585), .A(n183), .Z(n1583) );
  XOR U2607 ( .A(b[836]), .B(n1584), .Z(n1585) );
  XOR U2608 ( .A(n1586), .B(n1587), .Z(n1584) );
  ANDN U2609 ( .B(n1588), .A(n184), .Z(n1586) );
  XOR U2610 ( .A(b[835]), .B(n1587), .Z(n1588) );
  XOR U2611 ( .A(n1589), .B(n1590), .Z(n1587) );
  ANDN U2612 ( .B(n1591), .A(n185), .Z(n1589) );
  XOR U2613 ( .A(b[834]), .B(n1590), .Z(n1591) );
  XOR U2614 ( .A(n1592), .B(n1593), .Z(n1590) );
  ANDN U2615 ( .B(n1594), .A(n186), .Z(n1592) );
  XOR U2616 ( .A(b[833]), .B(n1593), .Z(n1594) );
  XOR U2617 ( .A(n1595), .B(n1596), .Z(n1593) );
  ANDN U2618 ( .B(n1597), .A(n187), .Z(n1595) );
  XOR U2619 ( .A(b[832]), .B(n1596), .Z(n1597) );
  XOR U2620 ( .A(n1598), .B(n1599), .Z(n1596) );
  ANDN U2621 ( .B(n1600), .A(n188), .Z(n1598) );
  XOR U2622 ( .A(b[831]), .B(n1599), .Z(n1600) );
  XOR U2623 ( .A(n1601), .B(n1602), .Z(n1599) );
  ANDN U2624 ( .B(n1603), .A(n189), .Z(n1601) );
  XOR U2625 ( .A(b[830]), .B(n1602), .Z(n1603) );
  XOR U2626 ( .A(n1604), .B(n1605), .Z(n1602) );
  ANDN U2627 ( .B(n1606), .A(n191), .Z(n1604) );
  XOR U2628 ( .A(b[829]), .B(n1605), .Z(n1606) );
  XOR U2629 ( .A(n1607), .B(n1608), .Z(n1605) );
  ANDN U2630 ( .B(n1609), .A(n192), .Z(n1607) );
  XOR U2631 ( .A(b[828]), .B(n1608), .Z(n1609) );
  XOR U2632 ( .A(n1610), .B(n1611), .Z(n1608) );
  ANDN U2633 ( .B(n1612), .A(n193), .Z(n1610) );
  XOR U2634 ( .A(b[827]), .B(n1611), .Z(n1612) );
  XOR U2635 ( .A(n1613), .B(n1614), .Z(n1611) );
  ANDN U2636 ( .B(n1615), .A(n194), .Z(n1613) );
  XOR U2637 ( .A(b[826]), .B(n1614), .Z(n1615) );
  XOR U2638 ( .A(n1616), .B(n1617), .Z(n1614) );
  ANDN U2639 ( .B(n1618), .A(n195), .Z(n1616) );
  XOR U2640 ( .A(b[825]), .B(n1617), .Z(n1618) );
  XOR U2641 ( .A(n1619), .B(n1620), .Z(n1617) );
  ANDN U2642 ( .B(n1621), .A(n196), .Z(n1619) );
  XOR U2643 ( .A(b[824]), .B(n1620), .Z(n1621) );
  XOR U2644 ( .A(n1622), .B(n1623), .Z(n1620) );
  ANDN U2645 ( .B(n1624), .A(n197), .Z(n1622) );
  XOR U2646 ( .A(b[823]), .B(n1623), .Z(n1624) );
  XOR U2647 ( .A(n1625), .B(n1626), .Z(n1623) );
  ANDN U2648 ( .B(n1627), .A(n198), .Z(n1625) );
  XOR U2649 ( .A(b[822]), .B(n1626), .Z(n1627) );
  XOR U2650 ( .A(n1628), .B(n1629), .Z(n1626) );
  ANDN U2651 ( .B(n1630), .A(n199), .Z(n1628) );
  XOR U2652 ( .A(b[821]), .B(n1629), .Z(n1630) );
  XOR U2653 ( .A(n1631), .B(n1632), .Z(n1629) );
  ANDN U2654 ( .B(n1633), .A(n200), .Z(n1631) );
  XOR U2655 ( .A(b[820]), .B(n1632), .Z(n1633) );
  XOR U2656 ( .A(n1634), .B(n1635), .Z(n1632) );
  ANDN U2657 ( .B(n1636), .A(n202), .Z(n1634) );
  XOR U2658 ( .A(b[819]), .B(n1635), .Z(n1636) );
  XOR U2659 ( .A(n1637), .B(n1638), .Z(n1635) );
  ANDN U2660 ( .B(n1639), .A(n203), .Z(n1637) );
  XOR U2661 ( .A(b[818]), .B(n1638), .Z(n1639) );
  XOR U2662 ( .A(n1640), .B(n1641), .Z(n1638) );
  ANDN U2663 ( .B(n1642), .A(n204), .Z(n1640) );
  XOR U2664 ( .A(b[817]), .B(n1641), .Z(n1642) );
  XOR U2665 ( .A(n1643), .B(n1644), .Z(n1641) );
  ANDN U2666 ( .B(n1645), .A(n205), .Z(n1643) );
  XOR U2667 ( .A(b[816]), .B(n1644), .Z(n1645) );
  XOR U2668 ( .A(n1646), .B(n1647), .Z(n1644) );
  ANDN U2669 ( .B(n1648), .A(n206), .Z(n1646) );
  XOR U2670 ( .A(b[815]), .B(n1647), .Z(n1648) );
  XOR U2671 ( .A(n1649), .B(n1650), .Z(n1647) );
  ANDN U2672 ( .B(n1651), .A(n207), .Z(n1649) );
  XOR U2673 ( .A(b[814]), .B(n1650), .Z(n1651) );
  XOR U2674 ( .A(n1652), .B(n1653), .Z(n1650) );
  ANDN U2675 ( .B(n1654), .A(n208), .Z(n1652) );
  XOR U2676 ( .A(b[813]), .B(n1653), .Z(n1654) );
  XOR U2677 ( .A(n1655), .B(n1656), .Z(n1653) );
  ANDN U2678 ( .B(n1657), .A(n209), .Z(n1655) );
  XOR U2679 ( .A(b[812]), .B(n1656), .Z(n1657) );
  XOR U2680 ( .A(n1658), .B(n1659), .Z(n1656) );
  ANDN U2681 ( .B(n1660), .A(n210), .Z(n1658) );
  XOR U2682 ( .A(b[811]), .B(n1659), .Z(n1660) );
  XOR U2683 ( .A(n1661), .B(n1662), .Z(n1659) );
  ANDN U2684 ( .B(n1663), .A(n211), .Z(n1661) );
  XOR U2685 ( .A(b[810]), .B(n1662), .Z(n1663) );
  XOR U2686 ( .A(n1664), .B(n1665), .Z(n1662) );
  ANDN U2687 ( .B(n1666), .A(n213), .Z(n1664) );
  XOR U2688 ( .A(b[809]), .B(n1665), .Z(n1666) );
  XOR U2689 ( .A(n1667), .B(n1668), .Z(n1665) );
  ANDN U2690 ( .B(n1669), .A(n214), .Z(n1667) );
  XOR U2691 ( .A(b[808]), .B(n1668), .Z(n1669) );
  XOR U2692 ( .A(n1670), .B(n1671), .Z(n1668) );
  ANDN U2693 ( .B(n1672), .A(n215), .Z(n1670) );
  XOR U2694 ( .A(b[807]), .B(n1671), .Z(n1672) );
  XOR U2695 ( .A(n1673), .B(n1674), .Z(n1671) );
  ANDN U2696 ( .B(n1675), .A(n216), .Z(n1673) );
  XOR U2697 ( .A(b[806]), .B(n1674), .Z(n1675) );
  XOR U2698 ( .A(n1676), .B(n1677), .Z(n1674) );
  ANDN U2699 ( .B(n1678), .A(n217), .Z(n1676) );
  XOR U2700 ( .A(b[805]), .B(n1677), .Z(n1678) );
  XOR U2701 ( .A(n1679), .B(n1680), .Z(n1677) );
  ANDN U2702 ( .B(n1681), .A(n218), .Z(n1679) );
  XOR U2703 ( .A(b[804]), .B(n1680), .Z(n1681) );
  XOR U2704 ( .A(n1682), .B(n1683), .Z(n1680) );
  ANDN U2705 ( .B(n1684), .A(n219), .Z(n1682) );
  XOR U2706 ( .A(b[803]), .B(n1683), .Z(n1684) );
  XOR U2707 ( .A(n1685), .B(n1686), .Z(n1683) );
  ANDN U2708 ( .B(n1687), .A(n220), .Z(n1685) );
  XOR U2709 ( .A(b[802]), .B(n1686), .Z(n1687) );
  XOR U2710 ( .A(n1688), .B(n1689), .Z(n1686) );
  ANDN U2711 ( .B(n1690), .A(n221), .Z(n1688) );
  XOR U2712 ( .A(b[801]), .B(n1689), .Z(n1690) );
  XOR U2713 ( .A(n1691), .B(n1692), .Z(n1689) );
  ANDN U2714 ( .B(n1693), .A(n222), .Z(n1691) );
  XOR U2715 ( .A(b[800]), .B(n1692), .Z(n1693) );
  XOR U2716 ( .A(n1694), .B(n1695), .Z(n1692) );
  ANDN U2717 ( .B(n1696), .A(n225), .Z(n1694) );
  XOR U2718 ( .A(b[799]), .B(n1695), .Z(n1696) );
  XOR U2719 ( .A(n1697), .B(n1698), .Z(n1695) );
  ANDN U2720 ( .B(n1699), .A(n226), .Z(n1697) );
  XOR U2721 ( .A(b[798]), .B(n1698), .Z(n1699) );
  XOR U2722 ( .A(n1700), .B(n1701), .Z(n1698) );
  ANDN U2723 ( .B(n1702), .A(n227), .Z(n1700) );
  XOR U2724 ( .A(b[797]), .B(n1701), .Z(n1702) );
  XOR U2725 ( .A(n1703), .B(n1704), .Z(n1701) );
  ANDN U2726 ( .B(n1705), .A(n228), .Z(n1703) );
  XOR U2727 ( .A(b[796]), .B(n1704), .Z(n1705) );
  XOR U2728 ( .A(n1706), .B(n1707), .Z(n1704) );
  ANDN U2729 ( .B(n1708), .A(n229), .Z(n1706) );
  XOR U2730 ( .A(b[795]), .B(n1707), .Z(n1708) );
  XOR U2731 ( .A(n1709), .B(n1710), .Z(n1707) );
  ANDN U2732 ( .B(n1711), .A(n230), .Z(n1709) );
  XOR U2733 ( .A(b[794]), .B(n1710), .Z(n1711) );
  XOR U2734 ( .A(n1712), .B(n1713), .Z(n1710) );
  ANDN U2735 ( .B(n1714), .A(n231), .Z(n1712) );
  XOR U2736 ( .A(b[793]), .B(n1713), .Z(n1714) );
  XOR U2737 ( .A(n1715), .B(n1716), .Z(n1713) );
  ANDN U2738 ( .B(n1717), .A(n232), .Z(n1715) );
  XOR U2739 ( .A(b[792]), .B(n1716), .Z(n1717) );
  XOR U2740 ( .A(n1718), .B(n1719), .Z(n1716) );
  ANDN U2741 ( .B(n1720), .A(n233), .Z(n1718) );
  XOR U2742 ( .A(b[791]), .B(n1719), .Z(n1720) );
  XOR U2743 ( .A(n1721), .B(n1722), .Z(n1719) );
  ANDN U2744 ( .B(n1723), .A(n234), .Z(n1721) );
  XOR U2745 ( .A(b[790]), .B(n1722), .Z(n1723) );
  XOR U2746 ( .A(n1724), .B(n1725), .Z(n1722) );
  ANDN U2747 ( .B(n1726), .A(n236), .Z(n1724) );
  XOR U2748 ( .A(b[789]), .B(n1725), .Z(n1726) );
  XOR U2749 ( .A(n1727), .B(n1728), .Z(n1725) );
  ANDN U2750 ( .B(n1729), .A(n237), .Z(n1727) );
  XOR U2751 ( .A(b[788]), .B(n1728), .Z(n1729) );
  XOR U2752 ( .A(n1730), .B(n1731), .Z(n1728) );
  ANDN U2753 ( .B(n1732), .A(n238), .Z(n1730) );
  XOR U2754 ( .A(b[787]), .B(n1731), .Z(n1732) );
  XOR U2755 ( .A(n1733), .B(n1734), .Z(n1731) );
  ANDN U2756 ( .B(n1735), .A(n239), .Z(n1733) );
  XOR U2757 ( .A(b[786]), .B(n1734), .Z(n1735) );
  XOR U2758 ( .A(n1736), .B(n1737), .Z(n1734) );
  ANDN U2759 ( .B(n1738), .A(n240), .Z(n1736) );
  XOR U2760 ( .A(b[785]), .B(n1737), .Z(n1738) );
  XOR U2761 ( .A(n1739), .B(n1740), .Z(n1737) );
  ANDN U2762 ( .B(n1741), .A(n241), .Z(n1739) );
  XOR U2763 ( .A(b[784]), .B(n1740), .Z(n1741) );
  XOR U2764 ( .A(n1742), .B(n1743), .Z(n1740) );
  ANDN U2765 ( .B(n1744), .A(n242), .Z(n1742) );
  XOR U2766 ( .A(b[783]), .B(n1743), .Z(n1744) );
  XOR U2767 ( .A(n1745), .B(n1746), .Z(n1743) );
  ANDN U2768 ( .B(n1747), .A(n243), .Z(n1745) );
  XOR U2769 ( .A(b[782]), .B(n1746), .Z(n1747) );
  XOR U2770 ( .A(n1748), .B(n1749), .Z(n1746) );
  ANDN U2771 ( .B(n1750), .A(n244), .Z(n1748) );
  XOR U2772 ( .A(b[781]), .B(n1749), .Z(n1750) );
  XOR U2773 ( .A(n1751), .B(n1752), .Z(n1749) );
  ANDN U2774 ( .B(n1753), .A(n245), .Z(n1751) );
  XOR U2775 ( .A(b[780]), .B(n1752), .Z(n1753) );
  XOR U2776 ( .A(n1754), .B(n1755), .Z(n1752) );
  ANDN U2777 ( .B(n1756), .A(n247), .Z(n1754) );
  XOR U2778 ( .A(b[779]), .B(n1755), .Z(n1756) );
  XOR U2779 ( .A(n1757), .B(n1758), .Z(n1755) );
  ANDN U2780 ( .B(n1759), .A(n248), .Z(n1757) );
  XOR U2781 ( .A(b[778]), .B(n1758), .Z(n1759) );
  XOR U2782 ( .A(n1760), .B(n1761), .Z(n1758) );
  ANDN U2783 ( .B(n1762), .A(n249), .Z(n1760) );
  XOR U2784 ( .A(b[777]), .B(n1761), .Z(n1762) );
  XOR U2785 ( .A(n1763), .B(n1764), .Z(n1761) );
  ANDN U2786 ( .B(n1765), .A(n250), .Z(n1763) );
  XOR U2787 ( .A(b[776]), .B(n1764), .Z(n1765) );
  XOR U2788 ( .A(n1766), .B(n1767), .Z(n1764) );
  ANDN U2789 ( .B(n1768), .A(n251), .Z(n1766) );
  XOR U2790 ( .A(b[775]), .B(n1767), .Z(n1768) );
  XOR U2791 ( .A(n1769), .B(n1770), .Z(n1767) );
  ANDN U2792 ( .B(n1771), .A(n252), .Z(n1769) );
  XOR U2793 ( .A(b[774]), .B(n1770), .Z(n1771) );
  XOR U2794 ( .A(n1772), .B(n1773), .Z(n1770) );
  ANDN U2795 ( .B(n1774), .A(n253), .Z(n1772) );
  XOR U2796 ( .A(b[773]), .B(n1773), .Z(n1774) );
  XOR U2797 ( .A(n1775), .B(n1776), .Z(n1773) );
  ANDN U2798 ( .B(n1777), .A(n254), .Z(n1775) );
  XOR U2799 ( .A(b[772]), .B(n1776), .Z(n1777) );
  XOR U2800 ( .A(n1778), .B(n1779), .Z(n1776) );
  ANDN U2801 ( .B(n1780), .A(n255), .Z(n1778) );
  XOR U2802 ( .A(b[771]), .B(n1779), .Z(n1780) );
  XOR U2803 ( .A(n1781), .B(n1782), .Z(n1779) );
  ANDN U2804 ( .B(n1783), .A(n256), .Z(n1781) );
  XOR U2805 ( .A(b[770]), .B(n1782), .Z(n1783) );
  XOR U2806 ( .A(n1784), .B(n1785), .Z(n1782) );
  ANDN U2807 ( .B(n1786), .A(n258), .Z(n1784) );
  XOR U2808 ( .A(b[769]), .B(n1785), .Z(n1786) );
  XOR U2809 ( .A(n1787), .B(n1788), .Z(n1785) );
  ANDN U2810 ( .B(n1789), .A(n259), .Z(n1787) );
  XOR U2811 ( .A(b[768]), .B(n1788), .Z(n1789) );
  XOR U2812 ( .A(n1790), .B(n1791), .Z(n1788) );
  ANDN U2813 ( .B(n1792), .A(n260), .Z(n1790) );
  XOR U2814 ( .A(b[767]), .B(n1791), .Z(n1792) );
  XOR U2815 ( .A(n1793), .B(n1794), .Z(n1791) );
  ANDN U2816 ( .B(n1795), .A(n261), .Z(n1793) );
  XOR U2817 ( .A(b[766]), .B(n1794), .Z(n1795) );
  XOR U2818 ( .A(n1796), .B(n1797), .Z(n1794) );
  ANDN U2819 ( .B(n1798), .A(n262), .Z(n1796) );
  XOR U2820 ( .A(b[765]), .B(n1797), .Z(n1798) );
  XOR U2821 ( .A(n1799), .B(n1800), .Z(n1797) );
  ANDN U2822 ( .B(n1801), .A(n263), .Z(n1799) );
  XOR U2823 ( .A(b[764]), .B(n1800), .Z(n1801) );
  XOR U2824 ( .A(n1802), .B(n1803), .Z(n1800) );
  ANDN U2825 ( .B(n1804), .A(n264), .Z(n1802) );
  XOR U2826 ( .A(b[763]), .B(n1803), .Z(n1804) );
  XOR U2827 ( .A(n1805), .B(n1806), .Z(n1803) );
  ANDN U2828 ( .B(n1807), .A(n265), .Z(n1805) );
  XOR U2829 ( .A(b[762]), .B(n1806), .Z(n1807) );
  XOR U2830 ( .A(n1808), .B(n1809), .Z(n1806) );
  ANDN U2831 ( .B(n1810), .A(n266), .Z(n1808) );
  XOR U2832 ( .A(b[761]), .B(n1809), .Z(n1810) );
  XOR U2833 ( .A(n1811), .B(n1812), .Z(n1809) );
  ANDN U2834 ( .B(n1813), .A(n267), .Z(n1811) );
  XOR U2835 ( .A(b[760]), .B(n1812), .Z(n1813) );
  XOR U2836 ( .A(n1814), .B(n1815), .Z(n1812) );
  ANDN U2837 ( .B(n1816), .A(n269), .Z(n1814) );
  XOR U2838 ( .A(b[759]), .B(n1815), .Z(n1816) );
  XOR U2839 ( .A(n1817), .B(n1818), .Z(n1815) );
  ANDN U2840 ( .B(n1819), .A(n270), .Z(n1817) );
  XOR U2841 ( .A(b[758]), .B(n1818), .Z(n1819) );
  XOR U2842 ( .A(n1820), .B(n1821), .Z(n1818) );
  ANDN U2843 ( .B(n1822), .A(n271), .Z(n1820) );
  XOR U2844 ( .A(b[757]), .B(n1821), .Z(n1822) );
  XOR U2845 ( .A(n1823), .B(n1824), .Z(n1821) );
  ANDN U2846 ( .B(n1825), .A(n272), .Z(n1823) );
  XOR U2847 ( .A(b[756]), .B(n1824), .Z(n1825) );
  XOR U2848 ( .A(n1826), .B(n1827), .Z(n1824) );
  ANDN U2849 ( .B(n1828), .A(n273), .Z(n1826) );
  XOR U2850 ( .A(b[755]), .B(n1827), .Z(n1828) );
  XOR U2851 ( .A(n1829), .B(n1830), .Z(n1827) );
  ANDN U2852 ( .B(n1831), .A(n274), .Z(n1829) );
  XOR U2853 ( .A(b[754]), .B(n1830), .Z(n1831) );
  XOR U2854 ( .A(n1832), .B(n1833), .Z(n1830) );
  ANDN U2855 ( .B(n1834), .A(n275), .Z(n1832) );
  XOR U2856 ( .A(b[753]), .B(n1833), .Z(n1834) );
  XOR U2857 ( .A(n1835), .B(n1836), .Z(n1833) );
  ANDN U2858 ( .B(n1837), .A(n276), .Z(n1835) );
  XOR U2859 ( .A(b[752]), .B(n1836), .Z(n1837) );
  XOR U2860 ( .A(n1838), .B(n1839), .Z(n1836) );
  ANDN U2861 ( .B(n1840), .A(n277), .Z(n1838) );
  XOR U2862 ( .A(b[751]), .B(n1839), .Z(n1840) );
  XOR U2863 ( .A(n1841), .B(n1842), .Z(n1839) );
  ANDN U2864 ( .B(n1843), .A(n278), .Z(n1841) );
  XOR U2865 ( .A(b[750]), .B(n1842), .Z(n1843) );
  XOR U2866 ( .A(n1844), .B(n1845), .Z(n1842) );
  ANDN U2867 ( .B(n1846), .A(n280), .Z(n1844) );
  XOR U2868 ( .A(b[749]), .B(n1845), .Z(n1846) );
  XOR U2869 ( .A(n1847), .B(n1848), .Z(n1845) );
  ANDN U2870 ( .B(n1849), .A(n281), .Z(n1847) );
  XOR U2871 ( .A(b[748]), .B(n1848), .Z(n1849) );
  XOR U2872 ( .A(n1850), .B(n1851), .Z(n1848) );
  ANDN U2873 ( .B(n1852), .A(n282), .Z(n1850) );
  XOR U2874 ( .A(b[747]), .B(n1851), .Z(n1852) );
  XOR U2875 ( .A(n1853), .B(n1854), .Z(n1851) );
  ANDN U2876 ( .B(n1855), .A(n283), .Z(n1853) );
  XOR U2877 ( .A(b[746]), .B(n1854), .Z(n1855) );
  XOR U2878 ( .A(n1856), .B(n1857), .Z(n1854) );
  ANDN U2879 ( .B(n1858), .A(n284), .Z(n1856) );
  XOR U2880 ( .A(b[745]), .B(n1857), .Z(n1858) );
  XOR U2881 ( .A(n1859), .B(n1860), .Z(n1857) );
  ANDN U2882 ( .B(n1861), .A(n285), .Z(n1859) );
  XOR U2883 ( .A(b[744]), .B(n1860), .Z(n1861) );
  XOR U2884 ( .A(n1862), .B(n1863), .Z(n1860) );
  ANDN U2885 ( .B(n1864), .A(n286), .Z(n1862) );
  XOR U2886 ( .A(b[743]), .B(n1863), .Z(n1864) );
  XOR U2887 ( .A(n1865), .B(n1866), .Z(n1863) );
  ANDN U2888 ( .B(n1867), .A(n287), .Z(n1865) );
  XOR U2889 ( .A(b[742]), .B(n1866), .Z(n1867) );
  XOR U2890 ( .A(n1868), .B(n1869), .Z(n1866) );
  ANDN U2891 ( .B(n1870), .A(n288), .Z(n1868) );
  XOR U2892 ( .A(b[741]), .B(n1869), .Z(n1870) );
  XOR U2893 ( .A(n1871), .B(n1872), .Z(n1869) );
  ANDN U2894 ( .B(n1873), .A(n289), .Z(n1871) );
  XOR U2895 ( .A(b[740]), .B(n1872), .Z(n1873) );
  XOR U2896 ( .A(n1874), .B(n1875), .Z(n1872) );
  ANDN U2897 ( .B(n1876), .A(n291), .Z(n1874) );
  XOR U2898 ( .A(b[739]), .B(n1875), .Z(n1876) );
  XOR U2899 ( .A(n1877), .B(n1878), .Z(n1875) );
  ANDN U2900 ( .B(n1879), .A(n292), .Z(n1877) );
  XOR U2901 ( .A(b[738]), .B(n1878), .Z(n1879) );
  XOR U2902 ( .A(n1880), .B(n1881), .Z(n1878) );
  ANDN U2903 ( .B(n1882), .A(n293), .Z(n1880) );
  XOR U2904 ( .A(b[737]), .B(n1881), .Z(n1882) );
  XOR U2905 ( .A(n1883), .B(n1884), .Z(n1881) );
  ANDN U2906 ( .B(n1885), .A(n294), .Z(n1883) );
  XOR U2907 ( .A(b[736]), .B(n1884), .Z(n1885) );
  XOR U2908 ( .A(n1886), .B(n1887), .Z(n1884) );
  ANDN U2909 ( .B(n1888), .A(n295), .Z(n1886) );
  XOR U2910 ( .A(b[735]), .B(n1887), .Z(n1888) );
  XOR U2911 ( .A(n1889), .B(n1890), .Z(n1887) );
  ANDN U2912 ( .B(n1891), .A(n296), .Z(n1889) );
  XOR U2913 ( .A(b[734]), .B(n1890), .Z(n1891) );
  XOR U2914 ( .A(n1892), .B(n1893), .Z(n1890) );
  ANDN U2915 ( .B(n1894), .A(n297), .Z(n1892) );
  XOR U2916 ( .A(b[733]), .B(n1893), .Z(n1894) );
  XOR U2917 ( .A(n1895), .B(n1896), .Z(n1893) );
  ANDN U2918 ( .B(n1897), .A(n298), .Z(n1895) );
  XOR U2919 ( .A(b[732]), .B(n1896), .Z(n1897) );
  XOR U2920 ( .A(n1898), .B(n1899), .Z(n1896) );
  ANDN U2921 ( .B(n1900), .A(n299), .Z(n1898) );
  XOR U2922 ( .A(b[731]), .B(n1899), .Z(n1900) );
  XOR U2923 ( .A(n1901), .B(n1902), .Z(n1899) );
  ANDN U2924 ( .B(n1903), .A(n300), .Z(n1901) );
  XOR U2925 ( .A(b[730]), .B(n1902), .Z(n1903) );
  XOR U2926 ( .A(n1904), .B(n1905), .Z(n1902) );
  ANDN U2927 ( .B(n1906), .A(n302), .Z(n1904) );
  XOR U2928 ( .A(b[729]), .B(n1905), .Z(n1906) );
  XOR U2929 ( .A(n1907), .B(n1908), .Z(n1905) );
  ANDN U2930 ( .B(n1909), .A(n303), .Z(n1907) );
  XOR U2931 ( .A(b[728]), .B(n1908), .Z(n1909) );
  XOR U2932 ( .A(n1910), .B(n1911), .Z(n1908) );
  ANDN U2933 ( .B(n1912), .A(n304), .Z(n1910) );
  XOR U2934 ( .A(b[727]), .B(n1911), .Z(n1912) );
  XOR U2935 ( .A(n1913), .B(n1914), .Z(n1911) );
  ANDN U2936 ( .B(n1915), .A(n305), .Z(n1913) );
  XOR U2937 ( .A(b[726]), .B(n1914), .Z(n1915) );
  XOR U2938 ( .A(n1916), .B(n1917), .Z(n1914) );
  ANDN U2939 ( .B(n1918), .A(n306), .Z(n1916) );
  XOR U2940 ( .A(b[725]), .B(n1917), .Z(n1918) );
  XOR U2941 ( .A(n1919), .B(n1920), .Z(n1917) );
  ANDN U2942 ( .B(n1921), .A(n307), .Z(n1919) );
  XOR U2943 ( .A(b[724]), .B(n1920), .Z(n1921) );
  XOR U2944 ( .A(n1922), .B(n1923), .Z(n1920) );
  ANDN U2945 ( .B(n1924), .A(n308), .Z(n1922) );
  XOR U2946 ( .A(b[723]), .B(n1923), .Z(n1924) );
  XOR U2947 ( .A(n1925), .B(n1926), .Z(n1923) );
  ANDN U2948 ( .B(n1927), .A(n309), .Z(n1925) );
  XOR U2949 ( .A(b[722]), .B(n1926), .Z(n1927) );
  XOR U2950 ( .A(n1928), .B(n1929), .Z(n1926) );
  ANDN U2951 ( .B(n1930), .A(n310), .Z(n1928) );
  XOR U2952 ( .A(b[721]), .B(n1929), .Z(n1930) );
  XOR U2953 ( .A(n1931), .B(n1932), .Z(n1929) );
  ANDN U2954 ( .B(n1933), .A(n311), .Z(n1931) );
  XOR U2955 ( .A(b[720]), .B(n1932), .Z(n1933) );
  XOR U2956 ( .A(n1934), .B(n1935), .Z(n1932) );
  ANDN U2957 ( .B(n1936), .A(n313), .Z(n1934) );
  XOR U2958 ( .A(b[719]), .B(n1935), .Z(n1936) );
  XOR U2959 ( .A(n1937), .B(n1938), .Z(n1935) );
  ANDN U2960 ( .B(n1939), .A(n314), .Z(n1937) );
  XOR U2961 ( .A(b[718]), .B(n1938), .Z(n1939) );
  XOR U2962 ( .A(n1940), .B(n1941), .Z(n1938) );
  ANDN U2963 ( .B(n1942), .A(n315), .Z(n1940) );
  XOR U2964 ( .A(b[717]), .B(n1941), .Z(n1942) );
  XOR U2965 ( .A(n1943), .B(n1944), .Z(n1941) );
  ANDN U2966 ( .B(n1945), .A(n316), .Z(n1943) );
  XOR U2967 ( .A(b[716]), .B(n1944), .Z(n1945) );
  XOR U2968 ( .A(n1946), .B(n1947), .Z(n1944) );
  ANDN U2969 ( .B(n1948), .A(n317), .Z(n1946) );
  XOR U2970 ( .A(b[715]), .B(n1947), .Z(n1948) );
  XOR U2971 ( .A(n1949), .B(n1950), .Z(n1947) );
  ANDN U2972 ( .B(n1951), .A(n318), .Z(n1949) );
  XOR U2973 ( .A(b[714]), .B(n1950), .Z(n1951) );
  XOR U2974 ( .A(n1952), .B(n1953), .Z(n1950) );
  ANDN U2975 ( .B(n1954), .A(n319), .Z(n1952) );
  XOR U2976 ( .A(b[713]), .B(n1953), .Z(n1954) );
  XOR U2977 ( .A(n1955), .B(n1956), .Z(n1953) );
  ANDN U2978 ( .B(n1957), .A(n320), .Z(n1955) );
  XOR U2979 ( .A(b[712]), .B(n1956), .Z(n1957) );
  XOR U2980 ( .A(n1958), .B(n1959), .Z(n1956) );
  ANDN U2981 ( .B(n1960), .A(n321), .Z(n1958) );
  XOR U2982 ( .A(b[711]), .B(n1959), .Z(n1960) );
  XOR U2983 ( .A(n1961), .B(n1962), .Z(n1959) );
  ANDN U2984 ( .B(n1963), .A(n322), .Z(n1961) );
  XOR U2985 ( .A(b[710]), .B(n1962), .Z(n1963) );
  XOR U2986 ( .A(n1964), .B(n1965), .Z(n1962) );
  ANDN U2987 ( .B(n1966), .A(n324), .Z(n1964) );
  XOR U2988 ( .A(b[709]), .B(n1965), .Z(n1966) );
  XOR U2989 ( .A(n1967), .B(n1968), .Z(n1965) );
  ANDN U2990 ( .B(n1969), .A(n325), .Z(n1967) );
  XOR U2991 ( .A(b[708]), .B(n1968), .Z(n1969) );
  XOR U2992 ( .A(n1970), .B(n1971), .Z(n1968) );
  ANDN U2993 ( .B(n1972), .A(n326), .Z(n1970) );
  XOR U2994 ( .A(b[707]), .B(n1971), .Z(n1972) );
  XOR U2995 ( .A(n1973), .B(n1974), .Z(n1971) );
  ANDN U2996 ( .B(n1975), .A(n327), .Z(n1973) );
  XOR U2997 ( .A(b[706]), .B(n1974), .Z(n1975) );
  XOR U2998 ( .A(n1976), .B(n1977), .Z(n1974) );
  ANDN U2999 ( .B(n1978), .A(n328), .Z(n1976) );
  XOR U3000 ( .A(b[705]), .B(n1977), .Z(n1978) );
  XOR U3001 ( .A(n1979), .B(n1980), .Z(n1977) );
  ANDN U3002 ( .B(n1981), .A(n329), .Z(n1979) );
  XOR U3003 ( .A(b[704]), .B(n1980), .Z(n1981) );
  XOR U3004 ( .A(n1982), .B(n1983), .Z(n1980) );
  ANDN U3005 ( .B(n1984), .A(n330), .Z(n1982) );
  XOR U3006 ( .A(b[703]), .B(n1983), .Z(n1984) );
  XOR U3007 ( .A(n1985), .B(n1986), .Z(n1983) );
  ANDN U3008 ( .B(n1987), .A(n331), .Z(n1985) );
  XOR U3009 ( .A(b[702]), .B(n1986), .Z(n1987) );
  XOR U3010 ( .A(n1988), .B(n1989), .Z(n1986) );
  ANDN U3011 ( .B(n1990), .A(n332), .Z(n1988) );
  XOR U3012 ( .A(b[701]), .B(n1989), .Z(n1990) );
  XOR U3013 ( .A(n1991), .B(n1992), .Z(n1989) );
  ANDN U3014 ( .B(n1993), .A(n333), .Z(n1991) );
  XOR U3015 ( .A(b[700]), .B(n1992), .Z(n1993) );
  XOR U3016 ( .A(n1994), .B(n1995), .Z(n1992) );
  ANDN U3017 ( .B(n1996), .A(n336), .Z(n1994) );
  XOR U3018 ( .A(b[699]), .B(n1995), .Z(n1996) );
  XOR U3019 ( .A(n1997), .B(n1998), .Z(n1995) );
  ANDN U3020 ( .B(n1999), .A(n337), .Z(n1997) );
  XOR U3021 ( .A(b[698]), .B(n1998), .Z(n1999) );
  XOR U3022 ( .A(n2000), .B(n2001), .Z(n1998) );
  ANDN U3023 ( .B(n2002), .A(n338), .Z(n2000) );
  XOR U3024 ( .A(b[697]), .B(n2001), .Z(n2002) );
  XOR U3025 ( .A(n2003), .B(n2004), .Z(n2001) );
  ANDN U3026 ( .B(n2005), .A(n339), .Z(n2003) );
  XOR U3027 ( .A(b[696]), .B(n2004), .Z(n2005) );
  XOR U3028 ( .A(n2006), .B(n2007), .Z(n2004) );
  ANDN U3029 ( .B(n2008), .A(n340), .Z(n2006) );
  XOR U3030 ( .A(b[695]), .B(n2007), .Z(n2008) );
  XOR U3031 ( .A(n2009), .B(n2010), .Z(n2007) );
  ANDN U3032 ( .B(n2011), .A(n341), .Z(n2009) );
  XOR U3033 ( .A(b[694]), .B(n2010), .Z(n2011) );
  XOR U3034 ( .A(n2012), .B(n2013), .Z(n2010) );
  ANDN U3035 ( .B(n2014), .A(n342), .Z(n2012) );
  XOR U3036 ( .A(b[693]), .B(n2013), .Z(n2014) );
  XOR U3037 ( .A(n2015), .B(n2016), .Z(n2013) );
  ANDN U3038 ( .B(n2017), .A(n343), .Z(n2015) );
  XOR U3039 ( .A(b[692]), .B(n2016), .Z(n2017) );
  XOR U3040 ( .A(n2018), .B(n2019), .Z(n2016) );
  ANDN U3041 ( .B(n2020), .A(n344), .Z(n2018) );
  XOR U3042 ( .A(b[691]), .B(n2019), .Z(n2020) );
  XOR U3043 ( .A(n2021), .B(n2022), .Z(n2019) );
  ANDN U3044 ( .B(n2023), .A(n345), .Z(n2021) );
  XOR U3045 ( .A(b[690]), .B(n2022), .Z(n2023) );
  XOR U3046 ( .A(n2024), .B(n2025), .Z(n2022) );
  ANDN U3047 ( .B(n2026), .A(n347), .Z(n2024) );
  XOR U3048 ( .A(b[689]), .B(n2025), .Z(n2026) );
  XOR U3049 ( .A(n2027), .B(n2028), .Z(n2025) );
  ANDN U3050 ( .B(n2029), .A(n348), .Z(n2027) );
  XOR U3051 ( .A(b[688]), .B(n2028), .Z(n2029) );
  XOR U3052 ( .A(n2030), .B(n2031), .Z(n2028) );
  ANDN U3053 ( .B(n2032), .A(n349), .Z(n2030) );
  XOR U3054 ( .A(b[687]), .B(n2031), .Z(n2032) );
  XOR U3055 ( .A(n2033), .B(n2034), .Z(n2031) );
  ANDN U3056 ( .B(n2035), .A(n350), .Z(n2033) );
  XOR U3057 ( .A(b[686]), .B(n2034), .Z(n2035) );
  XOR U3058 ( .A(n2036), .B(n2037), .Z(n2034) );
  ANDN U3059 ( .B(n2038), .A(n351), .Z(n2036) );
  XOR U3060 ( .A(b[685]), .B(n2037), .Z(n2038) );
  XOR U3061 ( .A(n2039), .B(n2040), .Z(n2037) );
  ANDN U3062 ( .B(n2041), .A(n352), .Z(n2039) );
  XOR U3063 ( .A(b[684]), .B(n2040), .Z(n2041) );
  XOR U3064 ( .A(n2042), .B(n2043), .Z(n2040) );
  ANDN U3065 ( .B(n2044), .A(n353), .Z(n2042) );
  XOR U3066 ( .A(b[683]), .B(n2043), .Z(n2044) );
  XOR U3067 ( .A(n2045), .B(n2046), .Z(n2043) );
  ANDN U3068 ( .B(n2047), .A(n354), .Z(n2045) );
  XOR U3069 ( .A(b[682]), .B(n2046), .Z(n2047) );
  XOR U3070 ( .A(n2048), .B(n2049), .Z(n2046) );
  ANDN U3071 ( .B(n2050), .A(n355), .Z(n2048) );
  XOR U3072 ( .A(b[681]), .B(n2049), .Z(n2050) );
  XOR U3073 ( .A(n2051), .B(n2052), .Z(n2049) );
  ANDN U3074 ( .B(n2053), .A(n356), .Z(n2051) );
  XOR U3075 ( .A(b[680]), .B(n2052), .Z(n2053) );
  XOR U3076 ( .A(n2054), .B(n2055), .Z(n2052) );
  ANDN U3077 ( .B(n2056), .A(n358), .Z(n2054) );
  XOR U3078 ( .A(b[679]), .B(n2055), .Z(n2056) );
  XOR U3079 ( .A(n2057), .B(n2058), .Z(n2055) );
  ANDN U3080 ( .B(n2059), .A(n359), .Z(n2057) );
  XOR U3081 ( .A(b[678]), .B(n2058), .Z(n2059) );
  XOR U3082 ( .A(n2060), .B(n2061), .Z(n2058) );
  ANDN U3083 ( .B(n2062), .A(n360), .Z(n2060) );
  XOR U3084 ( .A(b[677]), .B(n2061), .Z(n2062) );
  XOR U3085 ( .A(n2063), .B(n2064), .Z(n2061) );
  ANDN U3086 ( .B(n2065), .A(n361), .Z(n2063) );
  XOR U3087 ( .A(b[676]), .B(n2064), .Z(n2065) );
  XOR U3088 ( .A(n2066), .B(n2067), .Z(n2064) );
  ANDN U3089 ( .B(n2068), .A(n362), .Z(n2066) );
  XOR U3090 ( .A(b[675]), .B(n2067), .Z(n2068) );
  XOR U3091 ( .A(n2069), .B(n2070), .Z(n2067) );
  ANDN U3092 ( .B(n2071), .A(n363), .Z(n2069) );
  XOR U3093 ( .A(b[674]), .B(n2070), .Z(n2071) );
  XOR U3094 ( .A(n2072), .B(n2073), .Z(n2070) );
  ANDN U3095 ( .B(n2074), .A(n364), .Z(n2072) );
  XOR U3096 ( .A(b[673]), .B(n2073), .Z(n2074) );
  XOR U3097 ( .A(n2075), .B(n2076), .Z(n2073) );
  ANDN U3098 ( .B(n2077), .A(n365), .Z(n2075) );
  XOR U3099 ( .A(b[672]), .B(n2076), .Z(n2077) );
  XOR U3100 ( .A(n2078), .B(n2079), .Z(n2076) );
  ANDN U3101 ( .B(n2080), .A(n366), .Z(n2078) );
  XOR U3102 ( .A(b[671]), .B(n2079), .Z(n2080) );
  XOR U3103 ( .A(n2081), .B(n2082), .Z(n2079) );
  ANDN U3104 ( .B(n2083), .A(n367), .Z(n2081) );
  XOR U3105 ( .A(b[670]), .B(n2082), .Z(n2083) );
  XOR U3106 ( .A(n2084), .B(n2085), .Z(n2082) );
  ANDN U3107 ( .B(n2086), .A(n369), .Z(n2084) );
  XOR U3108 ( .A(b[669]), .B(n2085), .Z(n2086) );
  XOR U3109 ( .A(n2087), .B(n2088), .Z(n2085) );
  ANDN U3110 ( .B(n2089), .A(n370), .Z(n2087) );
  XOR U3111 ( .A(b[668]), .B(n2088), .Z(n2089) );
  XOR U3112 ( .A(n2090), .B(n2091), .Z(n2088) );
  ANDN U3113 ( .B(n2092), .A(n371), .Z(n2090) );
  XOR U3114 ( .A(b[667]), .B(n2091), .Z(n2092) );
  XOR U3115 ( .A(n2093), .B(n2094), .Z(n2091) );
  ANDN U3116 ( .B(n2095), .A(n372), .Z(n2093) );
  XOR U3117 ( .A(b[666]), .B(n2094), .Z(n2095) );
  XOR U3118 ( .A(n2096), .B(n2097), .Z(n2094) );
  ANDN U3119 ( .B(n2098), .A(n373), .Z(n2096) );
  XOR U3120 ( .A(b[665]), .B(n2097), .Z(n2098) );
  XOR U3121 ( .A(n2099), .B(n2100), .Z(n2097) );
  ANDN U3122 ( .B(n2101), .A(n374), .Z(n2099) );
  XOR U3123 ( .A(b[664]), .B(n2100), .Z(n2101) );
  XOR U3124 ( .A(n2102), .B(n2103), .Z(n2100) );
  ANDN U3125 ( .B(n2104), .A(n375), .Z(n2102) );
  XOR U3126 ( .A(b[663]), .B(n2103), .Z(n2104) );
  XOR U3127 ( .A(n2105), .B(n2106), .Z(n2103) );
  ANDN U3128 ( .B(n2107), .A(n376), .Z(n2105) );
  XOR U3129 ( .A(b[662]), .B(n2106), .Z(n2107) );
  XOR U3130 ( .A(n2108), .B(n2109), .Z(n2106) );
  ANDN U3131 ( .B(n2110), .A(n377), .Z(n2108) );
  XOR U3132 ( .A(b[661]), .B(n2109), .Z(n2110) );
  XOR U3133 ( .A(n2111), .B(n2112), .Z(n2109) );
  ANDN U3134 ( .B(n2113), .A(n378), .Z(n2111) );
  XOR U3135 ( .A(b[660]), .B(n2112), .Z(n2113) );
  XOR U3136 ( .A(n2114), .B(n2115), .Z(n2112) );
  ANDN U3137 ( .B(n2116), .A(n380), .Z(n2114) );
  XOR U3138 ( .A(b[659]), .B(n2115), .Z(n2116) );
  XOR U3139 ( .A(n2117), .B(n2118), .Z(n2115) );
  ANDN U3140 ( .B(n2119), .A(n381), .Z(n2117) );
  XOR U3141 ( .A(b[658]), .B(n2118), .Z(n2119) );
  XOR U3142 ( .A(n2120), .B(n2121), .Z(n2118) );
  ANDN U3143 ( .B(n2122), .A(n382), .Z(n2120) );
  XOR U3144 ( .A(b[657]), .B(n2121), .Z(n2122) );
  XOR U3145 ( .A(n2123), .B(n2124), .Z(n2121) );
  ANDN U3146 ( .B(n2125), .A(n383), .Z(n2123) );
  XOR U3147 ( .A(b[656]), .B(n2124), .Z(n2125) );
  XOR U3148 ( .A(n2126), .B(n2127), .Z(n2124) );
  ANDN U3149 ( .B(n2128), .A(n384), .Z(n2126) );
  XOR U3150 ( .A(b[655]), .B(n2127), .Z(n2128) );
  XOR U3151 ( .A(n2129), .B(n2130), .Z(n2127) );
  ANDN U3152 ( .B(n2131), .A(n385), .Z(n2129) );
  XOR U3153 ( .A(b[654]), .B(n2130), .Z(n2131) );
  XOR U3154 ( .A(n2132), .B(n2133), .Z(n2130) );
  ANDN U3155 ( .B(n2134), .A(n386), .Z(n2132) );
  XOR U3156 ( .A(b[653]), .B(n2133), .Z(n2134) );
  XOR U3157 ( .A(n2135), .B(n2136), .Z(n2133) );
  ANDN U3158 ( .B(n2137), .A(n387), .Z(n2135) );
  XOR U3159 ( .A(b[652]), .B(n2136), .Z(n2137) );
  XOR U3160 ( .A(n2138), .B(n2139), .Z(n2136) );
  ANDN U3161 ( .B(n2140), .A(n388), .Z(n2138) );
  XOR U3162 ( .A(b[651]), .B(n2139), .Z(n2140) );
  XOR U3163 ( .A(n2141), .B(n2142), .Z(n2139) );
  ANDN U3164 ( .B(n2143), .A(n389), .Z(n2141) );
  XOR U3165 ( .A(b[650]), .B(n2142), .Z(n2143) );
  XOR U3166 ( .A(n2144), .B(n2145), .Z(n2142) );
  ANDN U3167 ( .B(n2146), .A(n391), .Z(n2144) );
  XOR U3168 ( .A(b[649]), .B(n2145), .Z(n2146) );
  XOR U3169 ( .A(n2147), .B(n2148), .Z(n2145) );
  ANDN U3170 ( .B(n2149), .A(n392), .Z(n2147) );
  XOR U3171 ( .A(b[648]), .B(n2148), .Z(n2149) );
  XOR U3172 ( .A(n2150), .B(n2151), .Z(n2148) );
  ANDN U3173 ( .B(n2152), .A(n393), .Z(n2150) );
  XOR U3174 ( .A(b[647]), .B(n2151), .Z(n2152) );
  XOR U3175 ( .A(n2153), .B(n2154), .Z(n2151) );
  ANDN U3176 ( .B(n2155), .A(n394), .Z(n2153) );
  XOR U3177 ( .A(b[646]), .B(n2154), .Z(n2155) );
  XOR U3178 ( .A(n2156), .B(n2157), .Z(n2154) );
  ANDN U3179 ( .B(n2158), .A(n395), .Z(n2156) );
  XOR U3180 ( .A(b[645]), .B(n2157), .Z(n2158) );
  XOR U3181 ( .A(n2159), .B(n2160), .Z(n2157) );
  ANDN U3182 ( .B(n2161), .A(n396), .Z(n2159) );
  XOR U3183 ( .A(b[644]), .B(n2160), .Z(n2161) );
  XOR U3184 ( .A(n2162), .B(n2163), .Z(n2160) );
  ANDN U3185 ( .B(n2164), .A(n397), .Z(n2162) );
  XOR U3186 ( .A(b[643]), .B(n2163), .Z(n2164) );
  XOR U3187 ( .A(n2165), .B(n2166), .Z(n2163) );
  ANDN U3188 ( .B(n2167), .A(n398), .Z(n2165) );
  XOR U3189 ( .A(b[642]), .B(n2166), .Z(n2167) );
  XOR U3190 ( .A(n2168), .B(n2169), .Z(n2166) );
  ANDN U3191 ( .B(n2170), .A(n399), .Z(n2168) );
  XOR U3192 ( .A(b[641]), .B(n2169), .Z(n2170) );
  XOR U3193 ( .A(n2171), .B(n2172), .Z(n2169) );
  ANDN U3194 ( .B(n2173), .A(n400), .Z(n2171) );
  XOR U3195 ( .A(b[640]), .B(n2172), .Z(n2173) );
  XOR U3196 ( .A(n2174), .B(n2175), .Z(n2172) );
  ANDN U3197 ( .B(n2176), .A(n402), .Z(n2174) );
  XOR U3198 ( .A(b[639]), .B(n2175), .Z(n2176) );
  XOR U3199 ( .A(n2177), .B(n2178), .Z(n2175) );
  ANDN U3200 ( .B(n2179), .A(n403), .Z(n2177) );
  XOR U3201 ( .A(b[638]), .B(n2178), .Z(n2179) );
  XOR U3202 ( .A(n2180), .B(n2181), .Z(n2178) );
  ANDN U3203 ( .B(n2182), .A(n404), .Z(n2180) );
  XOR U3204 ( .A(b[637]), .B(n2181), .Z(n2182) );
  XOR U3205 ( .A(n2183), .B(n2184), .Z(n2181) );
  ANDN U3206 ( .B(n2185), .A(n405), .Z(n2183) );
  XOR U3207 ( .A(b[636]), .B(n2184), .Z(n2185) );
  XOR U3208 ( .A(n2186), .B(n2187), .Z(n2184) );
  ANDN U3209 ( .B(n2188), .A(n406), .Z(n2186) );
  XOR U3210 ( .A(b[635]), .B(n2187), .Z(n2188) );
  XOR U3211 ( .A(n2189), .B(n2190), .Z(n2187) );
  ANDN U3212 ( .B(n2191), .A(n407), .Z(n2189) );
  XOR U3213 ( .A(b[634]), .B(n2190), .Z(n2191) );
  XOR U3214 ( .A(n2192), .B(n2193), .Z(n2190) );
  ANDN U3215 ( .B(n2194), .A(n408), .Z(n2192) );
  XOR U3216 ( .A(b[633]), .B(n2193), .Z(n2194) );
  XOR U3217 ( .A(n2195), .B(n2196), .Z(n2193) );
  ANDN U3218 ( .B(n2197), .A(n409), .Z(n2195) );
  XOR U3219 ( .A(b[632]), .B(n2196), .Z(n2197) );
  XOR U3220 ( .A(n2198), .B(n2199), .Z(n2196) );
  ANDN U3221 ( .B(n2200), .A(n410), .Z(n2198) );
  XOR U3222 ( .A(b[631]), .B(n2199), .Z(n2200) );
  XOR U3223 ( .A(n2201), .B(n2202), .Z(n2199) );
  ANDN U3224 ( .B(n2203), .A(n411), .Z(n2201) );
  XOR U3225 ( .A(b[630]), .B(n2202), .Z(n2203) );
  XOR U3226 ( .A(n2204), .B(n2205), .Z(n2202) );
  ANDN U3227 ( .B(n2206), .A(n413), .Z(n2204) );
  XOR U3228 ( .A(b[629]), .B(n2205), .Z(n2206) );
  XOR U3229 ( .A(n2207), .B(n2208), .Z(n2205) );
  ANDN U3230 ( .B(n2209), .A(n414), .Z(n2207) );
  XOR U3231 ( .A(b[628]), .B(n2208), .Z(n2209) );
  XOR U3232 ( .A(n2210), .B(n2211), .Z(n2208) );
  ANDN U3233 ( .B(n2212), .A(n415), .Z(n2210) );
  XOR U3234 ( .A(b[627]), .B(n2211), .Z(n2212) );
  XOR U3235 ( .A(n2213), .B(n2214), .Z(n2211) );
  ANDN U3236 ( .B(n2215), .A(n416), .Z(n2213) );
  XOR U3237 ( .A(b[626]), .B(n2214), .Z(n2215) );
  XOR U3238 ( .A(n2216), .B(n2217), .Z(n2214) );
  ANDN U3239 ( .B(n2218), .A(n417), .Z(n2216) );
  XOR U3240 ( .A(b[625]), .B(n2217), .Z(n2218) );
  XOR U3241 ( .A(n2219), .B(n2220), .Z(n2217) );
  ANDN U3242 ( .B(n2221), .A(n418), .Z(n2219) );
  XOR U3243 ( .A(b[624]), .B(n2220), .Z(n2221) );
  XOR U3244 ( .A(n2222), .B(n2223), .Z(n2220) );
  ANDN U3245 ( .B(n2224), .A(n419), .Z(n2222) );
  XOR U3246 ( .A(b[623]), .B(n2223), .Z(n2224) );
  XOR U3247 ( .A(n2225), .B(n2226), .Z(n2223) );
  ANDN U3248 ( .B(n2227), .A(n420), .Z(n2225) );
  XOR U3249 ( .A(b[622]), .B(n2226), .Z(n2227) );
  XOR U3250 ( .A(n2228), .B(n2229), .Z(n2226) );
  ANDN U3251 ( .B(n2230), .A(n421), .Z(n2228) );
  XOR U3252 ( .A(b[621]), .B(n2229), .Z(n2230) );
  XOR U3253 ( .A(n2231), .B(n2232), .Z(n2229) );
  ANDN U3254 ( .B(n2233), .A(n422), .Z(n2231) );
  XOR U3255 ( .A(b[620]), .B(n2232), .Z(n2233) );
  XOR U3256 ( .A(n2234), .B(n2235), .Z(n2232) );
  ANDN U3257 ( .B(n2236), .A(n424), .Z(n2234) );
  XOR U3258 ( .A(b[619]), .B(n2235), .Z(n2236) );
  XOR U3259 ( .A(n2237), .B(n2238), .Z(n2235) );
  ANDN U3260 ( .B(n2239), .A(n425), .Z(n2237) );
  XOR U3261 ( .A(b[618]), .B(n2238), .Z(n2239) );
  XOR U3262 ( .A(n2240), .B(n2241), .Z(n2238) );
  ANDN U3263 ( .B(n2242), .A(n426), .Z(n2240) );
  XOR U3264 ( .A(b[617]), .B(n2241), .Z(n2242) );
  XOR U3265 ( .A(n2243), .B(n2244), .Z(n2241) );
  ANDN U3266 ( .B(n2245), .A(n427), .Z(n2243) );
  XOR U3267 ( .A(b[616]), .B(n2244), .Z(n2245) );
  XOR U3268 ( .A(n2246), .B(n2247), .Z(n2244) );
  ANDN U3269 ( .B(n2248), .A(n428), .Z(n2246) );
  XOR U3270 ( .A(b[615]), .B(n2247), .Z(n2248) );
  XOR U3271 ( .A(n2249), .B(n2250), .Z(n2247) );
  ANDN U3272 ( .B(n2251), .A(n429), .Z(n2249) );
  XOR U3273 ( .A(b[614]), .B(n2250), .Z(n2251) );
  XOR U3274 ( .A(n2252), .B(n2253), .Z(n2250) );
  ANDN U3275 ( .B(n2254), .A(n430), .Z(n2252) );
  XOR U3276 ( .A(b[613]), .B(n2253), .Z(n2254) );
  XOR U3277 ( .A(n2255), .B(n2256), .Z(n2253) );
  ANDN U3278 ( .B(n2257), .A(n431), .Z(n2255) );
  XOR U3279 ( .A(b[612]), .B(n2256), .Z(n2257) );
  XOR U3280 ( .A(n2258), .B(n2259), .Z(n2256) );
  ANDN U3281 ( .B(n2260), .A(n432), .Z(n2258) );
  XOR U3282 ( .A(b[611]), .B(n2259), .Z(n2260) );
  XOR U3283 ( .A(n2261), .B(n2262), .Z(n2259) );
  ANDN U3284 ( .B(n2263), .A(n433), .Z(n2261) );
  XOR U3285 ( .A(b[610]), .B(n2262), .Z(n2263) );
  XOR U3286 ( .A(n2264), .B(n2265), .Z(n2262) );
  ANDN U3287 ( .B(n2266), .A(n435), .Z(n2264) );
  XOR U3288 ( .A(b[609]), .B(n2265), .Z(n2266) );
  XOR U3289 ( .A(n2267), .B(n2268), .Z(n2265) );
  ANDN U3290 ( .B(n2269), .A(n436), .Z(n2267) );
  XOR U3291 ( .A(b[608]), .B(n2268), .Z(n2269) );
  XOR U3292 ( .A(n2270), .B(n2271), .Z(n2268) );
  ANDN U3293 ( .B(n2272), .A(n437), .Z(n2270) );
  XOR U3294 ( .A(b[607]), .B(n2271), .Z(n2272) );
  XOR U3295 ( .A(n2273), .B(n2274), .Z(n2271) );
  ANDN U3296 ( .B(n2275), .A(n438), .Z(n2273) );
  XOR U3297 ( .A(b[606]), .B(n2274), .Z(n2275) );
  XOR U3298 ( .A(n2276), .B(n2277), .Z(n2274) );
  ANDN U3299 ( .B(n2278), .A(n439), .Z(n2276) );
  XOR U3300 ( .A(b[605]), .B(n2277), .Z(n2278) );
  XOR U3301 ( .A(n2279), .B(n2280), .Z(n2277) );
  ANDN U3302 ( .B(n2281), .A(n440), .Z(n2279) );
  XOR U3303 ( .A(b[604]), .B(n2280), .Z(n2281) );
  XOR U3304 ( .A(n2282), .B(n2283), .Z(n2280) );
  ANDN U3305 ( .B(n2284), .A(n441), .Z(n2282) );
  XOR U3306 ( .A(b[603]), .B(n2283), .Z(n2284) );
  XOR U3307 ( .A(n2285), .B(n2286), .Z(n2283) );
  ANDN U3308 ( .B(n2287), .A(n442), .Z(n2285) );
  XOR U3309 ( .A(b[602]), .B(n2286), .Z(n2287) );
  XOR U3310 ( .A(n2288), .B(n2289), .Z(n2286) );
  ANDN U3311 ( .B(n2290), .A(n443), .Z(n2288) );
  XOR U3312 ( .A(b[601]), .B(n2289), .Z(n2290) );
  XOR U3313 ( .A(n2291), .B(n2292), .Z(n2289) );
  ANDN U3314 ( .B(n2293), .A(n444), .Z(n2291) );
  XOR U3315 ( .A(b[600]), .B(n2292), .Z(n2293) );
  XOR U3316 ( .A(n2294), .B(n2295), .Z(n2292) );
  ANDN U3317 ( .B(n2296), .A(n447), .Z(n2294) );
  XOR U3318 ( .A(b[599]), .B(n2295), .Z(n2296) );
  XOR U3319 ( .A(n2297), .B(n2298), .Z(n2295) );
  ANDN U3320 ( .B(n2299), .A(n448), .Z(n2297) );
  XOR U3321 ( .A(b[598]), .B(n2298), .Z(n2299) );
  XOR U3322 ( .A(n2300), .B(n2301), .Z(n2298) );
  ANDN U3323 ( .B(n2302), .A(n449), .Z(n2300) );
  XOR U3324 ( .A(b[597]), .B(n2301), .Z(n2302) );
  XOR U3325 ( .A(n2303), .B(n2304), .Z(n2301) );
  ANDN U3326 ( .B(n2305), .A(n450), .Z(n2303) );
  XOR U3327 ( .A(b[596]), .B(n2304), .Z(n2305) );
  XOR U3328 ( .A(n2306), .B(n2307), .Z(n2304) );
  ANDN U3329 ( .B(n2308), .A(n451), .Z(n2306) );
  XOR U3330 ( .A(b[595]), .B(n2307), .Z(n2308) );
  XOR U3331 ( .A(n2309), .B(n2310), .Z(n2307) );
  ANDN U3332 ( .B(n2311), .A(n452), .Z(n2309) );
  XOR U3333 ( .A(b[594]), .B(n2310), .Z(n2311) );
  XOR U3334 ( .A(n2312), .B(n2313), .Z(n2310) );
  ANDN U3335 ( .B(n2314), .A(n453), .Z(n2312) );
  XOR U3336 ( .A(b[593]), .B(n2313), .Z(n2314) );
  XOR U3337 ( .A(n2315), .B(n2316), .Z(n2313) );
  ANDN U3338 ( .B(n2317), .A(n454), .Z(n2315) );
  XOR U3339 ( .A(b[592]), .B(n2316), .Z(n2317) );
  XOR U3340 ( .A(n2318), .B(n2319), .Z(n2316) );
  ANDN U3341 ( .B(n2320), .A(n455), .Z(n2318) );
  XOR U3342 ( .A(b[591]), .B(n2319), .Z(n2320) );
  XOR U3343 ( .A(n2321), .B(n2322), .Z(n2319) );
  ANDN U3344 ( .B(n2323), .A(n456), .Z(n2321) );
  XOR U3345 ( .A(b[590]), .B(n2322), .Z(n2323) );
  XOR U3346 ( .A(n2324), .B(n2325), .Z(n2322) );
  ANDN U3347 ( .B(n2326), .A(n458), .Z(n2324) );
  XOR U3348 ( .A(b[589]), .B(n2325), .Z(n2326) );
  XOR U3349 ( .A(n2327), .B(n2328), .Z(n2325) );
  ANDN U3350 ( .B(n2329), .A(n459), .Z(n2327) );
  XOR U3351 ( .A(b[588]), .B(n2328), .Z(n2329) );
  XOR U3352 ( .A(n2330), .B(n2331), .Z(n2328) );
  ANDN U3353 ( .B(n2332), .A(n460), .Z(n2330) );
  XOR U3354 ( .A(b[587]), .B(n2331), .Z(n2332) );
  XOR U3355 ( .A(n2333), .B(n2334), .Z(n2331) );
  ANDN U3356 ( .B(n2335), .A(n461), .Z(n2333) );
  XOR U3357 ( .A(b[586]), .B(n2334), .Z(n2335) );
  XOR U3358 ( .A(n2336), .B(n2337), .Z(n2334) );
  ANDN U3359 ( .B(n2338), .A(n462), .Z(n2336) );
  XOR U3360 ( .A(b[585]), .B(n2337), .Z(n2338) );
  XOR U3361 ( .A(n2339), .B(n2340), .Z(n2337) );
  ANDN U3362 ( .B(n2341), .A(n463), .Z(n2339) );
  XOR U3363 ( .A(b[584]), .B(n2340), .Z(n2341) );
  XOR U3364 ( .A(n2342), .B(n2343), .Z(n2340) );
  ANDN U3365 ( .B(n2344), .A(n464), .Z(n2342) );
  XOR U3366 ( .A(b[583]), .B(n2343), .Z(n2344) );
  XOR U3367 ( .A(n2345), .B(n2346), .Z(n2343) );
  ANDN U3368 ( .B(n2347), .A(n465), .Z(n2345) );
  XOR U3369 ( .A(b[582]), .B(n2346), .Z(n2347) );
  XOR U3370 ( .A(n2348), .B(n2349), .Z(n2346) );
  ANDN U3371 ( .B(n2350), .A(n466), .Z(n2348) );
  XOR U3372 ( .A(b[581]), .B(n2349), .Z(n2350) );
  XOR U3373 ( .A(n2351), .B(n2352), .Z(n2349) );
  ANDN U3374 ( .B(n2353), .A(n467), .Z(n2351) );
  XOR U3375 ( .A(b[580]), .B(n2352), .Z(n2353) );
  XOR U3376 ( .A(n2354), .B(n2355), .Z(n2352) );
  ANDN U3377 ( .B(n2356), .A(n469), .Z(n2354) );
  XOR U3378 ( .A(b[579]), .B(n2355), .Z(n2356) );
  XOR U3379 ( .A(n2357), .B(n2358), .Z(n2355) );
  ANDN U3380 ( .B(n2359), .A(n470), .Z(n2357) );
  XOR U3381 ( .A(b[578]), .B(n2358), .Z(n2359) );
  XOR U3382 ( .A(n2360), .B(n2361), .Z(n2358) );
  ANDN U3383 ( .B(n2362), .A(n471), .Z(n2360) );
  XOR U3384 ( .A(b[577]), .B(n2361), .Z(n2362) );
  XOR U3385 ( .A(n2363), .B(n2364), .Z(n2361) );
  ANDN U3386 ( .B(n2365), .A(n472), .Z(n2363) );
  XOR U3387 ( .A(b[576]), .B(n2364), .Z(n2365) );
  XOR U3388 ( .A(n2366), .B(n2367), .Z(n2364) );
  ANDN U3389 ( .B(n2368), .A(n473), .Z(n2366) );
  XOR U3390 ( .A(b[575]), .B(n2367), .Z(n2368) );
  XOR U3391 ( .A(n2369), .B(n2370), .Z(n2367) );
  ANDN U3392 ( .B(n2371), .A(n474), .Z(n2369) );
  XOR U3393 ( .A(b[574]), .B(n2370), .Z(n2371) );
  XOR U3394 ( .A(n2372), .B(n2373), .Z(n2370) );
  ANDN U3395 ( .B(n2374), .A(n475), .Z(n2372) );
  XOR U3396 ( .A(b[573]), .B(n2373), .Z(n2374) );
  XOR U3397 ( .A(n2375), .B(n2376), .Z(n2373) );
  ANDN U3398 ( .B(n2377), .A(n476), .Z(n2375) );
  XOR U3399 ( .A(b[572]), .B(n2376), .Z(n2377) );
  XOR U3400 ( .A(n2378), .B(n2379), .Z(n2376) );
  ANDN U3401 ( .B(n2380), .A(n477), .Z(n2378) );
  XOR U3402 ( .A(b[571]), .B(n2379), .Z(n2380) );
  XOR U3403 ( .A(n2381), .B(n2382), .Z(n2379) );
  ANDN U3404 ( .B(n2383), .A(n478), .Z(n2381) );
  XOR U3405 ( .A(b[570]), .B(n2382), .Z(n2383) );
  XOR U3406 ( .A(n2384), .B(n2385), .Z(n2382) );
  ANDN U3407 ( .B(n2386), .A(n480), .Z(n2384) );
  XOR U3408 ( .A(b[569]), .B(n2385), .Z(n2386) );
  XOR U3409 ( .A(n2387), .B(n2388), .Z(n2385) );
  ANDN U3410 ( .B(n2389), .A(n481), .Z(n2387) );
  XOR U3411 ( .A(b[568]), .B(n2388), .Z(n2389) );
  XOR U3412 ( .A(n2390), .B(n2391), .Z(n2388) );
  ANDN U3413 ( .B(n2392), .A(n482), .Z(n2390) );
  XOR U3414 ( .A(b[567]), .B(n2391), .Z(n2392) );
  XOR U3415 ( .A(n2393), .B(n2394), .Z(n2391) );
  ANDN U3416 ( .B(n2395), .A(n483), .Z(n2393) );
  XOR U3417 ( .A(b[566]), .B(n2394), .Z(n2395) );
  XOR U3418 ( .A(n2396), .B(n2397), .Z(n2394) );
  ANDN U3419 ( .B(n2398), .A(n484), .Z(n2396) );
  XOR U3420 ( .A(b[565]), .B(n2397), .Z(n2398) );
  XOR U3421 ( .A(n2399), .B(n2400), .Z(n2397) );
  ANDN U3422 ( .B(n2401), .A(n485), .Z(n2399) );
  XOR U3423 ( .A(b[564]), .B(n2400), .Z(n2401) );
  XOR U3424 ( .A(n2402), .B(n2403), .Z(n2400) );
  ANDN U3425 ( .B(n2404), .A(n486), .Z(n2402) );
  XOR U3426 ( .A(b[563]), .B(n2403), .Z(n2404) );
  XOR U3427 ( .A(n2405), .B(n2406), .Z(n2403) );
  ANDN U3428 ( .B(n2407), .A(n487), .Z(n2405) );
  XOR U3429 ( .A(b[562]), .B(n2406), .Z(n2407) );
  XOR U3430 ( .A(n2408), .B(n2409), .Z(n2406) );
  ANDN U3431 ( .B(n2410), .A(n488), .Z(n2408) );
  XOR U3432 ( .A(b[561]), .B(n2409), .Z(n2410) );
  XOR U3433 ( .A(n2411), .B(n2412), .Z(n2409) );
  ANDN U3434 ( .B(n2413), .A(n489), .Z(n2411) );
  XOR U3435 ( .A(b[560]), .B(n2412), .Z(n2413) );
  XOR U3436 ( .A(n2414), .B(n2415), .Z(n2412) );
  ANDN U3437 ( .B(n2416), .A(n491), .Z(n2414) );
  XOR U3438 ( .A(b[559]), .B(n2415), .Z(n2416) );
  XOR U3439 ( .A(n2417), .B(n2418), .Z(n2415) );
  ANDN U3440 ( .B(n2419), .A(n492), .Z(n2417) );
  XOR U3441 ( .A(b[558]), .B(n2418), .Z(n2419) );
  XOR U3442 ( .A(n2420), .B(n2421), .Z(n2418) );
  ANDN U3443 ( .B(n2422), .A(n493), .Z(n2420) );
  XOR U3444 ( .A(b[557]), .B(n2421), .Z(n2422) );
  XOR U3445 ( .A(n2423), .B(n2424), .Z(n2421) );
  ANDN U3446 ( .B(n2425), .A(n494), .Z(n2423) );
  XOR U3447 ( .A(b[556]), .B(n2424), .Z(n2425) );
  XOR U3448 ( .A(n2426), .B(n2427), .Z(n2424) );
  ANDN U3449 ( .B(n2428), .A(n495), .Z(n2426) );
  XOR U3450 ( .A(b[555]), .B(n2427), .Z(n2428) );
  XOR U3451 ( .A(n2429), .B(n2430), .Z(n2427) );
  ANDN U3452 ( .B(n2431), .A(n496), .Z(n2429) );
  XOR U3453 ( .A(b[554]), .B(n2430), .Z(n2431) );
  XOR U3454 ( .A(n2432), .B(n2433), .Z(n2430) );
  ANDN U3455 ( .B(n2434), .A(n497), .Z(n2432) );
  XOR U3456 ( .A(b[553]), .B(n2433), .Z(n2434) );
  XOR U3457 ( .A(n2435), .B(n2436), .Z(n2433) );
  ANDN U3458 ( .B(n2437), .A(n498), .Z(n2435) );
  XOR U3459 ( .A(b[552]), .B(n2436), .Z(n2437) );
  XOR U3460 ( .A(n2438), .B(n2439), .Z(n2436) );
  ANDN U3461 ( .B(n2440), .A(n499), .Z(n2438) );
  XOR U3462 ( .A(b[551]), .B(n2439), .Z(n2440) );
  XOR U3463 ( .A(n2441), .B(n2442), .Z(n2439) );
  ANDN U3464 ( .B(n2443), .A(n500), .Z(n2441) );
  XOR U3465 ( .A(b[550]), .B(n2442), .Z(n2443) );
  XOR U3466 ( .A(n2444), .B(n2445), .Z(n2442) );
  ANDN U3467 ( .B(n2446), .A(n502), .Z(n2444) );
  XOR U3468 ( .A(b[549]), .B(n2445), .Z(n2446) );
  XOR U3469 ( .A(n2447), .B(n2448), .Z(n2445) );
  ANDN U3470 ( .B(n2449), .A(n503), .Z(n2447) );
  XOR U3471 ( .A(b[548]), .B(n2448), .Z(n2449) );
  XOR U3472 ( .A(n2450), .B(n2451), .Z(n2448) );
  ANDN U3473 ( .B(n2452), .A(n504), .Z(n2450) );
  XOR U3474 ( .A(b[547]), .B(n2451), .Z(n2452) );
  XOR U3475 ( .A(n2453), .B(n2454), .Z(n2451) );
  ANDN U3476 ( .B(n2455), .A(n505), .Z(n2453) );
  XOR U3477 ( .A(b[546]), .B(n2454), .Z(n2455) );
  XOR U3478 ( .A(n2456), .B(n2457), .Z(n2454) );
  ANDN U3479 ( .B(n2458), .A(n506), .Z(n2456) );
  XOR U3480 ( .A(b[545]), .B(n2457), .Z(n2458) );
  XOR U3481 ( .A(n2459), .B(n2460), .Z(n2457) );
  ANDN U3482 ( .B(n2461), .A(n507), .Z(n2459) );
  XOR U3483 ( .A(b[544]), .B(n2460), .Z(n2461) );
  XOR U3484 ( .A(n2462), .B(n2463), .Z(n2460) );
  ANDN U3485 ( .B(n2464), .A(n508), .Z(n2462) );
  XOR U3486 ( .A(b[543]), .B(n2463), .Z(n2464) );
  XOR U3487 ( .A(n2465), .B(n2466), .Z(n2463) );
  ANDN U3488 ( .B(n2467), .A(n509), .Z(n2465) );
  XOR U3489 ( .A(b[542]), .B(n2466), .Z(n2467) );
  XOR U3490 ( .A(n2468), .B(n2469), .Z(n2466) );
  ANDN U3491 ( .B(n2470), .A(n510), .Z(n2468) );
  XOR U3492 ( .A(b[541]), .B(n2469), .Z(n2470) );
  XOR U3493 ( .A(n2471), .B(n2472), .Z(n2469) );
  ANDN U3494 ( .B(n2473), .A(n511), .Z(n2471) );
  XOR U3495 ( .A(b[540]), .B(n2472), .Z(n2473) );
  XOR U3496 ( .A(n2474), .B(n2475), .Z(n2472) );
  ANDN U3497 ( .B(n2476), .A(n513), .Z(n2474) );
  XOR U3498 ( .A(b[539]), .B(n2475), .Z(n2476) );
  XOR U3499 ( .A(n2477), .B(n2478), .Z(n2475) );
  ANDN U3500 ( .B(n2479), .A(n514), .Z(n2477) );
  XOR U3501 ( .A(b[538]), .B(n2478), .Z(n2479) );
  XOR U3502 ( .A(n2480), .B(n2481), .Z(n2478) );
  ANDN U3503 ( .B(n2482), .A(n515), .Z(n2480) );
  XOR U3504 ( .A(b[537]), .B(n2481), .Z(n2482) );
  XOR U3505 ( .A(n2483), .B(n2484), .Z(n2481) );
  ANDN U3506 ( .B(n2485), .A(n516), .Z(n2483) );
  XOR U3507 ( .A(b[536]), .B(n2484), .Z(n2485) );
  XOR U3508 ( .A(n2486), .B(n2487), .Z(n2484) );
  ANDN U3509 ( .B(n2488), .A(n517), .Z(n2486) );
  XOR U3510 ( .A(b[535]), .B(n2487), .Z(n2488) );
  XOR U3511 ( .A(n2489), .B(n2490), .Z(n2487) );
  ANDN U3512 ( .B(n2491), .A(n518), .Z(n2489) );
  XOR U3513 ( .A(b[534]), .B(n2490), .Z(n2491) );
  XOR U3514 ( .A(n2492), .B(n2493), .Z(n2490) );
  ANDN U3515 ( .B(n2494), .A(n519), .Z(n2492) );
  XOR U3516 ( .A(b[533]), .B(n2493), .Z(n2494) );
  XOR U3517 ( .A(n2495), .B(n2496), .Z(n2493) );
  ANDN U3518 ( .B(n2497), .A(n520), .Z(n2495) );
  XOR U3519 ( .A(b[532]), .B(n2496), .Z(n2497) );
  XOR U3520 ( .A(n2498), .B(n2499), .Z(n2496) );
  ANDN U3521 ( .B(n2500), .A(n521), .Z(n2498) );
  XOR U3522 ( .A(b[531]), .B(n2499), .Z(n2500) );
  XOR U3523 ( .A(n2501), .B(n2502), .Z(n2499) );
  ANDN U3524 ( .B(n2503), .A(n522), .Z(n2501) );
  XOR U3525 ( .A(b[530]), .B(n2502), .Z(n2503) );
  XOR U3526 ( .A(n2504), .B(n2505), .Z(n2502) );
  ANDN U3527 ( .B(n2506), .A(n524), .Z(n2504) );
  XOR U3528 ( .A(b[529]), .B(n2505), .Z(n2506) );
  XOR U3529 ( .A(n2507), .B(n2508), .Z(n2505) );
  ANDN U3530 ( .B(n2509), .A(n525), .Z(n2507) );
  XOR U3531 ( .A(b[528]), .B(n2508), .Z(n2509) );
  XOR U3532 ( .A(n2510), .B(n2511), .Z(n2508) );
  ANDN U3533 ( .B(n2512), .A(n526), .Z(n2510) );
  XOR U3534 ( .A(b[527]), .B(n2511), .Z(n2512) );
  XOR U3535 ( .A(n2513), .B(n2514), .Z(n2511) );
  ANDN U3536 ( .B(n2515), .A(n527), .Z(n2513) );
  XOR U3537 ( .A(b[526]), .B(n2514), .Z(n2515) );
  XOR U3538 ( .A(n2516), .B(n2517), .Z(n2514) );
  ANDN U3539 ( .B(n2518), .A(n528), .Z(n2516) );
  XOR U3540 ( .A(b[525]), .B(n2517), .Z(n2518) );
  XOR U3541 ( .A(n2519), .B(n2520), .Z(n2517) );
  ANDN U3542 ( .B(n2521), .A(n529), .Z(n2519) );
  XOR U3543 ( .A(b[524]), .B(n2520), .Z(n2521) );
  XOR U3544 ( .A(n2522), .B(n2523), .Z(n2520) );
  ANDN U3545 ( .B(n2524), .A(n530), .Z(n2522) );
  XOR U3546 ( .A(b[523]), .B(n2523), .Z(n2524) );
  XOR U3547 ( .A(n2525), .B(n2526), .Z(n2523) );
  ANDN U3548 ( .B(n2527), .A(n531), .Z(n2525) );
  XOR U3549 ( .A(b[522]), .B(n2526), .Z(n2527) );
  XOR U3550 ( .A(n2528), .B(n2529), .Z(n2526) );
  ANDN U3551 ( .B(n2530), .A(n532), .Z(n2528) );
  XOR U3552 ( .A(b[521]), .B(n2529), .Z(n2530) );
  XOR U3553 ( .A(n2531), .B(n2532), .Z(n2529) );
  ANDN U3554 ( .B(n2533), .A(n533), .Z(n2531) );
  XOR U3555 ( .A(b[520]), .B(n2532), .Z(n2533) );
  XOR U3556 ( .A(n2534), .B(n2535), .Z(n2532) );
  ANDN U3557 ( .B(n2536), .A(n535), .Z(n2534) );
  XOR U3558 ( .A(b[519]), .B(n2535), .Z(n2536) );
  XOR U3559 ( .A(n2537), .B(n2538), .Z(n2535) );
  ANDN U3560 ( .B(n2539), .A(n536), .Z(n2537) );
  XOR U3561 ( .A(b[518]), .B(n2538), .Z(n2539) );
  XOR U3562 ( .A(n2540), .B(n2541), .Z(n2538) );
  ANDN U3563 ( .B(n2542), .A(n537), .Z(n2540) );
  XOR U3564 ( .A(b[517]), .B(n2541), .Z(n2542) );
  XOR U3565 ( .A(n2543), .B(n2544), .Z(n2541) );
  ANDN U3566 ( .B(n2545), .A(n538), .Z(n2543) );
  XOR U3567 ( .A(b[516]), .B(n2544), .Z(n2545) );
  XOR U3568 ( .A(n2546), .B(n2547), .Z(n2544) );
  ANDN U3569 ( .B(n2548), .A(n539), .Z(n2546) );
  XOR U3570 ( .A(b[515]), .B(n2547), .Z(n2548) );
  XOR U3571 ( .A(n2549), .B(n2550), .Z(n2547) );
  ANDN U3572 ( .B(n2551), .A(n540), .Z(n2549) );
  XOR U3573 ( .A(b[514]), .B(n2550), .Z(n2551) );
  XOR U3574 ( .A(n2552), .B(n2553), .Z(n2550) );
  ANDN U3575 ( .B(n2554), .A(n541), .Z(n2552) );
  XOR U3576 ( .A(b[513]), .B(n2553), .Z(n2554) );
  XOR U3577 ( .A(n2555), .B(n2556), .Z(n2553) );
  ANDN U3578 ( .B(n2557), .A(n542), .Z(n2555) );
  XOR U3579 ( .A(b[512]), .B(n2556), .Z(n2557) );
  XOR U3580 ( .A(n2558), .B(n2559), .Z(n2556) );
  ANDN U3581 ( .B(n2560), .A(n543), .Z(n2558) );
  XOR U3582 ( .A(b[511]), .B(n2559), .Z(n2560) );
  XOR U3583 ( .A(n2561), .B(n2562), .Z(n2559) );
  ANDN U3584 ( .B(n2563), .A(n544), .Z(n2561) );
  XOR U3585 ( .A(b[510]), .B(n2562), .Z(n2563) );
  XOR U3586 ( .A(n2564), .B(n2565), .Z(n2562) );
  ANDN U3587 ( .B(n2566), .A(n546), .Z(n2564) );
  XOR U3588 ( .A(b[509]), .B(n2565), .Z(n2566) );
  XOR U3589 ( .A(n2567), .B(n2568), .Z(n2565) );
  ANDN U3590 ( .B(n2569), .A(n547), .Z(n2567) );
  XOR U3591 ( .A(b[508]), .B(n2568), .Z(n2569) );
  XOR U3592 ( .A(n2570), .B(n2571), .Z(n2568) );
  ANDN U3593 ( .B(n2572), .A(n548), .Z(n2570) );
  XOR U3594 ( .A(b[507]), .B(n2571), .Z(n2572) );
  XOR U3595 ( .A(n2573), .B(n2574), .Z(n2571) );
  ANDN U3596 ( .B(n2575), .A(n549), .Z(n2573) );
  XOR U3597 ( .A(b[506]), .B(n2574), .Z(n2575) );
  XOR U3598 ( .A(n2576), .B(n2577), .Z(n2574) );
  ANDN U3599 ( .B(n2578), .A(n550), .Z(n2576) );
  XOR U3600 ( .A(b[505]), .B(n2577), .Z(n2578) );
  XOR U3601 ( .A(n2579), .B(n2580), .Z(n2577) );
  ANDN U3602 ( .B(n2581), .A(n551), .Z(n2579) );
  XOR U3603 ( .A(b[504]), .B(n2580), .Z(n2581) );
  XOR U3604 ( .A(n2582), .B(n2583), .Z(n2580) );
  ANDN U3605 ( .B(n2584), .A(n552), .Z(n2582) );
  XOR U3606 ( .A(b[503]), .B(n2583), .Z(n2584) );
  XOR U3607 ( .A(n2585), .B(n2586), .Z(n2583) );
  ANDN U3608 ( .B(n2587), .A(n553), .Z(n2585) );
  XOR U3609 ( .A(b[502]), .B(n2586), .Z(n2587) );
  XOR U3610 ( .A(n2588), .B(n2589), .Z(n2586) );
  ANDN U3611 ( .B(n2590), .A(n554), .Z(n2588) );
  XOR U3612 ( .A(b[501]), .B(n2589), .Z(n2590) );
  XOR U3613 ( .A(n2591), .B(n2592), .Z(n2589) );
  ANDN U3614 ( .B(n2593), .A(n555), .Z(n2591) );
  XOR U3615 ( .A(b[500]), .B(n2592), .Z(n2593) );
  XOR U3616 ( .A(n2594), .B(n2595), .Z(n2592) );
  ANDN U3617 ( .B(n2596), .A(n558), .Z(n2594) );
  XOR U3618 ( .A(b[499]), .B(n2595), .Z(n2596) );
  XOR U3619 ( .A(n2597), .B(n2598), .Z(n2595) );
  ANDN U3620 ( .B(n2599), .A(n559), .Z(n2597) );
  XOR U3621 ( .A(b[498]), .B(n2598), .Z(n2599) );
  XOR U3622 ( .A(n2600), .B(n2601), .Z(n2598) );
  ANDN U3623 ( .B(n2602), .A(n560), .Z(n2600) );
  XOR U3624 ( .A(b[497]), .B(n2601), .Z(n2602) );
  XOR U3625 ( .A(n2603), .B(n2604), .Z(n2601) );
  ANDN U3626 ( .B(n2605), .A(n561), .Z(n2603) );
  XOR U3627 ( .A(b[496]), .B(n2604), .Z(n2605) );
  XOR U3628 ( .A(n2606), .B(n2607), .Z(n2604) );
  ANDN U3629 ( .B(n2608), .A(n562), .Z(n2606) );
  XOR U3630 ( .A(b[495]), .B(n2607), .Z(n2608) );
  XOR U3631 ( .A(n2609), .B(n2610), .Z(n2607) );
  ANDN U3632 ( .B(n2611), .A(n563), .Z(n2609) );
  XOR U3633 ( .A(b[494]), .B(n2610), .Z(n2611) );
  XOR U3634 ( .A(n2612), .B(n2613), .Z(n2610) );
  ANDN U3635 ( .B(n2614), .A(n564), .Z(n2612) );
  XOR U3636 ( .A(b[493]), .B(n2613), .Z(n2614) );
  XOR U3637 ( .A(n2615), .B(n2616), .Z(n2613) );
  ANDN U3638 ( .B(n2617), .A(n565), .Z(n2615) );
  XOR U3639 ( .A(b[492]), .B(n2616), .Z(n2617) );
  XOR U3640 ( .A(n2618), .B(n2619), .Z(n2616) );
  ANDN U3641 ( .B(n2620), .A(n566), .Z(n2618) );
  XOR U3642 ( .A(b[491]), .B(n2619), .Z(n2620) );
  XOR U3643 ( .A(n2621), .B(n2622), .Z(n2619) );
  ANDN U3644 ( .B(n2623), .A(n567), .Z(n2621) );
  XOR U3645 ( .A(b[490]), .B(n2622), .Z(n2623) );
  XOR U3646 ( .A(n2624), .B(n2625), .Z(n2622) );
  ANDN U3647 ( .B(n2626), .A(n569), .Z(n2624) );
  XOR U3648 ( .A(b[489]), .B(n2625), .Z(n2626) );
  XOR U3649 ( .A(n2627), .B(n2628), .Z(n2625) );
  ANDN U3650 ( .B(n2629), .A(n570), .Z(n2627) );
  XOR U3651 ( .A(b[488]), .B(n2628), .Z(n2629) );
  XOR U3652 ( .A(n2630), .B(n2631), .Z(n2628) );
  ANDN U3653 ( .B(n2632), .A(n571), .Z(n2630) );
  XOR U3654 ( .A(b[487]), .B(n2631), .Z(n2632) );
  XOR U3655 ( .A(n2633), .B(n2634), .Z(n2631) );
  ANDN U3656 ( .B(n2635), .A(n572), .Z(n2633) );
  XOR U3657 ( .A(b[486]), .B(n2634), .Z(n2635) );
  XOR U3658 ( .A(n2636), .B(n2637), .Z(n2634) );
  ANDN U3659 ( .B(n2638), .A(n573), .Z(n2636) );
  XOR U3660 ( .A(b[485]), .B(n2637), .Z(n2638) );
  XOR U3661 ( .A(n2639), .B(n2640), .Z(n2637) );
  ANDN U3662 ( .B(n2641), .A(n574), .Z(n2639) );
  XOR U3663 ( .A(b[484]), .B(n2640), .Z(n2641) );
  XOR U3664 ( .A(n2642), .B(n2643), .Z(n2640) );
  ANDN U3665 ( .B(n2644), .A(n575), .Z(n2642) );
  XOR U3666 ( .A(b[483]), .B(n2643), .Z(n2644) );
  XOR U3667 ( .A(n2645), .B(n2646), .Z(n2643) );
  ANDN U3668 ( .B(n2647), .A(n576), .Z(n2645) );
  XOR U3669 ( .A(b[482]), .B(n2646), .Z(n2647) );
  XOR U3670 ( .A(n2648), .B(n2649), .Z(n2646) );
  ANDN U3671 ( .B(n2650), .A(n577), .Z(n2648) );
  XOR U3672 ( .A(b[481]), .B(n2649), .Z(n2650) );
  XOR U3673 ( .A(n2651), .B(n2652), .Z(n2649) );
  ANDN U3674 ( .B(n2653), .A(n578), .Z(n2651) );
  XOR U3675 ( .A(b[480]), .B(n2652), .Z(n2653) );
  XOR U3676 ( .A(n2654), .B(n2655), .Z(n2652) );
  ANDN U3677 ( .B(n2656), .A(n580), .Z(n2654) );
  XOR U3678 ( .A(b[479]), .B(n2655), .Z(n2656) );
  XOR U3679 ( .A(n2657), .B(n2658), .Z(n2655) );
  ANDN U3680 ( .B(n2659), .A(n581), .Z(n2657) );
  XOR U3681 ( .A(b[478]), .B(n2658), .Z(n2659) );
  XOR U3682 ( .A(n2660), .B(n2661), .Z(n2658) );
  ANDN U3683 ( .B(n2662), .A(n582), .Z(n2660) );
  XOR U3684 ( .A(b[477]), .B(n2661), .Z(n2662) );
  XOR U3685 ( .A(n2663), .B(n2664), .Z(n2661) );
  ANDN U3686 ( .B(n2665), .A(n583), .Z(n2663) );
  XOR U3687 ( .A(b[476]), .B(n2664), .Z(n2665) );
  XOR U3688 ( .A(n2666), .B(n2667), .Z(n2664) );
  ANDN U3689 ( .B(n2668), .A(n584), .Z(n2666) );
  XOR U3690 ( .A(b[475]), .B(n2667), .Z(n2668) );
  XOR U3691 ( .A(n2669), .B(n2670), .Z(n2667) );
  ANDN U3692 ( .B(n2671), .A(n585), .Z(n2669) );
  XOR U3693 ( .A(b[474]), .B(n2670), .Z(n2671) );
  XOR U3694 ( .A(n2672), .B(n2673), .Z(n2670) );
  ANDN U3695 ( .B(n2674), .A(n586), .Z(n2672) );
  XOR U3696 ( .A(b[473]), .B(n2673), .Z(n2674) );
  XOR U3697 ( .A(n2675), .B(n2676), .Z(n2673) );
  ANDN U3698 ( .B(n2677), .A(n587), .Z(n2675) );
  XOR U3699 ( .A(b[472]), .B(n2676), .Z(n2677) );
  XOR U3700 ( .A(n2678), .B(n2679), .Z(n2676) );
  ANDN U3701 ( .B(n2680), .A(n588), .Z(n2678) );
  XOR U3702 ( .A(b[471]), .B(n2679), .Z(n2680) );
  XOR U3703 ( .A(n2681), .B(n2682), .Z(n2679) );
  ANDN U3704 ( .B(n2683), .A(n589), .Z(n2681) );
  XOR U3705 ( .A(b[470]), .B(n2682), .Z(n2683) );
  XOR U3706 ( .A(n2684), .B(n2685), .Z(n2682) );
  ANDN U3707 ( .B(n2686), .A(n591), .Z(n2684) );
  XOR U3708 ( .A(b[469]), .B(n2685), .Z(n2686) );
  XOR U3709 ( .A(n2687), .B(n2688), .Z(n2685) );
  ANDN U3710 ( .B(n2689), .A(n592), .Z(n2687) );
  XOR U3711 ( .A(b[468]), .B(n2688), .Z(n2689) );
  XOR U3712 ( .A(n2690), .B(n2691), .Z(n2688) );
  ANDN U3713 ( .B(n2692), .A(n593), .Z(n2690) );
  XOR U3714 ( .A(b[467]), .B(n2691), .Z(n2692) );
  XOR U3715 ( .A(n2693), .B(n2694), .Z(n2691) );
  ANDN U3716 ( .B(n2695), .A(n594), .Z(n2693) );
  XOR U3717 ( .A(b[466]), .B(n2694), .Z(n2695) );
  XOR U3718 ( .A(n2696), .B(n2697), .Z(n2694) );
  ANDN U3719 ( .B(n2698), .A(n595), .Z(n2696) );
  XOR U3720 ( .A(b[465]), .B(n2697), .Z(n2698) );
  XOR U3721 ( .A(n2699), .B(n2700), .Z(n2697) );
  ANDN U3722 ( .B(n2701), .A(n596), .Z(n2699) );
  XOR U3723 ( .A(b[464]), .B(n2700), .Z(n2701) );
  XOR U3724 ( .A(n2702), .B(n2703), .Z(n2700) );
  ANDN U3725 ( .B(n2704), .A(n597), .Z(n2702) );
  XOR U3726 ( .A(b[463]), .B(n2703), .Z(n2704) );
  XOR U3727 ( .A(n2705), .B(n2706), .Z(n2703) );
  ANDN U3728 ( .B(n2707), .A(n598), .Z(n2705) );
  XOR U3729 ( .A(b[462]), .B(n2706), .Z(n2707) );
  XOR U3730 ( .A(n2708), .B(n2709), .Z(n2706) );
  ANDN U3731 ( .B(n2710), .A(n599), .Z(n2708) );
  XOR U3732 ( .A(b[461]), .B(n2709), .Z(n2710) );
  XOR U3733 ( .A(n2711), .B(n2712), .Z(n2709) );
  ANDN U3734 ( .B(n2713), .A(n600), .Z(n2711) );
  XOR U3735 ( .A(b[460]), .B(n2712), .Z(n2713) );
  XOR U3736 ( .A(n2714), .B(n2715), .Z(n2712) );
  ANDN U3737 ( .B(n2716), .A(n602), .Z(n2714) );
  XOR U3738 ( .A(b[459]), .B(n2715), .Z(n2716) );
  XOR U3739 ( .A(n2717), .B(n2718), .Z(n2715) );
  ANDN U3740 ( .B(n2719), .A(n603), .Z(n2717) );
  XOR U3741 ( .A(b[458]), .B(n2718), .Z(n2719) );
  XOR U3742 ( .A(n2720), .B(n2721), .Z(n2718) );
  ANDN U3743 ( .B(n2722), .A(n604), .Z(n2720) );
  XOR U3744 ( .A(b[457]), .B(n2721), .Z(n2722) );
  XOR U3745 ( .A(n2723), .B(n2724), .Z(n2721) );
  ANDN U3746 ( .B(n2725), .A(n605), .Z(n2723) );
  XOR U3747 ( .A(b[456]), .B(n2724), .Z(n2725) );
  XOR U3748 ( .A(n2726), .B(n2727), .Z(n2724) );
  ANDN U3749 ( .B(n2728), .A(n606), .Z(n2726) );
  XOR U3750 ( .A(b[455]), .B(n2727), .Z(n2728) );
  XOR U3751 ( .A(n2729), .B(n2730), .Z(n2727) );
  ANDN U3752 ( .B(n2731), .A(n607), .Z(n2729) );
  XOR U3753 ( .A(b[454]), .B(n2730), .Z(n2731) );
  XOR U3754 ( .A(n2732), .B(n2733), .Z(n2730) );
  ANDN U3755 ( .B(n2734), .A(n608), .Z(n2732) );
  XOR U3756 ( .A(b[453]), .B(n2733), .Z(n2734) );
  XOR U3757 ( .A(n2735), .B(n2736), .Z(n2733) );
  ANDN U3758 ( .B(n2737), .A(n609), .Z(n2735) );
  XOR U3759 ( .A(b[452]), .B(n2736), .Z(n2737) );
  XOR U3760 ( .A(n2738), .B(n2739), .Z(n2736) );
  ANDN U3761 ( .B(n2740), .A(n610), .Z(n2738) );
  XOR U3762 ( .A(b[451]), .B(n2739), .Z(n2740) );
  XOR U3763 ( .A(n2741), .B(n2742), .Z(n2739) );
  ANDN U3764 ( .B(n2743), .A(n611), .Z(n2741) );
  XOR U3765 ( .A(b[450]), .B(n2742), .Z(n2743) );
  XOR U3766 ( .A(n2744), .B(n2745), .Z(n2742) );
  ANDN U3767 ( .B(n2746), .A(n613), .Z(n2744) );
  XOR U3768 ( .A(b[449]), .B(n2745), .Z(n2746) );
  XOR U3769 ( .A(n2747), .B(n2748), .Z(n2745) );
  ANDN U3770 ( .B(n2749), .A(n614), .Z(n2747) );
  XOR U3771 ( .A(b[448]), .B(n2748), .Z(n2749) );
  XOR U3772 ( .A(n2750), .B(n2751), .Z(n2748) );
  ANDN U3773 ( .B(n2752), .A(n615), .Z(n2750) );
  XOR U3774 ( .A(b[447]), .B(n2751), .Z(n2752) );
  XOR U3775 ( .A(n2753), .B(n2754), .Z(n2751) );
  ANDN U3776 ( .B(n2755), .A(n616), .Z(n2753) );
  XOR U3777 ( .A(b[446]), .B(n2754), .Z(n2755) );
  XOR U3778 ( .A(n2756), .B(n2757), .Z(n2754) );
  ANDN U3779 ( .B(n2758), .A(n617), .Z(n2756) );
  XOR U3780 ( .A(b[445]), .B(n2757), .Z(n2758) );
  XOR U3781 ( .A(n2759), .B(n2760), .Z(n2757) );
  ANDN U3782 ( .B(n2761), .A(n618), .Z(n2759) );
  XOR U3783 ( .A(b[444]), .B(n2760), .Z(n2761) );
  XOR U3784 ( .A(n2762), .B(n2763), .Z(n2760) );
  ANDN U3785 ( .B(n2764), .A(n619), .Z(n2762) );
  XOR U3786 ( .A(b[443]), .B(n2763), .Z(n2764) );
  XOR U3787 ( .A(n2765), .B(n2766), .Z(n2763) );
  ANDN U3788 ( .B(n2767), .A(n620), .Z(n2765) );
  XOR U3789 ( .A(b[442]), .B(n2766), .Z(n2767) );
  XOR U3790 ( .A(n2768), .B(n2769), .Z(n2766) );
  ANDN U3791 ( .B(n2770), .A(n621), .Z(n2768) );
  XOR U3792 ( .A(b[441]), .B(n2769), .Z(n2770) );
  XOR U3793 ( .A(n2771), .B(n2772), .Z(n2769) );
  ANDN U3794 ( .B(n2773), .A(n622), .Z(n2771) );
  XOR U3795 ( .A(b[440]), .B(n2772), .Z(n2773) );
  XOR U3796 ( .A(n2774), .B(n2775), .Z(n2772) );
  ANDN U3797 ( .B(n2776), .A(n624), .Z(n2774) );
  XOR U3798 ( .A(b[439]), .B(n2775), .Z(n2776) );
  XOR U3799 ( .A(n2777), .B(n2778), .Z(n2775) );
  ANDN U3800 ( .B(n2779), .A(n625), .Z(n2777) );
  XOR U3801 ( .A(b[438]), .B(n2778), .Z(n2779) );
  XOR U3802 ( .A(n2780), .B(n2781), .Z(n2778) );
  ANDN U3803 ( .B(n2782), .A(n626), .Z(n2780) );
  XOR U3804 ( .A(b[437]), .B(n2781), .Z(n2782) );
  XOR U3805 ( .A(n2783), .B(n2784), .Z(n2781) );
  ANDN U3806 ( .B(n2785), .A(n627), .Z(n2783) );
  XOR U3807 ( .A(b[436]), .B(n2784), .Z(n2785) );
  XOR U3808 ( .A(n2786), .B(n2787), .Z(n2784) );
  ANDN U3809 ( .B(n2788), .A(n628), .Z(n2786) );
  XOR U3810 ( .A(b[435]), .B(n2787), .Z(n2788) );
  XOR U3811 ( .A(n2789), .B(n2790), .Z(n2787) );
  ANDN U3812 ( .B(n2791), .A(n629), .Z(n2789) );
  XOR U3813 ( .A(b[434]), .B(n2790), .Z(n2791) );
  XOR U3814 ( .A(n2792), .B(n2793), .Z(n2790) );
  ANDN U3815 ( .B(n2794), .A(n630), .Z(n2792) );
  XOR U3816 ( .A(b[433]), .B(n2793), .Z(n2794) );
  XOR U3817 ( .A(n2795), .B(n2796), .Z(n2793) );
  ANDN U3818 ( .B(n2797), .A(n631), .Z(n2795) );
  XOR U3819 ( .A(b[432]), .B(n2796), .Z(n2797) );
  XOR U3820 ( .A(n2798), .B(n2799), .Z(n2796) );
  ANDN U3821 ( .B(n2800), .A(n632), .Z(n2798) );
  XOR U3822 ( .A(b[431]), .B(n2799), .Z(n2800) );
  XOR U3823 ( .A(n2801), .B(n2802), .Z(n2799) );
  ANDN U3824 ( .B(n2803), .A(n633), .Z(n2801) );
  XOR U3825 ( .A(b[430]), .B(n2802), .Z(n2803) );
  XOR U3826 ( .A(n2804), .B(n2805), .Z(n2802) );
  ANDN U3827 ( .B(n2806), .A(n635), .Z(n2804) );
  XOR U3828 ( .A(b[429]), .B(n2805), .Z(n2806) );
  XOR U3829 ( .A(n2807), .B(n2808), .Z(n2805) );
  ANDN U3830 ( .B(n2809), .A(n636), .Z(n2807) );
  XOR U3831 ( .A(b[428]), .B(n2808), .Z(n2809) );
  XOR U3832 ( .A(n2810), .B(n2811), .Z(n2808) );
  ANDN U3833 ( .B(n2812), .A(n637), .Z(n2810) );
  XOR U3834 ( .A(b[427]), .B(n2811), .Z(n2812) );
  XOR U3835 ( .A(n2813), .B(n2814), .Z(n2811) );
  ANDN U3836 ( .B(n2815), .A(n638), .Z(n2813) );
  XOR U3837 ( .A(b[426]), .B(n2814), .Z(n2815) );
  XOR U3838 ( .A(n2816), .B(n2817), .Z(n2814) );
  ANDN U3839 ( .B(n2818), .A(n639), .Z(n2816) );
  XOR U3840 ( .A(b[425]), .B(n2817), .Z(n2818) );
  XOR U3841 ( .A(n2819), .B(n2820), .Z(n2817) );
  ANDN U3842 ( .B(n2821), .A(n640), .Z(n2819) );
  XOR U3843 ( .A(b[424]), .B(n2820), .Z(n2821) );
  XOR U3844 ( .A(n2822), .B(n2823), .Z(n2820) );
  ANDN U3845 ( .B(n2824), .A(n641), .Z(n2822) );
  XOR U3846 ( .A(b[423]), .B(n2823), .Z(n2824) );
  XOR U3847 ( .A(n2825), .B(n2826), .Z(n2823) );
  ANDN U3848 ( .B(n2827), .A(n642), .Z(n2825) );
  XOR U3849 ( .A(b[422]), .B(n2826), .Z(n2827) );
  XOR U3850 ( .A(n2828), .B(n2829), .Z(n2826) );
  ANDN U3851 ( .B(n2830), .A(n643), .Z(n2828) );
  XOR U3852 ( .A(b[421]), .B(n2829), .Z(n2830) );
  XOR U3853 ( .A(n2831), .B(n2832), .Z(n2829) );
  ANDN U3854 ( .B(n2833), .A(n644), .Z(n2831) );
  XOR U3855 ( .A(b[420]), .B(n2832), .Z(n2833) );
  XOR U3856 ( .A(n2834), .B(n2835), .Z(n2832) );
  ANDN U3857 ( .B(n2836), .A(n646), .Z(n2834) );
  XOR U3858 ( .A(b[419]), .B(n2835), .Z(n2836) );
  XOR U3859 ( .A(n2837), .B(n2838), .Z(n2835) );
  ANDN U3860 ( .B(n2839), .A(n647), .Z(n2837) );
  XOR U3861 ( .A(b[418]), .B(n2838), .Z(n2839) );
  XOR U3862 ( .A(n2840), .B(n2841), .Z(n2838) );
  ANDN U3863 ( .B(n2842), .A(n648), .Z(n2840) );
  XOR U3864 ( .A(b[417]), .B(n2841), .Z(n2842) );
  XOR U3865 ( .A(n2843), .B(n2844), .Z(n2841) );
  ANDN U3866 ( .B(n2845), .A(n649), .Z(n2843) );
  XOR U3867 ( .A(b[416]), .B(n2844), .Z(n2845) );
  XOR U3868 ( .A(n2846), .B(n2847), .Z(n2844) );
  ANDN U3869 ( .B(n2848), .A(n650), .Z(n2846) );
  XOR U3870 ( .A(b[415]), .B(n2847), .Z(n2848) );
  XOR U3871 ( .A(n2849), .B(n2850), .Z(n2847) );
  ANDN U3872 ( .B(n2851), .A(n651), .Z(n2849) );
  XOR U3873 ( .A(b[414]), .B(n2850), .Z(n2851) );
  XOR U3874 ( .A(n2852), .B(n2853), .Z(n2850) );
  ANDN U3875 ( .B(n2854), .A(n652), .Z(n2852) );
  XOR U3876 ( .A(b[413]), .B(n2853), .Z(n2854) );
  XOR U3877 ( .A(n2855), .B(n2856), .Z(n2853) );
  ANDN U3878 ( .B(n2857), .A(n653), .Z(n2855) );
  XOR U3879 ( .A(b[412]), .B(n2856), .Z(n2857) );
  XOR U3880 ( .A(n2858), .B(n2859), .Z(n2856) );
  ANDN U3881 ( .B(n2860), .A(n654), .Z(n2858) );
  XOR U3882 ( .A(b[411]), .B(n2859), .Z(n2860) );
  XOR U3883 ( .A(n2861), .B(n2862), .Z(n2859) );
  ANDN U3884 ( .B(n2863), .A(n655), .Z(n2861) );
  XOR U3885 ( .A(b[410]), .B(n2862), .Z(n2863) );
  XOR U3886 ( .A(n2864), .B(n2865), .Z(n2862) );
  ANDN U3887 ( .B(n2866), .A(n657), .Z(n2864) );
  XOR U3888 ( .A(b[409]), .B(n2865), .Z(n2866) );
  XOR U3889 ( .A(n2867), .B(n2868), .Z(n2865) );
  ANDN U3890 ( .B(n2869), .A(n658), .Z(n2867) );
  XOR U3891 ( .A(b[408]), .B(n2868), .Z(n2869) );
  XOR U3892 ( .A(n2870), .B(n2871), .Z(n2868) );
  ANDN U3893 ( .B(n2872), .A(n659), .Z(n2870) );
  XOR U3894 ( .A(b[407]), .B(n2871), .Z(n2872) );
  XOR U3895 ( .A(n2873), .B(n2874), .Z(n2871) );
  ANDN U3896 ( .B(n2875), .A(n660), .Z(n2873) );
  XOR U3897 ( .A(b[406]), .B(n2874), .Z(n2875) );
  XOR U3898 ( .A(n2876), .B(n2877), .Z(n2874) );
  ANDN U3899 ( .B(n2878), .A(n661), .Z(n2876) );
  XOR U3900 ( .A(b[405]), .B(n2877), .Z(n2878) );
  XOR U3901 ( .A(n2879), .B(n2880), .Z(n2877) );
  ANDN U3902 ( .B(n2881), .A(n662), .Z(n2879) );
  XOR U3903 ( .A(b[404]), .B(n2880), .Z(n2881) );
  XOR U3904 ( .A(n2882), .B(n2883), .Z(n2880) );
  ANDN U3905 ( .B(n2884), .A(n663), .Z(n2882) );
  XOR U3906 ( .A(b[403]), .B(n2883), .Z(n2884) );
  XOR U3907 ( .A(n2885), .B(n2886), .Z(n2883) );
  ANDN U3908 ( .B(n2887), .A(n664), .Z(n2885) );
  XOR U3909 ( .A(b[402]), .B(n2886), .Z(n2887) );
  XOR U3910 ( .A(n2888), .B(n2889), .Z(n2886) );
  ANDN U3911 ( .B(n2890), .A(n665), .Z(n2888) );
  XOR U3912 ( .A(b[401]), .B(n2889), .Z(n2890) );
  XOR U3913 ( .A(n2891), .B(n2892), .Z(n2889) );
  ANDN U3914 ( .B(n2893), .A(n666), .Z(n2891) );
  XOR U3915 ( .A(b[400]), .B(n2892), .Z(n2893) );
  XOR U3916 ( .A(n2894), .B(n2895), .Z(n2892) );
  ANDN U3917 ( .B(n2896), .A(n669), .Z(n2894) );
  XOR U3918 ( .A(b[399]), .B(n2895), .Z(n2896) );
  XOR U3919 ( .A(n2897), .B(n2898), .Z(n2895) );
  ANDN U3920 ( .B(n2899), .A(n670), .Z(n2897) );
  XOR U3921 ( .A(b[398]), .B(n2898), .Z(n2899) );
  XOR U3922 ( .A(n2900), .B(n2901), .Z(n2898) );
  ANDN U3923 ( .B(n2902), .A(n671), .Z(n2900) );
  XOR U3924 ( .A(b[397]), .B(n2901), .Z(n2902) );
  XOR U3925 ( .A(n2903), .B(n2904), .Z(n2901) );
  ANDN U3926 ( .B(n2905), .A(n672), .Z(n2903) );
  XOR U3927 ( .A(b[396]), .B(n2904), .Z(n2905) );
  XOR U3928 ( .A(n2906), .B(n2907), .Z(n2904) );
  ANDN U3929 ( .B(n2908), .A(n673), .Z(n2906) );
  XOR U3930 ( .A(b[395]), .B(n2907), .Z(n2908) );
  XOR U3931 ( .A(n2909), .B(n2910), .Z(n2907) );
  ANDN U3932 ( .B(n2911), .A(n674), .Z(n2909) );
  XOR U3933 ( .A(b[394]), .B(n2910), .Z(n2911) );
  XOR U3934 ( .A(n2912), .B(n2913), .Z(n2910) );
  ANDN U3935 ( .B(n2914), .A(n675), .Z(n2912) );
  XOR U3936 ( .A(b[393]), .B(n2913), .Z(n2914) );
  XOR U3937 ( .A(n2915), .B(n2916), .Z(n2913) );
  ANDN U3938 ( .B(n2917), .A(n676), .Z(n2915) );
  XOR U3939 ( .A(b[392]), .B(n2916), .Z(n2917) );
  XOR U3940 ( .A(n2918), .B(n2919), .Z(n2916) );
  ANDN U3941 ( .B(n2920), .A(n677), .Z(n2918) );
  XOR U3942 ( .A(b[391]), .B(n2919), .Z(n2920) );
  XOR U3943 ( .A(n2921), .B(n2922), .Z(n2919) );
  ANDN U3944 ( .B(n2923), .A(n678), .Z(n2921) );
  XOR U3945 ( .A(b[390]), .B(n2922), .Z(n2923) );
  XOR U3946 ( .A(n2924), .B(n2925), .Z(n2922) );
  ANDN U3947 ( .B(n2926), .A(n680), .Z(n2924) );
  XOR U3948 ( .A(b[389]), .B(n2925), .Z(n2926) );
  XOR U3949 ( .A(n2927), .B(n2928), .Z(n2925) );
  ANDN U3950 ( .B(n2929), .A(n681), .Z(n2927) );
  XOR U3951 ( .A(b[388]), .B(n2928), .Z(n2929) );
  XOR U3952 ( .A(n2930), .B(n2931), .Z(n2928) );
  ANDN U3953 ( .B(n2932), .A(n682), .Z(n2930) );
  XOR U3954 ( .A(b[387]), .B(n2931), .Z(n2932) );
  XOR U3955 ( .A(n2933), .B(n2934), .Z(n2931) );
  ANDN U3956 ( .B(n2935), .A(n683), .Z(n2933) );
  XOR U3957 ( .A(b[386]), .B(n2934), .Z(n2935) );
  XOR U3958 ( .A(n2936), .B(n2937), .Z(n2934) );
  ANDN U3959 ( .B(n2938), .A(n684), .Z(n2936) );
  XOR U3960 ( .A(b[385]), .B(n2937), .Z(n2938) );
  XOR U3961 ( .A(n2939), .B(n2940), .Z(n2937) );
  ANDN U3962 ( .B(n2941), .A(n685), .Z(n2939) );
  XOR U3963 ( .A(b[384]), .B(n2940), .Z(n2941) );
  XOR U3964 ( .A(n2942), .B(n2943), .Z(n2940) );
  ANDN U3965 ( .B(n2944), .A(n686), .Z(n2942) );
  XOR U3966 ( .A(b[383]), .B(n2943), .Z(n2944) );
  XOR U3967 ( .A(n2945), .B(n2946), .Z(n2943) );
  ANDN U3968 ( .B(n2947), .A(n687), .Z(n2945) );
  XOR U3969 ( .A(b[382]), .B(n2946), .Z(n2947) );
  XOR U3970 ( .A(n2948), .B(n2949), .Z(n2946) );
  ANDN U3971 ( .B(n2950), .A(n688), .Z(n2948) );
  XOR U3972 ( .A(b[381]), .B(n2949), .Z(n2950) );
  XOR U3973 ( .A(n2951), .B(n2952), .Z(n2949) );
  ANDN U3974 ( .B(n2953), .A(n689), .Z(n2951) );
  XOR U3975 ( .A(b[380]), .B(n2952), .Z(n2953) );
  XOR U3976 ( .A(n2954), .B(n2955), .Z(n2952) );
  ANDN U3977 ( .B(n2956), .A(n691), .Z(n2954) );
  XOR U3978 ( .A(b[379]), .B(n2955), .Z(n2956) );
  XOR U3979 ( .A(n2957), .B(n2958), .Z(n2955) );
  ANDN U3980 ( .B(n2959), .A(n692), .Z(n2957) );
  XOR U3981 ( .A(b[378]), .B(n2958), .Z(n2959) );
  XOR U3982 ( .A(n2960), .B(n2961), .Z(n2958) );
  ANDN U3983 ( .B(n2962), .A(n693), .Z(n2960) );
  XOR U3984 ( .A(b[377]), .B(n2961), .Z(n2962) );
  XOR U3985 ( .A(n2963), .B(n2964), .Z(n2961) );
  ANDN U3986 ( .B(n2965), .A(n694), .Z(n2963) );
  XOR U3987 ( .A(b[376]), .B(n2964), .Z(n2965) );
  XOR U3988 ( .A(n2966), .B(n2967), .Z(n2964) );
  ANDN U3989 ( .B(n2968), .A(n695), .Z(n2966) );
  XOR U3990 ( .A(b[375]), .B(n2967), .Z(n2968) );
  XOR U3991 ( .A(n2969), .B(n2970), .Z(n2967) );
  ANDN U3992 ( .B(n2971), .A(n696), .Z(n2969) );
  XOR U3993 ( .A(b[374]), .B(n2970), .Z(n2971) );
  XOR U3994 ( .A(n2972), .B(n2973), .Z(n2970) );
  ANDN U3995 ( .B(n2974), .A(n697), .Z(n2972) );
  XOR U3996 ( .A(b[373]), .B(n2973), .Z(n2974) );
  XOR U3997 ( .A(n2975), .B(n2976), .Z(n2973) );
  ANDN U3998 ( .B(n2977), .A(n698), .Z(n2975) );
  XOR U3999 ( .A(b[372]), .B(n2976), .Z(n2977) );
  XOR U4000 ( .A(n2978), .B(n2979), .Z(n2976) );
  ANDN U4001 ( .B(n2980), .A(n699), .Z(n2978) );
  XOR U4002 ( .A(b[371]), .B(n2979), .Z(n2980) );
  XOR U4003 ( .A(n2981), .B(n2982), .Z(n2979) );
  ANDN U4004 ( .B(n2983), .A(n700), .Z(n2981) );
  XOR U4005 ( .A(b[370]), .B(n2982), .Z(n2983) );
  XOR U4006 ( .A(n2984), .B(n2985), .Z(n2982) );
  ANDN U4007 ( .B(n2986), .A(n702), .Z(n2984) );
  XOR U4008 ( .A(b[369]), .B(n2985), .Z(n2986) );
  XOR U4009 ( .A(n2987), .B(n2988), .Z(n2985) );
  ANDN U4010 ( .B(n2989), .A(n703), .Z(n2987) );
  XOR U4011 ( .A(b[368]), .B(n2988), .Z(n2989) );
  XOR U4012 ( .A(n2990), .B(n2991), .Z(n2988) );
  ANDN U4013 ( .B(n2992), .A(n704), .Z(n2990) );
  XOR U4014 ( .A(b[367]), .B(n2991), .Z(n2992) );
  XOR U4015 ( .A(n2993), .B(n2994), .Z(n2991) );
  ANDN U4016 ( .B(n2995), .A(n705), .Z(n2993) );
  XOR U4017 ( .A(b[366]), .B(n2994), .Z(n2995) );
  XOR U4018 ( .A(n2996), .B(n2997), .Z(n2994) );
  ANDN U4019 ( .B(n2998), .A(n706), .Z(n2996) );
  XOR U4020 ( .A(b[365]), .B(n2997), .Z(n2998) );
  XOR U4021 ( .A(n2999), .B(n3000), .Z(n2997) );
  ANDN U4022 ( .B(n3001), .A(n707), .Z(n2999) );
  XOR U4023 ( .A(b[364]), .B(n3000), .Z(n3001) );
  XOR U4024 ( .A(n3002), .B(n3003), .Z(n3000) );
  ANDN U4025 ( .B(n3004), .A(n708), .Z(n3002) );
  XOR U4026 ( .A(b[363]), .B(n3003), .Z(n3004) );
  XOR U4027 ( .A(n3005), .B(n3006), .Z(n3003) );
  ANDN U4028 ( .B(n3007), .A(n709), .Z(n3005) );
  XOR U4029 ( .A(b[362]), .B(n3006), .Z(n3007) );
  XOR U4030 ( .A(n3008), .B(n3009), .Z(n3006) );
  ANDN U4031 ( .B(n3010), .A(n710), .Z(n3008) );
  XOR U4032 ( .A(b[361]), .B(n3009), .Z(n3010) );
  XOR U4033 ( .A(n3011), .B(n3012), .Z(n3009) );
  ANDN U4034 ( .B(n3013), .A(n711), .Z(n3011) );
  XOR U4035 ( .A(b[360]), .B(n3012), .Z(n3013) );
  XOR U4036 ( .A(n3014), .B(n3015), .Z(n3012) );
  ANDN U4037 ( .B(n3016), .A(n713), .Z(n3014) );
  XOR U4038 ( .A(b[359]), .B(n3015), .Z(n3016) );
  XOR U4039 ( .A(n3017), .B(n3018), .Z(n3015) );
  ANDN U4040 ( .B(n3019), .A(n714), .Z(n3017) );
  XOR U4041 ( .A(b[358]), .B(n3018), .Z(n3019) );
  XOR U4042 ( .A(n3020), .B(n3021), .Z(n3018) );
  ANDN U4043 ( .B(n3022), .A(n715), .Z(n3020) );
  XOR U4044 ( .A(b[357]), .B(n3021), .Z(n3022) );
  XOR U4045 ( .A(n3023), .B(n3024), .Z(n3021) );
  ANDN U4046 ( .B(n3025), .A(n716), .Z(n3023) );
  XOR U4047 ( .A(b[356]), .B(n3024), .Z(n3025) );
  XOR U4048 ( .A(n3026), .B(n3027), .Z(n3024) );
  ANDN U4049 ( .B(n3028), .A(n717), .Z(n3026) );
  XOR U4050 ( .A(b[355]), .B(n3027), .Z(n3028) );
  XOR U4051 ( .A(n3029), .B(n3030), .Z(n3027) );
  ANDN U4052 ( .B(n3031), .A(n718), .Z(n3029) );
  XOR U4053 ( .A(b[354]), .B(n3030), .Z(n3031) );
  XOR U4054 ( .A(n3032), .B(n3033), .Z(n3030) );
  ANDN U4055 ( .B(n3034), .A(n719), .Z(n3032) );
  XOR U4056 ( .A(b[353]), .B(n3033), .Z(n3034) );
  XOR U4057 ( .A(n3035), .B(n3036), .Z(n3033) );
  ANDN U4058 ( .B(n3037), .A(n720), .Z(n3035) );
  XOR U4059 ( .A(b[352]), .B(n3036), .Z(n3037) );
  XOR U4060 ( .A(n3038), .B(n3039), .Z(n3036) );
  ANDN U4061 ( .B(n3040), .A(n721), .Z(n3038) );
  XOR U4062 ( .A(b[351]), .B(n3039), .Z(n3040) );
  XOR U4063 ( .A(n3041), .B(n3042), .Z(n3039) );
  ANDN U4064 ( .B(n3043), .A(n722), .Z(n3041) );
  XOR U4065 ( .A(b[350]), .B(n3042), .Z(n3043) );
  XOR U4066 ( .A(n3044), .B(n3045), .Z(n3042) );
  ANDN U4067 ( .B(n3046), .A(n724), .Z(n3044) );
  XOR U4068 ( .A(b[349]), .B(n3045), .Z(n3046) );
  XOR U4069 ( .A(n3047), .B(n3048), .Z(n3045) );
  ANDN U4070 ( .B(n3049), .A(n725), .Z(n3047) );
  XOR U4071 ( .A(b[348]), .B(n3048), .Z(n3049) );
  XOR U4072 ( .A(n3050), .B(n3051), .Z(n3048) );
  ANDN U4073 ( .B(n3052), .A(n726), .Z(n3050) );
  XOR U4074 ( .A(b[347]), .B(n3051), .Z(n3052) );
  XOR U4075 ( .A(n3053), .B(n3054), .Z(n3051) );
  ANDN U4076 ( .B(n3055), .A(n727), .Z(n3053) );
  XOR U4077 ( .A(b[346]), .B(n3054), .Z(n3055) );
  XOR U4078 ( .A(n3056), .B(n3057), .Z(n3054) );
  ANDN U4079 ( .B(n3058), .A(n728), .Z(n3056) );
  XOR U4080 ( .A(b[345]), .B(n3057), .Z(n3058) );
  XOR U4081 ( .A(n3059), .B(n3060), .Z(n3057) );
  ANDN U4082 ( .B(n3061), .A(n729), .Z(n3059) );
  XOR U4083 ( .A(b[344]), .B(n3060), .Z(n3061) );
  XOR U4084 ( .A(n3062), .B(n3063), .Z(n3060) );
  ANDN U4085 ( .B(n3064), .A(n730), .Z(n3062) );
  XOR U4086 ( .A(b[343]), .B(n3063), .Z(n3064) );
  XOR U4087 ( .A(n3065), .B(n3066), .Z(n3063) );
  ANDN U4088 ( .B(n3067), .A(n731), .Z(n3065) );
  XOR U4089 ( .A(b[342]), .B(n3066), .Z(n3067) );
  XOR U4090 ( .A(n3068), .B(n3069), .Z(n3066) );
  ANDN U4091 ( .B(n3070), .A(n732), .Z(n3068) );
  XOR U4092 ( .A(b[341]), .B(n3069), .Z(n3070) );
  XOR U4093 ( .A(n3071), .B(n3072), .Z(n3069) );
  ANDN U4094 ( .B(n3073), .A(n733), .Z(n3071) );
  XOR U4095 ( .A(b[340]), .B(n3072), .Z(n3073) );
  XOR U4096 ( .A(n3074), .B(n3075), .Z(n3072) );
  ANDN U4097 ( .B(n3076), .A(n735), .Z(n3074) );
  XOR U4098 ( .A(b[339]), .B(n3075), .Z(n3076) );
  XOR U4099 ( .A(n3077), .B(n3078), .Z(n3075) );
  ANDN U4100 ( .B(n3079), .A(n736), .Z(n3077) );
  XOR U4101 ( .A(b[338]), .B(n3078), .Z(n3079) );
  XOR U4102 ( .A(n3080), .B(n3081), .Z(n3078) );
  ANDN U4103 ( .B(n3082), .A(n737), .Z(n3080) );
  XOR U4104 ( .A(b[337]), .B(n3081), .Z(n3082) );
  XOR U4105 ( .A(n3083), .B(n3084), .Z(n3081) );
  ANDN U4106 ( .B(n3085), .A(n738), .Z(n3083) );
  XOR U4107 ( .A(b[336]), .B(n3084), .Z(n3085) );
  XOR U4108 ( .A(n3086), .B(n3087), .Z(n3084) );
  ANDN U4109 ( .B(n3088), .A(n739), .Z(n3086) );
  XOR U4110 ( .A(b[335]), .B(n3087), .Z(n3088) );
  XOR U4111 ( .A(n3089), .B(n3090), .Z(n3087) );
  ANDN U4112 ( .B(n3091), .A(n740), .Z(n3089) );
  XOR U4113 ( .A(b[334]), .B(n3090), .Z(n3091) );
  XOR U4114 ( .A(n3092), .B(n3093), .Z(n3090) );
  ANDN U4115 ( .B(n3094), .A(n741), .Z(n3092) );
  XOR U4116 ( .A(b[333]), .B(n3093), .Z(n3094) );
  XOR U4117 ( .A(n3095), .B(n3096), .Z(n3093) );
  ANDN U4118 ( .B(n3097), .A(n742), .Z(n3095) );
  XOR U4119 ( .A(b[332]), .B(n3096), .Z(n3097) );
  XOR U4120 ( .A(n3098), .B(n3099), .Z(n3096) );
  ANDN U4121 ( .B(n3100), .A(n743), .Z(n3098) );
  XOR U4122 ( .A(b[331]), .B(n3099), .Z(n3100) );
  XOR U4123 ( .A(n3101), .B(n3102), .Z(n3099) );
  ANDN U4124 ( .B(n3103), .A(n744), .Z(n3101) );
  XOR U4125 ( .A(b[330]), .B(n3102), .Z(n3103) );
  XOR U4126 ( .A(n3104), .B(n3105), .Z(n3102) );
  ANDN U4127 ( .B(n3106), .A(n746), .Z(n3104) );
  XOR U4128 ( .A(b[329]), .B(n3105), .Z(n3106) );
  XOR U4129 ( .A(n3107), .B(n3108), .Z(n3105) );
  ANDN U4130 ( .B(n3109), .A(n747), .Z(n3107) );
  XOR U4131 ( .A(b[328]), .B(n3108), .Z(n3109) );
  XOR U4132 ( .A(n3110), .B(n3111), .Z(n3108) );
  ANDN U4133 ( .B(n3112), .A(n748), .Z(n3110) );
  XOR U4134 ( .A(b[327]), .B(n3111), .Z(n3112) );
  XOR U4135 ( .A(n3113), .B(n3114), .Z(n3111) );
  ANDN U4136 ( .B(n3115), .A(n749), .Z(n3113) );
  XOR U4137 ( .A(b[326]), .B(n3114), .Z(n3115) );
  XOR U4138 ( .A(n3116), .B(n3117), .Z(n3114) );
  ANDN U4139 ( .B(n3118), .A(n750), .Z(n3116) );
  XOR U4140 ( .A(b[325]), .B(n3117), .Z(n3118) );
  XOR U4141 ( .A(n3119), .B(n3120), .Z(n3117) );
  ANDN U4142 ( .B(n3121), .A(n751), .Z(n3119) );
  XOR U4143 ( .A(b[324]), .B(n3120), .Z(n3121) );
  XOR U4144 ( .A(n3122), .B(n3123), .Z(n3120) );
  ANDN U4145 ( .B(n3124), .A(n752), .Z(n3122) );
  XOR U4146 ( .A(b[323]), .B(n3123), .Z(n3124) );
  XOR U4147 ( .A(n3125), .B(n3126), .Z(n3123) );
  ANDN U4148 ( .B(n3127), .A(n753), .Z(n3125) );
  XOR U4149 ( .A(b[322]), .B(n3126), .Z(n3127) );
  XOR U4150 ( .A(n3128), .B(n3129), .Z(n3126) );
  ANDN U4151 ( .B(n3130), .A(n754), .Z(n3128) );
  XOR U4152 ( .A(b[321]), .B(n3129), .Z(n3130) );
  XOR U4153 ( .A(n3131), .B(n3132), .Z(n3129) );
  ANDN U4154 ( .B(n3133), .A(n755), .Z(n3131) );
  XOR U4155 ( .A(b[320]), .B(n3132), .Z(n3133) );
  XOR U4156 ( .A(n3134), .B(n3135), .Z(n3132) );
  ANDN U4157 ( .B(n3136), .A(n757), .Z(n3134) );
  XOR U4158 ( .A(b[319]), .B(n3135), .Z(n3136) );
  XOR U4159 ( .A(n3137), .B(n3138), .Z(n3135) );
  ANDN U4160 ( .B(n3139), .A(n758), .Z(n3137) );
  XOR U4161 ( .A(b[318]), .B(n3138), .Z(n3139) );
  XOR U4162 ( .A(n3140), .B(n3141), .Z(n3138) );
  ANDN U4163 ( .B(n3142), .A(n759), .Z(n3140) );
  XOR U4164 ( .A(b[317]), .B(n3141), .Z(n3142) );
  XOR U4165 ( .A(n3143), .B(n3144), .Z(n3141) );
  ANDN U4166 ( .B(n3145), .A(n760), .Z(n3143) );
  XOR U4167 ( .A(b[316]), .B(n3144), .Z(n3145) );
  XOR U4168 ( .A(n3146), .B(n3147), .Z(n3144) );
  ANDN U4169 ( .B(n3148), .A(n761), .Z(n3146) );
  XOR U4170 ( .A(b[315]), .B(n3147), .Z(n3148) );
  XOR U4171 ( .A(n3149), .B(n3150), .Z(n3147) );
  ANDN U4172 ( .B(n3151), .A(n762), .Z(n3149) );
  XOR U4173 ( .A(b[314]), .B(n3150), .Z(n3151) );
  XOR U4174 ( .A(n3152), .B(n3153), .Z(n3150) );
  ANDN U4175 ( .B(n3154), .A(n763), .Z(n3152) );
  XOR U4176 ( .A(b[313]), .B(n3153), .Z(n3154) );
  XOR U4177 ( .A(n3155), .B(n3156), .Z(n3153) );
  ANDN U4178 ( .B(n3157), .A(n764), .Z(n3155) );
  XOR U4179 ( .A(b[312]), .B(n3156), .Z(n3157) );
  XOR U4180 ( .A(n3158), .B(n3159), .Z(n3156) );
  ANDN U4181 ( .B(n3160), .A(n765), .Z(n3158) );
  XOR U4182 ( .A(b[311]), .B(n3159), .Z(n3160) );
  XOR U4183 ( .A(n3161), .B(n3162), .Z(n3159) );
  ANDN U4184 ( .B(n3163), .A(n766), .Z(n3161) );
  XOR U4185 ( .A(b[310]), .B(n3162), .Z(n3163) );
  XOR U4186 ( .A(n3164), .B(n3165), .Z(n3162) );
  ANDN U4187 ( .B(n3166), .A(n768), .Z(n3164) );
  XOR U4188 ( .A(b[309]), .B(n3165), .Z(n3166) );
  XOR U4189 ( .A(n3167), .B(n3168), .Z(n3165) );
  ANDN U4190 ( .B(n3169), .A(n769), .Z(n3167) );
  XOR U4191 ( .A(b[308]), .B(n3168), .Z(n3169) );
  XOR U4192 ( .A(n3170), .B(n3171), .Z(n3168) );
  ANDN U4193 ( .B(n3172), .A(n770), .Z(n3170) );
  XOR U4194 ( .A(b[307]), .B(n3171), .Z(n3172) );
  XOR U4195 ( .A(n3173), .B(n3174), .Z(n3171) );
  ANDN U4196 ( .B(n3175), .A(n771), .Z(n3173) );
  XOR U4197 ( .A(b[306]), .B(n3174), .Z(n3175) );
  XOR U4198 ( .A(n3176), .B(n3177), .Z(n3174) );
  ANDN U4199 ( .B(n3178), .A(n772), .Z(n3176) );
  XOR U4200 ( .A(b[305]), .B(n3177), .Z(n3178) );
  XOR U4201 ( .A(n3179), .B(n3180), .Z(n3177) );
  ANDN U4202 ( .B(n3181), .A(n773), .Z(n3179) );
  XOR U4203 ( .A(b[304]), .B(n3180), .Z(n3181) );
  XOR U4204 ( .A(n3182), .B(n3183), .Z(n3180) );
  ANDN U4205 ( .B(n3184), .A(n774), .Z(n3182) );
  XOR U4206 ( .A(b[303]), .B(n3183), .Z(n3184) );
  XOR U4207 ( .A(n3185), .B(n3186), .Z(n3183) );
  ANDN U4208 ( .B(n3187), .A(n775), .Z(n3185) );
  XOR U4209 ( .A(b[302]), .B(n3186), .Z(n3187) );
  XOR U4210 ( .A(n3188), .B(n3189), .Z(n3186) );
  ANDN U4211 ( .B(n3190), .A(n776), .Z(n3188) );
  XOR U4212 ( .A(b[301]), .B(n3189), .Z(n3190) );
  XOR U4213 ( .A(n3191), .B(n3192), .Z(n3189) );
  ANDN U4214 ( .B(n3193), .A(n777), .Z(n3191) );
  XOR U4215 ( .A(b[300]), .B(n3192), .Z(n3193) );
  XOR U4216 ( .A(n3194), .B(n3195), .Z(n3192) );
  ANDN U4217 ( .B(n3196), .A(n780), .Z(n3194) );
  XOR U4218 ( .A(b[299]), .B(n3195), .Z(n3196) );
  XOR U4219 ( .A(n3197), .B(n3198), .Z(n3195) );
  ANDN U4220 ( .B(n3199), .A(n781), .Z(n3197) );
  XOR U4221 ( .A(b[298]), .B(n3198), .Z(n3199) );
  XOR U4222 ( .A(n3200), .B(n3201), .Z(n3198) );
  ANDN U4223 ( .B(n3202), .A(n782), .Z(n3200) );
  XOR U4224 ( .A(b[297]), .B(n3201), .Z(n3202) );
  XOR U4225 ( .A(n3203), .B(n3204), .Z(n3201) );
  ANDN U4226 ( .B(n3205), .A(n783), .Z(n3203) );
  XOR U4227 ( .A(b[296]), .B(n3204), .Z(n3205) );
  XOR U4228 ( .A(n3206), .B(n3207), .Z(n3204) );
  ANDN U4229 ( .B(n3208), .A(n784), .Z(n3206) );
  XOR U4230 ( .A(b[295]), .B(n3207), .Z(n3208) );
  XOR U4231 ( .A(n3209), .B(n3210), .Z(n3207) );
  ANDN U4232 ( .B(n3211), .A(n785), .Z(n3209) );
  XOR U4233 ( .A(b[294]), .B(n3210), .Z(n3211) );
  XOR U4234 ( .A(n3212), .B(n3213), .Z(n3210) );
  ANDN U4235 ( .B(n3214), .A(n786), .Z(n3212) );
  XOR U4236 ( .A(b[293]), .B(n3213), .Z(n3214) );
  XOR U4237 ( .A(n3215), .B(n3216), .Z(n3213) );
  ANDN U4238 ( .B(n3217), .A(n787), .Z(n3215) );
  XOR U4239 ( .A(b[292]), .B(n3216), .Z(n3217) );
  XOR U4240 ( .A(n3218), .B(n3219), .Z(n3216) );
  ANDN U4241 ( .B(n3220), .A(n788), .Z(n3218) );
  XOR U4242 ( .A(b[291]), .B(n3219), .Z(n3220) );
  XOR U4243 ( .A(n3221), .B(n3222), .Z(n3219) );
  ANDN U4244 ( .B(n3223), .A(n789), .Z(n3221) );
  XOR U4245 ( .A(b[290]), .B(n3222), .Z(n3223) );
  XOR U4246 ( .A(n3224), .B(n3225), .Z(n3222) );
  ANDN U4247 ( .B(n3226), .A(n791), .Z(n3224) );
  XOR U4248 ( .A(b[289]), .B(n3225), .Z(n3226) );
  XOR U4249 ( .A(n3227), .B(n3228), .Z(n3225) );
  ANDN U4250 ( .B(n3229), .A(n792), .Z(n3227) );
  XOR U4251 ( .A(b[288]), .B(n3228), .Z(n3229) );
  XOR U4252 ( .A(n3230), .B(n3231), .Z(n3228) );
  ANDN U4253 ( .B(n3232), .A(n793), .Z(n3230) );
  XOR U4254 ( .A(b[287]), .B(n3231), .Z(n3232) );
  XOR U4255 ( .A(n3233), .B(n3234), .Z(n3231) );
  ANDN U4256 ( .B(n3235), .A(n794), .Z(n3233) );
  XOR U4257 ( .A(b[286]), .B(n3234), .Z(n3235) );
  XOR U4258 ( .A(n3236), .B(n3237), .Z(n3234) );
  ANDN U4259 ( .B(n3238), .A(n795), .Z(n3236) );
  XOR U4260 ( .A(b[285]), .B(n3237), .Z(n3238) );
  XOR U4261 ( .A(n3239), .B(n3240), .Z(n3237) );
  ANDN U4262 ( .B(n3241), .A(n796), .Z(n3239) );
  XOR U4263 ( .A(b[284]), .B(n3240), .Z(n3241) );
  XOR U4264 ( .A(n3242), .B(n3243), .Z(n3240) );
  ANDN U4265 ( .B(n3244), .A(n797), .Z(n3242) );
  XOR U4266 ( .A(b[283]), .B(n3243), .Z(n3244) );
  XOR U4267 ( .A(n3245), .B(n3246), .Z(n3243) );
  ANDN U4268 ( .B(n3247), .A(n798), .Z(n3245) );
  XOR U4269 ( .A(b[282]), .B(n3246), .Z(n3247) );
  XOR U4270 ( .A(n3248), .B(n3249), .Z(n3246) );
  ANDN U4271 ( .B(n3250), .A(n799), .Z(n3248) );
  XOR U4272 ( .A(b[281]), .B(n3249), .Z(n3250) );
  XOR U4273 ( .A(n3251), .B(n3252), .Z(n3249) );
  ANDN U4274 ( .B(n3253), .A(n800), .Z(n3251) );
  XOR U4275 ( .A(b[280]), .B(n3252), .Z(n3253) );
  XOR U4276 ( .A(n3254), .B(n3255), .Z(n3252) );
  ANDN U4277 ( .B(n3256), .A(n802), .Z(n3254) );
  XOR U4278 ( .A(b[279]), .B(n3255), .Z(n3256) );
  XOR U4279 ( .A(n3257), .B(n3258), .Z(n3255) );
  ANDN U4280 ( .B(n3259), .A(n803), .Z(n3257) );
  XOR U4281 ( .A(b[278]), .B(n3258), .Z(n3259) );
  XOR U4282 ( .A(n3260), .B(n3261), .Z(n3258) );
  ANDN U4283 ( .B(n3262), .A(n804), .Z(n3260) );
  XOR U4284 ( .A(b[277]), .B(n3261), .Z(n3262) );
  XOR U4285 ( .A(n3263), .B(n3264), .Z(n3261) );
  ANDN U4286 ( .B(n3265), .A(n805), .Z(n3263) );
  XOR U4287 ( .A(b[276]), .B(n3264), .Z(n3265) );
  XOR U4288 ( .A(n3266), .B(n3267), .Z(n3264) );
  ANDN U4289 ( .B(n3268), .A(n806), .Z(n3266) );
  XOR U4290 ( .A(b[275]), .B(n3267), .Z(n3268) );
  XOR U4291 ( .A(n3269), .B(n3270), .Z(n3267) );
  ANDN U4292 ( .B(n3271), .A(n807), .Z(n3269) );
  XOR U4293 ( .A(b[274]), .B(n3270), .Z(n3271) );
  XOR U4294 ( .A(n3272), .B(n3273), .Z(n3270) );
  ANDN U4295 ( .B(n3274), .A(n808), .Z(n3272) );
  XOR U4296 ( .A(b[273]), .B(n3273), .Z(n3274) );
  XOR U4297 ( .A(n3275), .B(n3276), .Z(n3273) );
  ANDN U4298 ( .B(n3277), .A(n809), .Z(n3275) );
  XOR U4299 ( .A(b[272]), .B(n3276), .Z(n3277) );
  XOR U4300 ( .A(n3278), .B(n3279), .Z(n3276) );
  ANDN U4301 ( .B(n3280), .A(n810), .Z(n3278) );
  XOR U4302 ( .A(b[271]), .B(n3279), .Z(n3280) );
  XOR U4303 ( .A(n3281), .B(n3282), .Z(n3279) );
  ANDN U4304 ( .B(n3283), .A(n811), .Z(n3281) );
  XOR U4305 ( .A(b[270]), .B(n3282), .Z(n3283) );
  XOR U4306 ( .A(n3284), .B(n3285), .Z(n3282) );
  ANDN U4307 ( .B(n3286), .A(n813), .Z(n3284) );
  XOR U4308 ( .A(b[269]), .B(n3285), .Z(n3286) );
  XOR U4309 ( .A(n3287), .B(n3288), .Z(n3285) );
  ANDN U4310 ( .B(n3289), .A(n814), .Z(n3287) );
  XOR U4311 ( .A(b[268]), .B(n3288), .Z(n3289) );
  XOR U4312 ( .A(n3290), .B(n3291), .Z(n3288) );
  ANDN U4313 ( .B(n3292), .A(n815), .Z(n3290) );
  XOR U4314 ( .A(b[267]), .B(n3291), .Z(n3292) );
  XOR U4315 ( .A(n3293), .B(n3294), .Z(n3291) );
  ANDN U4316 ( .B(n3295), .A(n816), .Z(n3293) );
  XOR U4317 ( .A(b[266]), .B(n3294), .Z(n3295) );
  XOR U4318 ( .A(n3296), .B(n3297), .Z(n3294) );
  ANDN U4319 ( .B(n3298), .A(n817), .Z(n3296) );
  XOR U4320 ( .A(b[265]), .B(n3297), .Z(n3298) );
  XOR U4321 ( .A(n3299), .B(n3300), .Z(n3297) );
  ANDN U4322 ( .B(n3301), .A(n818), .Z(n3299) );
  XOR U4323 ( .A(b[264]), .B(n3300), .Z(n3301) );
  XOR U4324 ( .A(n3302), .B(n3303), .Z(n3300) );
  ANDN U4325 ( .B(n3304), .A(n819), .Z(n3302) );
  XOR U4326 ( .A(b[263]), .B(n3303), .Z(n3304) );
  XOR U4327 ( .A(n3305), .B(n3306), .Z(n3303) );
  ANDN U4328 ( .B(n3307), .A(n820), .Z(n3305) );
  XOR U4329 ( .A(b[262]), .B(n3306), .Z(n3307) );
  XOR U4330 ( .A(n3308), .B(n3309), .Z(n3306) );
  ANDN U4331 ( .B(n3310), .A(n821), .Z(n3308) );
  XOR U4332 ( .A(b[261]), .B(n3309), .Z(n3310) );
  XOR U4333 ( .A(n3311), .B(n3312), .Z(n3309) );
  ANDN U4334 ( .B(n3313), .A(n822), .Z(n3311) );
  XOR U4335 ( .A(b[260]), .B(n3312), .Z(n3313) );
  XOR U4336 ( .A(n3314), .B(n3315), .Z(n3312) );
  ANDN U4337 ( .B(n3316), .A(n824), .Z(n3314) );
  XOR U4338 ( .A(b[259]), .B(n3315), .Z(n3316) );
  XOR U4339 ( .A(n3317), .B(n3318), .Z(n3315) );
  ANDN U4340 ( .B(n3319), .A(n825), .Z(n3317) );
  XOR U4341 ( .A(b[258]), .B(n3318), .Z(n3319) );
  XOR U4342 ( .A(n3320), .B(n3321), .Z(n3318) );
  ANDN U4343 ( .B(n3322), .A(n826), .Z(n3320) );
  XOR U4344 ( .A(b[257]), .B(n3321), .Z(n3322) );
  XOR U4345 ( .A(n3323), .B(n3324), .Z(n3321) );
  ANDN U4346 ( .B(n3325), .A(n827), .Z(n3323) );
  XOR U4347 ( .A(b[256]), .B(n3324), .Z(n3325) );
  XOR U4348 ( .A(n3326), .B(n3327), .Z(n3324) );
  ANDN U4349 ( .B(n3328), .A(n828), .Z(n3326) );
  XOR U4350 ( .A(b[255]), .B(n3327), .Z(n3328) );
  XOR U4351 ( .A(n3329), .B(n3330), .Z(n3327) );
  ANDN U4352 ( .B(n3331), .A(n829), .Z(n3329) );
  XOR U4353 ( .A(b[254]), .B(n3330), .Z(n3331) );
  XOR U4354 ( .A(n3332), .B(n3333), .Z(n3330) );
  ANDN U4355 ( .B(n3334), .A(n830), .Z(n3332) );
  XOR U4356 ( .A(b[253]), .B(n3333), .Z(n3334) );
  XOR U4357 ( .A(n3335), .B(n3336), .Z(n3333) );
  ANDN U4358 ( .B(n3337), .A(n831), .Z(n3335) );
  XOR U4359 ( .A(b[252]), .B(n3336), .Z(n3337) );
  XOR U4360 ( .A(n3338), .B(n3339), .Z(n3336) );
  ANDN U4361 ( .B(n3340), .A(n832), .Z(n3338) );
  XOR U4362 ( .A(b[251]), .B(n3339), .Z(n3340) );
  XOR U4363 ( .A(n3341), .B(n3342), .Z(n3339) );
  ANDN U4364 ( .B(n3343), .A(n833), .Z(n3341) );
  XOR U4365 ( .A(b[250]), .B(n3342), .Z(n3343) );
  XOR U4366 ( .A(n3344), .B(n3345), .Z(n3342) );
  ANDN U4367 ( .B(n3346), .A(n835), .Z(n3344) );
  XOR U4368 ( .A(b[249]), .B(n3345), .Z(n3346) );
  XOR U4369 ( .A(n3347), .B(n3348), .Z(n3345) );
  ANDN U4370 ( .B(n3349), .A(n836), .Z(n3347) );
  XOR U4371 ( .A(b[248]), .B(n3348), .Z(n3349) );
  XOR U4372 ( .A(n3350), .B(n3351), .Z(n3348) );
  ANDN U4373 ( .B(n3352), .A(n837), .Z(n3350) );
  XOR U4374 ( .A(b[247]), .B(n3351), .Z(n3352) );
  XOR U4375 ( .A(n3353), .B(n3354), .Z(n3351) );
  ANDN U4376 ( .B(n3355), .A(n838), .Z(n3353) );
  XOR U4377 ( .A(b[246]), .B(n3354), .Z(n3355) );
  XOR U4378 ( .A(n3356), .B(n3357), .Z(n3354) );
  ANDN U4379 ( .B(n3358), .A(n839), .Z(n3356) );
  XOR U4380 ( .A(b[245]), .B(n3357), .Z(n3358) );
  XOR U4381 ( .A(n3359), .B(n3360), .Z(n3357) );
  ANDN U4382 ( .B(n3361), .A(n840), .Z(n3359) );
  XOR U4383 ( .A(b[244]), .B(n3360), .Z(n3361) );
  XOR U4384 ( .A(n3362), .B(n3363), .Z(n3360) );
  ANDN U4385 ( .B(n3364), .A(n841), .Z(n3362) );
  XOR U4386 ( .A(b[243]), .B(n3363), .Z(n3364) );
  XOR U4387 ( .A(n3365), .B(n3366), .Z(n3363) );
  ANDN U4388 ( .B(n3367), .A(n842), .Z(n3365) );
  XOR U4389 ( .A(b[242]), .B(n3366), .Z(n3367) );
  XOR U4390 ( .A(n3368), .B(n3369), .Z(n3366) );
  ANDN U4391 ( .B(n3370), .A(n843), .Z(n3368) );
  XOR U4392 ( .A(b[241]), .B(n3369), .Z(n3370) );
  XOR U4393 ( .A(n3371), .B(n3372), .Z(n3369) );
  ANDN U4394 ( .B(n3373), .A(n844), .Z(n3371) );
  XOR U4395 ( .A(b[240]), .B(n3372), .Z(n3373) );
  XOR U4396 ( .A(n3374), .B(n3375), .Z(n3372) );
  ANDN U4397 ( .B(n3376), .A(n846), .Z(n3374) );
  XOR U4398 ( .A(b[239]), .B(n3375), .Z(n3376) );
  XOR U4399 ( .A(n3377), .B(n3378), .Z(n3375) );
  ANDN U4400 ( .B(n3379), .A(n847), .Z(n3377) );
  XOR U4401 ( .A(b[238]), .B(n3378), .Z(n3379) );
  XOR U4402 ( .A(n3380), .B(n3381), .Z(n3378) );
  ANDN U4403 ( .B(n3382), .A(n848), .Z(n3380) );
  XOR U4404 ( .A(b[237]), .B(n3381), .Z(n3382) );
  XOR U4405 ( .A(n3383), .B(n3384), .Z(n3381) );
  ANDN U4406 ( .B(n3385), .A(n849), .Z(n3383) );
  XOR U4407 ( .A(b[236]), .B(n3384), .Z(n3385) );
  XOR U4408 ( .A(n3386), .B(n3387), .Z(n3384) );
  ANDN U4409 ( .B(n3388), .A(n850), .Z(n3386) );
  XOR U4410 ( .A(b[235]), .B(n3387), .Z(n3388) );
  XOR U4411 ( .A(n3389), .B(n3390), .Z(n3387) );
  ANDN U4412 ( .B(n3391), .A(n851), .Z(n3389) );
  XOR U4413 ( .A(b[234]), .B(n3390), .Z(n3391) );
  XOR U4414 ( .A(n3392), .B(n3393), .Z(n3390) );
  ANDN U4415 ( .B(n3394), .A(n852), .Z(n3392) );
  XOR U4416 ( .A(b[233]), .B(n3393), .Z(n3394) );
  XOR U4417 ( .A(n3395), .B(n3396), .Z(n3393) );
  ANDN U4418 ( .B(n3397), .A(n853), .Z(n3395) );
  XOR U4419 ( .A(b[232]), .B(n3396), .Z(n3397) );
  XOR U4420 ( .A(n3398), .B(n3399), .Z(n3396) );
  ANDN U4421 ( .B(n3400), .A(n854), .Z(n3398) );
  XOR U4422 ( .A(b[231]), .B(n3399), .Z(n3400) );
  XOR U4423 ( .A(n3401), .B(n3402), .Z(n3399) );
  ANDN U4424 ( .B(n3403), .A(n855), .Z(n3401) );
  XOR U4425 ( .A(b[230]), .B(n3402), .Z(n3403) );
  XOR U4426 ( .A(n3404), .B(n3405), .Z(n3402) );
  ANDN U4427 ( .B(n3406), .A(n857), .Z(n3404) );
  XOR U4428 ( .A(b[229]), .B(n3405), .Z(n3406) );
  XOR U4429 ( .A(n3407), .B(n3408), .Z(n3405) );
  ANDN U4430 ( .B(n3409), .A(n858), .Z(n3407) );
  XOR U4431 ( .A(b[228]), .B(n3408), .Z(n3409) );
  XOR U4432 ( .A(n3410), .B(n3411), .Z(n3408) );
  ANDN U4433 ( .B(n3412), .A(n859), .Z(n3410) );
  XOR U4434 ( .A(b[227]), .B(n3411), .Z(n3412) );
  XOR U4435 ( .A(n3413), .B(n3414), .Z(n3411) );
  ANDN U4436 ( .B(n3415), .A(n860), .Z(n3413) );
  XOR U4437 ( .A(b[226]), .B(n3414), .Z(n3415) );
  XOR U4438 ( .A(n3416), .B(n3417), .Z(n3414) );
  ANDN U4439 ( .B(n3418), .A(n861), .Z(n3416) );
  XOR U4440 ( .A(b[225]), .B(n3417), .Z(n3418) );
  XOR U4441 ( .A(n3419), .B(n3420), .Z(n3417) );
  ANDN U4442 ( .B(n3421), .A(n862), .Z(n3419) );
  XOR U4443 ( .A(b[224]), .B(n3420), .Z(n3421) );
  XOR U4444 ( .A(n3422), .B(n3423), .Z(n3420) );
  ANDN U4445 ( .B(n3424), .A(n863), .Z(n3422) );
  XOR U4446 ( .A(b[223]), .B(n3423), .Z(n3424) );
  XOR U4447 ( .A(n3425), .B(n3426), .Z(n3423) );
  ANDN U4448 ( .B(n3427), .A(n864), .Z(n3425) );
  XOR U4449 ( .A(b[222]), .B(n3426), .Z(n3427) );
  XOR U4450 ( .A(n3428), .B(n3429), .Z(n3426) );
  ANDN U4451 ( .B(n3430), .A(n865), .Z(n3428) );
  XOR U4452 ( .A(b[221]), .B(n3429), .Z(n3430) );
  XOR U4453 ( .A(n3431), .B(n3432), .Z(n3429) );
  ANDN U4454 ( .B(n3433), .A(n866), .Z(n3431) );
  XOR U4455 ( .A(b[220]), .B(n3432), .Z(n3433) );
  XOR U4456 ( .A(n3434), .B(n3435), .Z(n3432) );
  ANDN U4457 ( .B(n3436), .A(n868), .Z(n3434) );
  XOR U4458 ( .A(b[219]), .B(n3435), .Z(n3436) );
  XOR U4459 ( .A(n3437), .B(n3438), .Z(n3435) );
  ANDN U4460 ( .B(n3439), .A(n869), .Z(n3437) );
  XOR U4461 ( .A(b[218]), .B(n3438), .Z(n3439) );
  XOR U4462 ( .A(n3440), .B(n3441), .Z(n3438) );
  ANDN U4463 ( .B(n3442), .A(n870), .Z(n3440) );
  XOR U4464 ( .A(b[217]), .B(n3441), .Z(n3442) );
  XOR U4465 ( .A(n3443), .B(n3444), .Z(n3441) );
  ANDN U4466 ( .B(n3445), .A(n871), .Z(n3443) );
  XOR U4467 ( .A(b[216]), .B(n3444), .Z(n3445) );
  XOR U4468 ( .A(n3446), .B(n3447), .Z(n3444) );
  ANDN U4469 ( .B(n3448), .A(n872), .Z(n3446) );
  XOR U4470 ( .A(b[215]), .B(n3447), .Z(n3448) );
  XOR U4471 ( .A(n3449), .B(n3450), .Z(n3447) );
  ANDN U4472 ( .B(n3451), .A(n873), .Z(n3449) );
  XOR U4473 ( .A(b[214]), .B(n3450), .Z(n3451) );
  XOR U4474 ( .A(n3452), .B(n3453), .Z(n3450) );
  ANDN U4475 ( .B(n3454), .A(n874), .Z(n3452) );
  XOR U4476 ( .A(b[213]), .B(n3453), .Z(n3454) );
  XOR U4477 ( .A(n3455), .B(n3456), .Z(n3453) );
  ANDN U4478 ( .B(n3457), .A(n875), .Z(n3455) );
  XOR U4479 ( .A(b[212]), .B(n3456), .Z(n3457) );
  XOR U4480 ( .A(n3458), .B(n3459), .Z(n3456) );
  ANDN U4481 ( .B(n3460), .A(n876), .Z(n3458) );
  XOR U4482 ( .A(b[211]), .B(n3459), .Z(n3460) );
  XOR U4483 ( .A(n3461), .B(n3462), .Z(n3459) );
  ANDN U4484 ( .B(n3463), .A(n877), .Z(n3461) );
  XOR U4485 ( .A(b[210]), .B(n3462), .Z(n3463) );
  XOR U4486 ( .A(n3464), .B(n3465), .Z(n3462) );
  ANDN U4487 ( .B(n3466), .A(n879), .Z(n3464) );
  XOR U4488 ( .A(b[209]), .B(n3465), .Z(n3466) );
  XOR U4489 ( .A(n3467), .B(n3468), .Z(n3465) );
  ANDN U4490 ( .B(n3469), .A(n880), .Z(n3467) );
  XOR U4491 ( .A(b[208]), .B(n3468), .Z(n3469) );
  XOR U4492 ( .A(n3470), .B(n3471), .Z(n3468) );
  ANDN U4493 ( .B(n3472), .A(n881), .Z(n3470) );
  XOR U4494 ( .A(b[207]), .B(n3471), .Z(n3472) );
  XOR U4495 ( .A(n3473), .B(n3474), .Z(n3471) );
  ANDN U4496 ( .B(n3475), .A(n882), .Z(n3473) );
  XOR U4497 ( .A(b[206]), .B(n3474), .Z(n3475) );
  XOR U4498 ( .A(n3476), .B(n3477), .Z(n3474) );
  ANDN U4499 ( .B(n3478), .A(n883), .Z(n3476) );
  XOR U4500 ( .A(b[205]), .B(n3477), .Z(n3478) );
  XOR U4501 ( .A(n3479), .B(n3480), .Z(n3477) );
  ANDN U4502 ( .B(n3481), .A(n884), .Z(n3479) );
  XOR U4503 ( .A(b[204]), .B(n3480), .Z(n3481) );
  XOR U4504 ( .A(n3482), .B(n3483), .Z(n3480) );
  ANDN U4505 ( .B(n3484), .A(n885), .Z(n3482) );
  XOR U4506 ( .A(b[203]), .B(n3483), .Z(n3484) );
  XOR U4507 ( .A(n3485), .B(n3486), .Z(n3483) );
  ANDN U4508 ( .B(n3487), .A(n886), .Z(n3485) );
  XOR U4509 ( .A(b[202]), .B(n3486), .Z(n3487) );
  XOR U4510 ( .A(n3488), .B(n3489), .Z(n3486) );
  ANDN U4511 ( .B(n3490), .A(n887), .Z(n3488) );
  XOR U4512 ( .A(b[201]), .B(n3489), .Z(n3490) );
  XOR U4513 ( .A(n3491), .B(n3492), .Z(n3489) );
  ANDN U4514 ( .B(n3493), .A(n888), .Z(n3491) );
  XOR U4515 ( .A(b[200]), .B(n3492), .Z(n3493) );
  XOR U4516 ( .A(n3494), .B(n3495), .Z(n3492) );
  ANDN U4517 ( .B(n3496), .A(n891), .Z(n3494) );
  XOR U4518 ( .A(b[199]), .B(n3495), .Z(n3496) );
  XOR U4519 ( .A(n3497), .B(n3498), .Z(n3495) );
  ANDN U4520 ( .B(n3499), .A(n892), .Z(n3497) );
  XOR U4521 ( .A(b[198]), .B(n3498), .Z(n3499) );
  XOR U4522 ( .A(n3500), .B(n3501), .Z(n3498) );
  ANDN U4523 ( .B(n3502), .A(n893), .Z(n3500) );
  XOR U4524 ( .A(b[197]), .B(n3501), .Z(n3502) );
  XOR U4525 ( .A(n3503), .B(n3504), .Z(n3501) );
  ANDN U4526 ( .B(n3505), .A(n894), .Z(n3503) );
  XOR U4527 ( .A(b[196]), .B(n3504), .Z(n3505) );
  XOR U4528 ( .A(n3506), .B(n3507), .Z(n3504) );
  ANDN U4529 ( .B(n3508), .A(n895), .Z(n3506) );
  XOR U4530 ( .A(b[195]), .B(n3507), .Z(n3508) );
  XOR U4531 ( .A(n3509), .B(n3510), .Z(n3507) );
  ANDN U4532 ( .B(n3511), .A(n896), .Z(n3509) );
  XOR U4533 ( .A(b[194]), .B(n3510), .Z(n3511) );
  XOR U4534 ( .A(n3512), .B(n3513), .Z(n3510) );
  ANDN U4535 ( .B(n3514), .A(n897), .Z(n3512) );
  XOR U4536 ( .A(b[193]), .B(n3513), .Z(n3514) );
  XOR U4537 ( .A(n3515), .B(n3516), .Z(n3513) );
  ANDN U4538 ( .B(n3517), .A(n898), .Z(n3515) );
  XOR U4539 ( .A(b[192]), .B(n3516), .Z(n3517) );
  XOR U4540 ( .A(n3518), .B(n3519), .Z(n3516) );
  ANDN U4541 ( .B(n3520), .A(n899), .Z(n3518) );
  XOR U4542 ( .A(b[191]), .B(n3519), .Z(n3520) );
  XOR U4543 ( .A(n3521), .B(n3522), .Z(n3519) );
  ANDN U4544 ( .B(n3523), .A(n900), .Z(n3521) );
  XOR U4545 ( .A(b[190]), .B(n3522), .Z(n3523) );
  XOR U4546 ( .A(n3524), .B(n3525), .Z(n3522) );
  ANDN U4547 ( .B(n3526), .A(n902), .Z(n3524) );
  XOR U4548 ( .A(b[189]), .B(n3525), .Z(n3526) );
  XOR U4549 ( .A(n3527), .B(n3528), .Z(n3525) );
  ANDN U4550 ( .B(n3529), .A(n903), .Z(n3527) );
  XOR U4551 ( .A(b[188]), .B(n3528), .Z(n3529) );
  XOR U4552 ( .A(n3530), .B(n3531), .Z(n3528) );
  ANDN U4553 ( .B(n3532), .A(n904), .Z(n3530) );
  XOR U4554 ( .A(b[187]), .B(n3531), .Z(n3532) );
  XOR U4555 ( .A(n3533), .B(n3534), .Z(n3531) );
  ANDN U4556 ( .B(n3535), .A(n905), .Z(n3533) );
  XOR U4557 ( .A(b[186]), .B(n3534), .Z(n3535) );
  XOR U4558 ( .A(n3536), .B(n3537), .Z(n3534) );
  ANDN U4559 ( .B(n3538), .A(n906), .Z(n3536) );
  XOR U4560 ( .A(b[185]), .B(n3537), .Z(n3538) );
  XOR U4561 ( .A(n3539), .B(n3540), .Z(n3537) );
  ANDN U4562 ( .B(n3541), .A(n907), .Z(n3539) );
  XOR U4563 ( .A(b[184]), .B(n3540), .Z(n3541) );
  XOR U4564 ( .A(n3542), .B(n3543), .Z(n3540) );
  ANDN U4565 ( .B(n3544), .A(n908), .Z(n3542) );
  XOR U4566 ( .A(b[183]), .B(n3543), .Z(n3544) );
  XOR U4567 ( .A(n3545), .B(n3546), .Z(n3543) );
  ANDN U4568 ( .B(n3547), .A(n909), .Z(n3545) );
  XOR U4569 ( .A(b[182]), .B(n3546), .Z(n3547) );
  XOR U4570 ( .A(n3548), .B(n3549), .Z(n3546) );
  ANDN U4571 ( .B(n3550), .A(n910), .Z(n3548) );
  XOR U4572 ( .A(b[181]), .B(n3549), .Z(n3550) );
  XOR U4573 ( .A(n3551), .B(n3552), .Z(n3549) );
  ANDN U4574 ( .B(n3553), .A(n911), .Z(n3551) );
  XOR U4575 ( .A(b[180]), .B(n3552), .Z(n3553) );
  XOR U4576 ( .A(n3554), .B(n3555), .Z(n3552) );
  ANDN U4577 ( .B(n3556), .A(n913), .Z(n3554) );
  XOR U4578 ( .A(b[179]), .B(n3555), .Z(n3556) );
  XOR U4579 ( .A(n3557), .B(n3558), .Z(n3555) );
  ANDN U4580 ( .B(n3559), .A(n914), .Z(n3557) );
  XOR U4581 ( .A(b[178]), .B(n3558), .Z(n3559) );
  XOR U4582 ( .A(n3560), .B(n3561), .Z(n3558) );
  ANDN U4583 ( .B(n3562), .A(n915), .Z(n3560) );
  XOR U4584 ( .A(b[177]), .B(n3561), .Z(n3562) );
  XOR U4585 ( .A(n3563), .B(n3564), .Z(n3561) );
  ANDN U4586 ( .B(n3565), .A(n916), .Z(n3563) );
  XOR U4587 ( .A(b[176]), .B(n3564), .Z(n3565) );
  XOR U4588 ( .A(n3566), .B(n3567), .Z(n3564) );
  ANDN U4589 ( .B(n3568), .A(n917), .Z(n3566) );
  XOR U4590 ( .A(b[175]), .B(n3567), .Z(n3568) );
  XOR U4591 ( .A(n3569), .B(n3570), .Z(n3567) );
  ANDN U4592 ( .B(n3571), .A(n918), .Z(n3569) );
  XOR U4593 ( .A(b[174]), .B(n3570), .Z(n3571) );
  XOR U4594 ( .A(n3572), .B(n3573), .Z(n3570) );
  ANDN U4595 ( .B(n3574), .A(n919), .Z(n3572) );
  XOR U4596 ( .A(b[173]), .B(n3573), .Z(n3574) );
  XOR U4597 ( .A(n3575), .B(n3576), .Z(n3573) );
  ANDN U4598 ( .B(n3577), .A(n920), .Z(n3575) );
  XOR U4599 ( .A(b[172]), .B(n3576), .Z(n3577) );
  XOR U4600 ( .A(n3578), .B(n3579), .Z(n3576) );
  ANDN U4601 ( .B(n3580), .A(n921), .Z(n3578) );
  XOR U4602 ( .A(b[171]), .B(n3579), .Z(n3580) );
  XOR U4603 ( .A(n3581), .B(n3582), .Z(n3579) );
  ANDN U4604 ( .B(n3583), .A(n922), .Z(n3581) );
  XOR U4605 ( .A(b[170]), .B(n3582), .Z(n3583) );
  XOR U4606 ( .A(n3584), .B(n3585), .Z(n3582) );
  ANDN U4607 ( .B(n3586), .A(n924), .Z(n3584) );
  XOR U4608 ( .A(b[169]), .B(n3585), .Z(n3586) );
  XOR U4609 ( .A(n3587), .B(n3588), .Z(n3585) );
  ANDN U4610 ( .B(n3589), .A(n925), .Z(n3587) );
  XOR U4611 ( .A(b[168]), .B(n3588), .Z(n3589) );
  XOR U4612 ( .A(n3590), .B(n3591), .Z(n3588) );
  ANDN U4613 ( .B(n3592), .A(n926), .Z(n3590) );
  XOR U4614 ( .A(b[167]), .B(n3591), .Z(n3592) );
  XOR U4615 ( .A(n3593), .B(n3594), .Z(n3591) );
  ANDN U4616 ( .B(n3595), .A(n927), .Z(n3593) );
  XOR U4617 ( .A(b[166]), .B(n3594), .Z(n3595) );
  XOR U4618 ( .A(n3596), .B(n3597), .Z(n3594) );
  ANDN U4619 ( .B(n3598), .A(n928), .Z(n3596) );
  XOR U4620 ( .A(b[165]), .B(n3597), .Z(n3598) );
  XOR U4621 ( .A(n3599), .B(n3600), .Z(n3597) );
  ANDN U4622 ( .B(n3601), .A(n929), .Z(n3599) );
  XOR U4623 ( .A(b[164]), .B(n3600), .Z(n3601) );
  XOR U4624 ( .A(n3602), .B(n3603), .Z(n3600) );
  ANDN U4625 ( .B(n3604), .A(n930), .Z(n3602) );
  XOR U4626 ( .A(b[163]), .B(n3603), .Z(n3604) );
  XOR U4627 ( .A(n3605), .B(n3606), .Z(n3603) );
  ANDN U4628 ( .B(n3607), .A(n931), .Z(n3605) );
  XOR U4629 ( .A(b[162]), .B(n3606), .Z(n3607) );
  XOR U4630 ( .A(n3608), .B(n3609), .Z(n3606) );
  ANDN U4631 ( .B(n3610), .A(n932), .Z(n3608) );
  XOR U4632 ( .A(b[161]), .B(n3609), .Z(n3610) );
  XOR U4633 ( .A(n3611), .B(n3612), .Z(n3609) );
  ANDN U4634 ( .B(n3613), .A(n933), .Z(n3611) );
  XOR U4635 ( .A(b[160]), .B(n3612), .Z(n3613) );
  XOR U4636 ( .A(n3614), .B(n3615), .Z(n3612) );
  ANDN U4637 ( .B(n3616), .A(n935), .Z(n3614) );
  XOR U4638 ( .A(b[159]), .B(n3615), .Z(n3616) );
  XOR U4639 ( .A(n3617), .B(n3618), .Z(n3615) );
  ANDN U4640 ( .B(n3619), .A(n936), .Z(n3617) );
  XOR U4641 ( .A(b[158]), .B(n3618), .Z(n3619) );
  XOR U4642 ( .A(n3620), .B(n3621), .Z(n3618) );
  ANDN U4643 ( .B(n3622), .A(n937), .Z(n3620) );
  XOR U4644 ( .A(b[157]), .B(n3621), .Z(n3622) );
  XOR U4645 ( .A(n3623), .B(n3624), .Z(n3621) );
  ANDN U4646 ( .B(n3625), .A(n938), .Z(n3623) );
  XOR U4647 ( .A(b[156]), .B(n3624), .Z(n3625) );
  XOR U4648 ( .A(n3626), .B(n3627), .Z(n3624) );
  ANDN U4649 ( .B(n3628), .A(n939), .Z(n3626) );
  XOR U4650 ( .A(b[155]), .B(n3627), .Z(n3628) );
  XOR U4651 ( .A(n3629), .B(n3630), .Z(n3627) );
  ANDN U4652 ( .B(n3631), .A(n940), .Z(n3629) );
  XOR U4653 ( .A(b[154]), .B(n3630), .Z(n3631) );
  XOR U4654 ( .A(n3632), .B(n3633), .Z(n3630) );
  ANDN U4655 ( .B(n3634), .A(n941), .Z(n3632) );
  XOR U4656 ( .A(b[153]), .B(n3633), .Z(n3634) );
  XOR U4657 ( .A(n3635), .B(n3636), .Z(n3633) );
  ANDN U4658 ( .B(n3637), .A(n942), .Z(n3635) );
  XOR U4659 ( .A(b[152]), .B(n3636), .Z(n3637) );
  XOR U4660 ( .A(n3638), .B(n3639), .Z(n3636) );
  ANDN U4661 ( .B(n3640), .A(n943), .Z(n3638) );
  XOR U4662 ( .A(b[151]), .B(n3639), .Z(n3640) );
  XOR U4663 ( .A(n3641), .B(n3642), .Z(n3639) );
  ANDN U4664 ( .B(n3643), .A(n944), .Z(n3641) );
  XOR U4665 ( .A(b[150]), .B(n3642), .Z(n3643) );
  XOR U4666 ( .A(n3644), .B(n3645), .Z(n3642) );
  ANDN U4667 ( .B(n3646), .A(n946), .Z(n3644) );
  XOR U4668 ( .A(b[149]), .B(n3645), .Z(n3646) );
  XOR U4669 ( .A(n3647), .B(n3648), .Z(n3645) );
  ANDN U4670 ( .B(n3649), .A(n947), .Z(n3647) );
  XOR U4671 ( .A(b[148]), .B(n3648), .Z(n3649) );
  XOR U4672 ( .A(n3650), .B(n3651), .Z(n3648) );
  ANDN U4673 ( .B(n3652), .A(n948), .Z(n3650) );
  XOR U4674 ( .A(b[147]), .B(n3651), .Z(n3652) );
  XOR U4675 ( .A(n3653), .B(n3654), .Z(n3651) );
  ANDN U4676 ( .B(n3655), .A(n949), .Z(n3653) );
  XOR U4677 ( .A(b[146]), .B(n3654), .Z(n3655) );
  XOR U4678 ( .A(n3656), .B(n3657), .Z(n3654) );
  ANDN U4679 ( .B(n3658), .A(n950), .Z(n3656) );
  XOR U4680 ( .A(b[145]), .B(n3657), .Z(n3658) );
  XOR U4681 ( .A(n3659), .B(n3660), .Z(n3657) );
  ANDN U4682 ( .B(n3661), .A(n951), .Z(n3659) );
  XOR U4683 ( .A(b[144]), .B(n3660), .Z(n3661) );
  XOR U4684 ( .A(n3662), .B(n3663), .Z(n3660) );
  ANDN U4685 ( .B(n3664), .A(n952), .Z(n3662) );
  XOR U4686 ( .A(b[143]), .B(n3663), .Z(n3664) );
  XOR U4687 ( .A(n3665), .B(n3666), .Z(n3663) );
  ANDN U4688 ( .B(n3667), .A(n953), .Z(n3665) );
  XOR U4689 ( .A(b[142]), .B(n3666), .Z(n3667) );
  XOR U4690 ( .A(n3668), .B(n3669), .Z(n3666) );
  ANDN U4691 ( .B(n3670), .A(n954), .Z(n3668) );
  XOR U4692 ( .A(b[141]), .B(n3669), .Z(n3670) );
  XOR U4693 ( .A(n3671), .B(n3672), .Z(n3669) );
  ANDN U4694 ( .B(n3673), .A(n955), .Z(n3671) );
  XOR U4695 ( .A(b[140]), .B(n3672), .Z(n3673) );
  XOR U4696 ( .A(n3674), .B(n3675), .Z(n3672) );
  ANDN U4697 ( .B(n3676), .A(n957), .Z(n3674) );
  XOR U4698 ( .A(b[139]), .B(n3675), .Z(n3676) );
  XOR U4699 ( .A(n3677), .B(n3678), .Z(n3675) );
  ANDN U4700 ( .B(n3679), .A(n958), .Z(n3677) );
  XOR U4701 ( .A(b[138]), .B(n3678), .Z(n3679) );
  XOR U4702 ( .A(n3680), .B(n3681), .Z(n3678) );
  ANDN U4703 ( .B(n3682), .A(n959), .Z(n3680) );
  XOR U4704 ( .A(b[137]), .B(n3681), .Z(n3682) );
  XOR U4705 ( .A(n3683), .B(n3684), .Z(n3681) );
  ANDN U4706 ( .B(n3685), .A(n960), .Z(n3683) );
  XOR U4707 ( .A(b[136]), .B(n3684), .Z(n3685) );
  XOR U4708 ( .A(n3686), .B(n3687), .Z(n3684) );
  ANDN U4709 ( .B(n3688), .A(n961), .Z(n3686) );
  XOR U4710 ( .A(b[135]), .B(n3687), .Z(n3688) );
  XOR U4711 ( .A(n3689), .B(n3690), .Z(n3687) );
  ANDN U4712 ( .B(n3691), .A(n962), .Z(n3689) );
  XOR U4713 ( .A(b[134]), .B(n3690), .Z(n3691) );
  XOR U4714 ( .A(n3692), .B(n3693), .Z(n3690) );
  ANDN U4715 ( .B(n3694), .A(n963), .Z(n3692) );
  XOR U4716 ( .A(b[133]), .B(n3693), .Z(n3694) );
  XOR U4717 ( .A(n3695), .B(n3696), .Z(n3693) );
  ANDN U4718 ( .B(n3697), .A(n964), .Z(n3695) );
  XOR U4719 ( .A(b[132]), .B(n3696), .Z(n3697) );
  XOR U4720 ( .A(n3698), .B(n3699), .Z(n3696) );
  ANDN U4721 ( .B(n3700), .A(n965), .Z(n3698) );
  XOR U4722 ( .A(b[131]), .B(n3699), .Z(n3700) );
  XOR U4723 ( .A(n3701), .B(n3702), .Z(n3699) );
  ANDN U4724 ( .B(n3703), .A(n966), .Z(n3701) );
  XOR U4725 ( .A(b[130]), .B(n3702), .Z(n3703) );
  XOR U4726 ( .A(n3704), .B(n3705), .Z(n3702) );
  ANDN U4727 ( .B(n3706), .A(n968), .Z(n3704) );
  XOR U4728 ( .A(b[129]), .B(n3705), .Z(n3706) );
  XOR U4729 ( .A(n3707), .B(n3708), .Z(n3705) );
  ANDN U4730 ( .B(n3709), .A(n969), .Z(n3707) );
  XOR U4731 ( .A(b[128]), .B(n3708), .Z(n3709) );
  XOR U4732 ( .A(n3710), .B(n3711), .Z(n3708) );
  ANDN U4733 ( .B(n3712), .A(n970), .Z(n3710) );
  XOR U4734 ( .A(b[127]), .B(n3711), .Z(n3712) );
  XOR U4735 ( .A(n3713), .B(n3714), .Z(n3711) );
  ANDN U4736 ( .B(n3715), .A(n971), .Z(n3713) );
  XOR U4737 ( .A(b[126]), .B(n3714), .Z(n3715) );
  XOR U4738 ( .A(n3716), .B(n3717), .Z(n3714) );
  ANDN U4739 ( .B(n3718), .A(n972), .Z(n3716) );
  XOR U4740 ( .A(b[125]), .B(n3717), .Z(n3718) );
  XOR U4741 ( .A(n3719), .B(n3720), .Z(n3717) );
  ANDN U4742 ( .B(n3721), .A(n973), .Z(n3719) );
  XOR U4743 ( .A(b[124]), .B(n3720), .Z(n3721) );
  XOR U4744 ( .A(n3722), .B(n3723), .Z(n3720) );
  ANDN U4745 ( .B(n3724), .A(n974), .Z(n3722) );
  XOR U4746 ( .A(b[123]), .B(n3723), .Z(n3724) );
  XOR U4747 ( .A(n3725), .B(n3726), .Z(n3723) );
  ANDN U4748 ( .B(n3727), .A(n975), .Z(n3725) );
  XOR U4749 ( .A(b[122]), .B(n3726), .Z(n3727) );
  XOR U4750 ( .A(n3728), .B(n3729), .Z(n3726) );
  ANDN U4751 ( .B(n3730), .A(n976), .Z(n3728) );
  XOR U4752 ( .A(b[121]), .B(n3729), .Z(n3730) );
  XOR U4753 ( .A(n3731), .B(n3732), .Z(n3729) );
  ANDN U4754 ( .B(n3733), .A(n977), .Z(n3731) );
  XOR U4755 ( .A(b[120]), .B(n3732), .Z(n3733) );
  XOR U4756 ( .A(n3734), .B(n3735), .Z(n3732) );
  ANDN U4757 ( .B(n3736), .A(n979), .Z(n3734) );
  XOR U4758 ( .A(b[119]), .B(n3735), .Z(n3736) );
  XOR U4759 ( .A(n3737), .B(n3738), .Z(n3735) );
  ANDN U4760 ( .B(n3739), .A(n980), .Z(n3737) );
  XOR U4761 ( .A(b[118]), .B(n3738), .Z(n3739) );
  XOR U4762 ( .A(n3740), .B(n3741), .Z(n3738) );
  ANDN U4763 ( .B(n3742), .A(n981), .Z(n3740) );
  XOR U4764 ( .A(b[117]), .B(n3741), .Z(n3742) );
  XOR U4765 ( .A(n3743), .B(n3744), .Z(n3741) );
  ANDN U4766 ( .B(n3745), .A(n982), .Z(n3743) );
  XOR U4767 ( .A(b[116]), .B(n3744), .Z(n3745) );
  XOR U4768 ( .A(n3746), .B(n3747), .Z(n3744) );
  ANDN U4769 ( .B(n3748), .A(n983), .Z(n3746) );
  XOR U4770 ( .A(b[115]), .B(n3747), .Z(n3748) );
  XOR U4771 ( .A(n3749), .B(n3750), .Z(n3747) );
  ANDN U4772 ( .B(n3751), .A(n984), .Z(n3749) );
  XOR U4773 ( .A(b[114]), .B(n3750), .Z(n3751) );
  XOR U4774 ( .A(n3752), .B(n3753), .Z(n3750) );
  ANDN U4775 ( .B(n3754), .A(n985), .Z(n3752) );
  XOR U4776 ( .A(b[113]), .B(n3753), .Z(n3754) );
  XOR U4777 ( .A(n3755), .B(n3756), .Z(n3753) );
  ANDN U4778 ( .B(n3757), .A(n986), .Z(n3755) );
  XOR U4779 ( .A(b[112]), .B(n3756), .Z(n3757) );
  XOR U4780 ( .A(n3758), .B(n3759), .Z(n3756) );
  ANDN U4781 ( .B(n3760), .A(n987), .Z(n3758) );
  XOR U4782 ( .A(b[111]), .B(n3759), .Z(n3760) );
  XOR U4783 ( .A(n3761), .B(n3762), .Z(n3759) );
  ANDN U4784 ( .B(n3763), .A(n988), .Z(n3761) );
  XOR U4785 ( .A(b[110]), .B(n3762), .Z(n3763) );
  XOR U4786 ( .A(n3764), .B(n3765), .Z(n3762) );
  ANDN U4787 ( .B(n3766), .A(n990), .Z(n3764) );
  XOR U4788 ( .A(b[109]), .B(n3765), .Z(n3766) );
  XOR U4789 ( .A(n3767), .B(n3768), .Z(n3765) );
  ANDN U4790 ( .B(n3769), .A(n991), .Z(n3767) );
  XOR U4791 ( .A(b[108]), .B(n3768), .Z(n3769) );
  XOR U4792 ( .A(n3770), .B(n3771), .Z(n3768) );
  ANDN U4793 ( .B(n3772), .A(n992), .Z(n3770) );
  XOR U4794 ( .A(b[107]), .B(n3771), .Z(n3772) );
  XOR U4795 ( .A(n3773), .B(n3774), .Z(n3771) );
  ANDN U4796 ( .B(n3775), .A(n993), .Z(n3773) );
  XOR U4797 ( .A(b[106]), .B(n3774), .Z(n3775) );
  XOR U4798 ( .A(n3776), .B(n3777), .Z(n3774) );
  ANDN U4799 ( .B(n3778), .A(n994), .Z(n3776) );
  XOR U4800 ( .A(b[105]), .B(n3777), .Z(n3778) );
  XOR U4801 ( .A(n3779), .B(n3780), .Z(n3777) );
  ANDN U4802 ( .B(n3781), .A(n995), .Z(n3779) );
  XOR U4803 ( .A(b[104]), .B(n3780), .Z(n3781) );
  XOR U4804 ( .A(n3782), .B(n3783), .Z(n3780) );
  ANDN U4805 ( .B(n3784), .A(n996), .Z(n3782) );
  XOR U4806 ( .A(b[103]), .B(n3783), .Z(n3784) );
  XOR U4807 ( .A(n3785), .B(n3786), .Z(n3783) );
  ANDN U4808 ( .B(n3787), .A(n997), .Z(n3785) );
  XOR U4809 ( .A(b[102]), .B(n3786), .Z(n3787) );
  XOR U4810 ( .A(n3788), .B(n3789), .Z(n3786) );
  ANDN U4811 ( .B(n3790), .A(n1016), .Z(n3788) );
  XOR U4812 ( .A(b[101]), .B(n3789), .Z(n3790) );
  XOR U4813 ( .A(n3791), .B(n3792), .Z(n3789) );
  ANDN U4814 ( .B(n3793), .A(n1057), .Z(n3791) );
  XOR U4815 ( .A(b[100]), .B(n3792), .Z(n3793) );
  XOR U4816 ( .A(n3794), .B(n3795), .Z(n3792) );
  ANDN U4817 ( .B(n3796), .A(n2), .Z(n3794) );
  XOR U4818 ( .A(b[99]), .B(n3795), .Z(n3796) );
  XOR U4819 ( .A(n3797), .B(n3798), .Z(n3795) );
  ANDN U4820 ( .B(n3799), .A(n13), .Z(n3797) );
  XOR U4821 ( .A(b[98]), .B(n3798), .Z(n3799) );
  XOR U4822 ( .A(n3800), .B(n3801), .Z(n3798) );
  ANDN U4823 ( .B(n3802), .A(n24), .Z(n3800) );
  XOR U4824 ( .A(b[97]), .B(n3801), .Z(n3802) );
  XOR U4825 ( .A(n3803), .B(n3804), .Z(n3801) );
  ANDN U4826 ( .B(n3805), .A(n35), .Z(n3803) );
  XOR U4827 ( .A(b[96]), .B(n3804), .Z(n3805) );
  XOR U4828 ( .A(n3806), .B(n3807), .Z(n3804) );
  ANDN U4829 ( .B(n3808), .A(n46), .Z(n3806) );
  XOR U4830 ( .A(b[95]), .B(n3807), .Z(n3808) );
  XOR U4831 ( .A(n3809), .B(n3810), .Z(n3807) );
  ANDN U4832 ( .B(n3811), .A(n57), .Z(n3809) );
  XOR U4833 ( .A(b[94]), .B(n3810), .Z(n3811) );
  XOR U4834 ( .A(n3812), .B(n3813), .Z(n3810) );
  ANDN U4835 ( .B(n3814), .A(n68), .Z(n3812) );
  XOR U4836 ( .A(b[93]), .B(n3813), .Z(n3814) );
  XOR U4837 ( .A(n3815), .B(n3816), .Z(n3813) );
  ANDN U4838 ( .B(n3817), .A(n79), .Z(n3815) );
  XOR U4839 ( .A(b[92]), .B(n3816), .Z(n3817) );
  XOR U4840 ( .A(n3818), .B(n3819), .Z(n3816) );
  ANDN U4841 ( .B(n3820), .A(n90), .Z(n3818) );
  XOR U4842 ( .A(b[91]), .B(n3819), .Z(n3820) );
  XOR U4843 ( .A(n3821), .B(n3822), .Z(n3819) );
  ANDN U4844 ( .B(n3823), .A(n101), .Z(n3821) );
  XOR U4845 ( .A(b[90]), .B(n3822), .Z(n3823) );
  XOR U4846 ( .A(n3824), .B(n3825), .Z(n3822) );
  ANDN U4847 ( .B(n3826), .A(n113), .Z(n3824) );
  XOR U4848 ( .A(b[89]), .B(n3825), .Z(n3826) );
  XOR U4849 ( .A(n3827), .B(n3828), .Z(n3825) );
  ANDN U4850 ( .B(n3829), .A(n124), .Z(n3827) );
  XOR U4851 ( .A(b[88]), .B(n3828), .Z(n3829) );
  XOR U4852 ( .A(n3830), .B(n3831), .Z(n3828) );
  ANDN U4853 ( .B(n3832), .A(n135), .Z(n3830) );
  XOR U4854 ( .A(b[87]), .B(n3831), .Z(n3832) );
  XOR U4855 ( .A(n3833), .B(n3834), .Z(n3831) );
  ANDN U4856 ( .B(n3835), .A(n146), .Z(n3833) );
  XOR U4857 ( .A(b[86]), .B(n3834), .Z(n3835) );
  XOR U4858 ( .A(n3836), .B(n3837), .Z(n3834) );
  ANDN U4859 ( .B(n3838), .A(n157), .Z(n3836) );
  XOR U4860 ( .A(b[85]), .B(n3837), .Z(n3838) );
  XOR U4861 ( .A(n3839), .B(n3840), .Z(n3837) );
  ANDN U4862 ( .B(n3841), .A(n168), .Z(n3839) );
  XOR U4863 ( .A(b[84]), .B(n3840), .Z(n3841) );
  XOR U4864 ( .A(n3842), .B(n3843), .Z(n3840) );
  ANDN U4865 ( .B(n3844), .A(n179), .Z(n3842) );
  XOR U4866 ( .A(b[83]), .B(n3843), .Z(n3844) );
  XOR U4867 ( .A(n3845), .B(n3846), .Z(n3843) );
  ANDN U4868 ( .B(n3847), .A(n190), .Z(n3845) );
  XOR U4869 ( .A(b[82]), .B(n3846), .Z(n3847) );
  XOR U4870 ( .A(n3848), .B(n3849), .Z(n3846) );
  ANDN U4871 ( .B(n3850), .A(n201), .Z(n3848) );
  XOR U4872 ( .A(b[81]), .B(n3849), .Z(n3850) );
  XOR U4873 ( .A(n3851), .B(n3852), .Z(n3849) );
  ANDN U4874 ( .B(n3853), .A(n212), .Z(n3851) );
  XOR U4875 ( .A(b[80]), .B(n3852), .Z(n3853) );
  XOR U4876 ( .A(n3854), .B(n3855), .Z(n3852) );
  ANDN U4877 ( .B(n3856), .A(n224), .Z(n3854) );
  XOR U4878 ( .A(b[79]), .B(n3855), .Z(n3856) );
  XOR U4879 ( .A(n3857), .B(n3858), .Z(n3855) );
  ANDN U4880 ( .B(n3859), .A(n235), .Z(n3857) );
  XOR U4881 ( .A(b[78]), .B(n3858), .Z(n3859) );
  XOR U4882 ( .A(n3860), .B(n3861), .Z(n3858) );
  ANDN U4883 ( .B(n3862), .A(n246), .Z(n3860) );
  XOR U4884 ( .A(b[77]), .B(n3861), .Z(n3862) );
  XOR U4885 ( .A(n3863), .B(n3864), .Z(n3861) );
  ANDN U4886 ( .B(n3865), .A(n257), .Z(n3863) );
  XOR U4887 ( .A(b[76]), .B(n3864), .Z(n3865) );
  XOR U4888 ( .A(n3866), .B(n3867), .Z(n3864) );
  ANDN U4889 ( .B(n3868), .A(n268), .Z(n3866) );
  XOR U4890 ( .A(b[75]), .B(n3867), .Z(n3868) );
  XOR U4891 ( .A(n3869), .B(n3870), .Z(n3867) );
  ANDN U4892 ( .B(n3871), .A(n279), .Z(n3869) );
  XOR U4893 ( .A(b[74]), .B(n3870), .Z(n3871) );
  XOR U4894 ( .A(n3872), .B(n3873), .Z(n3870) );
  ANDN U4895 ( .B(n3874), .A(n290), .Z(n3872) );
  XOR U4896 ( .A(b[73]), .B(n3873), .Z(n3874) );
  XOR U4897 ( .A(n3875), .B(n3876), .Z(n3873) );
  ANDN U4898 ( .B(n3877), .A(n301), .Z(n3875) );
  XOR U4899 ( .A(b[72]), .B(n3876), .Z(n3877) );
  XOR U4900 ( .A(n3878), .B(n3879), .Z(n3876) );
  ANDN U4901 ( .B(n3880), .A(n312), .Z(n3878) );
  XOR U4902 ( .A(b[71]), .B(n3879), .Z(n3880) );
  XOR U4903 ( .A(n3881), .B(n3882), .Z(n3879) );
  ANDN U4904 ( .B(n3883), .A(n323), .Z(n3881) );
  XOR U4905 ( .A(b[70]), .B(n3882), .Z(n3883) );
  XOR U4906 ( .A(n3884), .B(n3885), .Z(n3882) );
  ANDN U4907 ( .B(n3886), .A(n335), .Z(n3884) );
  XOR U4908 ( .A(b[69]), .B(n3885), .Z(n3886) );
  XOR U4909 ( .A(n3887), .B(n3888), .Z(n3885) );
  ANDN U4910 ( .B(n3889), .A(n346), .Z(n3887) );
  XOR U4911 ( .A(b[68]), .B(n3888), .Z(n3889) );
  XOR U4912 ( .A(n3890), .B(n3891), .Z(n3888) );
  ANDN U4913 ( .B(n3892), .A(n357), .Z(n3890) );
  XOR U4914 ( .A(b[67]), .B(n3891), .Z(n3892) );
  XOR U4915 ( .A(n3893), .B(n3894), .Z(n3891) );
  ANDN U4916 ( .B(n3895), .A(n368), .Z(n3893) );
  XOR U4917 ( .A(b[66]), .B(n3894), .Z(n3895) );
  XOR U4918 ( .A(n3896), .B(n3897), .Z(n3894) );
  ANDN U4919 ( .B(n3898), .A(n379), .Z(n3896) );
  XOR U4920 ( .A(b[65]), .B(n3897), .Z(n3898) );
  XOR U4921 ( .A(n3899), .B(n3900), .Z(n3897) );
  ANDN U4922 ( .B(n3901), .A(n390), .Z(n3899) );
  XOR U4923 ( .A(b[64]), .B(n3900), .Z(n3901) );
  XOR U4924 ( .A(n3902), .B(n3903), .Z(n3900) );
  ANDN U4925 ( .B(n3904), .A(n401), .Z(n3902) );
  XOR U4926 ( .A(b[63]), .B(n3903), .Z(n3904) );
  XOR U4927 ( .A(n3905), .B(n3906), .Z(n3903) );
  ANDN U4928 ( .B(n3907), .A(n412), .Z(n3905) );
  XOR U4929 ( .A(b[62]), .B(n3906), .Z(n3907) );
  XOR U4930 ( .A(n3908), .B(n3909), .Z(n3906) );
  ANDN U4931 ( .B(n3910), .A(n423), .Z(n3908) );
  XOR U4932 ( .A(b[61]), .B(n3909), .Z(n3910) );
  XOR U4933 ( .A(n3911), .B(n3912), .Z(n3909) );
  ANDN U4934 ( .B(n3913), .A(n434), .Z(n3911) );
  XOR U4935 ( .A(b[60]), .B(n3912), .Z(n3913) );
  XOR U4936 ( .A(n3914), .B(n3915), .Z(n3912) );
  ANDN U4937 ( .B(n3916), .A(n446), .Z(n3914) );
  XOR U4938 ( .A(b[59]), .B(n3915), .Z(n3916) );
  XOR U4939 ( .A(n3917), .B(n3918), .Z(n3915) );
  ANDN U4940 ( .B(n3919), .A(n457), .Z(n3917) );
  XOR U4941 ( .A(b[58]), .B(n3918), .Z(n3919) );
  XOR U4942 ( .A(n3920), .B(n3921), .Z(n3918) );
  ANDN U4943 ( .B(n3922), .A(n468), .Z(n3920) );
  XOR U4944 ( .A(b[57]), .B(n3921), .Z(n3922) );
  XOR U4945 ( .A(n3923), .B(n3924), .Z(n3921) );
  ANDN U4946 ( .B(n3925), .A(n479), .Z(n3923) );
  XOR U4947 ( .A(b[56]), .B(n3924), .Z(n3925) );
  XOR U4948 ( .A(n3926), .B(n3927), .Z(n3924) );
  ANDN U4949 ( .B(n3928), .A(n490), .Z(n3926) );
  XOR U4950 ( .A(b[55]), .B(n3927), .Z(n3928) );
  XOR U4951 ( .A(n3929), .B(n3930), .Z(n3927) );
  ANDN U4952 ( .B(n3931), .A(n501), .Z(n3929) );
  XOR U4953 ( .A(b[54]), .B(n3930), .Z(n3931) );
  XOR U4954 ( .A(n3932), .B(n3933), .Z(n3930) );
  ANDN U4955 ( .B(n3934), .A(n512), .Z(n3932) );
  XOR U4956 ( .A(b[53]), .B(n3933), .Z(n3934) );
  XOR U4957 ( .A(n3935), .B(n3936), .Z(n3933) );
  ANDN U4958 ( .B(n3937), .A(n523), .Z(n3935) );
  XOR U4959 ( .A(b[52]), .B(n3936), .Z(n3937) );
  XOR U4960 ( .A(n3938), .B(n3939), .Z(n3936) );
  ANDN U4961 ( .B(n3940), .A(n534), .Z(n3938) );
  XOR U4962 ( .A(b[51]), .B(n3939), .Z(n3940) );
  XOR U4963 ( .A(n3941), .B(n3942), .Z(n3939) );
  ANDN U4964 ( .B(n3943), .A(n545), .Z(n3941) );
  XOR U4965 ( .A(b[50]), .B(n3942), .Z(n3943) );
  XOR U4966 ( .A(n3944), .B(n3945), .Z(n3942) );
  ANDN U4967 ( .B(n3946), .A(n557), .Z(n3944) );
  XOR U4968 ( .A(b[49]), .B(n3945), .Z(n3946) );
  XOR U4969 ( .A(n3947), .B(n3948), .Z(n3945) );
  ANDN U4970 ( .B(n3949), .A(n568), .Z(n3947) );
  XOR U4971 ( .A(b[48]), .B(n3948), .Z(n3949) );
  XOR U4972 ( .A(n3950), .B(n3951), .Z(n3948) );
  ANDN U4973 ( .B(n3952), .A(n579), .Z(n3950) );
  XOR U4974 ( .A(b[47]), .B(n3951), .Z(n3952) );
  XOR U4975 ( .A(n3953), .B(n3954), .Z(n3951) );
  ANDN U4976 ( .B(n3955), .A(n590), .Z(n3953) );
  XOR U4977 ( .A(b[46]), .B(n3954), .Z(n3955) );
  XOR U4978 ( .A(n3956), .B(n3957), .Z(n3954) );
  ANDN U4979 ( .B(n3958), .A(n601), .Z(n3956) );
  XOR U4980 ( .A(b[45]), .B(n3957), .Z(n3958) );
  XOR U4981 ( .A(n3959), .B(n3960), .Z(n3957) );
  ANDN U4982 ( .B(n3961), .A(n612), .Z(n3959) );
  XOR U4983 ( .A(b[44]), .B(n3960), .Z(n3961) );
  XOR U4984 ( .A(n3962), .B(n3963), .Z(n3960) );
  ANDN U4985 ( .B(n3964), .A(n623), .Z(n3962) );
  XOR U4986 ( .A(b[43]), .B(n3963), .Z(n3964) );
  XOR U4987 ( .A(n3965), .B(n3966), .Z(n3963) );
  ANDN U4988 ( .B(n3967), .A(n634), .Z(n3965) );
  XOR U4989 ( .A(b[42]), .B(n3966), .Z(n3967) );
  XOR U4990 ( .A(n3968), .B(n3969), .Z(n3966) );
  ANDN U4991 ( .B(n3970), .A(n645), .Z(n3968) );
  XOR U4992 ( .A(b[41]), .B(n3969), .Z(n3970) );
  XOR U4993 ( .A(n3971), .B(n3972), .Z(n3969) );
  ANDN U4994 ( .B(n3973), .A(n656), .Z(n3971) );
  XOR U4995 ( .A(b[40]), .B(n3972), .Z(n3973) );
  XOR U4996 ( .A(n3974), .B(n3975), .Z(n3972) );
  ANDN U4997 ( .B(n3976), .A(n668), .Z(n3974) );
  XOR U4998 ( .A(b[39]), .B(n3975), .Z(n3976) );
  XOR U4999 ( .A(n3977), .B(n3978), .Z(n3975) );
  ANDN U5000 ( .B(n3979), .A(n679), .Z(n3977) );
  XOR U5001 ( .A(b[38]), .B(n3978), .Z(n3979) );
  XOR U5002 ( .A(n3980), .B(n3981), .Z(n3978) );
  ANDN U5003 ( .B(n3982), .A(n690), .Z(n3980) );
  XOR U5004 ( .A(b[37]), .B(n3981), .Z(n3982) );
  XOR U5005 ( .A(n3983), .B(n3984), .Z(n3981) );
  ANDN U5006 ( .B(n3985), .A(n701), .Z(n3983) );
  XOR U5007 ( .A(b[36]), .B(n3984), .Z(n3985) );
  XOR U5008 ( .A(n3986), .B(n3987), .Z(n3984) );
  ANDN U5009 ( .B(n3988), .A(n712), .Z(n3986) );
  XOR U5010 ( .A(b[35]), .B(n3987), .Z(n3988) );
  XOR U5011 ( .A(n3989), .B(n3990), .Z(n3987) );
  ANDN U5012 ( .B(n3991), .A(n723), .Z(n3989) );
  XOR U5013 ( .A(b[34]), .B(n3990), .Z(n3991) );
  XOR U5014 ( .A(n3992), .B(n3993), .Z(n3990) );
  ANDN U5015 ( .B(n3994), .A(n734), .Z(n3992) );
  XOR U5016 ( .A(b[33]), .B(n3993), .Z(n3994) );
  XOR U5017 ( .A(n3995), .B(n3996), .Z(n3993) );
  ANDN U5018 ( .B(n3997), .A(n745), .Z(n3995) );
  XOR U5019 ( .A(b[32]), .B(n3996), .Z(n3997) );
  XOR U5020 ( .A(n3998), .B(n3999), .Z(n3996) );
  ANDN U5021 ( .B(n4000), .A(n756), .Z(n3998) );
  XOR U5022 ( .A(b[31]), .B(n3999), .Z(n4000) );
  XOR U5023 ( .A(n4001), .B(n4002), .Z(n3999) );
  ANDN U5024 ( .B(n4003), .A(n767), .Z(n4001) );
  XOR U5025 ( .A(b[30]), .B(n4002), .Z(n4003) );
  XOR U5026 ( .A(n4004), .B(n4005), .Z(n4002) );
  ANDN U5027 ( .B(n4006), .A(n779), .Z(n4004) );
  XOR U5028 ( .A(b[29]), .B(n4005), .Z(n4006) );
  XOR U5029 ( .A(n4007), .B(n4008), .Z(n4005) );
  ANDN U5030 ( .B(n4009), .A(n790), .Z(n4007) );
  XOR U5031 ( .A(b[28]), .B(n4008), .Z(n4009) );
  XOR U5032 ( .A(n4010), .B(n4011), .Z(n4008) );
  ANDN U5033 ( .B(n4012), .A(n801), .Z(n4010) );
  XOR U5034 ( .A(b[27]), .B(n4011), .Z(n4012) );
  XOR U5035 ( .A(n4013), .B(n4014), .Z(n4011) );
  ANDN U5036 ( .B(n4015), .A(n812), .Z(n4013) );
  XOR U5037 ( .A(b[26]), .B(n4014), .Z(n4015) );
  XOR U5038 ( .A(n4016), .B(n4017), .Z(n4014) );
  ANDN U5039 ( .B(n4018), .A(n823), .Z(n4016) );
  XOR U5040 ( .A(b[25]), .B(n4017), .Z(n4018) );
  XOR U5041 ( .A(n4019), .B(n4020), .Z(n4017) );
  ANDN U5042 ( .B(n4021), .A(n834), .Z(n4019) );
  XOR U5043 ( .A(b[24]), .B(n4020), .Z(n4021) );
  XOR U5044 ( .A(n4022), .B(n4023), .Z(n4020) );
  ANDN U5045 ( .B(n4024), .A(n845), .Z(n4022) );
  XOR U5046 ( .A(b[23]), .B(n4023), .Z(n4024) );
  XOR U5047 ( .A(n4025), .B(n4026), .Z(n4023) );
  ANDN U5048 ( .B(n4027), .A(n856), .Z(n4025) );
  XOR U5049 ( .A(b[22]), .B(n4026), .Z(n4027) );
  XOR U5050 ( .A(n4028), .B(n4029), .Z(n4026) );
  ANDN U5051 ( .B(n4030), .A(n867), .Z(n4028) );
  XOR U5052 ( .A(b[21]), .B(n4029), .Z(n4030) );
  XOR U5053 ( .A(n4031), .B(n4032), .Z(n4029) );
  ANDN U5054 ( .B(n4033), .A(n878), .Z(n4031) );
  XOR U5055 ( .A(b[20]), .B(n4032), .Z(n4033) );
  XOR U5056 ( .A(n4034), .B(n4035), .Z(n4032) );
  ANDN U5057 ( .B(n4036), .A(n890), .Z(n4034) );
  XOR U5058 ( .A(b[19]), .B(n4035), .Z(n4036) );
  XOR U5059 ( .A(n4037), .B(n4038), .Z(n4035) );
  ANDN U5060 ( .B(n4039), .A(n901), .Z(n4037) );
  XOR U5061 ( .A(b[18]), .B(n4038), .Z(n4039) );
  XOR U5062 ( .A(n4040), .B(n4041), .Z(n4038) );
  ANDN U5063 ( .B(n4042), .A(n912), .Z(n4040) );
  XOR U5064 ( .A(b[17]), .B(n4041), .Z(n4042) );
  XOR U5065 ( .A(n4043), .B(n4044), .Z(n4041) );
  ANDN U5066 ( .B(n4045), .A(n923), .Z(n4043) );
  XOR U5067 ( .A(b[16]), .B(n4044), .Z(n4045) );
  XOR U5068 ( .A(n4046), .B(n4047), .Z(n4044) );
  ANDN U5069 ( .B(n4048), .A(n934), .Z(n4046) );
  XOR U5070 ( .A(b[15]), .B(n4047), .Z(n4048) );
  XOR U5071 ( .A(n4049), .B(n4050), .Z(n4047) );
  ANDN U5072 ( .B(n4051), .A(n945), .Z(n4049) );
  XOR U5073 ( .A(b[14]), .B(n4050), .Z(n4051) );
  XOR U5074 ( .A(n4052), .B(n4053), .Z(n4050) );
  ANDN U5075 ( .B(n4054), .A(n956), .Z(n4052) );
  XOR U5076 ( .A(b[13]), .B(n4053), .Z(n4054) );
  XOR U5077 ( .A(n4055), .B(n4056), .Z(n4053) );
  ANDN U5078 ( .B(n4057), .A(n967), .Z(n4055) );
  XOR U5079 ( .A(b[12]), .B(n4056), .Z(n4057) );
  XOR U5080 ( .A(n4058), .B(n4059), .Z(n4056) );
  ANDN U5081 ( .B(n4060), .A(n978), .Z(n4058) );
  XOR U5082 ( .A(b[11]), .B(n4059), .Z(n4060) );
  XOR U5083 ( .A(n4061), .B(n4062), .Z(n4059) );
  ANDN U5084 ( .B(n4063), .A(n989), .Z(n4061) );
  XOR U5085 ( .A(b[10]), .B(n4062), .Z(n4063) );
  XOR U5086 ( .A(n4064), .B(n4065), .Z(n4062) );
  ANDN U5087 ( .B(n4066), .A(n1), .Z(n4064) );
  XOR U5088 ( .A(b[9]), .B(n4065), .Z(n4066) );
  XOR U5089 ( .A(n4067), .B(n4068), .Z(n4065) );
  ANDN U5090 ( .B(n4069), .A(n112), .Z(n4067) );
  XOR U5091 ( .A(b[8]), .B(n4068), .Z(n4069) );
  XOR U5092 ( .A(n4070), .B(n4071), .Z(n4068) );
  ANDN U5093 ( .B(n4072), .A(n223), .Z(n4070) );
  XOR U5094 ( .A(b[7]), .B(n4071), .Z(n4072) );
  XOR U5095 ( .A(n4073), .B(n4074), .Z(n4071) );
  ANDN U5096 ( .B(n4075), .A(n334), .Z(n4073) );
  XOR U5097 ( .A(b[6]), .B(n4074), .Z(n4075) );
  XOR U5098 ( .A(n4076), .B(n4077), .Z(n4074) );
  ANDN U5099 ( .B(n4078), .A(n445), .Z(n4076) );
  XOR U5100 ( .A(b[5]), .B(n4077), .Z(n4078) );
  XOR U5101 ( .A(n4079), .B(n4080), .Z(n4077) );
  ANDN U5102 ( .B(n4081), .A(n556), .Z(n4079) );
  XOR U5103 ( .A(b[4]), .B(n4080), .Z(n4081) );
  XOR U5104 ( .A(n4082), .B(n4083), .Z(n4080) );
  ANDN U5105 ( .B(n4084), .A(n667), .Z(n4082) );
  XOR U5106 ( .A(b[3]), .B(n4083), .Z(n4084) );
  XOR U5107 ( .A(n4085), .B(n4086), .Z(n4083) );
  ANDN U5108 ( .B(n4087), .A(n778), .Z(n4085) );
  XOR U5109 ( .A(b[2]), .B(n4086), .Z(n4087) );
  XNOR U5110 ( .A(n4088), .B(n4089), .Z(n4086) );
  NANDN U5111 ( .A(n889), .B(n4090), .Z(n4089) );
  XOR U5112 ( .A(b[1]), .B(n4088), .Z(n4090) );
  XNOR U5113 ( .A(a[1]), .B(n4088), .Z(n889) );
  AND U5114 ( .A(b[0]), .B(a[0]), .Z(n4088) );
  XOR U5115 ( .A(b[0]), .B(a[0]), .Z(c[0]) );
endmodule

