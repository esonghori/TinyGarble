
module sha3_seq_CC3 ( clk, rst, in, out );
  input [575:0] in;
  output [1599:0] out;
  input clk, rst;
  wire   init, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
         n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
         n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
         n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
         n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
         n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
         n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
         n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
         n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
         n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
         n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
         n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
         n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
         n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966,
         n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974,
         n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982,
         n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990,
         n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
         n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006,
         n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014,
         n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
         n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
         n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038,
         n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046,
         n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054,
         n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062,
         n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
         n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078,
         n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
         n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
         n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
         n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110,
         n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118,
         n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
         n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134,
         n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
         n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150,
         n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158,
         n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
         n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
         n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182,
         n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
         n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198,
         n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
         n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
         n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
         n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
         n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238,
         n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
         n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254,
         n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262,
         n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270,
         n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278,
         n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286,
         n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294,
         n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302,
         n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310,
         n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318,
         n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326,
         n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334,
         n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
         n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350,
         n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358,
         n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
         n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
         n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382,
         n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390,
         n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398,
         n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406,
         n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
         n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422,
         n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430,
         n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438,
         n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446,
         n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454,
         n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462,
         n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
         n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
         n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486,
         n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494,
         n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502,
         n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510,
         n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518,
         n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526,
         n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534,
         n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542,
         n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550,
         n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558,
         n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566,
         n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
         n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582,
         n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590,
         n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598,
         n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606,
         n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614,
         n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622,
         n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630,
         n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638,
         n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646,
         n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654,
         n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662,
         n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670,
         n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678,
         n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686,
         n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694,
         n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702,
         n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710,
         n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718,
         n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726,
         n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734,
         n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742,
         n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750,
         n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758,
         n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766,
         n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774,
         n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782,
         n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790,
         n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798,
         n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806,
         n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814,
         n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822,
         n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830,
         n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838,
         n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846,
         n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854,
         n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862,
         n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870,
         n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878,
         n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886,
         n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894,
         n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902,
         n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910,
         n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918,
         n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926,
         n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934,
         n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942,
         n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950,
         n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958,
         n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966,
         n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974,
         n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982,
         n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990,
         n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998,
         n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006,
         n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014,
         n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022,
         n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030,
         n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038,
         n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046,
         n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054,
         n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062,
         n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070,
         n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078,
         n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086,
         n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094,
         n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102,
         n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110,
         n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118,
         n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126,
         n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134,
         n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142,
         n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150,
         n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158,
         n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166,
         n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174,
         n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182,
         n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190,
         n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198,
         n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206,
         n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214,
         n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222,
         n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230,
         n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238,
         n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246,
         n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254,
         n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262,
         n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270,
         n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278,
         n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286,
         n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294,
         n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302,
         n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310,
         n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318,
         n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
         n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334,
         n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342,
         n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350,
         n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358,
         n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366,
         n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374,
         n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
         n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
         n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
         n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406,
         n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
         n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
         n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430,
         n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
         n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
         n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
         n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
         n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
         n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
         n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
         n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
         n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502,
         n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
         n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
         n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
         n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
         n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
         n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
         n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
         n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
         n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598,
         n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
         n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
         n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622,
         n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630,
         n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638,
         n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646,
         n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
         n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
         n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670,
         n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
         n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
         n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
         n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
         n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
         n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
         n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
         n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
         n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
         n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
         n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
         n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
         n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854,
         n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862,
         n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870,
         n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
         n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886,
         n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
         n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902,
         n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910,
         n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918,
         n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926,
         n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934,
         n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942,
         n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
         n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,
         n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
         n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974,
         n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982,
         n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990,
         n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998,
         n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006,
         n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014,
         n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022,
         n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030,
         n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038,
         n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046,
         n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054,
         n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062,
         n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070,
         n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078,
         n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086,
         n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094,
         n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102,
         n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,
         n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118,
         n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126,
         n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134,
         n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142,
         n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150,
         n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158,
         n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,
         n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
         n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
         n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190,
         n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198,
         n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,
         n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214,
         n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222,
         n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230,
         n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238,
         n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246,
         n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254,
         n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262,
         n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270,
         n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278,
         n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286,
         n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294,
         n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302,
         n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310,
         n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318,
         n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326,
         n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334,
         n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342,
         n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350,
         n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358,
         n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366,
         n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374,
         n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382,
         n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390,
         n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398,
         n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406,
         n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414,
         n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422,
         n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430,
         n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438,
         n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446,
         n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454,
         n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462,
         n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470,
         n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478,
         n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486,
         n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494,
         n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502,
         n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510,
         n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518,
         n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526,
         n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534,
         n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542,
         n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550,
         n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558,
         n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566,
         n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574,
         n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582,
         n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590,
         n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598,
         n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606,
         n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614,
         n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622,
         n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630,
         n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638,
         n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646,
         n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654,
         n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662,
         n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670,
         n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678,
         n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686,
         n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694,
         n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702,
         n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710,
         n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718,
         n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726,
         n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734,
         n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742,
         n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750,
         n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758,
         n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766,
         n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774,
         n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782,
         n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790,
         n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798,
         n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806,
         n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814,
         n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822,
         n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830,
         n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838,
         n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846,
         n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854,
         n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862,
         n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870,
         n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878,
         n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886,
         n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894,
         n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902,
         n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910,
         n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918,
         n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926,
         n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934,
         n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942,
         n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950,
         n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958,
         n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966,
         n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974,
         n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982,
         n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990,
         n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998,
         n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006,
         n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014,
         n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022,
         n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030,
         n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038,
         n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046,
         n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054,
         n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062,
         n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070,
         n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078,
         n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086,
         n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094,
         n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102,
         n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110,
         n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118,
         n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126,
         n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134,
         n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142,
         n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150,
         n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158,
         n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166,
         n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174,
         n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182,
         n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190,
         n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198,
         n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206,
         n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214,
         n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222,
         n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230,
         n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238,
         n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246,
         n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254,
         n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262,
         n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270,
         n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278,
         n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286,
         n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294,
         n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302,
         n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310,
         n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318,
         n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326,
         n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334,
         n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342,
         n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350,
         n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358,
         n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366,
         n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374,
         n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382,
         n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390,
         n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398,
         n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406,
         n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414,
         n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422,
         n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430,
         n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438,
         n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446,
         n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454,
         n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462,
         n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470,
         n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478,
         n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486,
         n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494,
         n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502,
         n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510,
         n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518,
         n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526,
         n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534,
         n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542,
         n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550,
         n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558,
         n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566,
         n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574,
         n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582,
         n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590,
         n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598,
         n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606,
         n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614,
         n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622,
         n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630,
         n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638,
         n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646,
         n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654,
         n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662,
         n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670,
         n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678,
         n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686,
         n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694,
         n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702,
         n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710,
         n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718,
         n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726,
         n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734,
         n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742,
         n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750,
         n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758,
         n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766,
         n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774,
         n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782,
         n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790,
         n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798,
         n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806,
         n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814,
         n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822,
         n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830,
         n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838,
         n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846,
         n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854,
         n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862,
         n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870,
         n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878,
         n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886,
         n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894,
         n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902,
         n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910,
         n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918,
         n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926,
         n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934,
         n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942,
         n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950,
         n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958,
         n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966,
         n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974,
         n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982,
         n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990,
         n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998,
         n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006,
         n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014,
         n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022,
         n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030,
         n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038,
         n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046,
         n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054,
         n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062,
         n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070,
         n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078,
         n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086,
         n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094,
         n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102,
         n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110,
         n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118,
         n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126,
         n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134,
         n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142,
         n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150,
         n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158,
         n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166,
         n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174,
         n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182,
         n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190,
         n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198,
         n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206,
         n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214,
         n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222,
         n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230,
         n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238,
         n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246,
         n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254,
         n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262,
         n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270,
         n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278,
         n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286,
         n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294,
         n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302,
         n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310,
         n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318,
         n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326,
         n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334,
         n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342,
         n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350,
         n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358,
         n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366,
         n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374,
         n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382,
         n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390,
         n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398,
         n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406,
         n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414,
         n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422,
         n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430,
         n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438,
         n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446,
         n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454,
         n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462,
         n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470,
         n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478,
         n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486,
         n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494,
         n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502,
         n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510,
         n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518,
         n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526,
         n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534,
         n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542,
         n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550,
         n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558,
         n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566,
         n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574,
         n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582,
         n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590,
         n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598,
         n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606,
         n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614,
         n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622,
         n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630,
         n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638,
         n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646,
         n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654,
         n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662,
         n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670,
         n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678,
         n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686,
         n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694,
         n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702,
         n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710,
         n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718,
         n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726,
         n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734,
         n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742,
         n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750,
         n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758,
         n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766,
         n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774,
         n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782,
         n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790,
         n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798,
         n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806,
         n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814,
         n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822,
         n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830,
         n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838,
         n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846,
         n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854,
         n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862,
         n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870,
         n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878,
         n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886,
         n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894,
         n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902,
         n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910,
         n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918,
         n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926,
         n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934,
         n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942,
         n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950,
         n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958,
         n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966,
         n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974,
         n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982,
         n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990,
         n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998,
         n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006,
         n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014,
         n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022,
         n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030,
         n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038,
         n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046,
         n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054,
         n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062,
         n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070,
         n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078,
         n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086,
         n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094,
         n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102,
         n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110,
         n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118,
         n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126,
         n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134,
         n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142,
         n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150,
         n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158,
         n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166,
         n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174,
         n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182,
         n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190,
         n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198,
         n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206,
         n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214,
         n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222,
         n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230,
         n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238,
         n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246,
         n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254,
         n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262,
         n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270,
         n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278,
         n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286,
         n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294,
         n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302,
         n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310,
         n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318,
         n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326,
         n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334,
         n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342,
         n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350,
         n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358,
         n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366,
         n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374,
         n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382,
         n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390,
         n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398,
         n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406,
         n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414,
         n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422,
         n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430,
         n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438,
         n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446,
         n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454,
         n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462,
         n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470,
         n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478,
         n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486,
         n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494,
         n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502,
         n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510,
         n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518,
         n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526,
         n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534,
         n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542,
         n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550,
         n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558,
         n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566,
         n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574,
         n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582,
         n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590,
         n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598,
         n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606,
         n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614,
         n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622,
         n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630,
         n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638,
         n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646,
         n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654,
         n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662,
         n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670,
         n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678,
         n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686,
         n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694,
         n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702,
         n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710,
         n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718,
         n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726,
         n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734,
         n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742,
         n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750,
         n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758,
         n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766,
         n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774,
         n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782,
         n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790,
         n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798,
         n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806,
         n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814,
         n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822,
         n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830,
         n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838,
         n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846,
         n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854,
         n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862,
         n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870,
         n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878,
         n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886,
         n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894,
         n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902,
         n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910,
         n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918,
         n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926,
         n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934,
         n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942,
         n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950,
         n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958,
         n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966,
         n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974,
         n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982,
         n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990,
         n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998,
         n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006,
         n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014,
         n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022,
         n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030,
         n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038,
         n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046,
         n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054,
         n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062,
         n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070,
         n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078,
         n19079, n19080, n19081, n19082, n19083, n19084, n19085, n19086,
         n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094,
         n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102,
         n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110,
         n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118,
         n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126,
         n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134,
         n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142,
         n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150,
         n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158,
         n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166,
         n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174,
         n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182,
         n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190,
         n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198,
         n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206,
         n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214,
         n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222,
         n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19230,
         n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238,
         n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246,
         n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254,
         n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262,
         n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270,
         n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278,
         n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286,
         n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294,
         n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302,
         n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310,
         n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318,
         n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326,
         n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334,
         n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342,
         n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350,
         n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358,
         n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366,
         n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374,
         n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382,
         n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390,
         n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398,
         n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406,
         n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414,
         n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422,
         n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430,
         n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438,
         n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446,
         n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454,
         n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462,
         n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470,
         n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478,
         n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486,
         n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494,
         n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502,
         n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510,
         n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518,
         n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526,
         n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534,
         n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542,
         n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550,
         n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558,
         n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566,
         n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574,
         n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582,
         n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590,
         n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598,
         n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606,
         n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614,
         n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622,
         n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630,
         n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638,
         n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646,
         n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654,
         n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662,
         n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670,
         n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678,
         n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686,
         n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694,
         n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702,
         n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710,
         n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718,
         n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726,
         n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734,
         n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742,
         n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750,
         n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758,
         n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766,
         n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774,
         n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782,
         n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790,
         n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798,
         n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806,
         n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814,
         n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822,
         n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830,
         n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838,
         n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846,
         n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854,
         n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862,
         n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870,
         n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878,
         n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886,
         n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894,
         n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902,
         n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910,
         n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918,
         n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926,
         n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934,
         n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942,
         n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950,
         n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958,
         n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966,
         n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974,
         n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982,
         n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990,
         n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998,
         n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006,
         n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014,
         n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022,
         n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030,
         n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038,
         n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046,
         n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054,
         n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062,
         n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070,
         n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078,
         n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086,
         n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094,
         n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102,
         n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110,
         n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118,
         n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126,
         n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134,
         n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142,
         n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150,
         n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158,
         n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166,
         n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174,
         n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182,
         n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190,
         n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198,
         n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206,
         n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214,
         n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222,
         n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230,
         n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238,
         n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246,
         n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254,
         n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262,
         n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270,
         n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278,
         n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286,
         n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294,
         n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302,
         n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310,
         n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318,
         n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326,
         n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334,
         n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342,
         n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350,
         n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358,
         n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366,
         n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374,
         n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382,
         n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390,
         n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398,
         n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406,
         n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414,
         n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422,
         n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430,
         n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438,
         n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446,
         n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454,
         n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462,
         n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470,
         n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478,
         n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486,
         n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494,
         n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502,
         n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510,
         n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518,
         n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526,
         n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534,
         n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542,
         n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550,
         n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558,
         n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566,
         n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574,
         n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582,
         n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590,
         n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598,
         n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606,
         n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614,
         n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622,
         n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630,
         n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638,
         n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646,
         n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654,
         n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662,
         n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670,
         n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678,
         n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686,
         n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694,
         n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702,
         n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710,
         n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718,
         n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726,
         n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734,
         n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742,
         n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750,
         n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758,
         n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766,
         n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774,
         n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782,
         n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790,
         n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798,
         n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806,
         n20807, n20808, n20809, n20810, n20811, n20812, n20813, n20814,
         n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822,
         n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830,
         n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838,
         n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846,
         n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854,
         n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862,
         n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870,
         n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878,
         n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886,
         n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894,
         n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902,
         n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910,
         n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918,
         n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926,
         n20927, n20928, n20929, n20930, n20931, n20932, n20933, n20934,
         n20935, n20936, n20937, n20938, n20939, n20940, n20941, n20942,
         n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950,
         n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958,
         n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966,
         n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974,
         n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982,
         n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990,
         n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998,
         n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006,
         n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014,
         n21015, n21016, n21017, n21018, n21019, n21020, n21021, n21022,
         n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030,
         n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038,
         n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046,
         n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054,
         n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062,
         n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070,
         n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078,
         n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086,
         n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094,
         n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102,
         n21103, n21104, n21105, n21106, n21107, n21108, n21109, n21110,
         n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118,
         n21119, n21120, n21121, n21122, n21123, n21124, n21125, n21126,
         n21127, n21128, n21129, n21130, n21131, n21132, n21133, n21134,
         n21135, n21136, n21137, n21138, n21139, n21140, n21141, n21142,
         n21143, n21144, n21145, n21146, n21147, n21148, n21149, n21150,
         n21151, n21152, n21153, n21154, n21155, n21156, n21157, n21158,
         n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166,
         n21167, n21168, n21169, n21170, n21171, n21172, n21173, n21174,
         n21175, n21176, n21177, n21178, n21179, n21180, n21181, n21182,
         n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190,
         n21191, n21192, n21193, n21194, n21195, n21196, n21197, n21198,
         n21199, n21200, n21201, n21202, n21203, n21204, n21205, n21206,
         n21207, n21208, n21209, n21210, n21211, n21212, n21213, n21214,
         n21215, n21216, n21217, n21218, n21219, n21220, n21221, n21222,
         n21223, n21224, n21225, n21226, n21227, n21228, n21229, n21230,
         n21231, n21232, n21233, n21234, n21235, n21236, n21237, n21238,
         n21239, n21240, n21241, n21242, n21243, n21244, n21245, n21246,
         n21247, n21248, n21249, n21250, n21251, n21252, n21253, n21254,
         n21255, n21256, n21257, n21258, n21259, n21260, n21261, n21262,
         n21263, n21264, n21265, n21266, n21267, n21268, n21269, n21270,
         n21271, n21272, n21273, n21274, n21275, n21276, n21277, n21278,
         n21279, n21280, n21281, n21282, n21283, n21284, n21285, n21286,
         n21287, n21288, n21289, n21290, n21291, n21292, n21293, n21294,
         n21295, n21296, n21297, n21298, n21299, n21300, n21301, n21302,
         n21303, n21304, n21305, n21306, n21307, n21308, n21309, n21310,
         n21311, n21312, n21313, n21314, n21315, n21316, n21317, n21318,
         n21319, n21320, n21321, n21322, n21323, n21324, n21325, n21326,
         n21327, n21328, n21329, n21330, n21331, n21332, n21333, n21334,
         n21335, n21336, n21337, n21338, n21339, n21340, n21341, n21342,
         n21343, n21344, n21345, n21346, n21347, n21348, n21349, n21350,
         n21351, n21352, n21353, n21354, n21355, n21356, n21357, n21358,
         n21359, n21360, n21361, n21362, n21363, n21364, n21365, n21366,
         n21367, n21368, n21369, n21370, n21371, n21372, n21373, n21374,
         n21375, n21376, n21377, n21378, n21379, n21380, n21381, n21382,
         n21383, n21384, n21385, n21386, n21387, n21388, n21389, n21390,
         n21391, n21392, n21393, n21394, n21395, n21396, n21397, n21398,
         n21399, n21400, n21401, n21402, n21403, n21404, n21405, n21406,
         n21407, n21408, n21409, n21410, n21411, n21412, n21413, n21414,
         n21415, n21416, n21417, n21418, n21419, n21420, n21421, n21422,
         n21423, n21424, n21425, n21426, n21427, n21428, n21429, n21430,
         n21431, n21432, n21433, n21434, n21435, n21436, n21437, n21438,
         n21439, n21440, n21441, n21442, n21443, n21444, n21445, n21446,
         n21447, n21448, n21449, n21450, n21451, n21452, n21453, n21454,
         n21455, n21456, n21457, n21458, n21459, n21460, n21461, n21462,
         n21463, n21464, n21465, n21466, n21467, n21468, n21469, n21470,
         n21471, n21472, n21473, n21474, n21475, n21476, n21477, n21478,
         n21479, n21480, n21481, n21482, n21483, n21484, n21485, n21486,
         n21487, n21488, n21489, n21490, n21491, n21492, n21493, n21494,
         n21495, n21496, n21497, n21498, n21499, n21500, n21501, n21502,
         n21503, n21504, n21505, n21506, n21507, n21508, n21509, n21510,
         n21511, n21512, n21513, n21514, n21515, n21516, n21517, n21518,
         n21519, n21520, n21521, n21522, n21523, n21524, n21525, n21526,
         n21527, n21528, n21529, n21530, n21531, n21532, n21533, n21534,
         n21535, n21536, n21537, n21538, n21539, n21540, n21541, n21542,
         n21543, n21544, n21545, n21546, n21547, n21548, n21549, n21550,
         n21551, n21552, n21553, n21554, n21555, n21556, n21557, n21558,
         n21559, n21560, n21561, n21562, n21563, n21564, n21565, n21566,
         n21567, n21568, n21569, n21570, n21571, n21572, n21573, n21574,
         n21575, n21576, n21577, n21578, n21579, n21580, n21581, n21582,
         n21583, n21584, n21585, n21586, n21587, n21588, n21589, n21590,
         n21591, n21592, n21593, n21594, n21595, n21596, n21597, n21598,
         n21599, n21600, n21601, n21602, n21603, n21604, n21605, n21606,
         n21607, n21608, n21609, n21610, n21611, n21612, n21613, n21614,
         n21615, n21616, n21617, n21618, n21619, n21620, n21621, n21622,
         n21623, n21624, n21625, n21626, n21627, n21628, n21629, n21630,
         n21631, n21632, n21633, n21634, n21635, n21636, n21637, n21638,
         n21639, n21640, n21641, n21642, n21643, n21644, n21645, n21646,
         n21647, n21648, n21649, n21650, n21651, n21652, n21653, n21654,
         n21655, n21656, n21657, n21658, n21659, n21660, n21661, n21662,
         n21663, n21664, n21665, n21666, n21667, n21668, n21669, n21670,
         n21671, n21672, n21673, n21674, n21675, n21676, n21677, n21678,
         n21679, n21680, n21681, n21682, n21683, n21684, n21685, n21686,
         n21687, n21688, n21689, n21690, n21691, n21692, n21693, n21694,
         n21695, n21696, n21697, n21698, n21699, n21700, n21701, n21702,
         n21703, n21704, n21705, n21706, n21707, n21708, n21709, n21710,
         n21711, n21712, n21713, n21714, n21715, n21716, n21717, n21718,
         n21719, n21720, n21721, n21722, n21723, n21724, n21725, n21726,
         n21727, n21728, n21729, n21730, n21731, n21732, n21733, n21734,
         n21735, n21736, n21737, n21738, n21739, n21740, n21741, n21742,
         n21743, n21744, n21745, n21746, n21747, n21748, n21749, n21750,
         n21751, n21752, n21753, n21754, n21755, n21756, n21757, n21758,
         n21759, n21760, n21761, n21762, n21763, n21764, n21765, n21766,
         n21767, n21768, n21769, n21770, n21771, n21772, n21773, n21774,
         n21775, n21776, n21777, n21778, n21779, n21780, n21781, n21782,
         n21783, n21784, n21785, n21786, n21787, n21788, n21789, n21790,
         n21791, n21792, n21793, n21794, n21795, n21796, n21797, n21798,
         n21799, n21800, n21801, n21802, n21803, n21804, n21805, n21806,
         n21807, n21808, n21809, n21810, n21811, n21812, n21813, n21814,
         n21815, n21816, n21817, n21818, n21819, n21820, n21821, n21822,
         n21823, n21824, n21825, n21826, n21827, n21828, n21829, n21830,
         n21831, n21832, n21833, n21834, n21835, n21836, n21837, n21838,
         n21839, n21840, n21841, n21842, n21843, n21844, n21845, n21846,
         n21847, n21848, n21849, n21850, n21851, n21852, n21853, n21854,
         n21855, n21856, n21857, n21858, n21859, n21860, n21861, n21862,
         n21863, n21864, n21865, n21866, n21867, n21868, n21869, n21870,
         n21871, n21872, n21873, n21874, n21875, n21876, n21877, n21878,
         n21879, n21880, n21881, n21882, n21883, n21884, n21885, n21886,
         n21887, n21888, n21889, n21890, n21891, n21892, n21893, n21894,
         n21895, n21896, n21897, n21898, n21899, n21900, n21901, n21902,
         n21903, n21904, n21905, n21906, n21907, n21908, n21909, n21910,
         n21911, n21912, n21913, n21914, n21915, n21916, n21917, n21918,
         n21919, n21920, n21921, n21922, n21923, n21924, n21925, n21926,
         n21927, n21928, n21929, n21930, n21931, n21932, n21933, n21934,
         n21935, n21936, n21937, n21938, n21939, n21940, n21941, n21942,
         n21943, n21944, n21945, n21946, n21947, n21948, n21949, n21950,
         n21951, n21952, n21953, n21954, n21955, n21956, n21957, n21958,
         n21959, n21960, n21961, n21962, n21963, n21964, n21965, n21966,
         n21967, n21968, n21969, n21970, n21971, n21972, n21973, n21974,
         n21975, n21976, n21977, n21978, n21979, n21980, n21981, n21982,
         n21983, n21984, n21985, n21986, n21987, n21988, n21989, n21990,
         n21991, n21992, n21993, n21994, n21995, n21996, n21997, n21998,
         n21999, n22000, n22001, n22002, n22003, n22004, n22005, n22006,
         n22007, n22008, n22009, n22010, n22011, n22012, n22013, n22014,
         n22015, n22016, n22017, n22018, n22019, n22020, n22021, n22022,
         n22023, n22024, n22025, n22026, n22027, n22028, n22029, n22030,
         n22031, n22032, n22033, n22034, n22035, n22036, n22037, n22038,
         n22039, n22040, n22041, n22042, n22043, n22044, n22045, n22046,
         n22047, n22048, n22049, n22050, n22051, n22052, n22053, n22054,
         n22055, n22056, n22057, n22058, n22059, n22060, n22061, n22062,
         n22063, n22064, n22065, n22066, n22067, n22068, n22069, n22070,
         n22071, n22072, n22073, n22074, n22075, n22076, n22077, n22078,
         n22079, n22080, n22081, n22082, n22083, n22084, n22085, n22086,
         n22087, n22088, n22089, n22090, n22091, n22092, n22093, n22094,
         n22095, n22096, n22097, n22098, n22099, n22100, n22101, n22102,
         n22103, n22104, n22105, n22106, n22107, n22108, n22109, n22110,
         n22111, n22112, n22113, n22114, n22115, n22116, n22117, n22118,
         n22119, n22120, n22121, n22122, n22123, n22124, n22125, n22126,
         n22127, n22128, n22129, n22130, n22131, n22132, n22133, n22134,
         n22135, n22136, n22137, n22138, n22139, n22140, n22141, n22142,
         n22143, n22144, n22145, n22146, n22147, n22148, n22149, n22150,
         n22151, n22152, n22153, n22154, n22155, n22156, n22157, n22158,
         n22159, n22160, n22161, n22162, n22163, n22164, n22165, n22166,
         n22167, n22168, n22169, n22170, n22171, n22172, n22173, n22174,
         n22175, n22176, n22177, n22178, n22179, n22180, n22181, n22182,
         n22183, n22184, n22185, n22186, n22187, n22188, n22189, n22190,
         n22191, n22192, n22193, n22194, n22195, n22196, n22197, n22198,
         n22199, n22200, n22201, n22202, n22203, n22204, n22205, n22206,
         n22207, n22208, n22209, n22210, n22211, n22212, n22213, n22214,
         n22215, n22216, n22217, n22218, n22219, n22220, n22221, n22222,
         n22223, n22224, n22225, n22226, n22227, n22228, n22229, n22230,
         n22231, n22232, n22233, n22234, n22235, n22236, n22237, n22238,
         n22239, n22240, n22241, n22242, n22243, n22244, n22245, n22246,
         n22247, n22248, n22249, n22250, n22251, n22252, n22253, n22254,
         n22255, n22256, n22257, n22258, n22259, n22260, n22261, n22262,
         n22263, n22264, n22265, n22266, n22267, n22268, n22269, n22270,
         n22271, n22272, n22273, n22274, n22275, n22276, n22277, n22278,
         n22279, n22280, n22281, n22282, n22283, n22284, n22285, n22286,
         n22287, n22288, n22289, n22290, n22291, n22292, n22293, n22294,
         n22295, n22296, n22297, n22298, n22299, n22300, n22301, n22302,
         n22303, n22304, n22305, n22306, n22307, n22308, n22309, n22310,
         n22311, n22312, n22313, n22314, n22315, n22316, n22317, n22318,
         n22319, n22320, n22321, n22322, n22323, n22324, n22325, n22326,
         n22327, n22328, n22329, n22330, n22331, n22332, n22333, n22334,
         n22335, n22336, n22337, n22338, n22339, n22340, n22341, n22342,
         n22343, n22344, n22345, n22346, n22347, n22348, n22349, n22350,
         n22351, n22352, n22353, n22354, n22355, n22356, n22357, n22358,
         n22359, n22360, n22361, n22362, n22363, n22364, n22365, n22366,
         n22367, n22368, n22369, n22370, n22371, n22372, n22373, n22374,
         n22375, n22376, n22377, n22378, n22379, n22380, n22381, n22382,
         n22383, n22384, n22385, n22386, n22387, n22388, n22389, n22390,
         n22391, n22392, n22393, n22394, n22395, n22396, n22397, n22398,
         n22399, n22400, n22401, n22402, n22403, n22404, n22405, n22406,
         n22407, n22408, n22409, n22410, n22411, n22412, n22413, n22414,
         n22415, n22416, n22417, n22418, n22419, n22420, n22421, n22422,
         n22423, n22424, n22425, n22426, n22427, n22428, n22429, n22430,
         n22431, n22432, n22433, n22434, n22435, n22436, n22437, n22438,
         n22439, n22440, n22441, n22442, n22443, n22444, n22445, n22446,
         n22447, n22448, n22449, n22450, n22451, n22452, n22453, n22454,
         n22455, n22456, n22457, n22458, n22459, n22460, n22461, n22462,
         n22463, n22464, n22465, n22466, n22467, n22468, n22469, n22470,
         n22471, n22472, n22473, n22474, n22475, n22476, n22477, n22478,
         n22479, n22480, n22481, n22482, n22483, n22484, n22485, n22486,
         n22487, n22488, n22489, n22490, n22491, n22492, n22493, n22494,
         n22495, n22496, n22497, n22498, n22499, n22500, n22501, n22502,
         n22503, n22504, n22505, n22506, n22507, n22508, n22509, n22510,
         n22511, n22512, n22513, n22514, n22515, n22516, n22517, n22518,
         n22519, n22520, n22521, n22522, n22523, n22524, n22525, n22526,
         n22527, n22528, n22529, n22530, n22531, n22532, n22533, n22534,
         n22535, n22536, n22537, n22538, n22539, n22540, n22541, n22542,
         n22543, n22544, n22545, n22546, n22547, n22548, n22549, n22550,
         n22551, n22552, n22553, n22554, n22555, n22556, n22557, n22558,
         n22559, n22560, n22561, n22562, n22563, n22564, n22565, n22566,
         n22567, n22568, n22569, n22570, n22571, n22572, n22573, n22574,
         n22575, n22576, n22577, n22578, n22579, n22580, n22581, n22582,
         n22583, n22584, n22585, n22586, n22587, n22588, n22589, n22590,
         n22591, n22592, n22593, n22594, n22595, n22596, n22597, n22598,
         n22599, n22600, n22601, n22602, n22603, n22604, n22605, n22606,
         n22607, n22608, n22609, n22610, n22611, n22612, n22613, n22614,
         n22615, n22616, n22617, n22618, n22619, n22620, n22621, n22622,
         n22623, n22624, n22625, n22626, n22627, n22628, n22629, n22630,
         n22631, n22632, n22633, n22634, n22635, n22636, n22637, n22638,
         n22639, n22640, n22641, n22642, n22643, n22644, n22645, n22646,
         n22647, n22648, n22649, n22650, n22651, n22652, n22653, n22654,
         n22655, n22656, n22657, n22658, n22659, n22660, n22661, n22662,
         n22663, n22664, n22665, n22666, n22667, n22668, n22669, n22670,
         n22671, n22672, n22673, n22674, n22675, n22676, n22677, n22678,
         n22679, n22680, n22681, n22682, n22683, n22684, n22685, n22686,
         n22687, n22688, n22689, n22690, n22691, n22692, n22693, n22694,
         n22695, n22696, n22697, n22698, n22699, n22700, n22701, n22702,
         n22703, n22704, n22705, n22706, n22707, n22708, n22709, n22710,
         n22711, n22712, n22713, n22714, n22715, n22716, n22717, n22718,
         n22719, n22720, n22721, n22722, n22723, n22724, n22725, n22726,
         n22727, n22728, n22729, n22730, n22731, n22732, n22733, n22734,
         n22735, n22736, n22737, n22738, n22739, n22740, n22741, n22742,
         n22743, n22744, n22745, n22746, n22747, n22748, n22749, n22750,
         n22751, n22752, n22753, n22754, n22755, n22756, n22757, n22758,
         n22759, n22760, n22761, n22762, n22763, n22764, n22765, n22766,
         n22767, n22768, n22769, n22770, n22771, n22772, n22773, n22774,
         n22775, n22776, n22777, n22778, n22779, n22780, n22781, n22782,
         n22783, n22784, n22785, n22786, n22787, n22788, n22789, n22790,
         n22791, n22792, n22793, n22794, n22795, n22796, n22797, n22798,
         n22799, n22800, n22801, n22802, n22803, n22804, n22805, n22806,
         n22807, n22808, n22809, n22810, n22811, n22812, n22813, n22814,
         n22815, n22816, n22817, n22818, n22819, n22820, n22821, n22822,
         n22823, n22824, n22825, n22826, n22827, n22828, n22829, n22830,
         n22831, n22832, n22833, n22834, n22835, n22836, n22837, n22838,
         n22839, n22840, n22841, n22842, n22843, n22844, n22845, n22846,
         n22847, n22848, n22849, n22850, n22851, n22852, n22853, n22854,
         n22855, n22856, n22857, n22858, n22859, n22860, n22861, n22862,
         n22863, n22864, n22865, n22866, n22867, n22868, n22869, n22870,
         n22871, n22872, n22873, n22874, n22875, n22876, n22877, n22878,
         n22879, n22880, n22881, n22882, n22883, n22884, n22885, n22886,
         n22887, n22888, n22889, n22890, n22891, n22892, n22893, n22894,
         n22895, n22896, n22897, n22898, n22899, n22900, n22901, n22902,
         n22903, n22904, n22905, n22906, n22907, n22908, n22909, n22910,
         n22911, n22912, n22913, n22914, n22915, n22916, n22917, n22918,
         n22919, n22920, n22921, n22922, n22923, n22924, n22925, n22926,
         n22927, n22928, n22929, n22930, n22931, n22932, n22933, n22934,
         n22935, n22936, n22937, n22938, n22939, n22940, n22941, n22942,
         n22943, n22944, n22945, n22946, n22947, n22948, n22949, n22950,
         n22951, n22952, n22953, n22954, n22955, n22956, n22957, n22958,
         n22959, n22960, n22961, n22962, n22963, n22964, n22965, n22966,
         n22967, n22968, n22969, n22970, n22971, n22972, n22973, n22974,
         n22975, n22976, n22977, n22978, n22979, n22980, n22981, n22982,
         n22983, n22984, n22985, n22986, n22987, n22988, n22989, n22990,
         n22991, n22992, n22993, n22994, n22995, n22996, n22997, n22998,
         n22999, n23000, n23001, n23002, n23003, n23004, n23005, n23006,
         n23007, n23008, n23009, n23010, n23011, n23012, n23013, n23014,
         n23015, n23016, n23017, n23018, n23019, n23020, n23021, n23022,
         n23023, n23024, n23025, n23026, n23027, n23028, n23029, n23030,
         n23031, n23032, n23033, n23034, n23035, n23036, n23037, n23038,
         n23039, n23040, n23041, n23042, n23043, n23044, n23045, n23046,
         n23047, n23048, n23049, n23050, n23051, n23052, n23053, n23054,
         n23055, n23056, n23057, n23058, n23059, n23060, n23061, n23062,
         n23063, n23064, n23065, n23066, n23067, n23068, n23069, n23070,
         n23071, n23072, n23073, n23074, n23075, n23076, n23077, n23078,
         n23079, n23080, n23081, n23082, n23083, n23084, n23085, n23086,
         n23087, n23088, n23089, n23090, n23091, n23092, n23093, n23094,
         n23095, n23096, n23097, n23098, n23099, n23100, n23101, n23102,
         n23103, n23104, n23105, n23106, n23107, n23108, n23109, n23110,
         n23111, n23112, n23113, n23114, n23115, n23116, n23117, n23118,
         n23119, n23120, n23121, n23122, n23123, n23124, n23125, n23126,
         n23127, n23128, n23129, n23130, n23131, n23132, n23133, n23134,
         n23135, n23136, n23137, n23138, n23139, n23140, n23141, n23142,
         n23143, n23144, n23145, n23146, n23147, n23148, n23149, n23150,
         n23151, n23152, n23153, n23154, n23155, n23156, n23157, n23158,
         n23159, n23160, n23161, n23162, n23163, n23164, n23165, n23166,
         n23167, n23168, n23169, n23170, n23171, n23172, n23173, n23174,
         n23175, n23176, n23177, n23178, n23179, n23180, n23181, n23182,
         n23183, n23184, n23185, n23186, n23187, n23188, n23189, n23190,
         n23191, n23192, n23193, n23194, n23195, n23196, n23197, n23198,
         n23199, n23200, n23201, n23202, n23203, n23204, n23205, n23206,
         n23207, n23208, n23209, n23210, n23211, n23212, n23213, n23214,
         n23215, n23216, n23217, n23218, n23219, n23220, n23221, n23222,
         n23223, n23224, n23225, n23226, n23227, n23228, n23229, n23230,
         n23231, n23232, n23233, n23234, n23235, n23236, n23237, n23238,
         n23239, n23240, n23241, n23242, n23243, n23244, n23245, n23246,
         n23247, n23248, n23249, n23250, n23251, n23252, n23253, n23254,
         n23255, n23256, n23257, n23258, n23259, n23260, n23261, n23262,
         n23263, n23264, n23265, n23266, n23267, n23268, n23269, n23270,
         n23271, n23272, n23273, n23274, n23275, n23276, n23277, n23278,
         n23279, n23280, n23281, n23282, n23283, n23284, n23285, n23286,
         n23287, n23288, n23289, n23290, n23291, n23292, n23293, n23294,
         n23295, n23296, n23297, n23298, n23299, n23300, n23301, n23302,
         n23303, n23304, n23305, n23306, n23307, n23308, n23309, n23310,
         n23311, n23312, n23313, n23314, n23315, n23316, n23317, n23318,
         n23319, n23320, n23321, n23322, n23323, n23324, n23325, n23326,
         n23327, n23328, n23329, n23330, n23331, n23332, n23333, n23334,
         n23335, n23336, n23337, n23338, n23339, n23340, n23341, n23342,
         n23343, n23344, n23345, n23346, n23347, n23348, n23349, n23350,
         n23351, n23352, n23353, n23354, n23355, n23356, n23357, n23358,
         n23359, n23360, n23361, n23362, n23363, n23364, n23365, n23366,
         n23367, n23368, n23369, n23370, n23371, n23372, n23373, n23374,
         n23375, n23376, n23377, n23378, n23379, n23380, n23381, n23382,
         n23383, n23384, n23385, n23386, n23387, n23388, n23389, n23390,
         n23391, n23392, n23393, n23394, n23395, n23396, n23397, n23398,
         n23399, n23400, n23401, n23402, n23403, n23404, n23405, n23406,
         n23407, n23408, n23409, n23410, n23411, n23412, n23413, n23414,
         n23415, n23416, n23417, n23418, n23419, n23420, n23421, n23422,
         n23423, n23424, n23425, n23426, n23427, n23428, n23429, n23430,
         n23431, n23432, n23433, n23434, n23435, n23436, n23437, n23438,
         n23439, n23440, n23441, n23442, n23443, n23444, n23445, n23446,
         n23447, n23448, n23449, n23450, n23451, n23452, n23453, n23454,
         n23455, n23456, n23457, n23458, n23459, n23460, n23461, n23462,
         n23463, n23464, n23465, n23466, n23467, n23468, n23469, n23470,
         n23471, n23472, n23473, n23474, n23475, n23476, n23477, n23478,
         n23479, n23480, n23481, n23482, n23483, n23484, n23485, n23486,
         n23487, n23488, n23489, n23490, n23491, n23492, n23493, n23494,
         n23495, n23496, n23497, n23498, n23499, n23500, n23501, n23502,
         n23503, n23504, n23505, n23506, n23507, n23508, n23509, n23510,
         n23511, n23512, n23513, n23514, n23515, n23516, n23517, n23518,
         n23519, n23520, n23521, n23522, n23523, n23524, n23525, n23526,
         n23527, n23528, n23529, n23530, n23531, n23532, n23533, n23534,
         n23535, n23536, n23537, n23538, n23539, n23540, n23541, n23542,
         n23543, n23544, n23545, n23546, n23547, n23548, n23549, n23550,
         n23551, n23552, n23553, n23554, n23555, n23556, n23557, n23558,
         n23559, n23560, n23561, n23562, n23563, n23564, n23565, n23566,
         n23567, n23568, n23569, n23570, n23571, n23572, n23573, n23574,
         n23575, n23576, n23577, n23578, n23579, n23580, n23581, n23582,
         n23583, n23584, n23585, n23586, n23587, n23588, n23589, n23590,
         n23591, n23592, n23593, n23594, n23595, n23596, n23597, n23598,
         n23599, n23600, n23601, n23602, n23603, n23604, n23605, n23606,
         n23607, n23608, n23609, n23610, n23611, n23612, n23613, n23614,
         n23615, n23616, n23617, n23618, n23619, n23620, n23621, n23622,
         n23623, n23624, n23625, n23626, n23627, n23628, n23629, n23630,
         n23631, n23632, n23633, n23634, n23635, n23636, n23637, n23638,
         n23639, n23640, n23641, n23642, n23643, n23644, n23645, n23646,
         n23647, n23648, n23649, n23650, n23651, n23652, n23653, n23654,
         n23655, n23656, n23657, n23658, n23659, n23660, n23661, n23662,
         n23663, n23664, n23665, n23666, n23667, n23668, n23669, n23670,
         n23671, n23672, n23673, n23674, n23675, n23676, n23677, n23678,
         n23679, n23680, n23681, n23682, n23683, n23684, n23685, n23686,
         n23687, n23688, n23689, n23690, n23691, n23692, n23693, n23694,
         n23695, n23696, n23697, n23698, n23699, n23700, n23701, n23702,
         n23703, n23704, n23705, n23706, n23707, n23708, n23709, n23710,
         n23711, n23712, n23713, n23714, n23715, n23716, n23717, n23718,
         n23719, n23720, n23721, n23722, n23723, n23724, n23725, n23726,
         n23727, n23728, n23729, n23730, n23731, n23732, n23733, n23734,
         n23735, n23736, n23737, n23738, n23739, n23740, n23741, n23742,
         n23743, n23744, n23745, n23746, n23747, n23748, n23749, n23750,
         n23751, n23752, n23753, n23754, n23755, n23756, n23757, n23758,
         n23759, n23760, n23761, n23762, n23763, n23764, n23765, n23766,
         n23767, n23768, n23769, n23770, n23771, n23772, n23773, n23774,
         n23775, n23776, n23777, n23778, n23779, n23780, n23781, n23782,
         n23783, n23784, n23785, n23786, n23787, n23788, n23789, n23790,
         n23791, n23792, n23793, n23794, n23795, n23796, n23797, n23798,
         n23799, n23800, n23801, n23802, n23803, n23804, n23805, n23806,
         n23807, n23808, n23809, n23810, n23811, n23812, n23813, n23814,
         n23815, n23816, n23817, n23818, n23819, n23820, n23821, n23822,
         n23823, n23824, n23825, n23826, n23827, n23828, n23829, n23830,
         n23831, n23832, n23833, n23834, n23835, n23836, n23837, n23838,
         n23839, n23840, n23841, n23842, n23843, n23844, n23845, n23846,
         n23847, n23848, n23849, n23850, n23851, n23852, n23853, n23854,
         n23855, n23856, n23857, n23858, n23859, n23860, n23861, n23862,
         n23863, n23864, n23865, n23866, n23867, n23868, n23869, n23870,
         n23871, n23872, n23873, n23874, n23875, n23876, n23877, n23878,
         n23879, n23880, n23881, n23882, n23883, n23884, n23885, n23886,
         n23887, n23888, n23889, n23890, n23891, n23892, n23893, n23894,
         n23895, n23896, n23897, n23898, n23899, n23900, n23901, n23902,
         n23903, n23904, n23905, n23906, n23907, n23908, n23909, n23910,
         n23911, n23912, n23913, n23914, n23915, n23916, n23917, n23918,
         n23919, n23920, n23921, n23922, n23923, n23924, n23925, n23926,
         n23927, n23928, n23929, n23930, n23931, n23932, n23933, n23934,
         n23935, n23936, n23937, n23938, n23939, n23940, n23941, n23942,
         n23943, n23944, n23945, n23946, n23947, n23948, n23949, n23950,
         n23951, n23952, n23953, n23954, n23955, n23956, n23957, n23958,
         n23959, n23960, n23961, n23962, n23963, n23964, n23965, n23966,
         n23967, n23968, n23969, n23970, n23971, n23972, n23973, n23974,
         n23975, n23976, n23977, n23978, n23979, n23980, n23981, n23982,
         n23983, n23984, n23985, n23986, n23987, n23988, n23989, n23990,
         n23991, n23992, n23993, n23994, n23995, n23996, n23997, n23998,
         n23999, n24000, n24001, n24002, n24003, n24004, n24005, n24006,
         n24007, n24008, n24009, n24010, n24011, n24012, n24013, n24014,
         n24015, n24016, n24017, n24018, n24019, n24020, n24021, n24022,
         n24023, n24024, n24025, n24026, n24027, n24028, n24029, n24030,
         n24031, n24032, n24033, n24034, n24035, n24036, n24037, n24038,
         n24039, n24040, n24041, n24042, n24043, n24044, n24045, n24046,
         n24047, n24048, n24049, n24050, n24051, n24052, n24053, n24054,
         n24055, n24056, n24057, n24058, n24059, n24060, n24061, n24062,
         n24063, n24064, n24065, n24066, n24067, n24068, n24069, n24070,
         n24071, n24072, n24073, n24074, n24075, n24076, n24077, n24078,
         n24079, n24080, n24081, n24082, n24083, n24084, n24085, n24086,
         n24087, n24088, n24089, n24090, n24091, n24092, n24093, n24094,
         n24095, n24096, n24097, n24098, n24099, n24100, n24101, n24102,
         n24103, n24104, n24105, n24106, n24107, n24108, n24109, n24110,
         n24111, n24112, n24113, n24114, n24115, n24116, n24117, n24118,
         n24119, n24120, n24121, n24122, n24123, n24124, n24125, n24126,
         n24127, n24128, n24129, n24130, n24131, n24132, n24133, n24134,
         n24135, n24136, n24137, n24138, n24139, n24140, n24141, n24142,
         n24143, n24144, n24145, n24146, n24147, n24148, n24149, n24150,
         n24151, n24152, n24153, n24154, n24155, n24156, n24157, n24158,
         n24159, n24160, n24161, n24162, n24163, n24164, n24165, n24166,
         n24167, n24168, n24169, n24170, n24171, n24172, n24173, n24174,
         n24175, n24176, n24177, n24178, n24179, n24180, n24181, n24182,
         n24183, n24184, n24185, n24186, n24187, n24188, n24189, n24190,
         n24191, n24192, n24193, n24194, n24195, n24196, n24197, n24198,
         n24199, n24200, n24201, n24202, n24203, n24204, n24205, n24206,
         n24207, n24208, n24209, n24210, n24211, n24212, n24213, n24214,
         n24215, n24216, n24217, n24218, n24219, n24220, n24221, n24222,
         n24223, n24224, n24225, n24226, n24227, n24228, n24229, n24230,
         n24231, n24232, n24233, n24234, n24235, n24236, n24237, n24238,
         n24239, n24240, n24241, n24242, n24243, n24244, n24245, n24246,
         n24247, n24248, n24249, n24250, n24251, n24252, n24253, n24254,
         n24255, n24256, n24257, n24258, n24259, n24260, n24261, n24262,
         n24263, n24264, n24265, n24266, n24267, n24268, n24269, n24270,
         n24271, n24272, n24273, n24274, n24275, n24276, n24277, n24278,
         n24279, n24280, n24281, n24282, n24283, n24284, n24285, n24286,
         n24287, n24288, n24289, n24290, n24291, n24292, n24293, n24294,
         n24295, n24296, n24297, n24298, n24299, n24300, n24301, n24302,
         n24303, n24304, n24305, n24306, n24307, n24308, n24309, n24310,
         n24311, n24312, n24313, n24314, n24315, n24316, n24317, n24318,
         n24319, n24320, n24321, n24322, n24323, n24324, n24325, n24326,
         n24327, n24328, n24329, n24330, n24331, n24332, n24333, n24334,
         n24335, n24336, n24337, n24338, n24339, n24340, n24341, n24342,
         n24343, n24344, n24345, n24346, n24347, n24348, n24349, n24350,
         n24351, n24352, n24353, n24354, n24355, n24356, n24357, n24358,
         n24359, n24360, n24361, n24362, n24363, n24364, n24365, n24366,
         n24367, n24368, n24369, n24370, n24371, n24372, n24373, n24374,
         n24375, n24376, n24377, n24378, n24379, n24380, n24381, n24382,
         n24383, n24384, n24385, n24386, n24387, n24388, n24389, n24390,
         n24391, n24392, n24393, n24394, n24395, n24396, n24397, n24398,
         n24399, n24400, n24401, n24402, n24403, n24404, n24405, n24406,
         n24407, n24408, n24409, n24410, n24411, n24412, n24413, n24414,
         n24415, n24416, n24417, n24418, n24419, n24420, n24421, n24422,
         n24423, n24424, n24425, n24426, n24427, n24428, n24429, n24430,
         n24431, n24432, n24433, n24434, n24435, n24436, n24437, n24438,
         n24439, n24440, n24441, n24442, n24443, n24444, n24445, n24446,
         n24447, n24448, n24449, n24450, n24451, n24452, n24453, n24454,
         n24455, n24456, n24457, n24458, n24459, n24460, n24461, n24462,
         n24463, n24464, n24465, n24466, n24467, n24468, n24469, n24470,
         n24471, n24472, n24473, n24474, n24475, n24476, n24477, n24478,
         n24479, n24480, n24481, n24482, n24483, n24484, n24485, n24486,
         n24487, n24488, n24489, n24490, n24491, n24492, n24493, n24494,
         n24495, n24496, n24497, n24498, n24499, n24500, n24501, n24502,
         n24503, n24504, n24505, n24506, n24507, n24508, n24509, n24510,
         n24511, n24512, n24513, n24514, n24515, n24516, n24517, n24518,
         n24519, n24520, n24521, n24522, n24523, n24524, n24525, n24526,
         n24527, n24528, n24529, n24530, n24531, n24532, n24533, n24534,
         n24535, n24536, n24537, n24538, n24539, n24540, n24541, n24542,
         n24543, n24544, n24545, n24546, n24547, n24548, n24549, n24550,
         n24551, n24552, n24553, n24554, n24555, n24556, n24557, n24558,
         n24559, n24560, n24561, n24562, n24563, n24564, n24565, n24566,
         n24567, n24568, n24569, n24570, n24571, n24572, n24573, n24574,
         n24575, n24576, n24577, n24578, n24579, n24580, n24581, n24582,
         n24583, n24584, n24585, n24586, n24587, n24588, n24589, n24590,
         n24591, n24592, n24593, n24594, n24595, n24596, n24597, n24598,
         n24599, n24600, n24601, n24602, n24603, n24604, n24605, n24606,
         n24607, n24608, n24609, n24610, n24611, n24612, n24613, n24614,
         n24615, n24616, n24617, n24618, n24619, n24620, n24621, n24622,
         n24623, n24624, n24625, n24626, n24627, n24628, n24629, n24630,
         n24631, n24632, n24633, n24634, n24635, n24636, n24637, n24638,
         n24639, n24640, n24641, n24642, n24643, n24644, n24645, n24646,
         n24647, n24648, n24649, n24650, n24651, n24652, n24653, n24654,
         n24655, n24656, n24657, n24658, n24659, n24660, n24661, n24662,
         n24663, n24664, n24665, n24666, n24667, n24668, n24669, n24670,
         n24671, n24672, n24673, n24674, n24675, n24676, n24677, n24678,
         n24679, n24680, n24681, n24682, n24683, n24684, n24685, n24686,
         n24687, n24688, n24689, n24690, n24691, n24692, n24693, n24694,
         n24695, n24696, n24697, n24698, n24699, n24700, n24701, n24702,
         n24703, n24704, n24705, n24706, n24707, n24708, n24709, n24710,
         n24711, n24712, n24713, n24714, n24715, n24716, n24717, n24718,
         n24719, n24720, n24721, n24722, n24723, n24724, n24725, n24726,
         n24727, n24728, n24729, n24730, n24731, n24732, n24733, n24734,
         n24735, n24736, n24737, n24738, n24739, n24740, n24741, n24742,
         n24743, n24744, n24745, n24746, n24747, n24748, n24749, n24750,
         n24751, n24752, n24753, n24754, n24755, n24756, n24757, n24758,
         n24759, n24760, n24761, n24762, n24763, n24764, n24765, n24766,
         n24767, n24768, n24769, n24770, n24771, n24772, n24773, n24774,
         n24775, n24776, n24777, n24778, n24779, n24780, n24781, n24782,
         n24783, n24784, n24785, n24786, n24787, n24788, n24789, n24790,
         n24791, n24792, n24793, n24794, n24795, n24796, n24797, n24798,
         n24799, n24800, n24801, n24802, n24803, n24804, n24805, n24806,
         n24807, n24808, n24809, n24810, n24811, n24812, n24813, n24814,
         n24815, n24816, n24817, n24818, n24819, n24820, n24821, n24822,
         n24823, n24824, n24825, n24826, n24827, n24828, n24829, n24830,
         n24831, n24832, n24833, n24834, n24835, n24836, n24837, n24838,
         n24839, n24840, n24841, n24842, n24843, n24844, n24845, n24846,
         n24847, n24848, n24849, n24850, n24851, n24852, n24853, n24854,
         n24855, n24856, n24857, n24858, n24859, n24860, n24861, n24862,
         n24863, n24864, n24865, n24866, n24867, n24868, n24869, n24870,
         n24871, n24872, n24873, n24874, n24875, n24876, n24877, n24878,
         n24879, n24880, n24881, n24882, n24883, n24884, n24885, n24886,
         n24887, n24888, n24889, n24890, n24891, n24892, n24893, n24894,
         n24895, n24896, n24897, n24898, n24899, n24900, n24901, n24902,
         n24903, n24904, n24905, n24906, n24907, n24908, n24909, n24910,
         n24911, n24912, n24913, n24914, n24915, n24916, n24917, n24918,
         n24919, n24920, n24921, n24922, n24923, n24924, n24925, n24926,
         n24927, n24928, n24929, n24930, n24931, n24932, n24933, n24934,
         n24935, n24936, n24937, n24938, n24939, n24940, n24941, n24942,
         n24943, n24944, n24945, n24946, n24947, n24948, n24949, n24950,
         n24951, n24952, n24953, n24954, n24955, n24956, n24957, n24958,
         n24959, n24960, n24961, n24962, n24963, n24964, n24965, n24966,
         n24967, n24968, n24969, n24970, n24971, n24972, n24973, n24974,
         n24975, n24976, n24977, n24978, n24979, n24980, n24981, n24982,
         n24983, n24984, n24985, n24986, n24987, n24988, n24989, n24990,
         n24991, n24992, n24993, n24994, n24995, n24996, n24997, n24998,
         n24999, n25000, n25001, n25002, n25003, n25004, n25005, n25006,
         n25007, n25008, n25009, n25010, n25011, n25012, n25013, n25014,
         n25015, n25016, n25017, n25018, n25019, n25020, n25021, n25022,
         n25023, n25024, n25025, n25026, n25027, n25028, n25029, n25030,
         n25031, n25032, n25033, n25034, n25035, n25036, n25037, n25038,
         n25039, n25040, n25041, n25042, n25043, n25044, n25045, n25046,
         n25047, n25048, n25049, n25050, n25051, n25052, n25053, n25054,
         n25055, n25056, n25057, n25058, n25059, n25060, n25061, n25062,
         n25063, n25064, n25065, n25066, n25067, n25068, n25069, n25070,
         n25071, n25072, n25073, n25074, n25075, n25076, n25077, n25078,
         n25079, n25080, n25081, n25082, n25083, n25084, n25085, n25086,
         n25087, n25088, n25089, n25090, n25091, n25092, n25093, n25094,
         n25095, n25096, n25097, n25098, n25099, n25100, n25101, n25102,
         n25103, n25104, n25105, n25106, n25107, n25108, n25109, n25110,
         n25111, n25112, n25113, n25114, n25115, n25116, n25117, n25118,
         n25119, n25120, n25121, n25122, n25123, n25124, n25125, n25126,
         n25127, n25128, n25129, n25130, n25131, n25132, n25133, n25134,
         n25135, n25136, n25137, n25138, n25139, n25140, n25141, n25142,
         n25143, n25144, n25145, n25146, n25147, n25148, n25149, n25150,
         n25151, n25152, n25153, n25154, n25155, n25156, n25157, n25158,
         n25159, n25160, n25161, n25162, n25163, n25164, n25165, n25166,
         n25167, n25168, n25169, n25170, n25171, n25172, n25173, n25174,
         n25175, n25176, n25177, n25178, n25179, n25180, n25181, n25182,
         n25183, n25184, n25185, n25186, n25187, n25188, n25189, n25190,
         n25191, n25192, n25193, n25194, n25195, n25196, n25197, n25198,
         n25199, n25200, n25201, n25202, n25203, n25204, n25205, n25206,
         n25207, n25208, n25209, n25210, n25211, n25212, n25213, n25214,
         n25215, n25216, n25217, n25218, n25219, n25220, n25221, n25222,
         n25223, n25224, n25225, n25226, n25227, n25228, n25229, n25230,
         n25231, n25232, n25233, n25234, n25235, n25236, n25237, n25238,
         n25239, n25240, n25241, n25242, n25243, n25244, n25245, n25246,
         n25247, n25248, n25249, n25250, n25251, n25252, n25253, n25254,
         n25255, n25256, n25257, n25258, n25259, n25260, n25261, n25262,
         n25263, n25264, n25265, n25266, n25267, n25268, n25269, n25270,
         n25271, n25272, n25273, n25274, n25275, n25276, n25277, n25278,
         n25279, n25280, n25281, n25282, n25283, n25284, n25285, n25286,
         n25287, n25288, n25289, n25290, n25291, n25292, n25293, n25294,
         n25295, n25296, n25297, n25298, n25299, n25300, n25301, n25302,
         n25303, n25304, n25305, n25306, n25307, n25308, n25309, n25310,
         n25311, n25312, n25313, n25314, n25315, n25316, n25317, n25318,
         n25319, n25320, n25321, n25322, n25323, n25324, n25325, n25326,
         n25327, n25328, n25329, n25330, n25331, n25332, n25333, n25334,
         n25335, n25336, n25337, n25338, n25339, n25340, n25341, n25342,
         n25343, n25344, n25345, n25346, n25347, n25348, n25349, n25350,
         n25351, n25352, n25353, n25354, n25355, n25356, n25357, n25358,
         n25359, n25360, n25361, n25362, n25363, n25364, n25365, n25366,
         n25367, n25368, n25369, n25370, n25371, n25372, n25373, n25374,
         n25375, n25376, n25377, n25378, n25379, n25380, n25381, n25382,
         n25383, n25384, n25385, n25386, n25387, n25388, n25389, n25390,
         n25391, n25392, n25393, n25394, n25395, n25396, n25397, n25398,
         n25399, n25400, n25401, n25402, n25403, n25404, n25405, n25406,
         n25407, n25408, n25409, n25410, n25411, n25412, n25413, n25414,
         n25415, n25416, n25417, n25418, n25419, n25420, n25421, n25422,
         n25423, n25424, n25425, n25426, n25427, n25428, n25429, n25430,
         n25431, n25432, n25433, n25434, n25435, n25436, n25437, n25438,
         n25439, n25440, n25441, n25442, n25443, n25444, n25445, n25446,
         n25447, n25448, n25449, n25450, n25451, n25452, n25453, n25454,
         n25455, n25456, n25457, n25458, n25459, n25460, n25461, n25462,
         n25463, n25464, n25465, n25466, n25467, n25468, n25469, n25470,
         n25471, n25472, n25473, n25474, n25475, n25476, n25477, n25478,
         n25479, n25480, n25481, n25482, n25483, n25484, n25485, n25486,
         n25487, n25488, n25489, n25490, n25491, n25492, n25493, n25494,
         n25495, n25496, n25497, n25498, n25499, n25500, n25501, n25502,
         n25503, n25504, n25505, n25506, n25507, n25508, n25509, n25510,
         n25511, n25512, n25513, n25514, n25515, n25516, n25517, n25518,
         n25519, n25520, n25521, n25522, n25523, n25524, n25525, n25526,
         n25527, n25528, n25529, n25530, n25531, n25532, n25533, n25534,
         n25535, n25536, n25537, n25538, n25539, n25540, n25541, n25542,
         n25543, n25544, n25545, n25546, n25547, n25548, n25549, n25550,
         n25551, n25552, n25553, n25554, n25555, n25556, n25557, n25558,
         n25559, n25560, n25561, n25562, n25563, n25564, n25565, n25566,
         n25567, n25568, n25569, n25570, n25571, n25572, n25573, n25574,
         n25575, n25576, n25577, n25578, n25579, n25580, n25581, n25582,
         n25583, n25584, n25585, n25586, n25587, n25588, n25589, n25590,
         n25591, n25592, n25593, n25594, n25595, n25596, n25597, n25598,
         n25599, n25600, n25601, n25602, n25603, n25604, n25605, n25606,
         n25607, n25608, n25609, n25610, n25611, n25612, n25613, n25614,
         n25615, n25616, n25617, n25618, n25619, n25620, n25621, n25622,
         n25623, n25624, n25625, n25626, n25627, n25628, n25629, n25630,
         n25631, n25632, n25633, n25634, n25635, n25636, n25637, n25638,
         n25639, n25640, n25641, n25642, n25643, n25644, n25645, n25646,
         n25647, n25648, n25649, n25650, n25651, n25652, n25653, n25654,
         n25655, n25656, n25657, n25658, n25659, n25660, n25661, n25662,
         n25663, n25664, n25665, n25666, n25667, n25668, n25669, n25670,
         n25671, n25672, n25673, n25674, n25675, n25676, n25677, n25678,
         n25679, n25680, n25681, n25682, n25683, n25684, n25685, n25686,
         n25687, n25688, n25689, n25690, n25691, n25692, n25693, n25694,
         n25695, n25696, n25697, n25698, n25699, n25700, n25701, n25702,
         n25703, n25704, n25705, n25706, n25707, n25708, n25709, n25710,
         n25711, n25712, n25713, n25714, n25715, n25716, n25717, n25718,
         n25719, n25720, n25721, n25722, n25723, n25724, n25725, n25726,
         n25727, n25728, n25729, n25730, n25731, n25732, n25733, n25734,
         n25735, n25736, n25737, n25738, n25739, n25740, n25741, n25742,
         n25743, n25744, n25745, n25746, n25747, n25748, n25749, n25750,
         n25751, n25752, n25753, n25754, n25755, n25756, n25757, n25758,
         n25759, n25760, n25761, n25762, n25763, n25764, n25765, n25766,
         n25767, n25768, n25769, n25770, n25771, n25772, n25773, n25774,
         n25775, n25776, n25777, n25778, n25779, n25780, n25781, n25782,
         n25783, n25784, n25785, n25786, n25787, n25788, n25789, n25790,
         n25791, n25792, n25793, n25794, n25795, n25796, n25797, n25798,
         n25799, n25800, n25801, n25802, n25803, n25804, n25805, n25806,
         n25807, n25808, n25809, n25810, n25811, n25812, n25813, n25814,
         n25815, n25816, n25817, n25818, n25819, n25820, n25821, n25822,
         n25823, n25824, n25825, n25826, n25827, n25828, n25829, n25830,
         n25831, n25832, n25833, n25834, n25835, n25836, n25837, n25838,
         n25839, n25840, n25841, n25842, n25843, n25844, n25845, n25846,
         n25847, n25848, n25849, n25850, n25851, n25852, n25853, n25854,
         n25855, n25856, n25857, n25858, n25859, n25860, n25861, n25862,
         n25863, n25864, n25865, n25866, n25867, n25868, n25869, n25870,
         n25871, n25872, n25873, n25874, n25875, n25876, n25877, n25878,
         n25879, n25880, n25881, n25882, n25883, n25884, n25885, n25886,
         n25887, n25888, n25889, n25890, n25891, n25892, n25893, n25894,
         n25895, n25896, n25897, n25898, n25899, n25900, n25901, n25902,
         n25903, n25904, n25905, n25906, n25907, n25908, n25909, n25910,
         n25911, n25912, n25913, n25914, n25915, n25916, n25917, n25918,
         n25919, n25920, n25921, n25922, n25923, n25924, n25925, n25926,
         n25927, n25928, n25929, n25930, n25931, n25932, n25933, n25934,
         n25935, n25936, n25937, n25938, n25939, n25940, n25941, n25942,
         n25943, n25944, n25945, n25946, n25947, n25948, n25949, n25950,
         n25951, n25952, n25953, n25954, n25955, n25956, n25957, n25958,
         n25959, n25960, n25961, n25962, n25963, n25964, n25965, n25966,
         n25967, n25968, n25969, n25970, n25971, n25972, n25973, n25974,
         n25975, n25976, n25977, n25978, n25979, n25980, n25981, n25982,
         n25983, n25984, n25985, n25986, n25987, n25988, n25989, n25990,
         n25991, n25992, n25993, n25994, n25995, n25996, n25997, n25998,
         n25999, n26000, n26001, n26002, n26003, n26004, n26005, n26006,
         n26007, n26008, n26009, n26010, n26011, n26012, n26013, n26014,
         n26015, n26016, n26017, n26018, n26019, n26020, n26021, n26022,
         n26023, n26024, n26025, n26026, n26027, n26028, n26029, n26030,
         n26031, n26032, n26033, n26034, n26035, n26036, n26037, n26038,
         n26039, n26040, n26041, n26042, n26043, n26044, n26045, n26046,
         n26047, n26048, n26049, n26050, n26051, n26052, n26053, n26054,
         n26055, n26056, n26057, n26058, n26059, n26060, n26061, n26062,
         n26063, n26064, n26065, n26066, n26067, n26068, n26069, n26070,
         n26071, n26072, n26073, n26074, n26075, n26076, n26077, n26078,
         n26079, n26080, n26081, n26082, n26083, n26084, n26085, n26086,
         n26087, n26088, n26089, n26090, n26091, n26092, n26093, n26094,
         n26095, n26096, n26097, n26098, n26099, n26100, n26101, n26102,
         n26103, n26104, n26105, n26106, n26107, n26108, n26109, n26110,
         n26111, n26112, n26113, n26114, n26115, n26116, n26117, n26118,
         n26119, n26120, n26121, n26122, n26123, n26124, n26125, n26126,
         n26127, n26128, n26129, n26130, n26131, n26132, n26133, n26134,
         n26135, n26136, n26137, n26138, n26139, n26140, n26141, n26142,
         n26143, n26144, n26145, n26146, n26147, n26148, n26149, n26150,
         n26151, n26152, n26153, n26154, n26155, n26156, n26157, n26158,
         n26159, n26160, n26161, n26162, n26163, n26164, n26165, n26166,
         n26167, n26168, n26169, n26170, n26171, n26172, n26173, n26174,
         n26175, n26176, n26177, n26178, n26179, n26180, n26181, n26182,
         n26183, n26184, n26185, n26186, n26187, n26188, n26189, n26190,
         n26191, n26192, n26193, n26194, n26195, n26196, n26197, n26198,
         n26199, n26200, n26201, n26202, n26203, n26204, n26205, n26206,
         n26207, n26208, n26209, n26210, n26211, n26212, n26213, n26214,
         n26215, n26216, n26217, n26218, n26219, n26220, n26221, n26222,
         n26223, n26224, n26225, n26226, n26227, n26228, n26229, n26230,
         n26231, n26232, n26233, n26234, n26235, n26236, n26237, n26238,
         n26239, n26240, n26241, n26242, n26243, n26244, n26245, n26246,
         n26247, n26248, n26249, n26250, n26251, n26252, n26253, n26254,
         n26255, n26256, n26257, n26258, n26259, n26260, n26261, n26262,
         n26263, n26264, n26265, n26266, n26267, n26268, n26269, n26270,
         n26271, n26272, n26273, n26274, n26275, n26276, n26277, n26278,
         n26279, n26280, n26281, n26282, n26283, n26284, n26285, n26286,
         n26287, n26288, n26289, n26290, n26291, n26292, n26293, n26294,
         n26295, n26296, n26297, n26298, n26299, n26300, n26301, n26302,
         n26303, n26304, n26305, n26306, n26307, n26308, n26309, n26310,
         n26311, n26312, n26313, n26314, n26315, n26316, n26317, n26318,
         n26319, n26320, n26321, n26322, n26323, n26324, n26325, n26326,
         n26327, n26328, n26329, n26330, n26331, n26332, n26333, n26334,
         n26335, n26336, n26337, n26338, n26339, n26340, n26341, n26342,
         n26343, n26344, n26345, n26346, n26347, n26348, n26349, n26350,
         n26351, n26352, n26353, n26354, n26355, n26356, n26357, n26358,
         n26359, n26360, n26361, n26362, n26363, n26364, n26365, n26366,
         n26367, n26368, n26369, n26370, n26371, n26372, n26373, n26374,
         n26375, n26376, n26377, n26378, n26379, n26380, n26381, n26382,
         n26383, n26384, n26385, n26386, n26387, n26388, n26389, n26390,
         n26391, n26392, n26393, n26394, n26395, n26396, n26397, n26398,
         n26399, n26400, n26401, n26402, n26403, n26404, n26405, n26406,
         n26407, n26408, n26409, n26410, n26411, n26412, n26413, n26414,
         n26415, n26416, n26417, n26418, n26419, n26420, n26421, n26422,
         n26423, n26424, n26425, n26426, n26427, n26428, n26429, n26430,
         n26431, n26432, n26433, n26434, n26435, n26436, n26437, n26438,
         n26439, n26440, n26441, n26442, n26443, n26444, n26445, n26446,
         n26447, n26448, n26449, n26450, n26451, n26452, n26453, n26454,
         n26455, n26456, n26457, n26458, n26459, n26460, n26461, n26462,
         n26463, n26464, n26465, n26466, n26467, n26468, n26469, n26470,
         n26471, n26472, n26473, n26474, n26475, n26476, n26477, n26478,
         n26479, n26480, n26481, n26482, n26483, n26484, n26485, n26486,
         n26487, n26488, n26489, n26490, n26491, n26492, n26493, n26494,
         n26495, n26496, n26497, n26498, n26499, n26500, n26501, n26502,
         n26503, n26504, n26505, n26506, n26507, n26508, n26509, n26510,
         n26511, n26512, n26513, n26514, n26515, n26516, n26517, n26518,
         n26519, n26520, n26521, n26522, n26523, n26524, n26525, n26526,
         n26527, n26528, n26529, n26530, n26531, n26532, n26533, n26534,
         n26535, n26536, n26537, n26538, n26539, n26540, n26541, n26542,
         n26543, n26544, n26545, n26546, n26547, n26548, n26549, n26550,
         n26551, n26552, n26553, n26554, n26555, n26556, n26557, n26558,
         n26559, n26560, n26561, n26562, n26563, n26564, n26565, n26566,
         n26567, n26568, n26569, n26570, n26571, n26572, n26573, n26574,
         n26575, n26576, n26577, n26578, n26579, n26580, n26581, n26582,
         n26583, n26584, n26585, n26586, n26587, n26588, n26589, n26590,
         n26591, n26592, n26593, n26594, n26595, n26596, n26597, n26598,
         n26599, n26600, n26601, n26602, n26603, n26604, n26605, n26606,
         n26607, n26608, n26609, n26610, n26611, n26612, n26613, n26614,
         n26615, n26616, n26617, n26618, n26619, n26620, n26621, n26622,
         n26623, n26624, n26625, n26626, n26627, n26628, n26629, n26630,
         n26631, n26632, n26633, n26634, n26635, n26636, n26637, n26638,
         n26639, n26640, n26641, n26642, n26643, n26644, n26645, n26646,
         n26647, n26648, n26649, n26650, n26651, n26652, n26653, n26654,
         n26655, n26656, n26657, n26658, n26659, n26660, n26661, n26662,
         n26663, n26664, n26665, n26666, n26667, n26668, n26669, n26670,
         n26671, n26672, n26673, n26674, n26675, n26676, n26677, n26678,
         n26679, n26680, n26681, n26682, n26683, n26684, n26685, n26686,
         n26687, n26688, n26689, n26690, n26691, n26692, n26693, n26694,
         n26695, n26696, n26697, n26698, n26699, n26700, n26701, n26702,
         n26703, n26704, n26705, n26706, n26707, n26708, n26709, n26710,
         n26711, n26712, n26713, n26714, n26715, n26716, n26717, n26718,
         n26719, n26720, n26721, n26722, n26723, n26724, n26725, n26726,
         n26727, n26728, n26729, n26730, n26731, n26732, n26733, n26734,
         n26735, n26736, n26737, n26738, n26739, n26740, n26741, n26742,
         n26743, n26744, n26745, n26746, n26747, n26748, n26749, n26750,
         n26751, n26752, n26753, n26754, n26755, n26756, n26757, n26758,
         n26759, n26760, n26761, n26762, n26763, n26764, n26765, n26766,
         n26767, n26768, n26769, n26770, n26771, n26772, n26773, n26774,
         n26775, n26776, n26777, n26778, n26779, n26780, n26781, n26782,
         n26783, n26784, n26785, n26786, n26787, n26788, n26789, n26790,
         n26791, n26792, n26793, n26794, n26795, n26796, n26797, n26798,
         n26799, n26800, n26801, n26802, n26803, n26804, n26805, n26806,
         n26807, n26808, n26809, n26810, n26811, n26812, n26813, n26814,
         n26815, n26816, n26817, n26818, n26819, n26820, n26821, n26822,
         n26823, n26824, n26825, n26826, n26827, n26828, n26829, n26830,
         n26831, n26832, n26833, n26834, n26835, n26836, n26837, n26838,
         n26839, n26840, n26841, n26842, n26843, n26844, n26845, n26846,
         n26847, n26848, n26849, n26850, n26851, n26852, n26853, n26854,
         n26855, n26856, n26857, n26858, n26859, n26860, n26861, n26862,
         n26863, n26864, n26865, n26866, n26867, n26868, n26869, n26870,
         n26871, n26872, n26873, n26874, n26875, n26876, n26877, n26878,
         n26879, n26880, n26881, n26882, n26883, n26884, n26885, n26886,
         n26887, n26888, n26889, n26890, n26891, n26892, n26893, n26894,
         n26895, n26896, n26897, n26898, n26899, n26900, n26901, n26902,
         n26903, n26904, n26905, n26906, n26907, n26908, n26909, n26910,
         n26911, n26912, n26913, n26914, n26915, n26916, n26917, n26918,
         n26919, n26920, n26921, n26922, n26923, n26924, n26925, n26926,
         n26927, n26928, n26929, n26930, n26931, n26932, n26933, n26934,
         n26935, n26936, n26937, n26938, n26939, n26940, n26941, n26942,
         n26943, n26944, n26945, n26946, n26947, n26948, n26949, n26950,
         n26951, n26952, n26953, n26954, n26955, n26956, n26957, n26958,
         n26959, n26960, n26961, n26962, n26963, n26964, n26965, n26966,
         n26967, n26968, n26969, n26970, n26971, n26972, n26973, n26974,
         n26975, n26976, n26977, n26978, n26979, n26980, n26981, n26982,
         n26983, n26984, n26985, n26986, n26987, n26988, n26989, n26990,
         n26991, n26992, n26993, n26994, n26995, n26996, n26997, n26998,
         n26999, n27000, n27001, n27002, n27003, n27004, n27005, n27006,
         n27007, n27008, n27009, n27010, n27011, n27012, n27013, n27014,
         n27015, n27016, n27017, n27018, n27019, n27020, n27021, n27022,
         n27023, n27024, n27025, n27026, n27027, n27028, n27029, n27030,
         n27031, n27032, n27033, n27034, n27035, n27036, n27037, n27038,
         n27039, n27040, n27041, n27042, n27043, n27044, n27045, n27046,
         n27047, n27048, n27049, n27050, n27051, n27052, n27053, n27054,
         n27055, n27056, n27057, n27058, n27059, n27060, n27061, n27062,
         n27063, n27064, n27065, n27066, n27067, n27068, n27069, n27070,
         n27071, n27072, n27073, n27074, n27075, n27076, n27077, n27078,
         n27079, n27080, n27081, n27082, n27083, n27084, n27085, n27086,
         n27087, n27088, n27089, n27090, n27091, n27092, n27093, n27094,
         n27095, n27096, n27097, n27098, n27099, n27100, n27101, n27102,
         n27103, n27104, n27105, n27106, n27107, n27108, n27109, n27110,
         n27111, n27112, n27113, n27114, n27115, n27116, n27117, n27118,
         n27119, n27120, n27121, n27122, n27123, n27124, n27125, n27126,
         n27127, n27128, n27129, n27130, n27131, n27132, n27133, n27134,
         n27135, n27136, n27137, n27138, n27139, n27140, n27141, n27142,
         n27143, n27144, n27145, n27146, n27147, n27148, n27149, n27150,
         n27151, n27152, n27153, n27154, n27155, n27156, n27157, n27158,
         n27159, n27160, n27161, n27162, n27163, n27164, n27165, n27166,
         n27167, n27168, n27169, n27170, n27171, n27172, n27173, n27174,
         n27175, n27176, n27177, n27178, n27179, n27180, n27181, n27182,
         n27183, n27184, n27185, n27186, n27187, n27188, n27189, n27190,
         n27191, n27192, n27193, n27194, n27195, n27196, n27197, n27198,
         n27199, n27200, n27201, n27202, n27203, n27204, n27205, n27206,
         n27207, n27208, n27209, n27210, n27211, n27212, n27213, n27214,
         n27215, n27216, n27217, n27218, n27219, n27220, n27221, n27222,
         n27223, n27224, n27225, n27226, n27227, n27228, n27229, n27230,
         n27231, n27232, n27233, n27234, n27235, n27236, n27237, n27238,
         n27239, n27240, n27241, n27242, n27243, n27244, n27245, n27246,
         n27247, n27248, n27249, n27250, n27251, n27252, n27253, n27254,
         n27255, n27256, n27257, n27258, n27259, n27260, n27261, n27262,
         n27263, n27264, n27265, n27266, n27267, n27268, n27269, n27270,
         n27271, n27272, n27273, n27274, n27275, n27276, n27277, n27278,
         n27279, n27280, n27281, n27282, n27283, n27284, n27285, n27286,
         n27287, n27288, n27289, n27290, n27291, n27292, n27293, n27294,
         n27295, n27296, n27297, n27298, n27299, n27300, n27301, n27302,
         n27303, n27304, n27305, n27306, n27307, n27308, n27309, n27310,
         n27311, n27312, n27313, n27314, n27315, n27316, n27317, n27318,
         n27319, n27320, n27321, n27322, n27323, n27324, n27325, n27326,
         n27327, n27328, n27329, n27330, n27331, n27332, n27333, n27334,
         n27335, n27336, n27337, n27338, n27339, n27340, n27341, n27342,
         n27343, n27344, n27345, n27346, n27347, n27348, n27349, n27350,
         n27351, n27352, n27353, n27354, n27355, n27356, n27357, n27358,
         n27359, n27360, n27361, n27362, n27363, n27364, n27365, n27366,
         n27367, n27368, n27369, n27370, n27371, n27372, n27373, n27374,
         n27375, n27376, n27377, n27378, n27379, n27380, n27381, n27382,
         n27383, n27384, n27385, n27386, n27387, n27388, n27389, n27390,
         n27391, n27392, n27393, n27394, n27395, n27396, n27397, n27398,
         n27399, n27400, n27401, n27402, n27403, n27404, n27405, n27406,
         n27407, n27408, n27409, n27410, n27411, n27412, n27413, n27414,
         n27415, n27416, n27417, n27418, n27419, n27420, n27421, n27422,
         n27423, n27424, n27425, n27426, n27427, n27428, n27429, n27430,
         n27431, n27432, n27433, n27434, n27435, n27436, n27437, n27438,
         n27439, n27440, n27441, n27442, n27443, n27444, n27445, n27446,
         n27447, n27448, n27449, n27450, n27451, n27452, n27453, n27454,
         n27455, n27456, n27457, n27458, n27459, n27460, n27461, n27462,
         n27463, n27464, n27465, n27466, n27467, n27468, n27469, n27470,
         n27471, n27472, n27473, n27474, n27475, n27476, n27477, n27478,
         n27479, n27480, n27481, n27482, n27483, n27484, n27485, n27486,
         n27487, n27488, n27489, n27490, n27491, n27492, n27493, n27494,
         n27495, n27496, n27497, n27498, n27499, n27500, n27501, n27502,
         n27503, n27504, n27505, n27506, n27507, n27508, n27509, n27510,
         n27511, n27512, n27513, n27514, n27515, n27516, n27517, n27518,
         n27519, n27520, n27521, n27522, n27523, n27524, n27525, n27526,
         n27527, n27528, n27529, n27530, n27531, n27532, n27533, n27534,
         n27535, n27536, n27537, n27538, n27539, n27540, n27541, n27542,
         n27543, n27544, n27545, n27546, n27547, n27548, n27549, n27550,
         n27551, n27552, n27553, n27554, n27555, n27556, n27557, n27558,
         n27559, n27560, n27561, n27562, n27563, n27564, n27565, n27566,
         n27567, n27568, n27569, n27570, n27571, n27572, n27573, n27574,
         n27575, n27576, n27577, n27578, n27579, n27580, n27581, n27582,
         n27583, n27584, n27585, n27586, n27587, n27588, n27589, n27590,
         n27591, n27592, n27593, n27594, n27595, n27596, n27597, n27598,
         n27599, n27600, n27601, n27602, n27603, n27604, n27605, n27606,
         n27607, n27608, n27609, n27610, n27611, n27612, n27613, n27614,
         n27615, n27616, n27617, n27618, n27619, n27620, n27621, n27622,
         n27623, n27624, n27625, n27626, n27627, n27628, n27629, n27630,
         n27631, n27632, n27633, n27634, n27635, n27636, n27637, n27638,
         n27639, n27640, n27641, n27642, n27643, n27644, n27645, n27646,
         n27647, n27648, n27649, n27650, n27651, n27652, n27653, n27654,
         n27655, n27656, n27657, n27658, n27659, n27660, n27661, n27662,
         n27663, n27664, n27665, n27666, n27667, n27668, n27669, n27670,
         n27671, n27672, n27673, n27674, n27675, n27676, n27677, n27678,
         n27679, n27680, n27681, n27682, n27683, n27684, n27685, n27686,
         n27687, n27688, n27689, n27690, n27691, n27692, n27693, n27694,
         n27695, n27696, n27697, n27698, n27699, n27700, n27701, n27702,
         n27703, n27704, n27705, n27706, n27707, n27708, n27709, n27710,
         n27711, n27712, n27713, n27714, n27715, n27716, n27717, n27718,
         n27719, n27720, n27721, n27722, n27723, n27724, n27725, n27726,
         n27727, n27728, n27729, n27730, n27731, n27732, n27733, n27734,
         n27735, n27736, n27737, n27738, n27739, n27740, n27741, n27742,
         n27743, n27744, n27745, n27746, n27747, n27748, n27749, n27750,
         n27751, n27752, n27753, n27754, n27755, n27756, n27757, n27758,
         n27759, n27760, n27761, n27762, n27763, n27764, n27765, n27766,
         n27767, n27768, n27769, n27770, n27771, n27772, n27773, n27774,
         n27775, n27776, n27777, n27778, n27779, n27780, n27781, n27782,
         n27783, n27784, n27785, n27786, n27787, n27788, n27789, n27790,
         n27791, n27792, n27793, n27794, n27795, n27796, n27797, n27798,
         n27799, n27800, n27801, n27802, n27803, n27804, n27805, n27806,
         n27807, n27808, n27809, n27810, n27811, n27812, n27813, n27814,
         n27815, n27816, n27817, n27818, n27819, n27820, n27821, n27822,
         n27823, n27824, n27825, n27826, n27827, n27828, n27829, n27830,
         n27831, n27832, n27833, n27834, n27835, n27836, n27837, n27838,
         n27839, n27840, n27841, n27842, n27843, n27844, n27845, n27846,
         n27847, n27848, n27849, n27850, n27851, n27852, n27853, n27854,
         n27855, n27856, n27857, n27858, n27859, n27860, n27861, n27862,
         n27863, n27864, n27865, n27866, n27867, n27868, n27869, n27870,
         n27871, n27872, n27873, n27874, n27875, n27876, n27877, n27878,
         n27879, n27880, n27881, n27882, n27883, n27884, n27885, n27886,
         n27887, n27888, n27889, n27890, n27891, n27892, n27893, n27894,
         n27895, n27896, n27897, n27898, n27899, n27900, n27901, n27902,
         n27903, n27904, n27905, n27906, n27907, n27908, n27909, n27910,
         n27911, n27912, n27913, n27914, n27915, n27916, n27917, n27918,
         n27919, n27920, n27921, n27922, n27923, n27924, n27925, n27926,
         n27927, n27928, n27929, n27930, n27931, n27932, n27933, n27934,
         n27935, n27936, n27937, n27938, n27939, n27940, n27941, n27942,
         n27943, n27944, n27945, n27946, n27947, n27948, n27949, n27950,
         n27951, n27952, n27953, n27954, n27955, n27956, n27957, n27958,
         n27959, n27960, n27961, n27962, n27963, n27964, n27965, n27966,
         n27967, n27968, n27969, n27970, n27971, n27972, n27973, n27974,
         n27975, n27976, n27977, n27978, n27979, n27980, n27981, n27982,
         n27983, n27984, n27985, n27986, n27987, n27988, n27989, n27990,
         n27991, n27992, n27993, n27994, n27995, n27996, n27997, n27998,
         n27999, n28000, n28001, n28002, n28003, n28004, n28005, n28006,
         n28007, n28008, n28009, n28010, n28011, n28012, n28013, n28014,
         n28015, n28016, n28017, n28018, n28019, n28020, n28021, n28022,
         n28023, n28024, n28025, n28026, n28027, n28028, n28029, n28030,
         n28031, n28032, n28033, n28034, n28035, n28036, n28037, n28038,
         n28039, n28040, n28041, n28042, n28043, n28044, n28045, n28046,
         n28047, n28048, n28049, n28050, n28051, n28052, n28053, n28054,
         n28055, n28056, n28057, n28058, n28059, n28060, n28061, n28062,
         n28063, n28064, n28065, n28066, n28067, n28068, n28069, n28070,
         n28071, n28072, n28073, n28074, n28075, n28076, n28077, n28078,
         n28079, n28080, n28081, n28082, n28083, n28084, n28085, n28086,
         n28087, n28088, n28089, n28090, n28091, n28092, n28093, n28094,
         n28095, n28096, n28097, n28098, n28099, n28100, n28101, n28102,
         n28103, n28104, n28105, n28106, n28107, n28108, n28109, n28110,
         n28111, n28112, n28113, n28114, n28115, n28116, n28117, n28118,
         n28119, n28120, n28121, n28122, n28123, n28124, n28125, n28126,
         n28127, n28128, n28129, n28130, n28131, n28132, n28133, n28134,
         n28135, n28136, n28137, n28138, n28139, n28140, n28141, n28142,
         n28143, n28144, n28145, n28146, n28147, n28148, n28149, n28150,
         n28151, n28152, n28153, n28154, n28155, n28156, n28157, n28158,
         n28159, n28160, n28161, n28162, n28163, n28164, n28165, n28166,
         n28167, n28168, n28169, n28170, n28171, n28172, n28173, n28174,
         n28175, n28176, n28177, n28178, n28179, n28180, n28181, n28182,
         n28183, n28184, n28185, n28186, n28187, n28188, n28189, n28190,
         n28191, n28192, n28193, n28194, n28195, n28196, n28197, n28198,
         n28199, n28200, n28201, n28202, n28203, n28204, n28205, n28206,
         n28207, n28208, n28209, n28210, n28211, n28212, n28213, n28214,
         n28215, n28216, n28217, n28218, n28219, n28220, n28221, n28222,
         n28223, n28224, n28225, n28226, n28227, n28228, n28229, n28230,
         n28231, n28232, n28233, n28234, n28235, n28236, n28237, n28238,
         n28239, n28240, n28241, n28242, n28243, n28244, n28245, n28246,
         n28247, n28248, n28249, n28250, n28251, n28252, n28253, n28254,
         n28255, n28256, n28257, n28258, n28259, n28260, n28261, n28262,
         n28263, n28264, n28265, n28266, n28267, n28268, n28269, n28270,
         n28271, n28272, n28273, n28274, n28275, n28276, n28277, n28278,
         n28279, n28280, n28281, n28282, n28283, n28284, n28285, n28286,
         n28287, n28288, n28289, n28290, n28291, n28292, n28293, n28294,
         n28295, n28296, n28297, n28298, n28299, n28300, n28301, n28302,
         n28303, n28304, n28305, n28306, n28307, n28308, n28309, n28310,
         n28311, n28312, n28313, n28314, n28315, n28316, n28317, n28318,
         n28319, n28320, n28321, n28322, n28323, n28324, n28325, n28326,
         n28327, n28328, n28329, n28330, n28331, n28332, n28333, n28334,
         n28335, n28336, n28337, n28338, n28339, n28340, n28341, n28342,
         n28343, n28344, n28345, n28346, n28347, n28348, n28349, n28350,
         n28351, n28352, n28353, n28354, n28355, n28356, n28357, n28358,
         n28359, n28360, n28361, n28362, n28363, n28364, n28365, n28366,
         n28367, n28368, n28369, n28370, n28371, n28372, n28373, n28374,
         n28375, n28376, n28377, n28378, n28379, n28380, n28381, n28382,
         n28383, n28384, n28385, n28386, n28387, n28388, n28389, n28390,
         n28391, n28392, n28393, n28394, n28395, n28396, n28397, n28398,
         n28399, n28400, n28401, n28402, n28403, n28404, n28405, n28406,
         n28407, n28408, n28409, n28410, n28411, n28412, n28413, n28414,
         n28415, n28416, n28417, n28418, n28419, n28420, n28421, n28422,
         n28423, n28424, n28425, n28426, n28427, n28428, n28429, n28430,
         n28431, n28432, n28433, n28434, n28435, n28436, n28437, n28438,
         n28439, n28440, n28441, n28442, n28443, n28444, n28445, n28446,
         n28447, n28448, n28449, n28450, n28451, n28452, n28453, n28454,
         n28455, n28456, n28457, n28458, n28459, n28460, n28461, n28462,
         n28463, n28464, n28465, n28466, n28467, n28468, n28469, n28470,
         n28471, n28472, n28473, n28474, n28475, n28476, n28477, n28478,
         n28479, n28480, n28481, n28482, n28483, n28484, n28485, n28486,
         n28487, n28488, n28489, n28490, n28491, n28492, n28493, n28494,
         n28495, n28496, n28497, n28498, n28499, n28500, n28501, n28502,
         n28503, n28504, n28505, n28506, n28507, n28508, n28509, n28510,
         n28511, n28512, n28513, n28514, n28515, n28516, n28517, n28518,
         n28519, n28520, n28521, n28522, n28523, n28524, n28525, n28526,
         n28527, n28528, n28529, n28530, n28531, n28532, n28533, n28534,
         n28535, n28536, n28537, n28538, n28539, n28540, n28541, n28542,
         n28543, n28544, n28545, n28546, n28547, n28548, n28549, n28550,
         n28551, n28552, n28553, n28554, n28555, n28556, n28557, n28558,
         n28559, n28560, n28561, n28562, n28563, n28564, n28565, n28566,
         n28567, n28568, n28569, n28570, n28571, n28572, n28573, n28574,
         n28575, n28576, n28577, n28578, n28579, n28580, n28581, n28582,
         n28583, n28584, n28585, n28586, n28587, n28588, n28589, n28590,
         n28591, n28592, n28593, n28594, n28595, n28596, n28597, n28598,
         n28599, n28600, n28601, n28602, n28603, n28604, n28605, n28606,
         n28607, n28608, n28609, n28610, n28611, n28612, n28613, n28614,
         n28615, n28616, n28617, n28618, n28619, n28620, n28621, n28622,
         n28623, n28624, n28625, n28626, n28627, n28628, n28629, n28630,
         n28631, n28632, n28633, n28634, n28635, n28636, n28637, n28638,
         n28639, n28640, n28641, n28642, n28643, n28644, n28645, n28646,
         n28647, n28648, n28649, n28650, n28651, n28652, n28653, n28654,
         n28655, n28656, n28657, n28658, n28659, n28660, n28661, n28662,
         n28663, n28664, n28665, n28666, n28667, n28668, n28669, n28670,
         n28671, n28672, n28673, n28674, n28675, n28676, n28677, n28678,
         n28679, n28680, n28681, n28682, n28683, n28684, n28685, n28686,
         n28687, n28688, n28689, n28690, n28691, n28692, n28693, n28694,
         n28695, n28696, n28697, n28698, n28699, n28700, n28701, n28702,
         n28703, n28704, n28705, n28706, n28707, n28708, n28709, n28710,
         n28711, n28712, n28713, n28714, n28715, n28716, n28717, n28718,
         n28719, n28720, n28721, n28722, n28723, n28724, n28725, n28726,
         n28727, n28728, n28729, n28730, n28731, n28732, n28733, n28734,
         n28735, n28736, n28737, n28738, n28739, n28740, n28741, n28742,
         n28743, n28744, n28745, n28746, n28747, n28748, n28749, n28750,
         n28751, n28752, n28753, n28754, n28755, n28756, n28757, n28758,
         n28759, n28760, n28761, n28762, n28763, n28764, n28765, n28766,
         n28767, n28768, n28769, n28770, n28771, n28772, n28773, n28774,
         n28775, n28776, n28777, n28778, n28779, n28780, n28781, n28782,
         n28783, n28784, n28785, n28786, n28787, n28788, n28789, n28790,
         n28791, n28792, n28793, n28794, n28795, n28796, n28797, n28798,
         n28799, n28800, n28801, n28802, n28803, n28804, n28805, n28806,
         n28807, n28808, n28809, n28810, n28811, n28812, n28813, n28814,
         n28815, n28816, n28817, n28818, n28819, n28820, n28821, n28822,
         n28823, n28824, n28825, n28826, n28827, n28828, n28829, n28830,
         n28831, n28832, n28833, n28834, n28835, n28836, n28837, n28838,
         n28839, n28840, n28841, n28842, n28843, n28844, n28845, n28846,
         n28847, n28848, n28849, n28850, n28851, n28852, n28853, n28854,
         n28855, n28856, n28857, n28858, n28859, n28860, n28861, n28862,
         n28863, n28864, n28865, n28866, n28867, n28868, n28869, n28870,
         n28871, n28872, n28873, n28874, n28875, n28876, n28877, n28878,
         n28879, n28880, n28881, n28882, n28883, n28884, n28885, n28886,
         n28887, n28888, n28889, n28890, n28891, n28892, n28893, n28894,
         n28895, n28896, n28897, n28898, n28899, n28900, n28901, n28902,
         n28903, n28904, n28905, n28906, n28907, n28908, n28909, n28910,
         n28911, n28912, n28913, n28914, n28915, n28916, n28917, n28918,
         n28919, n28920, n28921, n28922, n28923, n28924, n28925, n28926,
         n28927, n28928, n28929, n28930, n28931, n28932, n28933, n28934,
         n28935, n28936, n28937, n28938, n28939, n28940, n28941, n28942,
         n28943, n28944, n28945, n28946, n28947, n28948, n28949, n28950,
         n28951, n28952, n28953, n28954, n28955, n28956, n28957, n28958,
         n28959, n28960, n28961, n28962, n28963, n28964, n28965, n28966,
         n28967, n28968, n28969, n28970, n28971, n28972, n28973, n28974,
         n28975, n28976, n28977, n28978, n28979, n28980, n28981, n28982,
         n28983, n28984, n28985, n28986, n28987, n28988, n28989, n28990,
         n28991, n28992, n28993, n28994, n28995, n28996, n28997, n28998,
         n28999, n29000, n29001, n29002, n29003, n29004, n29005, n29006,
         n29007, n29008, n29009, n29010, n29011, n29012, n29013, n29014,
         n29015, n29016, n29017, n29018, n29019, n29020, n29021, n29022,
         n29023, n29024, n29025, n29026, n29027, n29028, n29029, n29030,
         n29031, n29032, n29033, n29034, n29035, n29036, n29037, n29038,
         n29039, n29040, n29041, n29042, n29043, n29044, n29045, n29046,
         n29047, n29048, n29049, n29050, n29051, n29052, n29053, n29054,
         n29055, n29056, n29057, n29058, n29059, n29060, n29061, n29062,
         n29063, n29064, n29065, n29066, n29067, n29068, n29069, n29070,
         n29071, n29072, n29073, n29074, n29075, n29076, n29077, n29078,
         n29079, n29080, n29081, n29082, n29083, n29084, n29085, n29086,
         n29087, n29088, n29089, n29090, n29091, n29092, n29093, n29094,
         n29095, n29096, n29097, n29098, n29099, n29100, n29101, n29102,
         n29103, n29104, n29105, n29106, n29107, n29108, n29109, n29110,
         n29111, n29112, n29113, n29114, n29115, n29116, n29117, n29118,
         n29119, n29120, n29121, n29122, n29123, n29124, n29125, n29126,
         n29127, n29128, n29129, n29130, n29131, n29132, n29133, n29134,
         n29135, n29136, n29137, n29138, n29139, n29140, n29141, n29142,
         n29143, n29144, n29145, n29146, n29147, n29148, n29149, n29150,
         n29151, n29152, n29153, n29154, n29155, n29156, n29157, n29158,
         n29159, n29160, n29161, n29162, n29163, n29164, n29165, n29166,
         n29167, n29168, n29169, n29170, n29171, n29172, n29173, n29174,
         n29175, n29176, n29177, n29178, n29179, n29180, n29181, n29182,
         n29183, n29184, n29185, n29186, n29187, n29188, n29189, n29190,
         n29191, n29192, n29193, n29194, n29195, n29196, n29197, n29198,
         n29199, n29200, n29201, n29202, n29203, n29204, n29205, n29206,
         n29207, n29208, n29209, n29210, n29211, n29212, n29213, n29214,
         n29215, n29216, n29217, n29218, n29219, n29220, n29221, n29222,
         n29223, n29224, n29225, n29226, n29227, n29228, n29229, n29230,
         n29231, n29232, n29233, n29234, n29235, n29236, n29237, n29238,
         n29239, n29240, n29241, n29242, n29243, n29244, n29245, n29246,
         n29247, n29248, n29249, n29250, n29251, n29252, n29253, n29254,
         n29255, n29256, n29257, n29258, n29259, n29260, n29261, n29262,
         n29263, n29264, n29265, n29266, n29267, n29268, n29269, n29270,
         n29271, n29272, n29273, n29274, n29275, n29276, n29277, n29278,
         n29279, n29280, n29281, n29282, n29283, n29284, n29285, n29286,
         n29287, n29288, n29289, n29290, n29291, n29292, n29293, n29294,
         n29295, n29296, n29297, n29298, n29299, n29300, n29301, n29302,
         n29303, n29304, n29305, n29306, n29307, n29308, n29309, n29310,
         n29311, n29312, n29313, n29314, n29315, n29316, n29317, n29318,
         n29319, n29320, n29321, n29322, n29323, n29324, n29325, n29326,
         n29327, n29328, n29329, n29330, n29331, n29332, n29333, n29334,
         n29335, n29336, n29337, n29338, n29339, n29340, n29341, n29342,
         n29343, n29344, n29345, n29346, n29347, n29348, n29349, n29350,
         n29351, n29352, n29353, n29354, n29355, n29356, n29357, n29358,
         n29359, n29360, n29361, n29362, n29363, n29364, n29365, n29366,
         n29367, n29368, n29369, n29370, n29371, n29372, n29373, n29374,
         n29375, n29376, n29377, n29378, n29379, n29380, n29381, n29382,
         n29383, n29384, n29385, n29386, n29387, n29388, n29389, n29390,
         n29391, n29392, n29393, n29394, n29395, n29396, n29397, n29398,
         n29399, n29400, n29401, n29402, n29403, n29404, n29405, n29406,
         n29407, n29408, n29409, n29410, n29411, n29412, n29413, n29414,
         n29415, n29416, n29417, n29418, n29419, n29420, n29421, n29422,
         n29423, n29424, n29425, n29426, n29427, n29428, n29429, n29430,
         n29431, n29432, n29433, n29434, n29435, n29436, n29437, n29438,
         n29439, n29440, n29441, n29442, n29443, n29444, n29445, n29446,
         n29447, n29448, n29449, n29450, n29451, n29452, n29453, n29454,
         n29455, n29456, n29457, n29458, n29459, n29460, n29461, n29462,
         n29463, n29464, n29465, n29466, n29467, n29468, n29469, n29470,
         n29471, n29472, n29473, n29474, n29475, n29476, n29477, n29478,
         n29479, n29480, n29481, n29482, n29483, n29484, n29485, n29486,
         n29487, n29488, n29489, n29490, n29491, n29492, n29493, n29494,
         n29495, n29496, n29497, n29498, n29499, n29500, n29501, n29502,
         n29503, n29504, n29505, n29506, n29507, n29508, n29509, n29510,
         n29511, n29512, n29513, n29514, n29515, n29516, n29517, n29518,
         n29519, n29520, n29521, n29522, n29523, n29524, n29525, n29526,
         n29527, n29528, n29529, n29530, n29531, n29532, n29533, n29534,
         n29535, n29536, n29537, n29538, n29539, n29540, n29541, n29542,
         n29543, n29544, n29545, n29546, n29547, n29548, n29549, n29550,
         n29551, n29552, n29553, n29554, n29555, n29556, n29557, n29558,
         n29559, n29560, n29561, n29562, n29563, n29564, n29565, n29566,
         n29567, n29568, n29569, n29570, n29571, n29572, n29573, n29574,
         n29575, n29576, n29577, n29578, n29579, n29580, n29581, n29582,
         n29583, n29584, n29585, n29586, n29587, n29588, n29589, n29590,
         n29591, n29592, n29593, n29594, n29595, n29596, n29597, n29598,
         n29599, n29600, n29601, n29602, n29603, n29604, n29605, n29606,
         n29607, n29608, n29609, n29610, n29611, n29612, n29613, n29614,
         n29615, n29616, n29617, n29618, n29619, n29620, n29621, n29622,
         n29623, n29624, n29625, n29626, n29627, n29628, n29629, n29630,
         n29631, n29632, n29633, n29634, n29635, n29636, n29637, n29638,
         n29639, n29640, n29641, n29642, n29643, n29644, n29645, n29646,
         n29647, n29648, n29649, n29650, n29651, n29652, n29653, n29654,
         n29655, n29656, n29657, n29658, n29659, n29660, n29661, n29662,
         n29663, n29664, n29665, n29666, n29667, n29668, n29669, n29670,
         n29671, n29672, n29673, n29674, n29675, n29676, n29677, n29678,
         n29679, n29680, n29681, n29682, n29683, n29684, n29685, n29686,
         n29687, n29688, n29689, n29690, n29691, n29692, n29693, n29694,
         n29695, n29696, n29697, n29698, n29699, n29700, n29701, n29702,
         n29703, n29704, n29705, n29706, n29707, n29708, n29709, n29710,
         n29711, n29712, n29713, n29714, n29715, n29716, n29717, n29718,
         n29719, n29720, n29721, n29722, n29723, n29724, n29725, n29726,
         n29727, n29728, n29729, n29730, n29731, n29732, n29733, n29734,
         n29735, n29736, n29737, n29738, n29739, n29740, n29741, n29742,
         n29743, n29744, n29745, n29746, n29747, n29748, n29749, n29750,
         n29751, n29752, n29753, n29754, n29755, n29756, n29757, n29758,
         n29759, n29760, n29761, n29762, n29763, n29764, n29765, n29766,
         n29767, n29768, n29769, n29770, n29771, n29772, n29773, n29774,
         n29775, n29776, n29777, n29778, n29779, n29780, n29781, n29782,
         n29783, n29784, n29785, n29786, n29787, n29788, n29789, n29790,
         n29791, n29792, n29793, n29794, n29795, n29796, n29797, n29798,
         n29799, n29800, n29801, n29802, n29803, n29804, n29805, n29806,
         n29807, n29808, n29809, n29810, n29811, n29812, n29813, n29814,
         n29815, n29816, n29817, n29818, n29819, n29820, n29821, n29822,
         n29823, n29824, n29825, n29826, n29827, n29828, n29829, n29830,
         n29831, n29832, n29833, n29834, n29835, n29836, n29837, n29838,
         n29839, n29840, n29841, n29842, n29843, n29844, n29845, n29846,
         n29847, n29848, n29849, n29850, n29851, n29852, n29853, n29854,
         n29855, n29856, n29857, n29858, n29859, n29860, n29861, n29862,
         n29863, n29864, n29865, n29866, n29867, n29868, n29869, n29870,
         n29871, n29872, n29873, n29874, n29875, n29876, n29877, n29878,
         n29879, n29880, n29881, n29882, n29883, n29884, n29885, n29886,
         n29887, n29888, n29889, n29890, n29891, n29892, n29893, n29894,
         n29895, n29896, n29897, n29898, n29899, n29900, n29901, n29902,
         n29903, n29904, n29905, n29906, n29907, n29908, n29909, n29910,
         n29911, n29912, n29913, n29914, n29915, n29916, n29917, n29918,
         n29919, n29920, n29921, n29922, n29923, n29924, n29925, n29926,
         n29927, n29928, n29929, n29930, n29931, n29932, n29933, n29934,
         n29935, n29936, n29937, n29938, n29939, n29940, n29941, n29942,
         n29943, n29944, n29945, n29946, n29947, n29948, n29949, n29950,
         n29951, n29952, n29953, n29954, n29955, n29956, n29957, n29958,
         n29959, n29960, n29961, n29962, n29963, n29964, n29965, n29966,
         n29967, n29968, n29969, n29970, n29971, n29972, n29973, n29974,
         n29975, n29976, n29977, n29978, n29979, n29980, n29981, n29982,
         n29983, n29984, n29985, n29986, n29987, n29988, n29989, n29990,
         n29991, n29992, n29993, n29994, n29995, n29996, n29997, n29998,
         n29999, n30000, n30001, n30002, n30003, n30004, n30005, n30006,
         n30007, n30008, n30009, n30010, n30011, n30012, n30013, n30014,
         n30015, n30016, n30017, n30018, n30019, n30020, n30021, n30022,
         n30023, n30024, n30025, n30026, n30027, n30028, n30029, n30030,
         n30031, n30032, n30033, n30034, n30035, n30036, n30037, n30038,
         n30039, n30040, n30041, n30042, n30043, n30044, n30045, n30046,
         n30047, n30048, n30049, n30050, n30051, n30052, n30053, n30054,
         n30055, n30056, n30057, n30058, n30059, n30060, n30061, n30062,
         n30063, n30064, n30065, n30066, n30067, n30068, n30069, n30070,
         n30071, n30072, n30073, n30074, n30075, n30076, n30077, n30078,
         n30079, n30080, n30081, n30082, n30083, n30084, n30085, n30086,
         n30087, n30088, n30089, n30090, n30091, n30092, n30093, n30094,
         n30095, n30096, n30097, n30098, n30099, n30100, n30101, n30102,
         n30103, n30104, n30105, n30106, n30107, n30108, n30109, n30110,
         n30111, n30112, n30113, n30114, n30115, n30116, n30117, n30118,
         n30119, n30120, n30121, n30122, n30123, n30124, n30125, n30126,
         n30127, n30128, n30129, n30130, n30131, n30132, n30133, n30134,
         n30135, n30136, n30137, n30138, n30139, n30140, n30141, n30142,
         n30143, n30144, n30145, n30146, n30147, n30148, n30149, n30150,
         n30151, n30152, n30153, n30154, n30155, n30156, n30157, n30158,
         n30159, n30160, n30161, n30162, n30163, n30164, n30165, n30166,
         n30167, n30168, n30169, n30170, n30171, n30172, n30173, n30174,
         n30175, n30176, n30177, n30178, n30179, n30180, n30181, n30182,
         n30183, n30184, n30185, n30186, n30187, n30188, n30189, n30190,
         n30191, n30192, n30193, n30194, n30195, n30196, n30197, n30198,
         n30199, n30200, n30201, n30202, n30203, n30204, n30205, n30206,
         n30207, n30208, n30209, n30210, n30211, n30212, n30213, n30214,
         n30215, n30216, n30217, n30218, n30219, n30220, n30221, n30222,
         n30223, n30224, n30225, n30226, n30227, n30228, n30229, n30230,
         n30231, n30232, n30233, n30234, n30235, n30236, n30237, n30238,
         n30239, n30240, n30241, n30242, n30243, n30244, n30245, n30246,
         n30247, n30248, n30249, n30250, n30251, n30252, n30253, n30254,
         n30255, n30256, n30257, n30258, n30259, n30260, n30261, n30262,
         n30263, n30264, n30265, n30266, n30267, n30268, n30269, n30270,
         n30271, n30272, n30273, n30274, n30275, n30276, n30277, n30278,
         n30279, n30280, n30281, n30282, n30283, n30284, n30285, n30286,
         n30287, n30288, n30289, n30290, n30291, n30292, n30293, n30294,
         n30295, n30296, n30297, n30298, n30299, n30300, n30301, n30302,
         n30303, n30304, n30305, n30306, n30307, n30308, n30309, n30310,
         n30311, n30312, n30313, n30314, n30315, n30316, n30317, n30318,
         n30319, n30320, n30321, n30322, n30323, n30324, n30325, n30326,
         n30327, n30328, n30329, n30330, n30331, n30332, n30333, n30334,
         n30335, n30336, n30337, n30338, n30339, n30340, n30341, n30342,
         n30343, n30344, n30345, n30346, n30347, n30348, n30349, n30350,
         n30351, n30352, n30353, n30354, n30355, n30356, n30357, n30358,
         n30359, n30360, n30361, n30362, n30363, n30364, n30365, n30366,
         n30367, n30368, n30369, n30370, n30371, n30372, n30373, n30374,
         n30375, n30376, n30377, n30378, n30379, n30380, n30381, n30382,
         n30383, n30384, n30385, n30386, n30387, n30388, n30389, n30390,
         n30391, n30392, n30393, n30394, n30395, n30396, n30397, n30398,
         n30399, n30400, n30401, n30402, n30403, n30404, n30405, n30406,
         n30407, n30408, n30409, n30410, n30411, n30412, n30413, n30414,
         n30415, n30416, n30417, n30418, n30419, n30420, n30421, n30422,
         n30423, n30424, n30425, n30426, n30427, n30428, n30429, n30430,
         n30431, n30432, n30433, n30434, n30435, n30436, n30437, n30438,
         n30439, n30440, n30441, n30442, n30443, n30444, n30445, n30446,
         n30447, n30448, n30449, n30450, n30451, n30452, n30453, n30454,
         n30455, n30456, n30457, n30458, n30459, n30460, n30461, n30462,
         n30463, n30464, n30465, n30466, n30467, n30468, n30469, n30470,
         n30471, n30472, n30473, n30474, n30475, n30476, n30477, n30478,
         n30479, n30480, n30481, n30482, n30483, n30484, n30485, n30486,
         n30487, n30488, n30489, n30490, n30491, n30492, n30493, n30494,
         n30495, n30496, n30497, n30498, n30499, n30500, n30501, n30502,
         n30503, n30504, n30505, n30506, n30507, n30508, n30509, n30510,
         n30511, n30512, n30513, n30514, n30515, n30516, n30517, n30518,
         n30519, n30520, n30521, n30522, n30523, n30524, n30525, n30526,
         n30527, n30528, n30529, n30530, n30531, n30532, n30533, n30534,
         n30535, n30536, n30537, n30538, n30539, n30540, n30541, n30542,
         n30543, n30544, n30545, n30546, n30547, n30548, n30549, n30550,
         n30551, n30552, n30553, n30554, n30555, n30556, n30557, n30558,
         n30559, n30560, n30561, n30562, n30563, n30564, n30565, n30566,
         n30567, n30568, n30569, n30570, n30571, n30572, n30573, n30574,
         n30575, n30576, n30577, n30578, n30579, n30580, n30581, n30582,
         n30583, n30584, n30585, n30586, n30587, n30588, n30589, n30590,
         n30591, n30592, n30593, n30594, n30595, n30596, n30597, n30598,
         n30599, n30600, n30601, n30602, n30603, n30604, n30605, n30606,
         n30607, n30608, n30609, n30610, n30611, n30612, n30613, n30614,
         n30615, n30616, n30617, n30618, n30619, n30620, n30621, n30622,
         n30623, n30624, n30625, n30626, n30627, n30628, n30629, n30630,
         n30631, n30632, n30633, n30634, n30635, n30636, n30637, n30638,
         n30639, n30640, n30641, n30642, n30643, n30644, n30645, n30646,
         n30647, n30648, n30649, n30650, n30651, n30652, n30653, n30654,
         n30655, n30656, n30657, n30658, n30659, n30660, n30661, n30662,
         n30663, n30664, n30665, n30666, n30667, n30668, n30669, n30670,
         n30671, n30672, n30673, n30674, n30675, n30676, n30677, n30678,
         n30679, n30680, n30681, n30682, n30683, n30684, n30685, n30686,
         n30687, n30688, n30689, n30690, n30691, n30692, n30693, n30694,
         n30695, n30696, n30697, n30698, n30699, n30700, n30701, n30702,
         n30703, n30704, n30705, n30706, n30707, n30708, n30709, n30710,
         n30711, n30712, n30713, n30714, n30715, n30716, n30717, n30718,
         n30719, n30720, n30721, n30722, n30723, n30724, n30725, n30726,
         n30727, n30728, n30729, n30730, n30731, n30732, n30733, n30734,
         n30735, n30736, n30737, n30738, n30739, n30740, n30741, n30742,
         n30743, n30744, n30745, n30746, n30747, n30748, n30749, n30750,
         n30751, n30752, n30753, n30754, n30755, n30756, n30757, n30758,
         n30759, n30760, n30761, n30762, n30763, n30764, n30765, n30766,
         n30767, n30768, n30769, n30770, n30771, n30772, n30773, n30774,
         n30775, n30776, n30777, n30778, n30779, n30780, n30781, n30782,
         n30783, n30784, n30785, n30786, n30787, n30788, n30789, n30790,
         n30791, n30792, n30793, n30794, n30795, n30796, n30797, n30798,
         n30799, n30800, n30801, n30802, n30803, n30804, n30805, n30806,
         n30807, n30808, n30809, n30810, n30811, n30812, n30813, n30814,
         n30815, n30816, n30817, n30818, n30819, n30820, n30821, n30822,
         n30823, n30824, n30825, n30826, n30827, n30828, n30829, n30830,
         n30831, n30832, n30833, n30834, n30835, n30836, n30837, n30838,
         n30839, n30840, n30841, n30842, n30843, n30844, n30845, n30846,
         n30847, n30848, n30849, n30850, n30851, n30852, n30853, n30854,
         n30855, n30856, n30857, n30858, n30859, n30860, n30861, n30862,
         n30863, n30864, n30865, n30866, n30867, n30868, n30869, n30870,
         n30871, n30872, n30873, n30874, n30875, n30876, n30877, n30878,
         n30879, n30880, n30881, n30882, n30883, n30884, n30885, n30886,
         n30887, n30888, n30889, n30890, n30891, n30892, n30893, n30894,
         n30895, n30896, n30897, n30898, n30899, n30900, n30901, n30902,
         n30903, n30904, n30905, n30906, n30907, n30908, n30909, n30910,
         n30911, n30912, n30913, n30914, n30915, n30916, n30917, n30918,
         n30919, n30920, n30921, n30922, n30923, n30924, n30925, n30926,
         n30927, n30928, n30929, n30930, n30931, n30932, n30933, n30934,
         n30935, n30936, n30937, n30938, n30939, n30940, n30941, n30942,
         n30943, n30944, n30945, n30946, n30947, n30948, n30949, n30950,
         n30951, n30952, n30953, n30954, n30955, n30956, n30957, n30958,
         n30959, n30960, n30961, n30962, n30963, n30964, n30965, n30966,
         n30967, n30968, n30969, n30970, n30971, n30972, n30973, n30974,
         n30975, n30976, n30977, n30978, n30979, n30980, n30981, n30982,
         n30983, n30984, n30985, n30986, n30987, n30988, n30989, n30990,
         n30991, n30992, n30993, n30994, n30995, n30996, n30997, n30998,
         n30999, n31000, n31001, n31002, n31003, n31004, n31005, n31006,
         n31007, n31008, n31009, n31010, n31011, n31012, n31013, n31014,
         n31015, n31016, n31017, n31018, n31019, n31020, n31021, n31022,
         n31023, n31024, n31025, n31026, n31027, n31028, n31029, n31030,
         n31031, n31032, n31033, n31034, n31035, n31036, n31037, n31038,
         n31039, n31040, n31041, n31042, n31043, n31044, n31045, n31046,
         n31047, n31048, n31049, n31050, n31051, n31052, n31053, n31054,
         n31055, n31056, n31057, n31058, n31059, n31060, n31061, n31062,
         n31063, n31064, n31065, n31066, n31067, n31068, n31069, n31070,
         n31071, n31072, n31073, n31074, n31075, n31076, n31077, n31078,
         n31079, n31080, n31081, n31082, n31083, n31084, n31085, n31086,
         n31087, n31088, n31089, n31090, n31091, n31092, n31093, n31094,
         n31095, n31096, n31097, n31098, n31099, n31100, n31101, n31102,
         n31103, n31104, n31105, n31106, n31107, n31108, n31109, n31110,
         n31111, n31112, n31113, n31114, n31115, n31116, n31117, n31118,
         n31119, n31120, n31121, n31122, n31123, n31124, n31125, n31126,
         n31127, n31128, n31129, n31130, n31131, n31132, n31133, n31134,
         n31135, n31136, n31137, n31138, n31139, n31140, n31141, n31142,
         n31143, n31144, n31145, n31146, n31147, n31148, n31149, n31150,
         n31151, n31152, n31153, n31154, n31155, n31156, n31157, n31158,
         n31159, n31160, n31161, n31162, n31163, n31164, n31165, n31166,
         n31167, n31168, n31169, n31170, n31171, n31172, n31173, n31174,
         n31175, n31176, n31177, n31178, n31179, n31180, n31181, n31182,
         n31183, n31184, n31185, n31186, n31187, n31188, n31189, n31190,
         n31191, n31192, n31193, n31194, n31195, n31196, n31197, n31198,
         n31199, n31200, n31201, n31202, n31203, n31204, n31205, n31206,
         n31207, n31208, n31209, n31210, n31211, n31212, n31213, n31214,
         n31215, n31216, n31217, n31218, n31219, n31220, n31221, n31222,
         n31223, n31224, n31225, n31226, n31227, n31228, n31229, n31230,
         n31231, n31232, n31233, n31234, n31235, n31236, n31237, n31238,
         n31239, n31240, n31241, n31242, n31243, n31244, n31245, n31246,
         n31247, n31248, n31249, n31250, n31251, n31252, n31253, n31254,
         n31255, n31256, n31257, n31258, n31259, n31260, n31261, n31262,
         n31263, n31264, n31265, n31266, n31267, n31268, n31269, n31270,
         n31271, n31272, n31273, n31274, n31275, n31276, n31277, n31278,
         n31279, n31280, n31281, n31282, n31283, n31284, n31285, n31286,
         n31287, n31288, n31289, n31290, n31291, n31292, n31293, n31294,
         n31295, n31296, n31297, n31298, n31299, n31300, n31301, n31302,
         n31303, n31304, n31305, n31306, n31307, n31308, n31309, n31310,
         n31311, n31312, n31313, n31314, n31315, n31316, n31317, n31318,
         n31319, n31320, n31321, n31322, n31323, n31324, n31325, n31326,
         n31327, n31328, n31329, n31330, n31331, n31332, n31333, n31334,
         n31335, n31336, n31337, n31338, n31339, n31340, n31341, n31342,
         n31343, n31344, n31345, n31346, n31347, n31348, n31349, n31350,
         n31351, n31352, n31353, n31354, n31355, n31356, n31357, n31358,
         n31359, n31360, n31361, n31362, n31363, n31364, n31365, n31366,
         n31367, n31368, n31369, n31370, n31371, n31372, n31373, n31374,
         n31375, n31376, n31377, n31378, n31379, n31380, n31381, n31382,
         n31383, n31384, n31385, n31386, n31387, n31388, n31389, n31390,
         n31391, n31392, n31393, n31394, n31395, n31396, n31397, n31398,
         n31399, n31400, n31401, n31402, n31403, n31404, n31405, n31406,
         n31407, n31408, n31409, n31410, n31411, n31412, n31413, n31414,
         n31415, n31416, n31417, n31418, n31419, n31420, n31421, n31422,
         n31423, n31424, n31425, n31426, n31427, n31428, n31429, n31430,
         n31431, n31432, n31433, n31434, n31435, n31436, n31437, n31438,
         n31439, n31440, n31441, n31442, n31443, n31444, n31445, n31446,
         n31447, n31448, n31449, n31450, n31451, n31452, n31453, n31454,
         n31455, n31456, n31457, n31458, n31459, n31460, n31461, n31462,
         n31463, n31464, n31465, n31466, n31467, n31468, n31469, n31470,
         n31471, n31472, n31473, n31474, n31475, n31476, n31477, n31478,
         n31479, n31480, n31481, n31482, n31483, n31484, n31485, n31486,
         n31487, n31488, n31489, n31490, n31491, n31492, n31493, n31494,
         n31495, n31496, n31497, n31498, n31499, n31500, n31501, n31502,
         n31503, n31504, n31505, n31506, n31507, n31508, n31509, n31510,
         n31511, n31512, n31513, n31514, n31515, n31516, n31517, n31518,
         n31519, n31520, n31521, n31522, n31523, n31524, n31525, n31526,
         n31527, n31528, n31529, n31530, n31531, n31532, n31533, n31534,
         n31535, n31536, n31537, n31538, n31539, n31540, n31541, n31542,
         n31543, n31544, n31545, n31546, n31547, n31548, n31549, n31550,
         n31551, n31552, n31553, n31554, n31555, n31556, n31557, n31558,
         n31559, n31560, n31561, n31562, n31563, n31564, n31565, n31566,
         n31567, n31568, n31569, n31570, n31571, n31572, n31573, n31574,
         n31575, n31576, n31577, n31578, n31579, n31580, n31581, n31582,
         n31583, n31584, n31585, n31586, n31587, n31588, n31589, n31590,
         n31591, n31592, n31593, n31594, n31595, n31596, n31597, n31598,
         n31599, n31600, n31601, n31602, n31603, n31604, n31605, n31606,
         n31607, n31608, n31609, n31610, n31611, n31612, n31613, n31614,
         n31615, n31616, n31617, n31618, n31619, n31620, n31621, n31622,
         n31623, n31624, n31625, n31626, n31627, n31628, n31629, n31630,
         n31631, n31632, n31633, n31634, n31635, n31636, n31637, n31638,
         n31639, n31640, n31641, n31642, n31643, n31644, n31645, n31646,
         n31647, n31648, n31649, n31650, n31651, n31652, n31653, n31654,
         n31655, n31656, n31657, n31658, n31659, n31660, n31661, n31662,
         n31663, n31664, n31665, n31666, n31667, n31668, n31669, n31670,
         n31671, n31672, n31673, n31674, n31675, n31676, n31677, n31678,
         n31679, n31680, n31681, n31682, n31683, n31684, n31685, n31686,
         n31687, n31688, n31689, n31690, n31691, n31692, n31693, n31694,
         n31695, n31696, n31697, n31698, n31699, n31700, n31701, n31702,
         n31703, n31704, n31705, n31706, n31707, n31708, n31709, n31710,
         n31711, n31712, n31713, n31714, n31715, n31716, n31717, n31718,
         n31719, n31720, n31721, n31722, n31723, n31724, n31725, n31726,
         n31727, n31728, n31729, n31730, n31731, n31732, n31733, n31734,
         n31735, n31736, n31737, n31738, n31739, n31740, n31741, n31742,
         n31743, n31744, n31745, n31746, n31747, n31748, n31749, n31750,
         n31751, n31752, n31753, n31754, n31755, n31756, n31757, n31758,
         n31759, n31760, n31761, n31762, n31763, n31764, n31765, n31766,
         n31767, n31768, n31769, n31770, n31771, n31772, n31773, n31774,
         n31775, n31776, n31777, n31778, n31779, n31780, n31781, n31782,
         n31783, n31784, n31785, n31786, n31787, n31788, n31789, n31790,
         n31791, n31792, n31793, n31794, n31795, n31796, n31797, n31798,
         n31799, n31800, n31801, n31802, n31803, n31804, n31805, n31806,
         n31807, n31808, n31809, n31810, n31811, n31812, n31813, n31814,
         n31815, n31816, n31817, n31818, n31819, n31820, n31821, n31822,
         n31823, n31824, n31825, n31826, n31827, n31828, n31829, n31830,
         n31831, n31832, n31833, n31834, n31835, n31836, n31837, n31838,
         n31839, n31840, n31841, n31842, n31843, n31844, n31845, n31846,
         n31847, n31848, n31849, n31850, n31851, n31852, n31853, n31854,
         n31855, n31856, n31857, n31858, n31859, n31860, n31861, n31862,
         n31863, n31864, n31865, n31866, n31867, n31868, n31869, n31870,
         n31871, n31872, n31873, n31874, n31875, n31876, n31877, n31878,
         n31879, n31880, n31881, n31882, n31883, n31884, n31885, n31886,
         n31887, n31888, n31889, n31890, n31891, n31892, n31893, n31894,
         n31895, n31896, n31897, n31898, n31899, n31900, n31901, n31902,
         n31903, n31904, n31905, n31906, n31907, n31908, n31909, n31910,
         n31911, n31912, n31913, n31914, n31915, n31916, n31917, n31918,
         n31919, n31920, n31921, n31922, n31923, n31924, n31925, n31926,
         n31927, n31928, n31929, n31930, n31931, n31932, n31933, n31934,
         n31935, n31936, n31937, n31938, n31939, n31940, n31941, n31942,
         n31943, n31944, n31945, n31946, n31947, n31948, n31949, n31950,
         n31951, n31952, n31953, n31954, n31955, n31956, n31957, n31958,
         n31959, n31960, n31961, n31962, n31963, n31964, n31965, n31966,
         n31967, n31968, n31969, n31970, n31971, n31972, n31973, n31974,
         n31975, n31976, n31977, n31978, n31979, n31980, n31981, n31982,
         n31983, n31984, n31985, n31986, n31987, n31988, n31989, n31990,
         n31991, n31992, n31993, n31994, n31995, n31996, n31997, n31998,
         n31999, n32000, n32001, n32002, n32003, n32004, n32005, n32006,
         n32007, n32008, n32009, n32010, n32011, n32012, n32013, n32014,
         n32015, n32016, n32017, n32018, n32019, n32020, n32021, n32022,
         n32023, n32024, n32025, n32026, n32027, n32028, n32029, n32030,
         n32031, n32032, n32033, n32034, n32035, n32036, n32037, n32038,
         n32039, n32040, n32041, n32042, n32043, n32044, n32045, n32046,
         n32047, n32048, n32049, n32050, n32051, n32052, n32053, n32054,
         n32055, n32056, n32057, n32058, n32059, n32060, n32061, n32062,
         n32063, n32064, n32065, n32066, n32067, n32068, n32069, n32070,
         n32071, n32072, n32073, n32074, n32075, n32076, n32077, n32078,
         n32079, n32080, n32081, n32082, n32083, n32084, n32085, n32086,
         n32087, n32088, n32089, n32090, n32091, n32092, n32093, n32094,
         n32095, n32096, n32097, n32098, n32099, n32100, n32101, n32102,
         n32103, n32104, n32105, n32106, n32107, n32108, n32109, n32110,
         n32111, n32112, n32113, n32114, n32115, n32116, n32117, n32118,
         n32119, n32120, n32121, n32122, n32123, n32124, n32125, n32126,
         n32127, n32128, n32129, n32130, n32131, n32132, n32133, n32134,
         n32135, n32136, n32137, n32138, n32139, n32140, n32141, n32142,
         n32143, n32144, n32145, n32146, n32147, n32148, n32149, n32150,
         n32151, n32152, n32153, n32154, n32155, n32156, n32157, n32158,
         n32159, n32160, n32161, n32162, n32163, n32164, n32165, n32166,
         n32167, n32168, n32169, n32170, n32171, n32172, n32173, n32174,
         n32175, n32176, n32177, n32178, n32179, n32180, n32181, n32182,
         n32183, n32184, n32185, n32186, n32187, n32188, n32189, n32190,
         n32191, n32192, n32193, n32194, n32195, n32196, n32197, n32198,
         n32199, n32200, n32201, n32202, n32203, n32204, n32205, n32206,
         n32207, n32208, n32209, n32210, n32211, n32212, n32213, n32214,
         n32215, n32216, n32217, n32218, n32219, n32220, n32221, n32222,
         n32223, n32224, n32225, n32226, n32227, n32228, n32229, n32230,
         n32231, n32232, n32233, n32234, n32235, n32236, n32237, n32238,
         n32239, n32240, n32241, n32242, n32243, n32244, n32245, n32246,
         n32247, n32248, n32249, n32250, n32251, n32252, n32253, n32254,
         n32255, n32256, n32257, n32258, n32259, n32260, n32261, n32262,
         n32263, n32264, n32265, n32266, n32267, n32268, n32269, n32270,
         n32271, n32272, n32273, n32274, n32275, n32276, n32277, n32278,
         n32279, n32280, n32281, n32282, n32283, n32284, n32285, n32286,
         n32287, n32288, n32289, n32290, n32291, n32292, n32293, n32294,
         n32295, n32296, n32297, n32298, n32299, n32300, n32301, n32302,
         n32303, n32304, n32305, n32306, n32307, n32308, n32309, n32310,
         n32311, n32312, n32313, n32314, n32315, n32316, n32317, n32318,
         n32319, n32320, n32321, n32322, n32323, n32324, n32325, n32326,
         n32327, n32328, n32329, n32330, n32331, n32332, n32333, n32334,
         n32335, n32336, n32337, n32338, n32339, n32340, n32341, n32342,
         n32343, n32344, n32345, n32346, n32347, n32348, n32349, n32350,
         n32351, n32352, n32353, n32354, n32355, n32356, n32357, n32358,
         n32359, n32360, n32361, n32362, n32363, n32364, n32365, n32366,
         n32367, n32368, n32369, n32370, n32371, n32372, n32373, n32374,
         n32375, n32376, n32377, n32378, n32379, n32380, n32381, n32382,
         n32383, n32384, n32385, n32386, n32387, n32388, n32389, n32390,
         n32391, n32392, n32393, n32394, n32395, n32396, n32397, n32398,
         n32399, n32400, n32401, n32402, n32403, n32404, n32405, n32406,
         n32407, n32408, n32409, n32410, n32411, n32412, n32413, n32414,
         n32415, n32416, n32417, n32418, n32419, n32420, n32421, n32422,
         n32423, n32424, n32425, n32426, n32427, n32428, n32429, n32430,
         n32431, n32432, n32433, n32434, n32435, n32436, n32437, n32438,
         n32439, n32440, n32441, n32442, n32443, n32444, n32445, n32446,
         n32447, n32448, n32449, n32450, n32451, n32452, n32453, n32454,
         n32455, n32456, n32457, n32458, n32459, n32460, n32461, n32462,
         n32463, n32464, n32465, n32466, n32467, n32468, n32469, n32470,
         n32471, n32472, n32473, n32474, n32475, n32476, n32477, n32478,
         n32479, n32480, n32481, n32482, n32483, n32484, n32485, n32486,
         n32487, n32488, n32489, n32490, n32491, n32492, n32493, n32494,
         n32495, n32496, n32497, n32498, n32499, n32500, n32501, n32502,
         n32503, n32504, n32505, n32506, n32507, n32508, n32509, n32510,
         n32511, n32512, n32513, n32514, n32515, n32516, n32517, n32518,
         n32519, n32520, n32521, n32522, n32523, n32524, n32525, n32526,
         n32527, n32528, n32529, n32530, n32531, n32532, n32533, n32534,
         n32535, n32536, n32537, n32538, n32539, n32540, n32541, n32542,
         n32543, n32544, n32545, n32546, n32547, n32548, n32549, n32550,
         n32551, n32552, n32553, n32554, n32555, n32556, n32557, n32558,
         n32559, n32560, n32561, n32562, n32563, n32564, n32565, n32566,
         n32567, n32568, n32569, n32570, n32571, n32572, n32573, n32574,
         n32575, n32576, n32577, n32578, n32579, n32580, n32581, n32582,
         n32583, n32584, n32585, n32586, n32587, n32588, n32589, n32590,
         n32591, n32592, n32593, n32594, n32595, n32596, n32597, n32598,
         n32599, n32600, n32601, n32602, n32603, n32604, n32605, n32606,
         n32607, n32608, n32609, n32610, n32611, n32612, n32613, n32614,
         n32615, n32616, n32617, n32618, n32619, n32620, n32621, n32622,
         n32623, n32624, n32625, n32626, n32627, n32628, n32629, n32630,
         n32631, n32632, n32633, n32634, n32635, n32636, n32637, n32638,
         n32639, n32640, n32641, n32642, n32643, n32644, n32645, n32646,
         n32647, n32648, n32649, n32650, n32651, n32652, n32653, n32654,
         n32655, n32656, n32657, n32658, n32659, n32660, n32661, n32662,
         n32663, n32664, n32665, n32666, n32667, n32668, n32669, n32670,
         n32671, n32672, n32673, n32674, n32675, n32676, n32677, n32678,
         n32679, n32680, n32681, n32682, n32683, n32684, n32685, n32686,
         n32687, n32688, n32689, n32690, n32691, n32692, n32693, n32694,
         n32695, n32696, n32697, n32698, n32699, n32700, n32701, n32702,
         n32703, n32704, n32705, n32706, n32707, n32708, n32709, n32710,
         n32711, n32712, n32713, n32714, n32715, n32716, n32717, n32718,
         n32719, n32720, n32721, n32722, n32723, n32724, n32725, n32726,
         n32727, n32728, n32729, n32730, n32731, n32732, n32733, n32734,
         n32735, n32736, n32737, n32738, n32739, n32740, n32741, n32742,
         n32743, n32744, n32745, n32746, n32747, n32748, n32749, n32750,
         n32751, n32752, n32753, n32754, n32755, n32756, n32757, n32758,
         n32759, n32760, n32761, n32762, n32763, n32764, n32765, n32766,
         n32767, n32768, n32769, n32770, n32771, n32772, n32773, n32774,
         n32775, n32776, n32777, n32778, n32779, n32780, n32781, n32782,
         n32783, n32784, n32785, n32786, n32787, n32788, n32789, n32790,
         n32791, n32792, n32793, n32794, n32795, n32796, n32797, n32798,
         n32799, n32800, n32801, n32802, n32803, n32804, n32805, n32806,
         n32807, n32808, n32809, n32810, n32811, n32812, n32813, n32814,
         n32815, n32816, n32817, n32818, n32819, n32820, n32821, n32822,
         n32823, n32824, n32825, n32826, n32827, n32828, n32829, n32830,
         n32831, n32832, n32833, n32834, n32835, n32836, n32837, n32838,
         n32839, n32840, n32841, n32842, n32843, n32844, n32845, n32846,
         n32847, n32848, n32849, n32850, n32851, n32852, n32853, n32854,
         n32855, n32856, n32857, n32858, n32859, n32860, n32861, n32862,
         n32863, n32864, n32865, n32866, n32867, n32868, n32869, n32870,
         n32871, n32872, n32873, n32874, n32875, n32876, n32877, n32878,
         n32879, n32880, n32881, n32882, n32883, n32884, n32885, n32886,
         n32887, n32888, n32889, n32890, n32891, n32892, n32893, n32894,
         n32895, n32896, n32897, n32898, n32899, n32900, n32901, n32902,
         n32903, n32904, n32905, n32906, n32907, n32908, n32909, n32910,
         n32911, n32912, n32913, n32914, n32915, n32916, n32917, n32918,
         n32919, n32920, n32921, n32922, n32923, n32924, n32925, n32926,
         n32927, n32928, n32929, n32930, n32931, n32932, n32933, n32934,
         n32935, n32936, n32937, n32938, n32939, n32940, n32941, n32942,
         n32943, n32944, n32945, n32946, n32947, n32948, n32949, n32950,
         n32951, n32952, n32953, n32954, n32955, n32956, n32957, n32958,
         n32959, n32960, n32961, n32962, n32963, n32964, n32965, n32966,
         n32967, n32968, n32969, n32970, n32971, n32972, n32973, n32974,
         n32975, n32976, n32977, n32978, n32979, n32980, n32981, n32982,
         n32983, n32984, n32985, n32986, n32987, n32988, n32989, n32990,
         n32991, n32992, n32993, n32994, n32995, n32996, n32997, n32998,
         n32999, n33000, n33001, n33002, n33003, n33004, n33005, n33006,
         n33007, n33008, n33009, n33010, n33011, n33012, n33013, n33014,
         n33015, n33016, n33017, n33018, n33019, n33020, n33021, n33022,
         n33023, n33024, n33025, n33026, n33027, n33028, n33029, n33030,
         n33031, n33032, n33033, n33034, n33035, n33036, n33037, n33038,
         n33039, n33040, n33041, n33042, n33043, n33044, n33045, n33046,
         n33047, n33048, n33049, n33050, n33051, n33052, n33053, n33054,
         n33055, n33056, n33057, n33058, n33059, n33060, n33061, n33062,
         n33063, n33064, n33065, n33066, n33067, n33068, n33069, n33070,
         n33071, n33072, n33073, n33074, n33075, n33076, n33077, n33078,
         n33079, n33080, n33081, n33082, n33083, n33084, n33085, n33086,
         n33087, n33088, n33089, n33090, n33091, n33092, n33093, n33094,
         n33095, n33096, n33097, n33098, n33099, n33100, n33101, n33102,
         n33103, n33104, n33105, n33106, n33107, n33108, n33109, n33110,
         n33111, n33112, n33113, n33114, n33115, n33116, n33117, n33118,
         n33119, n33120, n33121, n33122, n33123, n33124, n33125, n33126,
         n33127, n33128, n33129, n33130, n33131, n33132, n33133, n33134,
         n33135, n33136, n33137, n33138, n33139, n33140, n33141, n33142,
         n33143, n33144, n33145, n33146, n33147, n33148, n33149, n33150,
         n33151, n33152, n33153, n33154, n33155, n33156, n33157, n33158,
         n33159, n33160, n33161, n33162, n33163, n33164, n33165, n33166,
         n33167, n33168, n33169, n33170, n33171, n33172, n33173, n33174,
         n33175, n33176, n33177, n33178, n33179, n33180, n33181, n33182,
         n33183, n33184, n33185, n33186, n33187, n33188, n33189, n33190,
         n33191, n33192, n33193, n33194, n33195, n33196, n33197, n33198,
         n33199, n33200, n33201, n33202, n33203, n33204, n33205, n33206,
         n33207, n33208, n33209, n33210, n33211, n33212, n33213, n33214,
         n33215, n33216, n33217, n33218, n33219, n33220, n33221, n33222,
         n33223, n33224, n33225, n33226, n33227, n33228, n33229, n33230,
         n33231, n33232, n33233, n33234, n33235, n33236, n33237, n33238,
         n33239, n33240, n33241, n33242, n33243, n33244, n33245, n33246,
         n33247, n33248, n33249, n33250, n33251, n33252, n33253, n33254,
         n33255, n33256, n33257, n33258, n33259, n33260, n33261, n33262,
         n33263, n33264, n33265, n33266, n33267, n33268, n33269, n33270,
         n33271, n33272, n33273, n33274, n33275, n33276, n33277, n33278,
         n33279, n33280, n33281, n33282, n33283, n33284, n33285, n33286,
         n33287, n33288, n33289, n33290, n33291, n33292, n33293, n33294,
         n33295, n33296, n33297, n33298, n33299, n33300, n33301, n33302,
         n33303, n33304, n33305, n33306, n33307, n33308, n33309, n33310,
         n33311, n33312, n33313, n33314, n33315, n33316, n33317, n33318,
         n33319, n33320, n33321, n33322, n33323, n33324, n33325, n33326,
         n33327, n33328, n33329, n33330, n33331, n33332, n33333, n33334,
         n33335, n33336, n33337, n33338, n33339, n33340, n33341, n33342,
         n33343, n33344, n33345, n33346, n33347, n33348, n33349, n33350,
         n33351, n33352, n33353, n33354, n33355, n33356, n33357, n33358,
         n33359, n33360, n33361, n33362, n33363, n33364, n33365, n33366,
         n33367, n33368, n33369, n33370, n33371, n33372, n33373, n33374,
         n33375, n33376, n33377, n33378, n33379, n33380, n33381, n33382,
         n33383, n33384, n33385, n33386, n33387, n33388, n33389, n33390,
         n33391, n33392, n33393, n33394, n33395, n33396, n33397, n33398,
         n33399, n33400, n33401, n33402, n33403, n33404, n33405, n33406,
         n33407, n33408, n33409, n33410, n33411, n33412, n33413, n33414,
         n33415, n33416, n33417, n33418, n33419, n33420, n33421, n33422,
         n33423, n33424, n33425, n33426, n33427, n33428, n33429, n33430,
         n33431, n33432, n33433, n33434, n33435, n33436, n33437, n33438,
         n33439, n33440, n33441, n33442, n33443, n33444, n33445, n33446,
         n33447, n33448, n33449, n33450, n33451, n33452, n33453, n33454,
         n33455, n33456, n33457, n33458, n33459, n33460, n33461, n33462,
         n33463, n33464, n33465, n33466, n33467, n33468, n33469, n33470,
         n33471, n33472, n33473, n33474, n33475, n33476, n33477, n33478,
         n33479, n33480, n33481, n33482, n33483, n33484, n33485, n33486,
         n33487, n33488, n33489, n33490, n33491, n33492, n33493, n33494,
         n33495, n33496, n33497, n33498, n33499, n33500, n33501, n33502,
         n33503, n33504, n33505, n33506, n33507, n33508, n33509, n33510,
         n33511, n33512, n33513, n33514, n33515, n33516, n33517, n33518,
         n33519, n33520, n33521, n33522, n33523, n33524, n33525, n33526,
         n33527, n33528, n33529, n33530, n33531, n33532, n33533, n33534,
         n33535, n33536, n33537, n33538, n33539, n33540, n33541, n33542,
         n33543, n33544, n33545, n33546, n33547, n33548, n33549, n33550,
         n33551, n33552, n33553, n33554, n33555, n33556, n33557, n33558,
         n33559, n33560, n33561, n33562, n33563, n33564, n33565, n33566,
         n33567, n33568, n33569, n33570, n33571, n33572, n33573, n33574,
         n33575, n33576, n33577, n33578, n33579, n33580, n33581, n33582,
         n33583, n33584, n33585, n33586, n33587, n33588, n33589, n33590,
         n33591, n33592, n33593, n33594, n33595, n33596, n33597, n33598,
         n33599, n33600, n33601, n33602, n33603, n33604, n33605, n33606,
         n33607, n33608, n33609, n33610, n33611, n33612, n33613, n33614,
         n33615, n33616, n33617, n33618, n33619, n33620, n33621, n33622,
         n33623, n33624, n33625, n33626, n33627, n33628, n33629, n33630,
         n33631, n33632, n33633, n33634, n33635, n33636, n33637, n33638,
         n33639, n33640, n33641, n33642, n33643, n33644, n33645, n33646,
         n33647, n33648, n33649, n33650, n33651, n33652, n33653, n33654,
         n33655, n33656, n33657, n33658, n33659, n33660, n33661, n33662,
         n33663, n33664, n33665, n33666, n33667, n33668, n33669, n33670,
         n33671, n33672, n33673, n33674, n33675, n33676, n33677, n33678,
         n33679, n33680, n33681, n33682, n33683, n33684, n33685, n33686,
         n33687, n33688, n33689, n33690, n33691, n33692, n33693, n33694,
         n33695, n33696, n33697, n33698, n33699, n33700, n33701, n33702,
         n33703, n33704, n33705, n33706, n33707, n33708, n33709, n33710,
         n33711, n33712, n33713, n33714, n33715, n33716, n33717, n33718,
         n33719, n33720, n33721, n33722, n33723, n33724, n33725, n33726,
         n33727, n33728, n33729, n33730, n33731, n33732, n33733, n33734,
         n33735, n33736, n33737, n33738, n33739, n33740, n33741, n33742,
         n33743, n33744, n33745, n33746, n33747, n33748, n33749, n33750,
         n33751, n33752, n33753, n33754, n33755, n33756, n33757, n33758,
         n33759, n33760, n33761, n33762, n33763, n33764, n33765, n33766,
         n33767, n33768, n33769, n33770, n33771, n33772, n33773, n33774,
         n33775, n33776, n33777, n33778, n33779, n33780, n33781, n33782,
         n33783, n33784, n33785, n33786, n33787, n33788, n33789, n33790,
         n33791, n33792, n33793, n33794, n33795, n33796, n33797, n33798,
         n33799, n33800, n33801, n33802, n33803, n33804, n33805, n33806,
         n33807, n33808, n33809, n33810, n33811, n33812, n33813, n33814,
         n33815, n33816, n33817, n33818, n33819, n33820, n33821, n33822,
         n33823, n33824, n33825, n33826, n33827, n33828, n33829, n33830,
         n33831, n33832, n33833, n33834, n33835, n33836, n33837, n33838,
         n33839, n33840, n33841, n33842, n33843, n33844, n33845, n33846,
         n33847, n33848, n33849, n33850, n33851, n33852, n33853, n33854,
         n33855, n33856, n33857, n33858, n33859, n33860, n33861, n33862,
         n33863, n33864, n33865, n33866, n33867, n33868, n33869, n33870,
         n33871, n33872, n33873, n33874, n33875, n33876, n33877, n33878,
         n33879, n33880, n33881, n33882, n33883, n33884, n33885, n33886,
         n33887, n33888, n33889, n33890, n33891, n33892, n33893, n33894,
         n33895, n33896, n33897, n33898, n33899, n33900, n33901, n33902,
         n33903, n33904, n33905, n33906, n33907, n33908, n33909, n33910,
         n33911, n33912, n33913, n33914, n33915, n33916, n33917, n33918,
         n33919, n33920, n33921, n33922, n33923, n33924, n33925, n33926,
         n33927, n33928, n33929, n33930, n33931, n33932, n33933, n33934,
         n33935, n33936, n33937, n33938, n33939, n33940, n33941, n33942,
         n33943, n33944, n33945, n33946, n33947, n33948, n33949, n33950,
         n33951, n33952, n33953, n33954, n33955, n33956, n33957, n33958,
         n33959, n33960, n33961, n33962, n33963, n33964, n33965, n33966,
         n33967, n33968, n33969, n33970, n33971, n33972, n33973, n33974,
         n33975, n33976, n33977, n33978, n33979, n33980, n33981, n33982,
         n33983, n33984, n33985, n33986, n33987, n33988, n33989, n33990,
         n33991, n33992, n33993, n33994, n33995, n33996, n33997, n33998,
         n33999, n34000, n34001, n34002, n34003, n34004, n34005, n34006,
         n34007, n34008, n34009, n34010, n34011, n34012, n34013, n34014,
         n34015, n34016, n34017, n34018, n34019, n34020, n34021, n34022,
         n34023, n34024, n34025, n34026, n34027, n34028, n34029, n34030,
         n34031, n34032, n34033, n34034, n34035, n34036, n34037, n34038,
         n34039, n34040, n34041, n34042, n34043, n34044, n34045, n34046,
         n34047, n34048, n34049, n34050, n34051, n34052, n34053, n34054,
         n34055, n34056, n34057, n34058, n34059, n34060, n34061, n34062,
         n34063, n34064, n34065, n34066, n34067, n34068, n34069, n34070,
         n34071, n34072, n34073, n34074, n34075, n34076, n34077, n34078,
         n34079, n34080, n34081, n34082, n34083, n34084, n34085, n34086,
         n34087, n34088, n34089, n34090, n34091, n34092, n34093, n34094,
         n34095, n34096, n34097, n34098, n34099, n34100, n34101, n34102,
         n34103, n34104, n34105, n34106, n34107, n34108, n34109, n34110,
         n34111, n34112, n34113, n34114, n34115, n34116, n34117, n34118,
         n34119, n34120, n34121, n34122, n34123, n34124, n34125, n34126,
         n34127, n34128, n34129, n34130, n34131, n34132, n34133, n34134,
         n34135, n34136, n34137, n34138, n34139, n34140, n34141, n34142,
         n34143, n34144, n34145, n34146, n34147, n34148, n34149, n34150,
         n34151, n34152, n34153, n34154, n34155, n34156, n34157, n34158,
         n34159, n34160, n34161, n34162, n34163, n34164, n34165, n34166,
         n34167, n34168, n34169, n34170, n34171, n34172, n34173, n34174,
         n34175, n34176, n34177, n34178, n34179, n34180, n34181, n34182,
         n34183, n34184, n34185, n34186, n34187, n34188, n34189, n34190,
         n34191, n34192, n34193, n34194, n34195, n34196, n34197, n34198,
         n34199, n34200, n34201, n34202, n34203, n34204, n34205, n34206,
         n34207, n34208, n34209, n34210, n34211, n34212, n34213, n34214,
         n34215, n34216, n34217, n34218, n34219, n34220, n34221, n34222,
         n34223, n34224, n34225, n34226, n34227, n34228, n34229, n34230,
         n34231, n34232, n34233, n34234, n34235, n34236, n34237, n34238,
         n34239, n34240, n34241, n34242, n34243, n34244, n34245, n34246,
         n34247, n34248, n34249, n34250, n34251, n34252, n34253, n34254,
         n34255, n34256, n34257, n34258, n34259, n34260, n34261, n34262,
         n34263, n34264, n34265, n34266, n34267, n34268, n34269, n34270,
         n34271, n34272, n34273, n34274, n34275, n34276, n34277, n34278,
         n34279, n34280, n34281, n34282, n34283, n34284, n34285, n34286,
         n34287, n34288, n34289, n34290, n34291, n34292, n34293, n34294,
         n34295, n34296, n34297, n34298, n34299, n34300, n34301, n34302,
         n34303, n34304, n34305, n34306, n34307, n34308, n34309, n34310,
         n34311, n34312, n34313, n34314, n34315, n34316, n34317, n34318,
         n34319, n34320, n34321, n34322, n34323, n34324, n34325, n34326,
         n34327, n34328, n34329, n34330, n34331, n34332, n34333, n34334,
         n34335, n34336, n34337, n34338, n34339, n34340, n34341, n34342,
         n34343, n34344, n34345, n34346, n34347, n34348, n34349, n34350,
         n34351, n34352, n34353, n34354, n34355, n34356, n34357, n34358,
         n34359, n34360, n34361, n34362, n34363, n34364, n34365, n34366,
         n34367, n34368, n34369, n34370, n34371, n34372, n34373, n34374,
         n34375, n34376, n34377, n34378, n34379, n34380, n34381, n34382,
         n34383, n34384, n34385, n34386, n34387, n34388, n34389, n34390,
         n34391, n34392, n34393, n34394, n34395, n34396, n34397, n34398,
         n34399, n34400, n34401, n34402, n34403, n34404, n34405, n34406,
         n34407, n34408, n34409, n34410, n34411, n34412, n34413, n34414,
         n34415, n34416, n34417, n34418, n34419, n34420, n34421, n34422,
         n34423, n34424, n34425, n34426, n34427, n34428, n34429, n34430,
         n34431, n34432, n34433, n34434, n34435, n34436, n34437, n34438,
         n34439, n34440, n34441, n34442, n34443, n34444, n34445, n34446,
         n34447, n34448, n34449, n34450, n34451, n34452, n34453, n34454,
         n34455, n34456, n34457, n34458, n34459, n34460, n34461, n34462,
         n34463, n34464, n34465, n34466, n34467, n34468, n34469, n34470,
         n34471, n34472, n34473, n34474, n34475, n34476, n34477, n34478,
         n34479, n34480, n34481, n34482, n34483, n34484, n34485, n34486,
         n34487, n34488, n34489, n34490, n34491, n34492, n34493, n34494,
         n34495, n34496, n34497, n34498, n34499, n34500, n34501, n34502,
         n34503, n34504, n34505, n34506, n34507, n34508, n34509, n34510,
         n34511, n34512, n34513, n34514, n34515, n34516, n34517, n34518,
         n34519, n34520, n34521, n34522, n34523, n34524, n34525, n34526,
         n34527, n34528, n34529, n34530, n34531, n34532, n34533, n34534,
         n34535, n34536, n34537, n34538, n34539, n34540, n34541, n34542,
         n34543, n34544, n34545, n34546, n34547, n34548, n34549, n34550,
         n34551, n34552, n34553, n34554, n34555, n34556, n34557, n34558,
         n34559, n34560, n34561, n34562, n34563, n34564, n34565, n34566,
         n34567, n34568, n34569, n34570, n34571, n34572, n34573, n34574,
         n34575, n34576, n34577, n34578, n34579, n34580, n34581, n34582,
         n34583, n34584, n34585, n34586, n34587, n34588, n34589, n34590,
         n34591, n34592, n34593, n34594, n34595, n34596, n34597, n34598,
         n34599, n34600, n34601, n34602, n34603, n34604, n34605, n34606,
         n34607, n34608, n34609, n34610, n34611, n34612, n34613, n34614,
         n34615, n34616, n34617, n34618, n34619, n34620, n34621, n34622,
         n34623, n34624, n34625, n34626, n34627, n34628, n34629, n34630,
         n34631, n34632, n34633, n34634, n34635, n34636, n34637, n34638,
         n34639, n34640, n34641, n34642, n34643, n34644, n34645, n34646,
         n34647, n34648, n34649, n34650, n34651, n34652, n34653, n34654,
         n34655, n34656, n34657, n34658, n34659, n34660, n34661, n34662,
         n34663, n34664, n34665, n34666, n34667, n34668, n34669, n34670,
         n34671, n34672, n34673, n34674, n34675, n34676, n34677, n34678,
         n34679, n34680, n34681, n34682, n34683, n34684, n34685, n34686,
         n34687, n34688, n34689, n34690, n34691, n34692, n34693, n34694,
         n34695, n34696, n34697, n34698, n34699, n34700, n34701, n34702,
         n34703, n34704, n34705, n34706, n34707, n34708, n34709, n34710,
         n34711, n34712, n34713, n34714, n34715, n34716, n34717, n34718,
         n34719, n34720, n34721, n34722, n34723, n34724, n34725, n34726,
         n34727, n34728, n34729, n34730, n34731, n34732, n34733, n34734,
         n34735, n34736, n34737, n34738, n34739, n34740, n34741, n34742,
         n34743, n34744, n34745, n34746, n34747, n34748, n34749, n34750,
         n34751, n34752, n34753, n34754, n34755, n34756, n34757, n34758,
         n34759, n34760, n34761, n34762, n34763, n34764, n34765, n34766,
         n34767, n34768, n34769, n34770, n34771, n34772, n34773, n34774,
         n34775, n34776, n34777, n34778, n34779, n34780, n34781, n34782,
         n34783, n34784, n34785, n34786, n34787, n34788, n34789, n34790,
         n34791, n34792, n34793, n34794, n34795, n34796, n34797, n34798,
         n34799, n34800, n34801, n34802, n34803, n34804, n34805, n34806,
         n34807, n34808, n34809, n34810, n34811, n34812, n34813, n34814,
         n34815, n34816, n34817, n34818, n34819, n34820, n34821, n34822,
         n34823, n34824, n34825, n34826, n34827, n34828, n34829, n34830,
         n34831, n34832, n34833, n34834, n34835, n34836, n34837, n34838,
         n34839, n34840, n34841, n34842, n34843, n34844, n34845, n34846,
         n34847, n34848, n34849, n34850, n34851, n34852, n34853, n34854,
         n34855, n34856, n34857, n34858, n34859, n34860, n34861, n34862,
         n34863, n34864, n34865, n34866, n34867, n34868, n34869, n34870,
         n34871, n34872, n34873, n34874, n34875, n34876, n34877, n34878,
         n34879, n34880, n34881, n34882, n34883, n34884, n34885, n34886,
         n34887, n34888, n34889, n34890, n34891, n34892, n34893, n34894,
         n34895, n34896, n34897, n34898, n34899, n34900, n34901, n34902,
         n34903, n34904, n34905, n34906, n34907, n34908, n34909, n34910,
         n34911, n34912, n34913, n34914, n34915, n34916, n34917, n34918,
         n34919, n34920, n34921, n34922, n34923, n34924, n34925, n34926,
         n34927, n34928, n34929, n34930, n34931, n34932, n34933, n34934,
         n34935, n34936, n34937, n34938, n34939, n34940, n34941, n34942,
         n34943, n34944, n34945, n34946, n34947, n34948, n34949, n34950,
         n34951, n34952, n34953, n34954, n34955, n34956, n34957, n34958,
         n34959, n34960, n34961, n34962, n34963, n34964, n34965, n34966,
         n34967, n34968, n34969, n34970, n34971, n34972, n34973, n34974,
         n34975, n34976, n34977, n34978, n34979, n34980, n34981, n34982,
         n34983, n34984, n34985, n34986, n34987, n34988, n34989, n34990,
         n34991, n34992, n34993, n34994, n34995, n34996, n34997, n34998,
         n34999, n35000, n35001, n35002, n35003, n35004, n35005, n35006,
         n35007, n35008, n35009, n35010, n35011, n35012, n35013, n35014,
         n35015, n35016, n35017, n35018, n35019, n35020, n35021, n35022,
         n35023, n35024, n35025, n35026, n35027, n35028, n35029, n35030,
         n35031, n35032, n35033, n35034, n35035, n35036, n35037, n35038,
         n35039, n35040, n35041, n35042, n35043, n35044, n35045, n35046,
         n35047, n35048, n35049, n35050, n35051, n35052, n35053, n35054,
         n35055, n35056, n35057, n35058, n35059, n35060, n35061, n35062,
         n35063, n35064, n35065, n35066, n35067, n35068, n35069, n35070,
         n35071, n35072, n35073, n35074, n35075, n35076, n35077, n35078,
         n35079, n35080, n35081, n35082, n35083, n35084, n35085, n35086,
         n35087, n35088, n35089, n35090, n35091, n35092, n35093, n35094,
         n35095, n35096, n35097, n35098, n35099, n35100, n35101, n35102,
         n35103, n35104, n35105, n35106, n35107, n35108, n35109, n35110,
         n35111, n35112, n35113, n35114, n35115, n35116, n35117, n35118,
         n35119, n35120, n35121, n35122, n35123, n35124, n35125, n35126,
         n35127, n35128, n35129, n35130, n35131, n35132, n35133, n35134,
         n35135, n35136, n35137, n35138, n35139, n35140, n35141, n35142,
         n35143, n35144, n35145, n35146, n35147, n35148, n35149, n35150,
         n35151, n35152, n35153, n35154, n35155, n35156, n35157, n35158,
         n35159, n35160, n35161, n35162, n35163, n35164, n35165, n35166,
         n35167, n35168, n35169, n35170, n35171, n35172, n35173, n35174,
         n35175, n35176, n35177, n35178, n35179, n35180, n35181, n35182,
         n35183, n35184, n35185, n35186, n35187, n35188, n35189, n35190,
         n35191, n35192, n35193, n35194, n35195, n35196, n35197, n35198,
         n35199, n35200, n35201, n35202, n35203, n35204, n35205, n35206,
         n35207, n35208, n35209, n35210, n35211, n35212, n35213, n35214,
         n35215, n35216, n35217, n35218, n35219, n35220, n35221, n35222,
         n35223, n35224, n35225, n35226, n35227, n35228, n35229, n35230,
         n35231, n35232, n35233, n35234, n35235, n35236, n35237, n35238,
         n35239, n35240, n35241, n35242, n35243, n35244, n35245, n35246,
         n35247, n35248, n35249, n35250, n35251, n35252, n35253, n35254,
         n35255, n35256, n35257, n35258, n35259, n35260, n35261, n35262,
         n35263, n35264, n35265, n35266, n35267, n35268, n35269, n35270,
         n35271, n35272, n35273, n35274, n35275, n35276, n35277, n35278,
         n35279, n35280, n35281, n35282, n35283, n35284, n35285, n35286,
         n35287, n35288, n35289, n35290, n35291, n35292, n35293, n35294,
         n35295, n35296, n35297, n35298, n35299, n35300, n35301, n35302,
         n35303, n35304, n35305, n35306, n35307, n35308, n35309, n35310,
         n35311, n35312, n35313, n35314, n35315, n35316, n35317, n35318,
         n35319, n35320, n35321, n35322, n35323, n35324, n35325, n35326,
         n35327, n35328, n35329, n35330, n35331, n35332, n35333, n35334,
         n35335, n35336, n35337, n35338, n35339, n35340, n35341, n35342,
         n35343, n35344, n35345, n35346, n35347, n35348, n35349, n35350,
         n35351, n35352, n35353, n35354, n35355, n35356, n35357, n35358,
         n35359, n35360, n35361, n35362, n35363, n35364, n35365, n35366,
         n35367, n35368, n35369, n35370, n35371, n35372, n35373, n35374,
         n35375, n35376, n35377, n35378, n35379, n35380, n35381, n35382,
         n35383, n35384, n35385, n35386, n35387, n35388, n35389, n35390,
         n35391, n35392, n35393, n35394, n35395, n35396, n35397, n35398,
         n35399, n35400, n35401, n35402, n35403, n35404, n35405, n35406,
         n35407, n35408, n35409, n35410, n35411, n35412, n35413, n35414,
         n35415, n35416, n35417, n35418, n35419, n35420, n35421, n35422,
         n35423, n35424, n35425, n35426, n35427, n35428, n35429, n35430,
         n35431, n35432, n35433, n35434, n35435, n35436, n35437, n35438,
         n35439, n35440, n35441, n35442, n35443, n35444, n35445, n35446,
         n35447, n35448, n35449, n35450, n35451, n35452, n35453, n35454,
         n35455, n35456, n35457, n35458, n35459, n35460, n35461, n35462,
         n35463, n35464, n35465, n35466, n35467, n35468, n35469, n35470,
         n35471, n35472, n35473, n35474, n35475, n35476, n35477, n35478,
         n35479, n35480, n35481, n35482, n35483, n35484, n35485, n35486,
         n35487, n35488, n35489, n35490, n35491, n35492, n35493, n35494,
         n35495, n35496, n35497, n35498, n35499, n35500, n35501, n35502,
         n35503, n35504, n35505, n35506, n35507, n35508, n35509, n35510,
         n35511, n35512, n35513, n35514, n35515, n35516, n35517, n35518,
         n35519, n35520, n35521, n35522, n35523, n35524, n35525, n35526,
         n35527, n35528, n35529, n35530, n35531, n35532, n35533, n35534,
         n35535, n35536, n35537, n35538, n35539, n35540, n35541, n35542,
         n35543, n35544, n35545, n35546, n35547, n35548, n35549, n35550,
         n35551, n35552, n35553, n35554, n35555, n35556, n35557, n35558,
         n35559, n35560, n35561, n35562, n35563, n35564, n35565, n35566,
         n35567, n35568, n35569, n35570, n35571, n35572, n35573, n35574,
         n35575, n35576, n35577, n35578, n35579, n35580, n35581, n35582,
         n35583, n35584, n35585, n35586, n35587, n35588, n35589, n35590,
         n35591, n35592, n35593, n35594, n35595, n35596, n35597, n35598,
         n35599, n35600, n35601, n35602, n35603, n35604, n35605, n35606,
         n35607, n35608, n35609, n35610, n35611, n35612, n35613, n35614,
         n35615, n35616, n35617, n35618, n35619, n35620, n35621, n35622,
         n35623, n35624, n35625, n35626, n35627, n35628, n35629, n35630,
         n35631, n35632, n35633, n35634, n35635, n35636, n35637, n35638,
         n35639, n35640, n35641, n35642, n35643, n35644, n35645, n35646,
         n35647, n35648, n35649, n35650, n35651, n35652, n35653, n35654,
         n35655, n35656, n35657, n35658, n35659, n35660, n35661, n35662,
         n35663, n35664, n35665, n35666, n35667, n35668, n35669, n35670,
         n35671, n35672, n35673, n35674, n35675, n35676, n35677, n35678,
         n35679, n35680, n35681, n35682, n35683, n35684, n35685, n35686,
         n35687, n35688, n35689, n35690, n35691, n35692, n35693, n35694,
         n35695, n35696, n35697, n35698, n35699, n35700, n35701, n35702,
         n35703, n35704, n35705, n35706, n35707, n35708, n35709, n35710,
         n35711, n35712, n35713, n35714, n35715, n35716, n35717, n35718,
         n35719, n35720, n35721, n35722, n35723, n35724, n35725, n35726,
         n35727, n35728, n35729, n35730, n35731, n35732, n35733, n35734,
         n35735, n35736, n35737, n35738, n35739, n35740, n35741, n35742,
         n35743, n35744, n35745, n35746, n35747, n35748, n35749, n35750,
         n35751, n35752, n35753, n35754, n35755, n35756, n35757, n35758,
         n35759, n35760, n35761, n35762, n35763, n35764, n35765, n35766,
         n35767, n35768, n35769, n35770, n35771, n35772, n35773, n35774,
         n35775, n35776, n35777, n35778, n35779, n35780, n35781, n35782,
         n35783, n35784, n35785, n35786, n35787, n35788, n35789, n35790,
         n35791, n35792, n35793, n35794, n35795, n35796, n35797, n35798,
         n35799, n35800, n35801, n35802, n35803, n35804, n35805, n35806,
         n35807, n35808, n35809, n35810, n35811, n35812, n35813, n35814,
         n35815, n35816, n35817, n35818, n35819, n35820, n35821, n35822,
         n35823, n35824, n35825, n35826, n35827, n35828, n35829, n35830,
         n35831, n35832, n35833, n35834, n35835, n35836, n35837, n35838,
         n35839, n35840, n35841, n35842, n35843, n35844, n35845, n35846,
         n35847, n35848, n35849, n35850, n35851, n35852, n35853, n35854,
         n35855, n35856, n35857, n35858, n35859, n35860, n35861, n35862,
         n35863, n35864, n35865, n35866, n35867, n35868, n35869, n35870,
         n35871, n35872, n35873, n35874, n35875, n35876, n35877, n35878,
         n35879, n35880, n35881, n35882, n35883, n35884, n35885, n35886,
         n35887, n35888, n35889, n35890, n35891, n35892, n35893, n35894,
         n35895, n35896, n35897, n35898, n35899, n35900, n35901, n35902,
         n35903, n35904, n35905, n35906, n35907, n35908, n35909, n35910,
         n35911, n35912, n35913, n35914, n35915, n35916, n35917, n35918,
         n35919, n35920, n35921, n35922, n35923, n35924, n35925, n35926,
         n35927, n35928, n35929, n35930, n35931, n35932, n35933, n35934,
         n35935, n35936, n35937, n35938, n35939, n35940, n35941, n35942,
         n35943, n35944, n35945, n35946, n35947, n35948, n35949, n35950,
         n35951, n35952, n35953, n35954, n35955, n35956, n35957, n35958,
         n35959, n35960, n35961, n35962, n35963, n35964, n35965, n35966,
         n35967, n35968, n35969, n35970, n35971, n35972, n35973, n35974,
         n35975, n35976, n35977, n35978, n35979, n35980, n35981, n35982,
         n35983, n35984, n35985, n35986, n35987, n35988, n35989, n35990,
         n35991, n35992, n35993, n35994, n35995, n35996, n35997, n35998,
         n35999, n36000, n36001, n36002, n36003, n36004, n36005, n36006,
         n36007, n36008, n36009, n36010, n36011, n36012, n36013, n36014,
         n36015, n36016, n36017, n36018, n36019, n36020, n36021, n36022,
         n36023, n36024, n36025, n36026, n36027, n36028, n36029, n36030,
         n36031, n36032, n36033, n36034, n36035, n36036, n36037, n36038,
         n36039, n36040, n36041, n36042, n36043, n36044, n36045, n36046,
         n36047, n36048, n36049, n36050, n36051, n36052, n36053, n36054,
         n36055, n36056, n36057, n36058, n36059, n36060, n36061, n36062,
         n36063, n36064, n36065, n36066, n36067, n36068, n36069, n36070,
         n36071, n36072, n36073, n36074, n36075, n36076, n36077, n36078,
         n36079, n36080, n36081, n36082, n36083, n36084, n36085, n36086,
         n36087, n36088, n36089, n36090, n36091, n36092, n36093, n36094,
         n36095, n36096, n36097, n36098, n36099, n36100, n36101, n36102,
         n36103, n36104, n36105, n36106, n36107, n36108, n36109, n36110,
         n36111, n36112, n36113, n36114, n36115, n36116, n36117, n36118,
         n36119, n36120, n36121, n36122, n36123, n36124, n36125, n36126,
         n36127, n36128, n36129, n36130, n36131, n36132, n36133, n36134,
         n36135, n36136, n36137, n36138, n36139, n36140, n36141, n36142,
         n36143, n36144, n36145, n36146, n36147, n36148, n36149, n36150,
         n36151, n36152, n36153, n36154, n36155, n36156, n36157, n36158,
         n36159, n36160, n36161, n36162, n36163, n36164, n36165, n36166,
         n36167, n36168, n36169, n36170, n36171, n36172, n36173, n36174,
         n36175, n36176, n36177, n36178, n36179, n36180, n36181, n36182,
         n36183, n36184, n36185, n36186, n36187, n36188, n36189, n36190,
         n36191, n36192, n36193, n36194, n36195, n36196, n36197, n36198,
         n36199, n36200, n36201, n36202, n36203, n36204, n36205, n36206,
         n36207, n36208, n36209, n36210, n36211, n36212, n36213, n36214,
         n36215, n36216, n36217, n36218, n36219, n36220, n36221, n36222,
         n36223, n36224, n36225, n36226, n36227, n36228, n36229, n36230,
         n36231, n36232, n36233, n36234, n36235, n36236, n36237, n36238,
         n36239, n36240, n36241, n36242, n36243, n36244, n36245, n36246,
         n36247, n36248, n36249, n36250, n36251, n36252, n36253, n36254,
         n36255, n36256, n36257, n36258, n36259, n36260, n36261, n36262,
         n36263, n36264, n36265, n36266, n36267, n36268, n36269, n36270,
         n36271, n36272, n36273, n36274, n36275, n36276, n36277, n36278,
         n36279, n36280, n36281, n36282, n36283, n36284, n36285, n36286,
         n36287, n36288, n36289, n36290, n36291, n36292, n36293, n36294,
         n36295, n36296, n36297, n36298, n36299, n36300, n36301, n36302,
         n36303, n36304, n36305, n36306, n36307, n36308, n36309, n36310,
         n36311, n36312, n36313, n36314, n36315, n36316, n36317, n36318,
         n36319, n36320, n36321, n36322, n36323, n36324, n36325, n36326,
         n36327, n36328, n36329, n36330, n36331, n36332, n36333, n36334,
         n36335, n36336, n36337, n36338, n36339, n36340, n36341, n36342,
         n36343, n36344, n36345, n36346, n36347, n36348, n36349, n36350,
         n36351, n36352, n36353, n36354, n36355, n36356, n36357, n36358,
         n36359, n36360, n36361, n36362, n36363, n36364, n36365, n36366,
         n36367, n36368, n36369, n36370, n36371, n36372, n36373, n36374,
         n36375, n36376, n36377, n36378, n36379, n36380, n36381, n36382,
         n36383, n36384, n36385, n36386, n36387, n36388, n36389, n36390,
         n36391, n36392, n36393, n36394, n36395, n36396, n36397, n36398,
         n36399, n36400, n36401, n36402, n36403, n36404, n36405, n36406,
         n36407, n36408, n36409, n36410, n36411, n36412, n36413, n36414,
         n36415, n36416, n36417, n36418, n36419, n36420, n36421, n36422,
         n36423, n36424, n36425, n36426, n36427, n36428, n36429, n36430,
         n36431, n36432, n36433, n36434, n36435, n36436, n36437, n36438,
         n36439, n36440, n36441, n36442, n36443, n36444, n36445, n36446,
         n36447, n36448, n36449, n36450, n36451, n36452, n36453, n36454,
         n36455, n36456, n36457, n36458, n36459, n36460, n36461, n36462,
         n36463, n36464, n36465, n36466, n36467, n36468, n36469, n36470,
         n36471, n36472, n36473, n36474, n36475, n36476, n36477, n36478,
         n36479, n36480, n36481, n36482, n36483, n36484, n36485, n36486,
         n36487, n36488, n36489, n36490, n36491, n36492, n36493, n36494,
         n36495, n36496, n36497, n36498, n36499, n36500, n36501, n36502,
         n36503, n36504, n36505, n36506, n36507, n36508, n36509, n36510,
         n36511, n36512, n36513, n36514, n36515, n36516, n36517, n36518,
         n36519, n36520, n36521, n36522, n36523, n36524, n36525, n36526,
         n36527, n36528, n36529, n36530, n36531, n36532, n36533, n36534,
         n36535, n36536, n36537, n36538, n36539, n36540, n36541, n36542,
         n36543, n36544, n36545, n36546, n36547, n36548, n36549, n36550,
         n36551, n36552, n36553, n36554, n36555, n36556, n36557, n36558,
         n36559, n36560, n36561, n36562, n36563, n36564, n36565, n36566,
         n36567, n36568, n36569, n36570, n36571, n36572, n36573, n36574,
         n36575, n36576, n36577, n36578, n36579, n36580, n36581, n36582,
         n36583, n36584, n36585, n36586, n36587, n36588, n36589, n36590,
         n36591, n36592, n36593, n36594, n36595, n36596, n36597, n36598,
         n36599, n36600, n36601, n36602, n36603, n36604, n36605, n36606,
         n36607, n36608, n36609, n36610, n36611, n36612, n36613, n36614,
         n36615, n36616, n36617, n36618, n36619, n36620, n36621, n36622,
         n36623, n36624, n36625, n36626, n36627, n36628, n36629, n36630,
         n36631, n36632, n36633, n36634, n36635, n36636, n36637, n36638,
         n36639, n36640, n36641, n36642, n36643, n36644, n36645, n36646,
         n36647, n36648, n36649, n36650, n36651, n36652, n36653, n36654,
         n36655, n36656, n36657, n36658, n36659, n36660, n36661, n36662,
         n36663, n36664, n36665, n36666, n36667, n36668, n36669, n36670,
         n36671, n36672, n36673, n36674, n36675, n36676, n36677, n36678,
         n36679, n36680, n36681, n36682, n36683, n36684, n36685, n36686,
         n36687, n36688, n36689, n36690, n36691, n36692, n36693, n36694,
         n36695, n36696, n36697, n36698, n36699, n36700, n36701, n36702,
         n36703, n36704, n36705, n36706, n36707, n36708, n36709, n36710,
         n36711, n36712, n36713, n36714, n36715, n36716, n36717, n36718,
         n36719, n36720, n36721, n36722, n36723, n36724, n36725, n36726,
         n36727, n36728, n36729, n36730, n36731, n36732, n36733, n36734,
         n36735, n36736, n36737, n36738, n36739, n36740, n36741, n36742,
         n36743, n36744, n36745, n36746, n36747, n36748, n36749, n36750,
         n36751, n36752, n36753, n36754, n36755, n36756, n36757, n36758,
         n36759, n36760, n36761, n36762, n36763, n36764, n36765, n36766,
         n36767, n36768, n36769, n36770, n36771, n36772, n36773, n36774,
         n36775, n36776, n36777, n36778, n36779, n36780, n36781, n36782,
         n36783, n36784, n36785, n36786, n36787, n36788, n36789, n36790,
         n36791, n36792, n36793, n36794, n36795, n36796, n36797, n36798,
         n36799, n36800, n36801, n36802, n36803, n36804, n36805, n36806,
         n36807, n36808, n36809, n36810, n36811, n36812, n36813, n36814,
         n36815, n36816, n36817, n36818, n36819, n36820, n36821, n36822,
         n36823, n36824, n36825, n36826, n36827, n36828, n36829, n36830,
         n36831, n36832, n36833, n36834, n36835, n36836, n36837, n36838,
         n36839, n36840, n36841, n36842, n36843, n36844, n36845, n36846,
         n36847, n36848, n36849, n36850, n36851, n36852, n36853, n36854,
         n36855, n36856, n36857, n36858, n36859, n36860, n36861, n36862,
         n36863, n36864, n36865, n36866, n36867, n36868, n36869, n36870,
         n36871, n36872, n36873, n36874, n36875, n36876, n36877, n36878,
         n36879, n36880, n36881, n36882, n36883, n36884, n36885, n36886,
         n36887, n36888, n36889, n36890, n36891, n36892, n36893, n36894,
         n36895, n36896, n36897, n36898, n36899, n36900, n36901, n36902,
         n36903, n36904, n36905, n36906, n36907, n36908, n36909, n36910,
         n36911, n36912, n36913, n36914, n36915, n36916, n36917, n36918,
         n36919, n36920, n36921, n36922, n36923, n36924, n36925, n36926,
         n36927, n36928, n36929, n36930, n36931, n36932, n36933, n36934,
         n36935, n36936, n36937, n36938, n36939, n36940, n36941, n36942,
         n36943, n36944, n36945, n36946, n36947, n36948, n36949, n36950,
         n36951, n36952, n36953, n36954, n36955, n36956, n36957, n36958,
         n36959, n36960, n36961, n36962, n36963, n36964, n36965, n36966,
         n36967, n36968, n36969, n36970, n36971, n36972, n36973, n36974,
         n36975, n36976, n36977, n36978, n36979, n36980, n36981, n36982,
         n36983, n36984, n36985, n36986, n36987, n36988, n36989, n36990,
         n36991, n36992, n36993, n36994, n36995, n36996, n36997, n36998,
         n36999, n37000, n37001, n37002, n37003, n37004, n37005, n37006,
         n37007, n37008, n37009, n37010, n37011, n37012, n37013, n37014,
         n37015, n37016, n37017, n37018, n37019, n37020, n37021, n37022,
         n37023, n37024, n37025, n37026, n37027, n37028, n37029, n37030,
         n37031, n37032, n37033, n37034, n37035, n37036, n37037, n37038,
         n37039, n37040, n37041, n37042, n37043, n37044, n37045, n37046,
         n37047, n37048, n37049, n37050, n37051, n37052, n37053, n37054,
         n37055, n37056, n37057, n37058, n37059, n37060, n37061, n37062,
         n37063, n37064, n37065, n37066, n37067, n37068, n37069, n37070,
         n37071, n37072, n37073, n37074, n37075, n37076, n37077, n37078,
         n37079, n37080, n37081, n37082, n37083, n37084, n37085, n37086,
         n37087, n37088, n37089, n37090, n37091, n37092, n37093, n37094,
         n37095, n37096, n37097, n37098, n37099, n37100, n37101, n37102,
         n37103, n37104, n37105, n37106, n37107, n37108, n37109, n37110,
         n37111, n37112, n37113, n37114, n37115, n37116, n37117, n37118,
         n37119, n37120, n37121, n37122, n37123, n37124, n37125, n37126,
         n37127, n37128, n37129, n37130, n37131, n37132, n37133, n37134,
         n37135, n37136, n37137, n37138, n37139, n37140, n37141, n37142,
         n37143, n37144, n37145, n37146, n37147, n37148, n37149, n37150,
         n37151, n37152, n37153, n37154, n37155, n37156, n37157, n37158,
         n37159, n37160, n37161, n37162, n37163, n37164, n37165, n37166,
         n37167, n37168, n37169, n37170, n37171, n37172, n37173, n37174,
         n37175, n37176, n37177, n37178, n37179, n37180, n37181, n37182,
         n37183, n37184, n37185, n37186, n37187, n37188, n37189, n37190,
         n37191, n37192, n37193, n37194, n37195, n37196, n37197, n37198,
         n37199, n37200, n37201, n37202, n37203, n37204, n37205, n37206,
         n37207, n37208, n37209, n37210, n37211, n37212, n37213, n37214,
         n37215, n37216, n37217, n37218, n37219, n37220, n37221, n37222,
         n37223, n37224, n37225, n37226, n37227, n37228, n37229, n37230,
         n37231, n37232, n37233, n37234, n37235, n37236, n37237, n37238,
         n37239, n37240, n37241, n37242, n37243, n37244, n37245, n37246,
         n37247, n37248, n37249, n37250, n37251, n37252, n37253, n37254,
         n37255, n37256, n37257, n37258, n37259, n37260, n37261, n37262,
         n37263, n37264, n37265, n37266, n37267, n37268, n37269, n37270,
         n37271, n37272, n37273, n37274, n37275, n37276, n37277, n37278,
         n37279, n37280, n37281, n37282, n37283, n37284, n37285, n37286,
         n37287, n37288, n37289, n37290, n37291, n37292, n37293, n37294,
         n37295, n37296, n37297, n37298, n37299, n37300, n37301, n37302,
         n37303, n37304, n37305, n37306, n37307, n37308, n37309, n37310,
         n37311, n37312, n37313, n37314, n37315, n37316, n37317, n37318,
         n37319, n37320, n37321, n37322, n37323, n37324, n37325, n37326,
         n37327, n37328, n37329, n37330, n37331, n37332, n37333, n37334,
         n37335, n37336, n37337, n37338, n37339, n37340, n37341, n37342,
         n37343, n37344, n37345, n37346, n37347, n37348, n37349, n37350,
         n37351, n37352, n37353, n37354, n37355, n37356, n37357, n37358,
         n37359, n37360, n37361, n37362, n37363, n37364, n37365, n37366,
         n37367, n37368, n37369, n37370, n37371, n37372, n37373, n37374,
         n37375, n37376, n37377, n37378, n37379, n37380, n37381, n37382,
         n37383, n37384, n37385, n37386, n37387, n37388, n37389, n37390,
         n37391, n37392, n37393, n37394, n37395, n37396, n37397, n37398,
         n37399, n37400, n37401, n37402, n37403, n37404, n37405, n37406,
         n37407, n37408, n37409, n37410, n37411, n37412, n37413, n37414,
         n37415, n37416, n37417, n37418, n37419, n37420, n37421, n37422,
         n37423, n37424, n37425, n37426, n37427, n37428, n37429, n37430,
         n37431, n37432, n37433, n37434, n37435, n37436, n37437, n37438,
         n37439, n37440, n37441, n37442, n37443, n37444, n37445, n37446,
         n37447, n37448, n37449, n37450, n37451, n37452, n37453, n37454,
         n37455, n37456, n37457, n37458, n37459, n37460, n37461, n37462,
         n37463, n37464, n37465, n37466, n37467, n37468, n37469, n37470,
         n37471, n37472, n37473, n37474, n37475, n37476, n37477, n37478,
         n37479, n37480, n37481, n37482, n37483, n37484, n37485, n37486,
         n37487, n37488, n37489, n37490, n37491, n37492, n37493, n37494,
         n37495, n37496, n37497, n37498, n37499, n37500, n37501, n37502,
         n37503, n37504, n37505, n37506, n37507, n37508, n37509, n37510,
         n37511, n37512, n37513, n37514, n37515, n37516, n37517, n37518,
         n37519, n37520, n37521, n37522, n37523, n37524, n37525, n37526,
         n37527, n37528, n37529, n37530, n37531, n37532, n37533, n37534,
         n37535, n37536, n37537, n37538, n37539, n37540, n37541, n37542,
         n37543, n37544, n37545, n37546, n37547, n37548, n37549, n37550,
         n37551, n37552, n37553, n37554, n37555, n37556, n37557, n37558,
         n37559, n37560, n37561, n37562, n37563, n37564, n37565, n37566,
         n37567, n37568, n37569, n37570, n37571, n37572, n37573, n37574,
         n37575, n37576, n37577, n37578, n37579, n37580, n37581, n37582,
         n37583, n37584, n37585, n37586, n37587, n37588, n37589, n37590,
         n37591, n37592, n37593, n37594, n37595, n37596, n37597, n37598,
         n37599, n37600, n37601, n37602, n37603, n37604, n37605, n37606,
         n37607, n37608, n37609, n37610, n37611, n37612, n37613, n37614,
         n37615, n37616, n37617, n37618, n37619, n37620, n37621, n37622,
         n37623, n37624, n37625, n37626, n37627, n37628, n37629, n37630,
         n37631, n37632, n37633, n37634, n37635, n37636, n37637, n37638,
         n37639, n37640, n37641, n37642, n37643, n37644, n37645, n37646,
         n37647, n37648, n37649, n37650, n37651, n37652, n37653, n37654,
         n37655, n37656, n37657, n37658, n37659, n37660, n37661, n37662,
         n37663, n37664, n37665, n37666, n37667, n37668, n37669, n37670,
         n37671, n37672, n37673, n37674, n37675, n37676, n37677, n37678,
         n37679, n37680, n37681, n37682, n37683, n37684, n37685, n37686,
         n37687, n37688, n37689, n37690, n37691, n37692, n37693, n37694,
         n37695, n37696, n37697, n37698, n37699, n37700, n37701, n37702,
         n37703, n37704, n37705, n37706, n37707, n37708, n37709, n37710,
         n37711, n37712, n37713, n37714, n37715, n37716, n37717, n37718,
         n37719, n37720, n37721, n37722, n37723, n37724, n37725, n37726,
         n37727, n37728, n37729, n37730, n37731, n37732, n37733, n37734,
         n37735, n37736, n37737, n37738, n37739, n37740, n37741, n37742,
         n37743, n37744, n37745, n37746, n37747, n37748, n37749, n37750,
         n37751, n37752, n37753, n37754, n37755, n37756, n37757, n37758,
         n37759, n37760, n37761, n37762, n37763, n37764, n37765, n37766,
         n37767, n37768, n37769, n37770, n37771, n37772, n37773, n37774,
         n37775, n37776, n37777, n37778, n37779, n37780, n37781, n37782,
         n37783, n37784, n37785, n37786, n37787, n37788, n37789, n37790,
         n37791, n37792, n37793, n37794, n37795, n37796, n37797, n37798,
         n37799, n37800, n37801, n37802, n37803, n37804, n37805, n37806,
         n37807, n37808, n37809, n37810, n37811, n37812, n37813, n37814,
         n37815, n37816, n37817, n37818, n37819, n37820, n37821, n37822,
         n37823, n37824, n37825, n37826, n37827, n37828, n37829, n37830,
         n37831, n37832, n37833, n37834, n37835, n37836, n37837, n37838,
         n37839, n37840, n37841, n37842, n37843, n37844, n37845, n37846,
         n37847, n37848, n37849, n37850, n37851, n37852, n37853, n37854,
         n37855, n37856, n37857, n37858, n37859, n37860, n37861, n37862,
         n37863, n37864, n37865, n37866, n37867, n37868, n37869, n37870,
         n37871, n37872, n37873, n37874, n37875, n37876, n37877, n37878,
         n37879, n37880, n37881, n37882, n37883, n37884, n37885, n37886,
         n37887, n37888, n37889, n37890, n37891, n37892, n37893, n37894,
         n37895, n37896, n37897, n37898, n37899, n37900, n37901, n37902,
         n37903, n37904, n37905, n37906, n37907, n37908, n37909, n37910,
         n37911, n37912, n37913, n37914, n37915, n37916, n37917, n37918,
         n37919, n37920, n37921, n37922, n37923, n37924, n37925, n37926,
         n37927, n37928, n37929, n37930, n37931, n37932, n37933, n37934,
         n37935, n37936, n37937, n37938, n37939, n37940, n37941, n37942,
         n37943, n37944, n37945, n37946, n37947, n37948, n37949, n37950,
         n37951, n37952, n37953, n37954, n37955, n37956, n37957, n37958,
         n37959, n37960, n37961, n37962, n37963, n37964, n37965, n37966,
         n37967, n37968, n37969, n37970, n37971, n37972, n37973, n37974,
         n37975, n37976, n37977, n37978, n37979, n37980, n37981, n37982,
         n37983, n37984, n37985, n37986, n37987, n37988, n37989, n37990,
         n37991, n37992, n37993, n37994, n37995, n37996, n37997, n37998,
         n37999, n38000, n38001, n38002, n38003, n38004, n38005, n38006,
         n38007, n38008, n38009, n38010, n38011, n38012, n38013, n38014,
         n38015, n38016, n38017, n38018, n38019, n38020, n38021, n38022,
         n38023, n38024, n38025, n38026, n38027, n38028, n38029, n38030,
         n38031, n38032, n38033, n38034, n38035, n38036, n38037, n38038,
         n38039, n38040, n38041, n38042, n38043, n38044, n38045, n38046,
         n38047, n38048, n38049, n38050, n38051, n38052, n38053, n38054,
         n38055, n38056, n38057, n38058, n38059, n38060, n38061, n38062,
         n38063, n38064, n38065, n38066, n38067, n38068, n38069, n38070,
         n38071, n38072, n38073, n38074, n38075, n38076, n38077, n38078,
         n38079, n38080, n38081, n38082, n38083, n38084, n38085, n38086,
         n38087, n38088, n38089, n38090, n38091, n38092, n38093, n38094,
         n38095, n38096, n38097, n38098, n38099, n38100, n38101, n38102,
         n38103, n38104, n38105, n38106, n38107, n38108, n38109, n38110,
         n38111, n38112, n38113, n38114, n38115, n38116, n38117, n38118,
         n38119, n38120, n38121, n38122, n38123, n38124, n38125, n38126,
         n38127, n38128, n38129, n38130, n38131, n38132, n38133, n38134,
         n38135, n38136, n38137, n38138, n38139, n38140, n38141, n38142,
         n38143, n38144, n38145, n38146, n38147, n38148, n38149, n38150,
         n38151, n38152, n38153, n38154, n38155, n38156, n38157, n38158,
         n38159, n38160, n38161, n38162, n38163, n38164, n38165, n38166,
         n38167, n38168, n38169, n38170, n38171, n38172, n38173, n38174,
         n38175, n38176, n38177, n38178, n38179, n38180, n38181, n38182,
         n38183, n38184, n38185, n38186, n38187, n38188, n38189, n38190,
         n38191, n38192, n38193, n38194, n38195, n38196, n38197, n38198,
         n38199, n38200, n38201, n38202, n38203, n38204, n38205, n38206,
         n38207, n38208, n38209, n38210, n38211, n38212, n38213, n38214,
         n38215, n38216, n38217, n38218, n38219, n38220, n38221, n38222,
         n38223, n38224, n38225, n38226, n38227, n38228, n38229, n38230,
         n38231, n38232, n38233, n38234, n38235, n38236, n38237, n38238,
         n38239, n38240, n38241, n38242, n38243, n38244, n38245, n38246,
         n38247, n38248, n38249, n38250, n38251, n38252, n38253, n38254,
         n38255, n38256, n38257, n38258, n38259, n38260, n38261, n38262,
         n38263, n38264, n38265, n38266, n38267, n38268, n38269, n38270,
         n38271, n38272, n38273, n38274, n38275, n38276, n38277, n38278,
         n38279, n38280, n38281, n38282, n38283, n38284, n38285, n38286,
         n38287, n38288, n38289, n38290, n38291, n38292, n38293, n38294,
         n38295, n38296, n38297, n38298, n38299, n38300, n38301, n38302,
         n38303, n38304, n38305, n38306, n38307, n38308, n38309, n38310,
         n38311, n38312, n38313, n38314, n38315, n38316, n38317, n38318,
         n38319, n38320, n38321, n38322, n38323, n38324, n38325, n38326,
         n38327, n38328, n38329, n38330, n38331, n38332, n38333, n38334,
         n38335, n38336, n38337, n38338, n38339, n38340, n38341, n38342,
         n38343, n38344, n38345, n38346, n38347, n38348, n38349, n38350,
         n38351, n38352, n38353, n38354, n38355, n38356, n38357, n38358,
         n38359, n38360, n38361, n38362, n38363, n38364, n38365, n38366,
         n38367, n38368, n38369, n38370, n38371, n38372, n38373, n38374,
         n38375, n38376, n38377, n38378, n38379, n38380, n38381, n38382,
         n38383, n38384, n38385, n38386, n38387, n38388, n38389, n38390,
         n38391, n38392, n38393, n38394, n38395, n38396, n38397, n38398,
         n38399, n38400, n38401, n38402, n38403, n38404, n38405, n38406,
         n38407, n38408, n38409, n38410, n38411, n38412, n38413, n38414,
         n38415, n38416, n38417, n38418, n38419, n38420, n38421, n38422,
         n38423, n38424, n38425, n38426, n38427, n38428, n38429, n38430,
         n38431, n38432, n38433, n38434, n38435, n38436, n38437, n38438,
         n38439, n38440, n38441, n38442, n38443, n38444, n38445, n38446,
         n38447, n38448, n38449, n38450, n38451, n38452, n38453, n38454,
         n38455, n38456, n38457, n38458, n38459, n38460, n38461, n38462,
         n38463, n38464, n38465, n38466, n38467, n38468, n38469, n38470,
         n38471, n38472, n38473, n38474, n38475, n38476, n38477, n38478,
         n38479, n38480, n38481, n38482, n38483, n38484, n38485, n38486,
         n38487, n38488, n38489, n38490, n38491, n38492, n38493, n38494,
         n38495, n38496, n38497, n38498, n38499, n38500, n38501, n38502,
         n38503, n38504, n38505, n38506, n38507, n38508, n38509, n38510,
         n38511, n38512, n38513, n38514, n38515, n38516, n38517, n38518,
         n38519, n38520, n38521, n38522, n38523, n38524, n38525, n38526,
         n38527, n38528, n38529, n38530, n38531, n38532, n38533, n38534,
         n38535, n38536, n38537, n38538, n38539, n38540, n38541, n38542,
         n38543, n38544, n38545, n38546, n38547, n38548, n38549, n38550,
         n38551, n38552, n38553, n38554, n38555, n38556, n38557, n38558,
         n38559, n38560, n38561, n38562, n38563, n38564, n38565, n38566,
         n38567, n38568, n38569, n38570, n38571, n38572, n38573, n38574,
         n38575, n38576, n38577, n38578, n38579, n38580, n38581, n38582,
         n38583, n38584, n38585, n38586, n38587, n38588, n38589, n38590,
         n38591, n38592, n38593, n38594, n38595, n38596, n38597, n38598,
         n38599, n38600, n38601, n38602, n38603, n38604, n38605, n38606,
         n38607, n38608, n38609, n38610, n38611, n38612, n38613, n38614,
         n38615, n38616, n38617, n38618, n38619, n38620, n38621, n38622,
         n38623, n38624, n38625, n38626, n38627, n38628, n38629, n38630,
         n38631, n38632, n38633, n38634, n38635, n38636, n38637, n38638,
         n38639, n38640, n38641, n38642, n38643, n38644, n38645, n38646,
         n38647, n38648, n38649, n38650, n38651, n38652, n38653, n38654,
         n38655, n38656, n38657, n38658, n38659, n38660, n38661, n38662,
         n38663, n38664, n38665, n38666, n38667, n38668, n38669, n38670,
         n38671, n38672, n38673, n38674, n38675, n38676, n38677, n38678,
         n38679, n38680, n38681, n38682, n38683, n38684, n38685, n38686,
         n38687, n38688, n38689, n38690, n38691, n38692, n38693, n38694,
         n38695, n38696, n38697, n38698, n38699, n38700, n38701, n38702,
         n38703, n38704, n38705, n38706, n38707, n38708, n38709, n38710,
         n38711, n38712, n38713, n38714, n38715, n38716, n38717, n38718,
         n38719, n38720, n38721, n38722, n38723, n38724, n38725, n38726,
         n38727, n38728, n38729, n38730, n38731, n38732, n38733, n38734,
         n38735, n38736, n38737, n38738, n38739, n38740, n38741, n38742,
         n38743, n38744, n38745, n38746, n38747, n38748, n38749, n38750,
         n38751, n38752, n38753, n38754, n38755, n38756, n38757, n38758,
         n38759, n38760, n38761, n38762, n38763, n38764, n38765, n38766,
         n38767, n38768, n38769, n38770, n38771, n38772, n38773, n38774,
         n38775, n38776, n38777, n38778, n38779, n38780, n38781, n38782,
         n38783, n38784, n38785, n38786, n38787, n38788, n38789, n38790,
         n38791, n38792, n38793, n38794, n38795, n38796, n38797, n38798,
         n38799, n38800, n38801, n38802, n38803, n38804, n38805, n38806,
         n38807, n38808, n38809, n38810, n38811, n38812, n38813, n38814,
         n38815, n38816, n38817, n38818, n38819, n38820, n38821, n38822,
         n38823, n38824, n38825, n38826, n38827, n38828, n38829, n38830,
         n38831, n38832, n38833, n38834, n38835, n38836, n38837, n38838,
         n38839, n38840, n38841, n38842, n38843, n38844, n38845, n38846,
         n38847, n38848, n38849, n38850, n38851, n38852, n38853, n38854,
         n38855, n38856, n38857, n38858, n38859, n38860, n38861, n38862,
         n38863, n38864, n38865, n38866, n38867, n38868, n38869, n38870,
         n38871, n38872, n38873, n38874, n38875, n38876, n38877, n38878,
         n38879, n38880, n38881, n38882, n38883, n38884, n38885, n38886,
         n38887, n38888, n38889, n38890, n38891, n38892, n38893, n38894,
         n38895, n38896, n38897, n38898, n38899, n38900, n38901, n38902,
         n38903, n38904, n38905, n38906, n38907, n38908, n38909, n38910,
         n38911, n38912, n38913, n38914, n38915, n38916, n38917, n38918,
         n38919, n38920, n38921, n38922, n38923, n38924, n38925, n38926,
         n38927, n38928, n38929, n38930, n38931, n38932, n38933, n38934,
         n38935, n38936, n38937, n38938, n38939, n38940, n38941, n38942,
         n38943, n38944, n38945, n38946, n38947, n38948, n38949, n38950,
         n38951, n38952, n38953, n38954, n38955, n38956, n38957, n38958,
         n38959, n38960, n38961, n38962, n38963, n38964, n38965, n38966,
         n38967, n38968, n38969, n38970, n38971, n38972, n38973, n38974,
         n38975, n38976, n38977, n38978, n38979, n38980, n38981, n38982,
         n38983, n38984, n38985, n38986, n38987, n38988, n38989, n38990,
         n38991, n38992, n38993, n38994, n38995, n38996, n38997, n38998,
         n38999, n39000, n39001, n39002, n39003, n39004, n39005, n39006,
         n39007, n39008, n39009, n39010, n39011, n39012, n39013, n39014,
         n39015, n39016, n39017, n39018, n39019, n39020, n39021, n39022,
         n39023, n39024, n39025, n39026, n39027, n39028, n39029, n39030,
         n39031, n39032, n39033, n39034, n39035, n39036, n39037, n39038,
         n39039, n39040, n39041, n39042, n39043, n39044, n39045, n39046,
         n39047, n39048, n39049, n39050, n39051, n39052, n39053, n39054,
         n39055, n39056, n39057, n39058, n39059, n39060, n39061, n39062,
         n39063, n39064, n39065, n39066, n39067, n39068, n39069, n39070,
         n39071, n39072, n39073, n39074, n39075, n39076, n39077, n39078,
         n39079, n39080, n39081, n39082, n39083, n39084, n39085, n39086,
         n39087, n39088, n39089, n39090, n39091, n39092, n39093, n39094,
         n39095, n39096, n39097, n39098, n39099, n39100, n39101, n39102,
         n39103, n39104, n39105, n39106, n39107, n39108, n39109, n39110,
         n39111, n39112, n39113, n39114, n39115, n39116, n39117, n39118,
         n39119, n39120, n39121, n39122, n39123, n39124, n39125, n39126,
         n39127, n39128, n39129, n39130, n39131, n39132, n39133, n39134,
         n39135, n39136, n39137, n39138, n39139, n39140, n39141, n39142,
         n39143, n39144, n39145, n39146, n39147, n39148, n39149, n39150,
         n39151, n39152, n39153, n39154, n39155, n39156, n39157, n39158,
         n39159, n39160, n39161, n39162, n39163, n39164, n39165, n39166,
         n39167, n39168, n39169, n39170, n39171, n39172, n39173, n39174,
         n39175, n39176, n39177, n39178, n39179, n39180, n39181, n39182,
         n39183, n39184, n39185, n39186, n39187, n39188, n39189, n39190,
         n39191, n39192, n39193, n39194, n39195, n39196, n39197, n39198,
         n39199, n39200, n39201, n39202, n39203, n39204, n39205, n39206,
         n39207, n39208, n39209, n39210, n39211, n39212, n39213, n39214,
         n39215, n39216, n39217, n39218, n39219, n39220, n39221, n39222,
         n39223, n39224, n39225, n39226, n39227, n39228, n39229, n39230,
         n39231, n39232, n39233, n39234, n39235, n39236, n39237, n39238,
         n39239, n39240, n39241, n39242, n39243, n39244, n39245, n39246,
         n39247, n39248, n39249, n39250, n39251, n39252, n39253, n39254,
         n39255, n39256, n39257, n39258, n39259, n39260, n39261, n39262,
         n39263, n39264, n39265, n39266, n39267, n39268, n39269, n39270,
         n39271, n39272, n39273, n39274, n39275, n39276, n39277, n39278,
         n39279, n39280, n39281, n39282, n39283, n39284, n39285, n39286,
         n39287, n39288, n39289, n39290, n39291, n39292, n39293, n39294,
         n39295, n39296, n39297, n39298, n39299, n39300, n39301, n39302,
         n39303, n39304, n39305, n39306, n39307, n39308, n39309, n39310,
         n39311, n39312, n39313, n39314, n39315, n39316, n39317, n39318,
         n39319, n39320, n39321, n39322, n39323, n39324, n39325, n39326,
         n39327, n39328, n39329, n39330, n39331, n39332, n39333, n39334,
         n39335, n39336, n39337, n39338, n39339, n39340, n39341, n39342,
         n39343, n39344, n39345, n39346, n39347, n39348, n39349, n39350,
         n39351, n39352, n39353, n39354, n39355, n39356, n39357, n39358,
         n39359, n39360, n39361, n39362, n39363, n39364, n39365, n39366,
         n39367, n39368, n39369, n39370, n39371, n39372, n39373, n39374,
         n39375, n39376, n39377, n39378, n39379, n39380, n39381, n39382,
         n39383, n39384, n39385, n39386, n39387, n39388, n39389, n39390,
         n39391, n39392, n39393, n39394, n39395, n39396, n39397, n39398,
         n39399, n39400, n39401, n39402, n39403, n39404, n39405, n39406,
         n39407, n39408, n39409, n39410, n39411, n39412, n39413, n39414,
         n39415, n39416, n39417, n39418, n39419, n39420, n39421, n39422,
         n39423, n39424, n39425, n39426, n39427, n39428, n39429, n39430,
         n39431, n39432, n39433, n39434, n39435, n39436, n39437, n39438,
         n39439, n39440, n39441, n39442, n39443, n39444, n39445, n39446,
         n39447, n39448, n39449, n39450, n39451, n39452, n39453, n39454,
         n39455, n39456, n39457, n39458, n39459, n39460, n39461, n39462,
         n39463, n39464, n39465, n39466, n39467, n39468, n39469, n39470,
         n39471, n39472, n39473, n39474, n39475, n39476, n39477, n39478,
         n39479, n39480, n39481, n39482, n39483, n39484, n39485, n39486,
         n39487, n39488, n39489, n39490, n39491, n39492, n39493, n39494,
         n39495, n39496, n39497, n39498, n39499, n39500, n39501, n39502,
         n39503, n39504, n39505, n39506, n39507, n39508, n39509, n39510,
         n39511, n39512, n39513, n39514, n39515, n39516, n39517, n39518,
         n39519, n39520, n39521, n39522, n39523, n39524, n39525, n39526,
         n39527, n39528, n39529, n39530, n39531, n39532, n39533, n39534,
         n39535, n39536, n39537, n39538, n39539, n39540, n39541, n39542,
         n39543, n39544, n39545, n39546, n39547, n39548, n39549, n39550,
         n39551, n39552, n39553, n39554, n39555, n39556, n39557, n39558,
         n39559, n39560, n39561, n39562, n39563, n39564, n39565, n39566,
         n39567, n39568, n39569, n39570, n39571, n39572, n39573, n39574,
         n39575, n39576, n39577, n39578, n39579, n39580, n39581, n39582,
         n39583, n39584, n39585, n39586, n39587, n39588, n39589, n39590,
         n39591, n39592, n39593, n39594, n39595, n39596, n39597, n39598,
         n39599, n39600, n39601, n39602, n39603, n39604, n39605, n39606,
         n39607, n39608, n39609, n39610, n39611, n39612, n39613, n39614,
         n39615, n39616, n39617, n39618, n39619, n39620, n39621, n39622,
         n39623, n39624, n39625, n39626, n39627, n39628, n39629, n39630,
         n39631, n39632, n39633, n39634, n39635, n39636, n39637, n39638,
         n39639, n39640, n39641, n39642, n39643, n39644, n39645, n39646,
         n39647, n39648, n39649, n39650, n39651, n39652, n39653, n39654,
         n39655, n39656, n39657, n39658, n39659, n39660, n39661, n39662,
         n39663, n39664, n39665, n39666, n39667, n39668, n39669, n39670,
         n39671, n39672, n39673, n39674, n39675, n39676, n39677, n39678,
         n39679, n39680, n39681, n39682, n39683, n39684, n39685, n39686,
         n39687, n39688, n39689, n39690, n39691, n39692, n39693, n39694,
         n39695, n39696, n39697, n39698, n39699, n39700, n39701, n39702,
         n39703, n39704, n39705, n39706, n39707, n39708, n39709, n39710,
         n39711, n39712, n39713, n39714, n39715, n39716, n39717, n39718,
         n39719, n39720, n39721, n39722, n39723, n39724, n39725, n39726,
         n39727, n39728, n39729, n39730, n39731, n39732, n39733, n39734,
         n39735, n39736, n39737, n39738, n39739, n39740, n39741, n39742,
         n39743, n39744, n39745, n39746, n39747, n39748, n39749, n39750,
         n39751, n39752, n39753, n39754, n39755, n39756, n39757, n39758,
         n39759, n39760, n39761, n39762, n39763, n39764, n39765, n39766,
         n39767, n39768, n39769, n39770, n39771, n39772, n39773, n39774,
         n39775, n39776, n39777, n39778, n39779, n39780, n39781, n39782,
         n39783, n39784, n39785, n39786, n39787, n39788, n39789, n39790,
         n39791, n39792, n39793, n39794, n39795, n39796, n39797, n39798,
         n39799, n39800, n39801, n39802, n39803, n39804, n39805, n39806,
         n39807, n39808, n39809, n39810, n39811, n39812, n39813, n39814,
         n39815, n39816, n39817, n39818, n39819, n39820, n39821, n39822,
         n39823, n39824, n39825, n39826, n39827, n39828, n39829, n39830,
         n39831, n39832, n39833, n39834, n39835, n39836, n39837, n39838,
         n39839, n39840, n39841, n39842, n39843, n39844, n39845, n39846,
         n39847, n39848, n39849, n39850, n39851, n39852, n39853, n39854,
         n39855, n39856, n39857, n39858, n39859, n39860, n39861, n39862,
         n39863, n39864, n39865, n39866, n39867, n39868, n39869, n39870,
         n39871, n39872, n39873, n39874, n39875, n39876, n39877, n39878,
         n39879, n39880, n39881, n39882, n39883, n39884, n39885, n39886,
         n39887, n39888, n39889, n39890, n39891, n39892, n39893, n39894,
         n39895, n39896, n39897, n39898, n39899, n39900, n39901, n39902,
         n39903, n39904, n39905, n39906, n39907, n39908, n39909, n39910,
         n39911, n39912, n39913, n39914, n39915, n39916, n39917, n39918,
         n39919, n39920, n39921, n39922, n39923, n39924, n39925, n39926,
         n39927, n39928, n39929, n39930, n39931, n39932, n39933, n39934,
         n39935, n39936, n39937, n39938, n39939, n39940, n39941, n39942,
         n39943, n39944, n39945, n39946, n39947, n39948, n39949, n39950,
         n39951, n39952, n39953, n39954, n39955, n39956, n39957, n39958,
         n39959, n39960, n39961, n39962, n39963, n39964, n39965, n39966,
         n39967, n39968, n39969, n39970, n39971, n39972, n39973, n39974,
         n39975, n39976, n39977, n39978, n39979, n39980, n39981, n39982,
         n39983, n39984, n39985, n39986, n39987, n39988, n39989, n39990,
         n39991, n39992, n39993, n39994, n39995, n39996, n39997, n39998,
         n39999, n40000, n40001, n40002, n40003, n40004, n40005, n40006,
         n40007, n40008, n40009, n40010, n40011, n40012, n40013, n40014,
         n40015, n40016, n40017, n40018, n40019, n40020, n40021, n40022,
         n40023, n40024, n40025, n40026, n40027, n40028, n40029, n40030,
         n40031, n40032, n40033, n40034, n40035, n40036, n40037, n40038,
         n40039, n40040, n40041, n40042, n40043, n40044, n40045, n40046,
         n40047, n40048, n40049, n40050, n40051, n40052, n40053, n40054,
         n40055, n40056, n40057, n40058, n40059, n40060, n40061, n40062,
         n40063, n40064, n40065, n40066, n40067, n40068, n40069, n40070,
         n40071, n40072, n40073, n40074, n40075, n40076, n40077, n40078,
         n40079, n40080, n40081, n40082, n40083, n40084, n40085, n40086,
         n40087, n40088, n40089, n40090, n40091, n40092, n40093, n40094,
         n40095, n40096, n40097, n40098, n40099, n40100, n40101, n40102,
         n40103, n40104, n40105, n40106, n40107, n40108, n40109, n40110,
         n40111, n40112, n40113, n40114, n40115, n40116, n40117, n40118,
         n40119, n40120, n40121, n40122, n40123, n40124, n40125, n40126,
         n40127, n40128, n40129, n40130, n40131, n40132, n40133, n40134,
         n40135, n40136, n40137, n40138, n40139, n40140, n40141, n40142,
         n40143, n40144, n40145, n40146, n40147, n40148, n40149, n40150,
         n40151, n40152, n40153, n40154, n40155, n40156, n40157, n40158,
         n40159, n40160, n40161, n40162, n40163, n40164, n40165, n40166,
         n40167, n40168, n40169, n40170, n40171, n40172, n40173, n40174,
         n40175, n40176, n40177, n40178, n40179, n40180, n40181, n40182,
         n40183, n40184, n40185, n40186, n40187, n40188, n40189, n40190,
         n40191, n40192, n40193, n40194, n40195, n40196, n40197, n40198,
         n40199, n40200, n40201, n40202, n40203, n40204, n40205, n40206,
         n40207, n40208, n40209, n40210, n40211, n40212, n40213, n40214,
         n40215, n40216, n40217, n40218, n40219, n40220, n40221, n40222,
         n40223, n40224, n40225, n40226, n40227, n40228, n40229, n40230,
         n40231, n40232, n40233, n40234, n40235, n40236, n40237, n40238,
         n40239, n40240, n40241, n40242, n40243, n40244, n40245, n40246,
         n40247, n40248, n40249, n40250, n40251, n40252, n40253, n40254,
         n40255, n40256, n40257, n40258, n40259, n40260, n40261, n40262,
         n40263, n40264, n40265, n40266, n40267, n40268, n40269, n40270,
         n40271, n40272, n40273, n40274, n40275, n40276, n40277, n40278,
         n40279, n40280, n40281, n40282, n40283, n40284, n40285, n40286,
         n40287, n40288, n40289, n40290, n40291, n40292, n40293, n40294,
         n40295, n40296, n40297, n40298, n40299, n40300, n40301, n40302,
         n40303, n40304, n40305, n40306, n40307, n40308, n40309, n40310,
         n40311, n40312, n40313, n40314, n40315, n40316, n40317, n40318,
         n40319, n40320, n40321, n40322, n40323, n40324, n40325, n40326,
         n40327, n40328, n40329, n40330, n40331, n40332, n40333, n40334,
         n40335, n40336, n40337, n40338, n40339, n40340, n40341, n40342,
         n40343, n40344, n40345, n40346, n40347, n40348, n40349, n40350,
         n40351, n40352, n40353, n40354, n40355, n40356, n40357, n40358,
         n40359, n40360, n40361, n40362, n40363, n40364, n40365, n40366,
         n40367, n40368, n40369, n40370, n40371, n40372, n40373, n40374,
         n40375, n40376, n40377, n40378, n40379, n40380, n40381, n40382,
         n40383, n40384, n40385, n40386, n40387, n40388, n40389, n40390,
         n40391, n40392, n40393, n40394, n40395, n40396, n40397, n40398,
         n40399, n40400, n40401, n40402, n40403, n40404, n40405, n40406,
         n40407, n40408, n40409, n40410, n40411, n40412, n40413, n40414,
         n40415, n40416, n40417, n40418, n40419, n40420, n40421, n40422,
         n40423, n40424, n40425, n40426, n40427, n40428, n40429, n40430,
         n40431, n40432, n40433, n40434, n40435, n40436, n40437, n40438,
         n40439, n40440, n40441, n40442, n40443, n40444, n40445, n40446,
         n40447, n40448, n40449, n40450, n40451, n40452, n40453, n40454,
         n40455, n40456, n40457, n40458, n40459, n40460, n40461, n40462,
         n40463, n40464, n40465, n40466, n40467, n40468, n40469, n40470,
         n40471, n40472, n40473, n40474, n40475, n40476, n40477, n40478,
         n40479, n40480, n40481, n40482, n40483, n40484, n40485, n40486,
         n40487, n40488, n40489, n40490, n40491, n40492, n40493, n40494,
         n40495, n40496, n40497, n40498, n40499, n40500, n40501, n40502,
         n40503, n40504, n40505, n40506, n40507, n40508, n40509, n40510,
         n40511, n40512, n40513, n40514, n40515, n40516, n40517, n40518,
         n40519, n40520, n40521, n40522, n40523, n40524, n40525, n40526,
         n40527, n40528, n40529, n40530, n40531, n40532, n40533, n40534,
         n40535, n40536, n40537, n40538, n40539, n40540, n40541, n40542,
         n40543, n40544, n40545, n40546, n40547, n40548, n40549, n40550,
         n40551, n40552, n40553, n40554, n40555, n40556, n40557, n40558,
         n40559, n40560, n40561, n40562, n40563, n40564, n40565, n40566,
         n40567, n40568, n40569, n40570, n40571, n40572, n40573, n40574,
         n40575, n40576, n40577, n40578, n40579, n40580, n40581, n40582,
         n40583, n40584, n40585, n40586, n40587, n40588, n40589, n40590,
         n40591, n40592, n40593, n40594, n40595, n40596, n40597, n40598,
         n40599, n40600, n40601, n40602, n40603, n40604, n40605, n40606,
         n40607, n40608, n40609, n40610, n40611, n40612, n40613, n40614,
         n40615, n40616, n40617, n40618, n40619, n40620, n40621, n40622,
         n40623, n40624, n40625, n40626, n40627, n40628, n40629, n40630,
         n40631, n40632, n40633, n40634, n40635, n40636, n40637, n40638,
         n40639, n40640, n40641, n40642, n40643, n40644, n40645, n40646,
         n40647, n40648, n40649, n40650, n40651, n40652, n40653, n40654,
         n40655, n40656, n40657, n40658, n40659, n40660, n40661, n40662,
         n40663, n40664, n40665, n40666, n40667, n40668, n40669, n40670,
         n40671, n40672, n40673, n40674, n40675, n40676, n40677, n40678,
         n40679, n40680, n40681, n40682, n40683, n40684, n40685, n40686,
         n40687, n40688, n40689, n40690, n40691, n40692, n40693, n40694,
         n40695, n40696, n40697, n40698, n40699, n40700, n40701, n40702,
         n40703, n40704, n40705, n40706, n40707, n40708, n40709, n40710,
         n40711, n40712, n40713, n40714, n40715, n40716, n40717, n40718,
         n40719, n40720, n40721, n40722, n40723, n40724, n40725, n40726,
         n40727, n40728, n40729, n40730, n40731, n40732, n40733, n40734,
         n40735, n40736, n40737, n40738, n40739, n40740, n40741, n40742,
         n40743, n40744, n40745, n40746, n40747, n40748, n40749, n40750,
         n40751, n40752, n40753, n40754, n40755, n40756, n40757, n40758,
         n40759, n40760, n40761, n40762, n40763, n40764, n40765, n40766,
         n40767, n40768, n40769, n40770, n40771, n40772, n40773, n40774,
         n40775, n40776, n40777, n40778, n40779, n40780, n40781, n40782,
         n40783, n40784, n40785, n40786, n40787, n40788, n40789, n40790,
         n40791, n40792, n40793, n40794, n40795, n40796, n40797, n40798,
         n40799, n40800, n40801, n40802, n40803, n40804, n40805, n40806,
         n40807, n40808, n40809, n40810, n40811, n40812, n40813, n40814,
         n40815, n40816, n40817, n40818, n40819, n40820, n40821, n40822,
         n40823, n40824, n40825, n40826, n40827, n40828, n40829, n40830,
         n40831, n40832, n40833, n40834, n40835, n40836, n40837, n40838,
         n40839, n40840, n40841, n40842, n40843, n40844, n40845, n40846,
         n40847, n40848, n40849, n40850, n40851, n40852, n40853, n40854,
         n40855, n40856, n40857, n40858, n40859, n40860, n40861, n40862,
         n40863, n40864, n40865, n40866, n40867, n40868, n40869, n40870,
         n40871, n40872, n40873, n40874, n40875, n40876, n40877, n40878,
         n40879, n40880, n40881, n40882, n40883, n40884, n40885, n40886,
         n40887, n40888, n40889, n40890, n40891, n40892, n40893, n40894,
         n40895, n40896, n40897, n40898, n40899, n40900, n40901, n40902,
         n40903, n40904, n40905, n40906, n40907, n40908, n40909, n40910,
         n40911, n40912, n40913, n40914, n40915, n40916, n40917, n40918,
         n40919, n40920, n40921, n40922, n40923, n40924, n40925, n40926,
         n40927, n40928, n40929, n40930, n40931, n40932, n40933, n40934,
         n40935, n40936, n40937, n40938, n40939, n40940, n40941, n40942,
         n40943, n40944, n40945, n40946, n40947, n40948, n40949, n40950,
         n40951, n40952, n40953, n40954, n40955, n40956, n40957, n40958,
         n40959, n40960, n40961, n40962, n40963, n40964, n40965, n40966,
         n40967, n40968, n40969, n40970, n40971, n40972, n40973, n40974,
         n40975, n40976, n40977, n40978, n40979, n40980, n40981, n40982,
         n40983, n40984, n40985, n40986, n40987, n40988, n40989, n40990,
         n40991, n40992, n40993, n40994, n40995, n40996, n40997, n40998,
         n40999, n41000, n41001, n41002, n41003, n41004, n41005, n41006,
         n41007, n41008, n41009, n41010, n41011, n41012, n41013, n41014,
         n41015, n41016, n41017, n41018, n41019, n41020, n41021, n41022,
         n41023, n41024, n41025, n41026, n41027, n41028, n41029, n41030,
         n41031, n41032, n41033, n41034, n41035, n41036, n41037, n41038,
         n41039, n41040, n41041, n41042, n41043, n41044, n41045, n41046,
         n41047, n41048, n41049, n41050, n41051, n41052, n41053, n41054,
         n41055, n41056, n41057, n41058, n41059, n41060, n41061, n41062,
         n41063, n41064, n41065, n41066, n41067, n41068, n41069, n41070,
         n41071, n41072, n41073, n41074, n41075, n41076, n41077, n41078,
         n41079, n41080, n41081, n41082, n41083, n41084, n41085, n41086,
         n41087, n41088, n41089, n41090, n41091, n41092, n41093, n41094,
         n41095, n41096, n41097, n41098, n41099, n41100, n41101, n41102,
         n41103, n41104, n41105, n41106, n41107, n41108, n41109, n41110,
         n41111, n41112, n41113, n41114, n41115, n41116, n41117, n41118,
         n41119, n41120, n41121, n41122, n41123, n41124, n41125, n41126,
         n41127, n41128, n41129, n41130, n41131, n41132, n41133, n41134,
         n41135, n41136, n41137, n41138, n41139, n41140, n41141, n41142,
         n41143, n41144, n41145, n41146, n41147, n41148, n41149, n41150,
         n41151, n41152, n41153, n41154, n41155, n41156, n41157, n41158,
         n41159, n41160, n41161, n41162, n41163, n41164, n41165, n41166,
         n41167, n41168, n41169, n41170, n41171, n41172, n41173, n41174,
         n41175, n41176, n41177, n41178, n41179, n41180, n41181, n41182,
         n41183, n41184, n41185, n41186, n41187, n41188, n41189, n41190,
         n41191, n41192, n41193, n41194, n41195, n41196, n41197, n41198,
         n41199, n41200, n41201, n41202, n41203, n41204, n41205, n41206,
         n41207, n41208, n41209, n41210, n41211, n41212, n41213, n41214,
         n41215, n41216, n41217, n41218, n41219, n41220, n41221, n41222,
         n41223, n41224, n41225, n41226, n41227, n41228, n41229, n41230,
         n41231, n41232, n41233, n41234, n41235, n41236, n41237, n41238,
         n41239, n41240, n41241, n41242, n41243, n41244, n41245, n41246,
         n41247, n41248, n41249, n41250, n41251, n41252, n41253, n41254,
         n41255, n41256, n41257, n41258, n41259, n41260, n41261, n41262,
         n41263, n41264, n41265, n41266, n41267, n41268, n41269, n41270,
         n41271, n41272, n41273, n41274, n41275, n41276, n41277, n41278,
         n41279, n41280, n41281, n41282, n41283, n41284, n41285, n41286,
         n41287, n41288, n41289, n41290, n41291, n41292, n41293, n41294,
         n41295, n41296, n41297, n41298, n41299, n41300, n41301, n41302,
         n41303, n41304, n41305, n41306, n41307, n41308, n41309, n41310,
         n41311, n41312, n41313, n41314, n41315, n41316, n41317, n41318,
         n41319, n41320, n41321, n41322, n41323, n41324, n41325, n41326,
         n41327, n41328, n41329, n41330, n41331, n41332, n41333, n41334,
         n41335, n41336, n41337, n41338, n41339, n41340, n41341, n41342,
         n41343, n41344, n41345, n41346, n41347, n41348, n41349, n41350,
         n41351, n41352, n41353, n41354, n41355, n41356, n41357, n41358,
         n41359, n41360, n41361, n41362, n41363, n41364, n41365, n41366,
         n41367, n41368, n41369, n41370, n41371, n41372, n41373, n41374,
         n41375, n41376, n41377, n41378, n41379, n41380, n41381, n41382,
         n41383, n41384, n41385, n41386, n41387, n41388, n41389, n41390,
         n41391, n41392, n41393, n41394, n41395, n41396, n41397, n41398,
         n41399, n41400, n41401, n41402, n41403, n41404, n41405, n41406,
         n41407, n41408, n41409, n41410, n41411, n41412, n41413, n41414,
         n41415, n41416, n41417, n41418, n41419, n41420, n41421, n41422,
         n41423, n41424, n41425, n41426, n41427, n41428, n41429, n41430,
         n41431, n41432, n41433, n41434, n41435, n41436, n41437, n41438,
         n41439, n41440, n41441, n41442, n41443, n41444, n41445, n41446,
         n41447, n41448, n41449, n41450, n41451, n41452, n41453, n41454,
         n41455, n41456, n41457, n41458, n41459, n41460, n41461, n41462,
         n41463, n41464, n41465, n41466, n41467, n41468, n41469, n41470,
         n41471, n41472, n41473, n41474, n41475, n41476, n41477, n41478,
         n41479, n41480, n41481, n41482, n41483, n41484, n41485, n41486,
         n41487, n41488, n41489, n41490, n41491, n41492, n41493, n41494,
         n41495, n41496, n41497, n41498, n41499, n41500, n41501, n41502,
         n41503, n41504, n41505, n41506, n41507, n41508, n41509, n41510,
         n41511, n41512, n41513, n41514, n41515, n41516, n41517, n41518,
         n41519, n41520, n41521, n41522, n41523, n41524, n41525, n41526,
         n41527, n41528, n41529, n41530, n41531, n41532, n41533, n41534,
         n41535, n41536, n41537, n41538, n41539, n41540, n41541, n41542,
         n41543, n41544, n41545, n41546, n41547, n41548, n41549, n41550,
         n41551, n41552, n41553, n41554, n41555, n41556, n41557, n41558,
         n41559, n41560, n41561, n41562, n41563, n41564, n41565, n41566,
         n41567, n41568, n41569, n41570, n41571, n41572, n41573, n41574,
         n41575, n41576, n41577, n41578, n41579, n41580, n41581, n41582,
         n41583, n41584, n41585, n41586, n41587, n41588, n41589, n41590,
         n41591, n41592, n41593, n41594, n41595, n41596, n41597, n41598,
         n41599, n41600, n41601, n41602, n41603, n41604, n41605, n41606,
         n41607, n41608, n41609, n41610, n41611, n41612, n41613, n41614,
         n41615, n41616, n41617, n41618, n41619, n41620, n41621, n41622,
         n41623, n41624, n41625, n41626, n41627, n41628, n41629, n41630,
         n41631, n41632, n41633, n41634, n41635, n41636, n41637, n41638,
         n41639, n41640, n41641, n41642, n41643, n41644, n41645, n41646,
         n41647, n41648, n41649, n41650, n41651, n41652, n41653, n41654,
         n41655, n41656, n41657, n41658, n41659, n41660, n41661, n41662,
         n41663, n41664, n41665, n41666, n41667, n41668, n41669, n41670,
         n41671, n41672, n41673, n41674, n41675, n41676, n41677, n41678,
         n41679, n41680, n41681, n41682, n41683, n41684, n41685, n41686,
         n41687, n41688, n41689, n41690, n41691, n41692, n41693, n41694,
         n41695, n41696, n41697, n41698, n41699, n41700, n41701, n41702,
         n41703, n41704, n41705, n41706, n41707, n41708, n41709, n41710,
         n41711, n41712, n41713, n41714, n41715, n41716, n41717, n41718,
         n41719, n41720, n41721, n41722, n41723, n41724, n41725, n41726,
         n41727, n41728, n41729, n41730, n41731, n41732, n41733, n41734,
         n41735, n41736, n41737, n41738, n41739, n41740, n41741, n41742,
         n41743, n41744, n41745, n41746, n41747, n41748, n41749, n41750,
         n41751, n41752, n41753, n41754, n41755, n41756, n41757, n41758,
         n41759, n41760, n41761, n41762, n41763, n41764, n41765, n41766,
         n41767, n41768, n41769, n41770, n41771, n41772, n41773, n41774,
         n41775, n41776, n41777, n41778, n41779, n41780, n41781, n41782,
         n41783, n41784, n41785, n41786, n41787, n41788, n41789, n41790,
         n41791, n41792, n41793, n41794, n41795, n41796, n41797, n41798,
         n41799, n41800, n41801, n41802, n41803, n41804, n41805, n41806,
         n41807, n41808, n41809, n41810, n41811, n41812, n41813, n41814,
         n41815, n41816, n41817, n41818, n41819, n41820, n41821, n41822,
         n41823, n41824, n41825, n41826, n41827, n41828, n41829, n41830,
         n41831, n41832, n41833, n41834, n41835, n41836, n41837, n41838,
         n41839, n41840, n41841, n41842, n41843, n41844, n41845, n41846,
         n41847, n41848, n41849, n41850, n41851, n41852, n41853, n41854,
         n41855, n41856, n41857, n41858, n41859, n41860, n41861, n41862,
         n41863, n41864, n41865, n41866, n41867, n41868, n41869, n41870,
         n41871, n41872, n41873, n41874, n41875, n41876, n41877, n41878,
         n41879, n41880, n41881, n41882, n41883, n41884, n41885, n41886,
         n41887, n41888, n41889, n41890, n41891, n41892, n41893, n41894,
         n41895, n41896, n41897, n41898, n41899, n41900, n41901, n41902,
         n41903, n41904, n41905, n41906, n41907, n41908, n41909, n41910,
         n41911, n41912, n41913, n41914, n41915, n41916, n41917, n41918,
         n41919, n41920, n41921, n41922, n41923, n41924, n41925, n41926,
         n41927, n41928, n41929, n41930, n41931, n41932, n41933, n41934,
         n41935, n41936, n41937, n41938, n41939, n41940, n41941, n41942,
         n41943, n41944, n41945, n41946, n41947, n41948, n41949, n41950,
         n41951, n41952, n41953, n41954, n41955, n41956, n41957, n41958,
         n41959, n41960, n41961, n41962, n41963, n41964, n41965, n41966,
         n41967, n41968, n41969, n41970, n41971, n41972, n41973, n41974,
         n41975, n41976, n41977, n41978, n41979, n41980, n41981, n41982,
         n41983, n41984, n41985, n41986, n41987, n41988, n41989, n41990,
         n41991, n41992, n41993, n41994, n41995, n41996, n41997, n41998,
         n41999, n42000, n42001, n42002, n42003, n42004, n42005, n42006,
         n42007, n42008, n42009, n42010, n42011, n42012, n42013, n42014,
         n42015, n42016, n42017, n42018, n42019, n42020, n42021, n42022,
         n42023, n42024, n42025, n42026, n42027, n42028, n42029, n42030,
         n42031, n42032, n42033, n42034, n42035, n42036, n42037, n42038,
         n42039, n42040, n42041, n42042, n42043, n42044, n42045, n42046,
         n42047, n42048, n42049, n42050, n42051, n42052, n42053, n42054,
         n42055, n42056, n42057, n42058, n42059, n42060, n42061, n42062,
         n42063, n42064, n42065, n42066, n42067, n42068, n42069, n42070,
         n42071, n42072, n42073, n42074, n42075, n42076, n42077, n42078,
         n42079, n42080, n42081, n42082, n42083, n42084, n42085, n42086,
         n42087, n42088, n42089, n42090, n42091, n42092, n42093, n42094,
         n42095, n42096, n42097, n42098, n42099, n42100, n42101, n42102,
         n42103, n42104, n42105, n42106, n42107, n42108, n42109, n42110,
         n42111, n42112, n42113, n42114, n42115, n42116, n42117, n42118,
         n42119, n42120, n42121, n42122, n42123, n42124, n42125, n42126,
         n42127, n42128, n42129, n42130, n42131, n42132, n42133, n42134,
         n42135, n42136, n42137, n42138, n42139, n42140, n42141, n42142,
         n42143, n42144, n42145, n42146, n42147, n42148, n42149, n42150,
         n42151, n42152, n42153, n42154, n42155, n42156, n42157, n42158,
         n42159, n42160, n42161, n42162, n42163, n42164, n42165, n42166,
         n42167, n42168, n42169, n42170, n42171, n42172, n42173, n42174,
         n42175, n42176, n42177, n42178, n42179, n42180, n42181, n42182,
         n42183, n42184, n42185, n42186, n42187, n42188, n42189, n42190,
         n42191, n42192, n42193, n42194, n42195, n42196, n42197, n42198,
         n42199, n42200, n42201, n42202, n42203, n42204, n42205, n42206,
         n42207, n42208, n42209, n42210, n42211, n42212, n42213, n42214,
         n42215, n42216, n42217, n42218, n42219, n42220, n42221, n42222,
         n42223, n42224, n42225, n42226, n42227, n42228, n42229, n42230,
         n42231, n42232, n42233, n42234, n42235, n42236, n42237, n42238,
         n42239, n42240, n42241, n42242, n42243, n42244, n42245, n42246,
         n42247, n42248, n42249, n42250, n42251, n42252, n42253, n42254,
         n42255, n42256, n42257, n42258, n42259, n42260, n42261, n42262,
         n42263, n42264, n42265, n42266, n42267, n42268, n42269, n42270,
         n42271, n42272, n42273, n42274, n42275, n42276, n42277, n42278,
         n42279, n42280, n42281, n42282, n42283, n42284, n42285, n42286,
         n42287, n42288, n42289, n42290, n42291, n42292, n42293, n42294,
         n42295, n42296, n42297, n42298, n42299, n42300, n42301, n42302,
         n42303, n42304, n42305, n42306, n42307, n42308, n42309, n42310,
         n42311, n42312, n42313, n42314, n42315, n42316, n42317, n42318,
         n42319, n42320, n42321, n42322, n42323, n42324, n42325, n42326,
         n42327, n42328, n42329, n42330, n42331, n42332, n42333, n42334,
         n42335, n42336, n42337, n42338, n42339, n42340, n42341, n42342,
         n42343, n42344, n42345, n42346, n42347, n42348, n42349, n42350,
         n42351, n42352, n42353, n42354, n42355, n42356, n42357, n42358,
         n42359, n42360, n42361, n42362, n42363, n42364, n42365, n42366,
         n42367, n42368, n42369, n42370, n42371, n42372, n42373, n42374,
         n42375, n42376, n42377, n42378, n42379, n42380, n42381, n42382,
         n42383, n42384, n42385, n42386, n42387, n42388, n42389, n42390,
         n42391, n42392, n42393, n42394, n42395, n42396, n42397, n42398,
         n42399, n42400, n42401, n42402, n42403, n42404, n42405, n42406,
         n42407, n42408, n42409, n42410, n42411, n42412, n42413, n42414,
         n42415, n42416, n42417, n42418, n42419, n42420, n42421, n42422,
         n42423, n42424, n42425, n42426, n42427, n42428, n42429, n42430,
         n42431, n42432, n42433, n42434, n42435, n42436, n42437, n42438,
         n42439, n42440, n42441, n42442, n42443, n42444, n42445, n42446,
         n42447, n42448, n42449, n42450, n42451, n42452, n42453, n42454,
         n42455, n42456, n42457, n42458, n42459, n42460, n42461, n42462,
         n42463, n42464, n42465, n42466, n42467, n42468, n42469, n42470,
         n42471, n42472, n42473, n42474, n42475, n42476, n42477, n42478,
         n42479, n42480, n42481, n42482, n42483, n42484, n42485, n42486,
         n42487, n42488, n42489, n42490, n42491, n42492, n42493, n42494,
         n42495, n42496, n42497, n42498, n42499, n42500, n42501, n42502,
         n42503, n42504, n42505, n42506, n42507, n42508, n42509, n42510,
         n42511, n42512, n42513, n42514, n42515, n42516, n42517, n42518,
         n42519, n42520, n42521, n42522, n42523, n42524, n42525, n42526,
         n42527, n42528, n42529, n42530, n42531, n42532, n42533, n42534,
         n42535, n42536, n42537, n42538, n42539, n42540, n42541, n42542,
         n42543, n42544, n42545, n42546, n42547, n42548, n42549, n42550,
         n42551, n42552, n42553, n42554, n42555, n42556, n42557, n42558,
         n42559, n42560, n42561, n42562, n42563, n42564, n42565, n42566,
         n42567, n42568, n42569, n42570, n42571, n42572, n42573, n42574,
         n42575, n42576, n42577, n42578, n42579, n42580, n42581, n42582,
         n42583, n42584, n42585, n42586, n42587, n42588, n42589, n42590,
         n42591, n42592, n42593, n42594, n42595, n42596, n42597, n42598,
         n42599, n42600, n42601, n42602, n42603, n42604, n42605, n42606,
         n42607, n42608, n42609, n42610, n42611, n42612, n42613, n42614,
         n42615, n42616, n42617, n42618, n42619, n42620, n42621, n42622,
         n42623, n42624, n42625, n42626, n42627, n42628, n42629, n42630,
         n42631, n42632, n42633, n42634, n42635, n42636, n42637, n42638,
         n42639, n42640, n42641, n42642, n42643, n42644, n42645, n42646,
         n42647, n42648, n42649, n42650, n42651, n42652, n42653, n42654,
         n42655, n42656, n42657, n42658, n42659, n42660, n42661, n42662,
         n42663, n42664, n42665, n42666, n42667, n42668, n42669, n42670,
         n42671, n42672, n42673, n42674, n42675, n42676, n42677, n42678,
         n42679, n42680, n42681, n42682, n42683, n42684, n42685, n42686,
         n42687, n42688, n42689, n42690, n42691, n42692, n42693, n42694,
         n42695, n42696, n42697, n42698, n42699, n42700, n42701, n42702,
         n42703, n42704, n42705, n42706, n42707, n42708, n42709, n42710,
         n42711, n42712, n42713, n42714, n42715, n42716, n42717, n42718,
         n42719, n42720, n42721, n42722, n42723, n42724, n42725, n42726,
         n42727, n42728, n42729, n42730, n42731, n42732, n42733, n42734,
         n42735, n42736, n42737, n42738, n42739, n42740, n42741, n42742,
         n42743, n42744, n42745, n42746, n42747, n42748, n42749, n42750,
         n42751, n42752, n42753, n42754, n42755, n42756, n42757, n42758,
         n42759, n42760, n42761, n42762, n42763, n42764, n42765, n42766,
         n42767, n42768, n42769, n42770, n42771, n42772, n42773, n42774,
         n42775, n42776, n42777, n42778, n42779, n42780, n42781, n42782,
         n42783, n42784, n42785, n42786, n42787, n42788, n42789, n42790,
         n42791, n42792, n42793, n42794, n42795, n42796, n42797, n42798,
         n42799, n42800, n42801, n42802, n42803, n42804, n42805, n42806,
         n42807, n42808, n42809, n42810, n42811, n42812, n42813, n42814,
         n42815, n42816, n42817, n42818, n42819, n42820, n42821, n42822,
         n42823, n42824, n42825, n42826, n42827, n42828, n42829, n42830,
         n42831, n42832, n42833, n42834, n42835, n42836, n42837, n42838,
         n42839, n42840, n42841, n42842, n42843, n42844, n42845, n42846,
         n42847, n42848, n42849, n42850, n42851, n42852, n42853, n42854,
         n42855, n42856, n42857, n42858, n42859, n42860, n42861, n42862,
         n42863, n42864, n42865, n42866, n42867, n42868, n42869, n42870,
         n42871, n42872, n42873, n42874, n42875, n42876, n42877, n42878,
         n42879, n42880, n42881, n42882, n42883, n42884, n42885, n42886,
         n42887, n42888, n42889, n42890, n42891, n42892, n42893, n42894,
         n42895, n42896, n42897, n42898, n42899, n42900, n42901, n42902,
         n42903, n42904, n42905, n42906, n42907, n42908, n42909, n42910,
         n42911, n42912, n42913, n42914, n42915, n42916, n42917, n42918,
         n42919, n42920, n42921, n42922, n42923, n42924, n42925, n42926,
         n42927, n42928, n42929, n42930, n42931, n42932, n42933, n42934,
         n42935, n42936, n42937, n42938, n42939, n42940, n42941, n42942,
         n42943, n42944, n42945, n42946, n42947, n42948, n42949, n42950,
         n42951, n42952, n42953, n42954, n42955, n42956, n42957, n42958,
         n42959, n42960, n42961, n42962, n42963, n42964, n42965, n42966,
         n42967, n42968, n42969, n42970, n42971, n42972, n42973, n42974,
         n42975, n42976, n42977, n42978, n42979, n42980, n42981, n42982,
         n42983, n42984, n42985, n42986, n42987, n42988, n42989, n42990,
         n42991, n42992, n42993, n42994, n42995, n42996, n42997, n42998,
         n42999, n43000, n43001, n43002, n43003, n43004, n43005, n43006,
         n43007, n43008, n43009, n43010, n43011, n43012, n43013, n43014,
         n43015, n43016, n43017, n43018, n43019, n43020, n43021, n43022,
         n43023, n43024, n43025, n43026, n43027, n43028, n43029, n43030,
         n43031, n43032, n43033, n43034, n43035, n43036, n43037, n43038,
         n43039, n43040, n43041, n43042, n43043, n43044, n43045, n43046,
         n43047, n43048, n43049, n43050, n43051, n43052, n43053, n43054,
         n43055, n43056, n43057, n43058, n43059, n43060, n43061, n43062,
         n43063, n43064, n43065, n43066, n43067, n43068, n43069, n43070,
         n43071, n43072, n43073, n43074, n43075, n43076, n43077, n43078,
         n43079, n43080, n43081, n43082, n43083, n43084, n43085, n43086,
         n43087, n43088, n43089, n43090, n43091, n43092, n43093, n43094,
         n43095, n43096, n43097, n43098, n43099, n43100, n43101, n43102,
         n43103, n43104, n43105, n43106, n43107, n43108, n43109, n43110,
         n43111, n43112, n43113, n43114, n43115, n43116, n43117, n43118,
         n43119, n43120, n43121, n43122, n43123, n43124, n43125, n43126,
         n43127, n43128, n43129, n43130, n43131, n43132, n43133, n43134,
         n43135, n43136, n43137, n43138, n43139, n43140, n43141, n43142,
         n43143, n43144, n43145, n43146, n43147, n43148, n43149, n43150,
         n43151, n43152, n43153, n43154, n43155, n43156, n43157, n43158,
         n43159, n43160, n43161, n43162, n43163, n43164, n43165, n43166,
         n43167, n43168, n43169, n43170, n43171, n43172, n43173, n43174,
         n43175, n43176, n43177, n43178, n43179, n43180, n43181, n43182,
         n43183, n43184, n43185, n43186, n43187, n43188, n43189, n43190,
         n43191, n43192, n43193, n43194, n43195, n43196, n43197, n43198,
         n43199, n43200, n43201, n43202, n43203, n43204, n43205, n43206,
         n43207, n43208, n43209, n43210, n43211, n43212, n43213, n43214,
         n43215, n43216, n43217, n43218, n43219, n43220, n43221, n43222,
         n43223, n43224, n43225, n43226, n43227, n43228, n43229, n43230,
         n43231, n43232, n43233, n43234, n43235, n43236, n43237, n43238,
         n43239, n43240, n43241, n43242, n43243, n43244, n43245, n43246,
         n43247, n43248, n43249, n43250, n43251, n43252, n43253, n43254,
         n43255, n43256, n43257, n43258, n43259, n43260, n43261, n43262,
         n43263, n43264, n43265, n43266, n43267, n43268, n43269, n43270,
         n43271, n43272, n43273, n43274, n43275, n43276, n43277, n43278,
         n43279, n43280, n43281, n43282, n43283, n43284, n43285, n43286,
         n43287, n43288, n43289, n43290, n43291, n43292, n43293, n43294,
         n43295, n43296, n43297, n43298, n43299, n43300, n43301, n43302,
         n43303, n43304, n43305, n43306, n43307, n43308, n43309, n43310,
         n43311, n43312, n43313, n43314, n43315, n43316, n43317, n43318,
         n43319, n43320, n43321, n43322, n43323, n43324, n43325, n43326,
         n43327, n43328, n43329, n43330, n43331, n43332, n43333, n43334,
         n43335, n43336, n43337, n43338, n43339, n43340, n43341, n43342,
         n43343, n43344, n43345, n43346, n43347, n43348, n43349, n43350,
         n43351, n43352, n43353, n43354, n43355, n43356, n43357, n43358,
         n43359, n43360, n43361, n43362, n43363, n43364, n43365, n43366,
         n43367, n43368, n43369, n43370, n43371, n43372, n43373, n43374,
         n43375, n43376, n43377, n43378, n43379, n43380, n43381, n43382,
         n43383, n43384, n43385, n43386, n43387, n43388, n43389, n43390,
         n43391, n43392, n43393, n43394, n43395, n43396, n43397, n43398,
         n43399, n43400, n43401, n43402, n43403, n43404, n43405, n43406,
         n43407, n43408, n43409, n43410, n43411, n43412, n43413, n43414,
         n43415, n43416, n43417, n43418, n43419, n43420, n43421, n43422,
         n43423, n43424, n43425, n43426, n43427, n43428, n43429, n43430,
         n43431, n43432, n43433, n43434, n43435, n43436, n43437, n43438,
         n43439, n43440, n43441, n43442, n43443, n43444, n43445, n43446,
         n43447, n43448, n43449, n43450, n43451, n43452, n43453, n43454,
         n43455, n43456, n43457, n43458, n43459, n43460, n43461, n43462,
         n43463, n43464, n43465, n43466, n43467, n43468, n43469, n43470,
         n43471, n43472, n43473, n43474, n43475, n43476, n43477, n43478,
         n43479, n43480, n43481, n43482, n43483, n43484, n43485, n43486,
         n43487, n43488, n43489, n43490, n43491, n43492, n43493, n43494,
         n43495, n43496, n43497, n43498, n43499, n43500, n43501, n43502,
         n43503, n43504, n43505, n43506, n43507, n43508, n43509, n43510,
         n43511, n43512, n43513, n43514, n43515, n43516, n43517, n43518,
         n43519, n43520, n43521, n43522, n43523, n43524, n43525, n43526,
         n43527, n43528, n43529, n43530, n43531, n43532, n43533, n43534,
         n43535, n43536, n43537, n43538, n43539, n43540, n43541, n43542,
         n43543, n43544, n43545, n43546, n43547, n43548, n43549, n43550,
         n43551, n43552, n43553, n43554, n43555, n43556, n43557, n43558,
         n43559, n43560, n43561, n43562, n43563, n43564, n43565, n43566,
         n43567, n43568, n43569, n43570, n43571, n43572, n43573, n43574,
         n43575, n43576, n43577, n43578, n43579, n43580, n43581, n43582,
         n43583, n43584, n43585, n43586, n43587, n43588, n43589, n43590,
         n43591, n43592, n43593, n43594, n43595, n43596, n43597, n43598,
         n43599, n43600, n43601, n43602, n43603, n43604, n43605, n43606,
         n43607, n43608, n43609, n43610, n43611, n43612, n43613, n43614,
         n43615, n43616, n43617, n43618, n43619, n43620, n43621, n43622,
         n43623, n43624, n43625, n43626, n43627, n43628, n43629, n43630,
         n43631, n43632, n43633, n43634, n43635, n43636, n43637, n43638,
         n43639, n43640, n43641, n43642, n43643, n43644, n43645, n43646,
         n43647, n43648, n43649, n43650, n43651, n43652, n43653, n43654,
         n43655, n43656, n43657, n43658, n43659, n43660, n43661, n43662,
         n43663, n43664, n43665, n43666, n43667, n43668, n43669, n43670,
         n43671, n43672, n43673, n43674, n43675, n43676, n43677, n43678,
         n43679, n43680, n43681, n43682, n43683, n43684, n43685, n43686,
         n43687, n43688, n43689, n43690, n43691, n43692, n43693, n43694,
         n43695, n43696, n43697, n43698, n43699, n43700, n43701, n43702,
         n43703, n43704, n43705, n43706, n43707, n43708, n43709, n43710,
         n43711, n43712, n43713, n43714, n43715, n43716, n43717, n43718,
         n43719, n43720, n43721, n43722, n43723, n43724, n43725, n43726,
         n43727, n43728, n43729, n43730, n43731, n43732, n43733, n43734,
         n43735, n43736, n43737, n43738, n43739, n43740, n43741, n43742,
         n43743, n43744, n43745, n43746, n43747, n43748, n43749, n43750,
         n43751, n43752, n43753, n43754, n43755, n43756, n43757, n43758,
         n43759, n43760, n43761, n43762, n43763, n43764, n43765, n43766,
         n43767, n43768, n43769, n43770, n43771, n43772, n43773, n43774,
         n43775, n43776, n43777, n43778, n43779, n43780, n43781, n43782,
         n43783, n43784, n43785, n43786, n43787, n43788, n43789, n43790,
         n43791, n43792, n43793, n43794, n43795, n43796, n43797, n43798,
         n43799, n43800, n43801, n43802, n43803, n43804, n43805, n43806,
         n43807, n43808, n43809, n43810, n43811, n43812, n43813, n43814,
         n43815, n43816, n43817, n43818, n43819, n43820, n43821, n43822,
         n43823, n43824, n43825, n43826, n43827, n43828, n43829, n43830,
         n43831, n43832, n43833, n43834, n43835, n43836, n43837, n43838,
         n43839, n43840, n43841, n43842, n43843, n43844, n43845, n43846,
         n43847, n43848, n43849, n43850, n43851, n43852, n43853, n43854,
         n43855, n43856, n43857, n43858, n43859, n43860, n43861, n43862,
         n43863, n43864, n43865, n43866, n43867, n43868, n43869, n43870,
         n43871, n43872, n43873, n43874, n43875, n43876, n43877, n43878,
         n43879, n43880, n43881, n43882, n43883, n43884, n43885, n43886,
         n43887, n43888, n43889, n43890, n43891, n43892, n43893, n43894,
         n43895, n43896, n43897, n43898, n43899, n43900, n43901, n43902,
         n43903, n43904, n43905, n43906, n43907, n43908, n43909, n43910,
         n43911, n43912, n43913, n43914, n43915, n43916, n43917, n43918,
         n43919, n43920, n43921, n43922, n43923, n43924, n43925, n43926,
         n43927, n43928, n43929, n43930, n43931, n43932, n43933, n43934,
         n43935, n43936, n43937, n43938, n43939, n43940, n43941, n43942,
         n43943, n43944, n43945, n43946, n43947, n43948, n43949, n43950,
         n43951, n43952, n43953, n43954, n43955, n43956, n43957, n43958,
         n43959, n43960, n43961, n43962, n43963, n43964, n43965, n43966,
         n43967, n43968, n43969, n43970, n43971, n43972, n43973, n43974,
         n43975, n43976, n43977, n43978, n43979, n43980, n43981, n43982,
         n43983, n43984, n43985, n43986, n43987, n43988, n43989, n43990,
         n43991, n43992, n43993, n43994, n43995, n43996, n43997, n43998,
         n43999, n44000, n44001, n44002, n44003, n44004, n44005, n44006,
         n44007, n44008, n44009, n44010, n44011, n44012, n44013, n44014,
         n44015, n44016, n44017, n44018, n44019, n44020, n44021, n44022,
         n44023, n44024, n44025, n44026, n44027, n44028, n44029, n44030,
         n44031, n44032, n44033, n44034, n44035, n44036, n44037, n44038,
         n44039, n44040, n44041, n44042, n44043, n44044, n44045, n44046,
         n44047, n44048, n44049, n44050, n44051, n44052, n44053, n44054,
         n44055, n44056, n44057, n44058, n44059, n44060, n44061, n44062,
         n44063, n44064, n44065, n44066, n44067, n44068, n44069, n44070,
         n44071, n44072, n44073, n44074, n44075, n44076, n44077, n44078,
         n44079, n44080, n44081, n44082, n44083, n44084, n44085, n44086,
         n44087, n44088, n44089, n44090, n44091, n44092, n44093, n44094,
         n44095, n44096, n44097, n44098, n44099, n44100, n44101, n44102,
         n44103, n44104, n44105, n44106, n44107, n44108, n44109, n44110,
         n44111, n44112, n44113, n44114, n44115, n44116, n44117, n44118,
         n44119, n44120, n44121, n44122, n44123, n44124, n44125, n44126,
         n44127, n44128, n44129, n44130, n44131, n44132, n44133, n44134,
         n44135, n44136, n44137, n44138, n44139, n44140, n44141, n44142,
         n44143, n44144, n44145, n44146, n44147, n44148, n44149, n44150,
         n44151, n44152, n44153, n44154, n44155, n44156, n44157, n44158,
         n44159, n44160, n44161, n44162, n44163, n44164, n44165, n44166,
         n44167, n44168, n44169, n44170, n44171, n44172, n44173, n44174,
         n44175, n44176, n44177, n44178, n44179, n44180, n44181, n44182,
         n44183, n44184, n44185, n44186, n44187, n44188, n44189, n44190,
         n44191, n44192, n44193, n44194, n44195, n44196, n44197, n44198,
         n44199, n44200, n44201, n44202, n44203, n44204, n44205, n44206,
         n44207, n44208, n44209, n44210, n44211, n44212, n44213, n44214,
         n44215, n44216, n44217, n44218, n44219, n44220, n44221, n44222,
         n44223, n44224, n44225, n44226, n44227, n44228, n44229, n44230,
         n44231, n44232, n44233, n44234, n44235, n44236, n44237, n44238,
         n44239, n44240, n44241, n44242, n44243, n44244, n44245, n44246,
         n44247, n44248, n44249, n44250, n44251, n44252, n44253, n44254,
         n44255, n44256, n44257, n44258, n44259, n44260, n44261, n44262,
         n44263, n44264, n44265, n44266, n44267, n44268, n44269, n44270,
         n44271, n44272, n44273, n44274, n44275, n44276, n44277, n44278,
         n44279, n44280, n44281, n44282, n44283, n44284, n44285, n44286,
         n44287, n44288, n44289, n44290, n44291, n44292, n44293, n44294,
         n44295, n44296, n44297, n44298, n44299, n44300, n44301, n44302,
         n44303, n44304, n44305, n44306, n44307, n44308, n44309, n44310,
         n44311, n44312, n44313, n44314, n44315, n44316, n44317, n44318,
         n44319, n44320, n44321, n44322, n44323, n44324, n44325, n44326,
         n44327, n44328, n44329, n44330, n44331, n44332, n44333, n44334,
         n44335, n44336, n44337, n44338, n44339, n44340, n44341, n44342,
         n44343, n44344, n44345, n44346, n44347, n44348, n44349, n44350,
         n44351, n44352, n44353, n44354, n44355, n44356, n44357, n44358,
         n44359, n44360, n44361, n44362, n44363, n44364, n44365, n44366,
         n44367, n44368, n44369, n44370, n44371, n44372, n44373, n44374,
         n44375, n44376, n44377, n44378, n44379, n44380, n44381, n44382,
         n44383, n44384, n44385, n44386, n44387, n44388, n44389, n44390,
         n44391, n44392, n44393, n44394, n44395, n44396, n44397, n44398,
         n44399, n44400, n44401, n44402, n44403, n44404, n44405, n44406,
         n44407, n44408, n44409, n44410, n44411, n44412, n44413, n44414,
         n44415, n44416, n44417, n44418, n44419, n44420, n44421, n44422,
         n44423, n44424, n44425, n44426, n44427, n44428, n44429, n44430,
         n44431, n44432, n44433, n44434, n44435, n44436, n44437, n44438,
         n44439, n44440, n44441, n44442, n44443, n44444, n44445, n44446,
         n44447, n44448, n44449, n44450, n44451, n44452, n44453, n44454,
         n44455, n44456, n44457, n44458, n44459, n44460, n44461, n44462,
         n44463, n44464, n44465, n44466, n44467, n44468, n44469, n44470,
         n44471, n44472, n44473, n44474, n44475, n44476, n44477, n44478,
         n44479, n44480, n44481, n44482, n44483, n44484, n44485, n44486,
         n44487, n44488, n44489, n44490, n44491, n44492, n44493, n44494,
         n44495, n44496, n44497, n44498, n44499, n44500, n44501, n44502,
         n44503, n44504, n44505, n44506, n44507, n44508, n44509, n44510,
         n44511, n44512, n44513, n44514, n44515, n44516, n44517, n44518,
         n44519, n44520, n44521, n44522, n44523, n44524, n44525, n44526,
         n44527, n44528, n44529, n44530, n44531, n44532, n44533, n44534,
         n44535, n44536, n44537, n44538, n44539, n44540, n44541, n44542,
         n44543, n44544, n44545, n44546, n44547, n44548, n44549, n44550,
         n44551, n44552, n44553, n44554, n44555, n44556, n44557, n44558,
         n44559, n44560, n44561, n44562, n44563, n44564, n44565, n44566,
         n44567, n44568, n44569, n44570, n44571, n44572, n44573, n44574,
         n44575, n44576, n44577, n44578, n44579, n44580, n44581, n44582,
         n44583, n44584, n44585, n44586, n44587, n44588, n44589, n44590,
         n44591, n44592, n44593, n44594, n44595, n44596, n44597, n44598,
         n44599, n44600, n44601, n44602, n44603, n44604, n44605, n44606,
         n44607, n44608, n44609, n44610, n44611, n44612, n44613, n44614,
         n44615, n44616, n44617, n44618, n44619, n44620, n44621, n44622,
         n44623, n44624, n44625, n44626, n44627, n44628, n44629, n44630,
         n44631, n44632, n44633, n44634, n44635, n44636, n44637, n44638,
         n44639, n44640, n44641, n44642, n44643, n44644, n44645, n44646,
         n44647, n44648, n44649, n44650, n44651, n44652, n44653, n44654,
         n44655, n44656, n44657, n44658, n44659, n44660, n44661, n44662,
         n44663, n44664, n44665, n44666, n44667, n44668, n44669, n44670,
         n44671, n44672, n44673, n44674, n44675, n44676, n44677, n44678,
         n44679, n44680, n44681, n44682, n44683, n44684, n44685, n44686,
         n44687, n44688, n44689, n44690, n44691, n44692, n44693, n44694,
         n44695, n44696, n44697, n44698, n44699, n44700, n44701, n44702,
         n44703, n44704, n44705, n44706, n44707, n44708, n44709, n44710,
         n44711, n44712, n44713, n44714, n44715, n44716, n44717, n44718,
         n44719, n44720, n44721, n44722, n44723, n44724, n44725, n44726,
         n44727, n44728, n44729, n44730, n44731, n44732, n44733, n44734,
         n44735, n44736, n44737, n44738, n44739, n44740, n44741, n44742,
         n44743, n44744, n44745, n44746, n44747, n44748, n44749, n44750,
         n44751, n44752, n44753, n44754, n44755, n44756, n44757, n44758,
         n44759, n44760, n44761, n44762, n44763, n44764, n44765, n44766,
         n44767, n44768, n44769, n44770, n44771, n44772, n44773, n44774,
         n44775, n44776, n44777, n44778, n44779, n44780, n44781, n44782,
         n44783, n44784, n44785, n44786, n44787, n44788, n44789, n44790,
         n44791, n44792, n44793, n44794, n44795, n44796, n44797, n44798,
         n44799, n44800, n44801, n44802, n44803, n44804, n44805, n44806,
         n44807, n44808, n44809, n44810, n44811, n44812, n44813, n44814,
         n44815, n44816, n44817, n44818, n44819, n44820, n44821, n44822,
         n44823, n44824, n44825, n44826, n44827, n44828, n44829, n44830,
         n44831, n44832, n44833, n44834, n44835, n44836, n44837, n44838,
         n44839, n44840, n44841, n44842, n44843, n44844, n44845, n44846,
         n44847, n44848, n44849, n44850, n44851, n44852, n44853, n44854,
         n44855, n44856, n44857, n44858, n44859, n44860, n44861, n44862,
         n44863, n44864, n44865, n44866, n44867, n44868, n44869, n44870,
         n44871, n44872, n44873, n44874, n44875, n44876, n44877, n44878,
         n44879, n44880, n44881, n44882, n44883, n44884, n44885, n44886,
         n44887, n44888, n44889, n44890, n44891, n44892, n44893, n44894,
         n44895, n44896, n44897, n44898, n44899, n44900, n44901, n44902,
         n44903, n44904, n44905, n44906, n44907, n44908, n44909, n44910,
         n44911, n44912, n44913, n44914, n44915, n44916, n44917, n44918,
         n44919, n44920, n44921, n44922, n44923, n44924, n44925, n44926,
         n44927, n44928, n44929, n44930, n44931, n44932, n44933, n44934,
         n44935, n44936, n44937, n44938, n44939, n44940, n44941, n44942,
         n44943, n44944, n44945, n44946, n44947, n44948, n44949, n44950,
         n44951, n44952, n44953, n44954, n44955, n44956, n44957, n44958,
         n44959, n44960, n44961, n44962, n44963, n44964, n44965, n44966,
         n44967, n44968, n44969, n44970, n44971, n44972, n44973, n44974,
         n44975, n44976, n44977, n44978, n44979, n44980, n44981, n44982,
         n44983, n44984, n44985, n44986, n44987, n44988, n44989, n44990,
         n44991, n44992, n44993, n44994, n44995, n44996, n44997, n44998,
         n44999, n45000, n45001, n45002, n45003, n45004, n45005, n45006,
         n45007, n45008, n45009, n45010, n45011, n45012, n45013, n45014,
         n45015, n45016, n45017, n45018, n45019, n45020, n45021, n45022,
         n45023, n45024, n45025, n45026, n45027, n45028, n45029, n45030,
         n45031, n45032, n45033, n45034, n45035, n45036, n45037, n45038,
         n45039, n45040, n45041, n45042, n45043, n45044, n45045, n45046,
         n45047, n45048, n45049, n45050, n45051, n45052, n45053, n45054,
         n45055, n45056, n45057, n45058, n45059, n45060, n45061, n45062,
         n45063, n45064, n45065, n45066, n45067, n45068, n45069, n45070,
         n45071, n45072, n45073, n45074, n45075, n45076, n45077, n45078,
         n45079, n45080, n45081, n45082, n45083, n45084, n45085, n45086,
         n45087, n45088, n45089, n45090, n45091, n45092, n45093, n45094,
         n45095, n45096, n45097, n45098, n45099, n45100, n45101, n45102,
         n45103, n45104, n45105, n45106, n45107, n45108, n45109, n45110,
         n45111, n45112, n45113, n45114, n45115, n45116, n45117, n45118,
         n45119, n45120, n45121, n45122, n45123, n45124, n45125, n45126,
         n45127, n45128, n45129, n45130, n45131, n45132, n45133, n45134,
         n45135, n45136, n45137, n45138, n45139, n45140, n45141, n45142,
         n45143, n45144, n45145, n45146, n45147, n45148, n45149, n45150,
         n45151, n45152, n45153, n45154, n45155, n45156, n45157, n45158,
         n45159, n45160, n45161, n45162, n45163, n45164, n45165, n45166,
         n45167, n45168, n45169, n45170, n45171, n45172, n45173, n45174,
         n45175, n45176, n45177, n45178, n45179, n45180, n45181, n45182,
         n45183, n45184, n45185, n45186, n45187, n45188, n45189, n45190,
         n45191, n45192, n45193, n45194, n45195, n45196, n45197, n45198,
         n45199, n45200, n45201, n45202, n45203, n45204, n45205, n45206,
         n45207, n45208, n45209, n45210, n45211, n45212, n45213, n45214,
         n45215, n45216, n45217, n45218, n45219, n45220, n45221, n45222,
         n45223, n45224, n45225, n45226, n45227, n45228, n45229, n45230,
         n45231, n45232, n45233, n45234, n45235, n45236, n45237, n45238,
         n45239, n45240, n45241, n45242, n45243, n45244, n45245, n45246,
         n45247, n45248, n45249, n45250, n45251, n45252, n45253, n45254,
         n45255, n45256, n45257, n45258, n45259, n45260, n45261, n45262,
         n45263, n45264, n45265, n45266, n45267, n45268, n45269, n45270,
         n45271, n45272, n45273, n45274, n45275, n45276, n45277, n45278,
         n45279, n45280, n45281, n45282, n45283, n45284, n45285, n45286,
         n45287, n45288, n45289, n45290, n45291, n45292, n45293, n45294,
         n45295, n45296, n45297, n45298, n45299, n45300, n45301, n45302,
         n45303, n45304, n45305, n45306, n45307, n45308, n45309, n45310,
         n45311, n45312, n45313, n45314, n45315, n45316, n45317, n45318,
         n45319, n45320, n45321, n45322, n45323, n45324, n45325, n45326,
         n45327, n45328, n45329, n45330, n45331, n45332, n45333, n45334,
         n45335, n45336, n45337, n45338, n45339, n45340, n45341, n45342,
         n45343, n45344, n45345, n45346, n45347, n45348, n45349, n45350,
         n45351, n45352, n45353, n45354, n45355, n45356, n45357, n45358,
         n45359, n45360, n45361, n45362, n45363, n45364, n45365, n45366,
         n45367, n45368, n45369, n45370, n45371, n45372, n45373, n45374,
         n45375, n45376, n45377, n45378, n45379, n45380, n45381, n45382,
         n45383, n45384, n45385, n45386, n45387, n45388, n45389, n45390,
         n45391, n45392, n45393, n45394, n45395, n45396, n45397, n45398,
         n45399, n45400, n45401, n45402, n45403, n45404, n45405, n45406,
         n45407, n45408, n45409, n45410, n45411, n45412, n45413, n45414,
         n45415, n45416, n45417, n45418, n45419, n45420, n45421, n45422,
         n45423, n45424, n45425, n45426, n45427, n45428, n45429, n45430,
         n45431, n45432, n45433, n45434, n45435, n45436, n45437, n45438,
         n45439, n45440, n45441, n45442, n45443, n45444, n45445, n45446,
         n45447, n45448, n45449, n45450, n45451, n45452, n45453, n45454,
         n45455, n45456, n45457, n45458, n45459, n45460, n45461, n45462,
         n45463, n45464, n45465, n45466, n45467, n45468, n45469, n45470,
         n45471, n45472, n45473, n45474, n45475, n45476, n45477, n45478,
         n45479, n45480, n45481, n45482, n45483, n45484, n45485, n45486,
         n45487, n45488, n45489, n45490, n45491, n45492, n45493, n45494,
         n45495, n45496, n45497, n45498, n45499, n45500, n45501, n45502,
         n45503, n45504, n45505, n45506, n45507, n45508, n45509, n45510,
         n45511, n45512, n45513, n45514, n45515, n45516, n45517, n45518,
         n45519, n45520, n45521, n45522, n45523, n45524, n45525, n45526,
         n45527, n45528, n45529, n45530, n45531, n45532, n45533, n45534,
         n45535, n45536, n45537, n45538, n45539, n45540, n45541, n45542,
         n45543, n45544, n45545, n45546, n45547, n45548, n45549, n45550,
         n45551, n45552, n45553, n45554, n45555, n45556, n45557, n45558,
         n45559, n45560, n45561, n45562, n45563, n45564, n45565, n45566,
         n45567, n45568, n45569, n45570, n45571, n45572, n45573, n45574,
         n45575, n45576, n45577, n45578, n45579, n45580, n45581, n45582,
         n45583, n45584, n45585, n45586, n45587, n45588, n45589, n45590,
         n45591, n45592, n45593, n45594, n45595, n45596, n45597, n45598,
         n45599, n45600, n45601, n45602, n45603, n45604, n45605, n45606,
         n45607, n45608, n45609, n45610, n45611, n45612, n45613, n45614,
         n45615, n45616, n45617, n45618, n45619, n45620, n45621, n45622,
         n45623, n45624, n45625, n45626, n45627, n45628, n45629, n45630,
         n45631, n45632, n45633, n45634, n45635, n45636, n45637, n45638,
         n45639, n45640, n45641, n45642, n45643, n45644, n45645, n45646,
         n45647, n45648, n45649, n45650, n45651, n45652, n45653, n45654,
         n45655, n45656, n45657, n45658, n45659, n45660, n45661, n45662,
         n45663, n45664, n45665, n45666, n45667, n45668, n45669, n45670,
         n45671, n45672, n45673, n45674, n45675, n45676, n45677, n45678,
         n45679, n45680, n45681, n45682, n45683, n45684, n45685, n45686,
         n45687, n45688, n45689, n45690, n45691, n45692, n45693, n45694,
         n45695, n45696, n45697, n45698, n45699, n45700, n45701, n45702,
         n45703, n45704, n45705, n45706, n45707, n45708, n45709, n45710,
         n45711, n45712, n45713, n45714, n45715, n45716, n45717, n45718,
         n45719, n45720, n45721, n45722, n45723, n45724, n45725, n45726,
         n45727, n45728, n45729, n45730, n45731, n45732, n45733, n45734,
         n45735, n45736, n45737, n45738, n45739, n45740, n45741, n45742,
         n45743, n45744, n45745, n45746, n45747, n45748, n45749, n45750,
         n45751, n45752, n45753, n45754, n45755, n45756, n45757, n45758,
         n45759, n45760, n45761, n45762, n45763, n45764, n45765, n45766,
         n45767, n45768, n45769, n45770, n45771, n45772, n45773, n45774,
         n45775, n45776, n45777, n45778, n45779, n45780, n45781, n45782,
         n45783, n45784, n45785, n45786, n45787, n45788, n45789, n45790,
         n45791, n45792, n45793, n45794, n45795, n45796, n45797, n45798,
         n45799, n45800, n45801, n45802, n45803, n45804, n45805, n45806,
         n45807, n45808, n45809, n45810, n45811, n45812, n45813, n45814,
         n45815, n45816, n45817, n45818, n45819, n45820, n45821, n45822,
         n45823, n45824, n45825, n45826, n45827, n45828, n45829, n45830,
         n45831, n45832, n45833, n45834, n45835, n45836, n45837, n45838,
         n45839, n45840, n45841, n45842, n45843, n45844, n45845, n45846,
         n45847, n45848, n45849, n45850, n45851, n45852, n45853, n45854,
         n45855, n45856, n45857, n45858, n45859, n45860, n45861, n45862,
         n45863, n45864, n45865, n45866, n45867, n45868, n45869, n45870,
         n45871, n45872, n45873, n45874, n45875, n45876, n45877, n45878,
         n45879, n45880, n45881, n45882, n45883, n45884, n45885, n45886,
         n45887, n45888, n45889, n45890, n45891, n45892, n45893, n45894,
         n45895, n45896, n45897, n45898, n45899, n45900, n45901, n45902,
         n45903, n45904, n45905, n45906, n45907, n45908, n45909, n45910,
         n45911, n45912, n45913, n45914, n45915, n45916, n45917, n45918,
         n45919, n45920, n45921, n45922, n45923, n45924, n45925, n45926,
         n45927, n45928, n45929, n45930, n45931, n45932, n45933, n45934,
         n45935, n45936, n45937, n45938, n45939, n45940, n45941, n45942,
         n45943, n45944, n45945, n45946, n45947, n45948, n45949, n45950,
         n45951, n45952, n45953, n45954, n45955, n45956, n45957, n45958,
         n45959, n45960, n45961, n45962, n45963, n45964, n45965, n45966,
         n45967, n45968, n45969, n45970, n45971, n45972, n45973, n45974,
         n45975, n45976, n45977, n45978, n45979, n45980, n45981, n45982,
         n45983, n45984, n45985, n45986, n45987, n45988, n45989, n45990,
         n45991, n45992, n45993, n45994, n45995, n45996, n45997, n45998,
         n45999, n46000, n46001, n46002, n46003, n46004, n46005, n46006,
         n46007, n46008, n46009, n46010, n46011, n46012, n46013, n46014,
         n46015, n46016, n46017, n46018, n46019, n46020, n46021, n46022,
         n46023, n46024, n46025, n46026, n46027, n46028, n46029, n46030,
         n46031, n46032, n46033, n46034, n46035, n46036, n46037, n46038,
         n46039, n46040, n46041, n46042, n46043, n46044, n46045, n46046,
         n46047, n46048, n46049, n46050, n46051, n46052, n46053, n46054,
         n46055, n46056, n46057, n46058, n46059, n46060, n46061, n46062,
         n46063, n46064, n46065, n46066, n46067, n46068, n46069, n46070,
         n46071, n46072, n46073, n46074, n46075, n46076, n46077, n46078,
         n46079, n46080, n46081, n46082, n46083, n46084, n46085, n46086,
         n46087, n46088, n46089, n46090, n46091, n46092, n46093, n46094,
         n46095, n46096, n46097, n46098, n46099, n46100, n46101, n46102,
         n46103, n46104, n46105, n46106, n46107, n46108, n46109, n46110,
         n46111, n46112, n46113, n46114, n46115, n46116, n46117, n46118,
         n46119, n46120, n46121, n46122, n46123, n46124, n46125, n46126,
         n46127, n46128, n46129, n46130, n46131, n46132, n46133, n46134,
         n46135, n46136, n46137, n46138, n46139, n46140, n46141, n46142,
         n46143, n46144, n46145, n46146, n46147, n46148, n46149, n46150,
         n46151, n46152, n46153, n46154, n46155, n46156, n46157, n46158,
         n46159, n46160, n46161, n46162, n46163, n46164, n46165, n46166,
         n46167, n46168, n46169, n46170, n46171, n46172, n46173, n46174,
         n46175, n46176, n46177, n46178, n46179, n46180, n46181, n46182,
         n46183, n46184, n46185, n46186, n46187, n46188, n46189, n46190,
         n46191, n46192, n46193, n46194, n46195, n46196, n46197, n46198,
         n46199, n46200, n46201, n46202, n46203, n46204, n46205, n46206,
         n46207, n46208, n46209, n46210, n46211, n46212, n46213, n46214,
         n46215, n46216, n46217, n46218, n46219, n46220, n46221, n46222,
         n46223, n46224, n46225, n46226, n46227, n46228, n46229, n46230,
         n46231, n46232, n46233, n46234, n46235, n46236, n46237, n46238,
         n46239, n46240, n46241, n46242, n46243, n46244, n46245, n46246,
         n46247, n46248, n46249, n46250, n46251, n46252, n46253, n46254,
         n46255, n46256, n46257, n46258, n46259, n46260, n46261, n46262,
         n46263, n46264, n46265, n46266, n46267, n46268, n46269, n46270,
         n46271, n46272, n46273, n46274, n46275, n46276, n46277, n46278,
         n46279, n46280, n46281, n46282, n46283, n46284, n46285, n46286,
         n46287, n46288, n46289, n46290, n46291, n46292, n46293, n46294,
         n46295, n46296, n46297, n46298, n46299, n46300, n46301, n46302,
         n46303, n46304, n46305, n46306, n46307, n46308, n46309, n46310,
         n46311, n46312, n46313, n46314, n46315, n46316, n46317, n46318,
         n46319, n46320, n46321, n46322, n46323, n46324, n46325, n46326,
         n46327, n46328, n46329, n46330, n46331, n46332, n46333, n46334,
         n46335, n46336, n46337, n46338, n46339, n46340, n46341, n46342,
         n46343, n46344, n46345, n46346, n46347, n46348, n46349, n46350,
         n46351, n46352, n46353, n46354, n46355, n46356, n46357, n46358,
         n46359, n46360, n46361, n46362, n46363, n46364, n46365, n46366,
         n46367, n46368, n46369, n46370, n46371, n46372, n46373, n46374,
         n46375, n46376, n46377, n46378, n46379, n46380, n46381, n46382,
         n46383, n46384, n46385, n46386, n46387, n46388, n46389, n46390,
         n46391, n46392, n46393, n46394, n46395, n46396, n46397, n46398,
         n46399, n46400, n46401, n46402, n46403, n46404, n46405, n46406,
         n46407, n46408, n46409, n46410, n46411, n46412, n46413, n46414,
         n46415, n46416, n46417, n46418, n46419, n46420, n46421, n46422,
         n46423, n46424, n46425, n46426, n46427, n46428, n46429, n46430,
         n46431, n46432, n46433, n46434, n46435, n46436, n46437, n46438,
         n46439, n46440, n46441, n46442, n46443, n46444, n46445, n46446,
         n46447, n46448, n46449, n46450, n46451, n46452, n46453, n46454,
         n46455, n46456, n46457, n46458, n46459, n46460, n46461, n46462,
         n46463, n46464, n46465, n46466, n46467, n46468, n46469, n46470,
         n46471, n46472, n46473, n46474, n46475, n46476, n46477, n46478,
         n46479, n46480, n46481, n46482, n46483, n46484, n46485, n46486,
         n46487, n46488, n46489, n46490, n46491, n46492, n46493, n46494,
         n46495, n46496, n46497, n46498, n46499, n46500, n46501, n46502,
         n46503, n46504, n46505, n46506, n46507, n46508, n46509, n46510,
         n46511, n46512, n46513, n46514, n46515, n46516, n46517, n46518,
         n46519, n46520, n46521, n46522, n46523, n46524, n46525, n46526,
         n46527, n46528, n46529, n46530, n46531, n46532, n46533, n46534,
         n46535, n46536, n46537, n46538, n46539, n46540, n46541, n46542,
         n46543, n46544, n46545, n46546, n46547, n46548, n46549, n46550,
         n46551, n46552, n46553, n46554, n46555, n46556, n46557, n46558,
         n46559, n46560, n46561, n46562, n46563, n46564, n46565, n46566,
         n46567, n46568, n46569, n46570, n46571, n46572, n46573, n46574,
         n46575, n46576, n46577, n46578, n46579, n46580, n46581, n46582,
         n46583, n46584, n46585, n46586, n46587, n46588, n46589, n46590,
         n46591, n46592, n46593, n46594, n46595, n46596, n46597, n46598,
         n46599, n46600, n46601, n46602, n46603, n46604, n46605, n46606,
         n46607, n46608, n46609, n46610, n46611, n46612, n46613, n46614,
         n46615, n46616, n46617, n46618, n46619, n46620, n46621, n46622,
         n46623, n46624, n46625, n46626, n46627, n46628, n46629, n46630,
         n46631, n46632, n46633, n46634, n46635, n46636, n46637, n46638,
         n46639, n46640, n46641, n46642, n46643, n46644, n46645, n46646,
         n46647, n46648, n46649, n46650, n46651, n46652, n46653, n46654,
         n46655, n46656, n46657, n46658, n46659, n46660, n46661, n46662,
         n46663, n46664, n46665, n46666, n46667, n46668, n46669, n46670,
         n46671, n46672, n46673, n46674, n46675, n46676, n46677, n46678,
         n46679, n46680, n46681, n46682, n46683, n46684, n46685, n46686,
         n46687, n46688, n46689, n46690, n46691, n46692, n46693, n46694,
         n46695, n46696, n46697, n46698, n46699, n46700, n46701, n46702,
         n46703, n46704, n46705, n46706, n46707, n46708, n46709, n46710,
         n46711, n46712, n46713, n46714, n46715, n46716, n46717, n46718,
         n46719, n46720, n46721, n46722, n46723, n46724, n46725, n46726,
         n46727, n46728, n46729, n46730, n46731, n46732, n46733, n46734,
         n46735, n46736, n46737, n46738, n46739, n46740, n46741, n46742,
         n46743, n46744, n46745, n46746, n46747, n46748, n46749, n46750,
         n46751, n46752, n46753, n46754, n46755, n46756, n46757, n46758,
         n46759, n46760, n46761, n46762, n46763, n46764, n46765, n46766,
         n46767, n46768, n46769, n46770, n46771, n46772, n46773, n46774,
         n46775, n46776, n46777, n46778, n46779, n46780, n46781, n46782,
         n46783, n46784, n46785, n46786, n46787, n46788, n46789, n46790,
         n46791, n46792, n46793, n46794, n46795, n46796, n46797, n46798,
         n46799, n46800, n46801, n46802, n46803, n46804, n46805, n46806,
         n46807, n46808, n46809, n46810, n46811, n46812, n46813, n46814,
         n46815, n46816, n46817, n46818, n46819, n46820, n46821, n46822,
         n46823, n46824, n46825, n46826, n46827, n46828, n46829, n46830,
         n46831, n46832, n46833, n46834, n46835, n46836, n46837, n46838,
         n46839, n46840, n46841, n46842, n46843, n46844, n46845, n46846,
         n46847, n46848, n46849, n46850, n46851, n46852, n46853, n46854,
         n46855, n46856, n46857, n46858, n46859, n46860, n46861, n46862,
         n46863, n46864, n46865, n46866, n46867, n46868, n46869, n46870,
         n46871, n46872, n46873, n46874, n46875, n46876, n46877, n46878,
         n46879, n46880, n46881, n46882, n46883, n46884, n46885, n46886,
         n46887, n46888, n46889, n46890, n46891, n46892, n46893, n46894,
         n46895, n46896, n46897, n46898, n46899, n46900, n46901, n46902,
         n46903, n46904, n46905, n46906, n46907, n46908, n46909, n46910,
         n46911, n46912, n46913, n46914, n46915, n46916, n46917, n46918,
         n46919, n46920, n46921, n46922, n46923, n46924, n46925, n46926,
         n46927, n46928, n46929, n46930, n46931, n46932, n46933, n46934,
         n46935, n46936, n46937, n46938, n46939, n46940, n46941, n46942,
         n46943, n46944, n46945, n46946, n46947, n46948, n46949, n46950,
         n46951, n46952, n46953, n46954, n46955, n46956, n46957, n46958,
         n46959, n46960, n46961, n46962, n46963, n46964, n46965, n46966,
         n46967, n46968, n46969, n46970, n46971, n46972, n46973, n46974,
         n46975, n46976, n46977, n46978, n46979, n46980, n46981, n46982,
         n46983, n46984, n46985, n46986, n46987, n46988, n46989, n46990,
         n46991, n46992, n46993, n46994, n46995, n46996, n46997, n46998,
         n46999, n47000, n47001, n47002, n47003, n47004, n47005, n47006,
         n47007, n47008, n47009, n47010, n47011, n47012, n47013, n47014,
         n47015, n47016, n47017, n47018, n47019, n47020, n47021, n47022,
         n47023, n47024, n47025, n47026, n47027, n47028, n47029, n47030,
         n47031, n47032, n47033, n47034, n47035, n47036, n47037, n47038,
         n47039, n47040, n47041, n47042, n47043, n47044, n47045, n47046,
         n47047, n47048, n47049, n47050, n47051, n47052, n47053, n47054,
         n47055, n47056, n47057, n47058, n47059, n47060, n47061, n47062,
         n47063, n47064, n47065, n47066, n47067, n47068, n47069, n47070,
         n47071, n47072, n47073, n47074, n47075, n47076, n47077, n47078,
         n47079, n47080, n47081, n47082, n47083, n47084, n47085, n47086,
         n47087, n47088, n47089, n47090, n47091, n47092, n47093, n47094,
         n47095, n47096, n47097, n47098, n47099, n47100, n47101, n47102,
         n47103, n47104, n47105, n47106, n47107, n47108, n47109, n47110,
         n47111, n47112, n47113, n47114, n47115, n47116, n47117, n47118,
         n47119, n47120, n47121, n47122, n47123, n47124, n47125, n47126,
         n47127, n47128, n47129, n47130, n47131, n47132, n47133, n47134,
         n47135, n47136, n47137, n47138, n47139, n47140, n47141, n47142,
         n47143, n47144, n47145, n47146, n47147, n47148, n47149, n47150,
         n47151, n47152, n47153, n47154, n47155, n47156, n47157, n47158,
         n47159, n47160, n47161, n47162, n47163, n47164, n47165, n47166,
         n47167, n47168, n47169, n47170, n47171, n47172, n47173, n47174,
         n47175, n47176, n47177, n47178, n47179, n47180, n47181, n47182,
         n47183, n47184, n47185, n47186, n47187, n47188, n47189, n47190,
         n47191, n47192, n47193, n47194, n47195, n47196, n47197, n47198,
         n47199, n47200, n47201, n47202, n47203, n47204, n47205, n47206,
         n47207, n47208, n47209, n47210, n47211, n47212, n47213, n47214,
         n47215, n47216, n47217, n47218, n47219, n47220, n47221, n47222,
         n47223, n47224, n47225, n47226, n47227, n47228, n47229, n47230,
         n47231, n47232, n47233, n47234, n47235, n47236, n47237, n47238,
         n47239, n47240, n47241, n47242, n47243, n47244, n47245, n47246,
         n47247, n47248, n47249, n47250, n47251, n47252, n47253, n47254,
         n47255, n47256, n47257, n47258, n47259, n47260, n47261, n47262,
         n47263, n47264, n47265, n47266, n47267, n47268, n47269, n47270,
         n47271, n47272, n47273, n47274, n47275, n47276, n47277, n47278,
         n47279, n47280, n47281, n47282, n47283, n47284, n47285, n47286,
         n47287, n47288, n47289, n47290, n47291, n47292, n47293, n47294,
         n47295, n47296, n47297, n47298, n47299, n47300, n47301, n47302,
         n47303, n47304, n47305, n47306, n47307, n47308, n47309, n47310,
         n47311, n47312, n47313, n47314, n47315, n47316, n47317, n47318,
         n47319, n47320, n47321, n47322, n47323, n47324, n47325, n47326,
         n47327, n47328, n47329, n47330, n47331, n47332, n47333, n47334,
         n47335, n47336, n47337, n47338, n47339, n47340, n47341, n47342,
         n47343, n47344, n47345, n47346, n47347, n47348, n47349, n47350,
         n47351, n47352, n47353, n47354, n47355, n47356, n47357, n47358,
         n47359, n47360, n47361, n47362, n47363, n47364, n47365, n47366,
         n47367, n47368, n47369, n47370, n47371, n47372, n47373, n47374,
         n47375, n47376, n47377, n47378, n47379, n47380, n47381, n47382,
         n47383, n47384, n47385, n47386, n47387, n47388, n47389, n47390,
         n47391, n47392, n47393, n47394, n47395, n47396, n47397, n47398,
         n47399, n47400, n47401, n47402, n47403, n47404, n47405, n47406,
         n47407, n47408, n47409, n47410, n47411, n47412, n47413, n47414,
         n47415, n47416, n47417, n47418, n47419, n47420, n47421, n47422,
         n47423, n47424, n47425, n47426, n47427, n47428, n47429, n47430,
         n47431, n47432, n47433, n47434, n47435, n47436, n47437, n47438,
         n47439, n47440, n47441, n47442, n47443, n47444, n47445, n47446,
         n47447, n47448, n47449, n47450, n47451, n47452, n47453, n47454,
         n47455, n47456, n47457, n47458, n47459, n47460, n47461, n47462,
         n47463, n47464, n47465, n47466, n47467, n47468, n47469, n47470,
         n47471, n47472, n47473, n47474, n47475, n47476, n47477, n47478,
         n47479, n47480, n47481, n47482, n47483, n47484, n47485, n47486,
         n47487, n47488, n47489, n47490, n47491, n47492, n47493, n47494,
         n47495, n47496, n47497, n47498, n47499, n47500, n47501, n47502,
         n47503, n47504, n47505, n47506, n47507, n47508, n47509, n47510,
         n47511, n47512, n47513, n47514, n47515, n47516, n47517, n47518,
         n47519, n47520, n47521, n47522, n47523, n47524, n47525, n47526,
         n47527, n47528, n47529, n47530, n47531, n47532, n47533, n47534,
         n47535, n47536, n47537, n47538, n47539, n47540, n47541, n47542,
         n47543, n47544, n47545, n47546, n47547, n47548, n47549, n47550,
         n47551, n47552, n47553, n47554, n47555, n47556, n47557, n47558,
         n47559, n47560, n47561, n47562, n47563, n47564, n47565, n47566,
         n47567, n47568, n47569, n47570, n47571, n47572, n47573, n47574,
         n47575, n47576, n47577, n47578, n47579, n47580, n47581, n47582,
         n47583, n47584, n47585, n47586, n47587, n47588, n47589, n47590,
         n47591, n47592, n47593, n47594, n47595, n47596, n47597, n47598,
         n47599, n47600, n47601, n47602, n47603, n47604, n47605, n47606,
         n47607, n47608, n47609, n47610, n47611, n47612, n47613, n47614,
         n47615, n47616, n47617, n47618, n47619, n47620, n47621, n47622,
         n47623, n47624, n47625, n47626, n47627, n47628, n47629, n47630,
         n47631, n47632, n47633, n47634, n47635, n47636, n47637, n47638,
         n47639, n47640, n47641, n47642, n47643, n47644, n47645, n47646,
         n47647, n47648, n47649, n47650, n47651, n47652, n47653, n47654,
         n47655, n47656, n47657, n47658, n47659, n47660, n47661, n47662,
         n47663, n47664, n47665, n47666, n47667, n47668, n47669, n47670,
         n47671, n47672, n47673, n47674, n47675, n47676, n47677, n47678,
         n47679, n47680, n47681, n47682, n47683, n47684, n47685, n47686,
         n47687, n47688, n47689, n47690, n47691, n47692, n47693, n47694,
         n47695, n47696, n47697, n47698, n47699, n47700, n47701, n47702,
         n47703, n47704, n47705, n47706, n47707, n47708, n47709, n47710,
         n47711, n47712, n47713, n47714, n47715, n47716, n47717, n47718,
         n47719, n47720, n47721, n47722, n47723, n47724, n47725, n47726,
         n47727, n47728, n47729, n47730, n47731, n47732, n47733, n47734,
         n47735, n47736, n47737, n47738, n47739, n47740, n47741, n47742,
         n47743, n47744, n47745, n47746, n47747, n47748, n47749, n47750,
         n47751, n47752, n47753, n47754, n47755, n47756, n47757, n47758,
         n47759, n47760, n47761, n47762, n47763, n47764, n47765, n47766,
         n47767, n47768, n47769, n47770, n47771, n47772, n47773, n47774,
         n47775, n47776, n47777, n47778, n47779, n47780, n47781, n47782,
         n47783, n47784, n47785, n47786, n47787, n47788, n47789, n47790,
         n47791, n47792, n47793, n47794, n47795, n47796, n47797, n47798,
         n47799, n47800, n47801, n47802, n47803, n47804, n47805, n47806,
         n47807, n47808, n47809, n47810, n47811, n47812, n47813, n47814,
         n47815, n47816, n47817, n47818, n47819, n47820, n47821, n47822,
         n47823, n47824, n47825, n47826, n47827, n47828, n47829, n47830,
         n47831, n47832, n47833, n47834, n47835, n47836, n47837, n47838,
         n47839, n47840, n47841, n47842, n47843, n47844, n47845, n47846,
         n47847, n47848, n47849, n47850, n47851, n47852, n47853, n47854,
         n47855, n47856, n47857, n47858, n47859, n47860, n47861, n47862,
         n47863, n47864, n47865, n47866, n47867, n47868, n47869, n47870,
         n47871, n47872, n47873, n47874, n47875, n47876, n47877, n47878,
         n47879, n47880, n47881, n47882, n47883, n47884, n47885, n47886,
         n47887, n47888, n47889, n47890, n47891, n47892, n47893, n47894,
         n47895, n47896, n47897, n47898, n47899, n47900, n47901, n47902,
         n47903, n47904, n47905, n47906, n47907, n47908, n47909, n47910,
         n47911, n47912, n47913, n47914, n47915, n47916, n47917, n47918,
         n47919, n47920, n47921, n47922, n47923, n47924, n47925, n47926,
         n47927, n47928, n47929, n47930, n47931, n47932, n47933, n47934,
         n47935, n47936, n47937, n47938, n47939, n47940, n47941, n47942,
         n47943, n47944, n47945, n47946, n47947, n47948, n47949, n47950,
         n47951, n47952, n47953, n47954, n47955, n47956, n47957, n47958,
         n47959, n47960, n47961, n47962, n47963, n47964, n47965, n47966,
         n47967, n47968, n47969, n47970, n47971, n47972, n47973, n47974,
         n47975, n47976, n47977, n47978, n47979, n47980, n47981, n47982,
         n47983, n47984, n47985, n47986, n47987, n47988, n47989, n47990,
         n47991, n47992, n47993, n47994, n47995, n47996, n47997, n47998,
         n47999, n48000, n48001, n48002, n48003, n48004, n48005, n48006,
         n48007, n48008, n48009, n48010, n48011, n48012, n48013, n48014,
         n48015, n48016, n48017, n48018, n48019, n48020, n48021, n48022,
         n48023, n48024, n48025, n48026, n48027, n48028, n48029, n48030,
         n48031, n48032, n48033, n48034, n48035, n48036, n48037, n48038,
         n48039, n48040, n48041, n48042, n48043, n48044, n48045, n48046,
         n48047, n48048, n48049, n48050, n48051, n48052, n48053, n48054,
         n48055, n48056, n48057, n48058, n48059, n48060, n48061, n48062,
         n48063, n48064, n48065, n48066, n48067, n48068, n48069, n48070,
         n48071, n48072, n48073, n48074, n48075, n48076, n48077, n48078,
         n48079, n48080, n48081, n48082, n48083, n48084, n48085, n48086,
         n48087, n48088, n48089, n48090, n48091, n48092, n48093, n48094,
         n48095, n48096, n48097, n48098, n48099, n48100, n48101, n48102,
         n48103, n48104, n48105, n48106, n48107, n48108, n48109, n48110,
         n48111, n48112, n48113, n48114, n48115, n48116, n48117, n48118,
         n48119, n48120, n48121, n48122, n48123, n48124, n48125, n48126,
         n48127, n48128, n48129, n48130, n48131, n48132, n48133, n48134,
         n48135, n48136, n48137, n48138, n48139, n48140, n48141, n48142,
         n48143, n48144, n48145, n48146, n48147, n48148, n48149, n48150,
         n48151, n48152, n48153, n48154, n48155, n48156, n48157, n48158,
         n48159, n48160, n48161, n48162, n48163, n48164, n48165, n48166,
         n48167, n48168, n48169, n48170, n48171, n48172, n48173, n48174,
         n48175, n48176, n48177, n48178, n48179, n48180, n48181, n48182,
         n48183, n48184, n48185, n48186, n48187, n48188, n48189, n48190,
         n48191, n48192, n48193, n48194, n48195, n48196, n48197, n48198,
         n48199, n48200, n48201, n48202, n48203, n48204, n48205, n48206,
         n48207, n48208, n48209, n48210, n48211, n48212, n48213, n48214,
         n48215, n48216, n48217, n48218, n48219, n48220, n48221, n48222,
         n48223, n48224, n48225, n48226, n48227, n48228, n48229, n48230,
         n48231, n48232, n48233, n48234, n48235, n48236, n48237, n48238,
         n48239, n48240, n48241, n48242, n48243, n48244, n48245, n48246,
         n48247, n48248, n48249, n48250, n48251, n48252, n48253, n48254,
         n48255, n48256, n48257, n48258, n48259, n48260, n48261, n48262,
         n48263, n48264, n48265, n48266, n48267, n48268, n48269, n48270,
         n48271, n48272, n48273, n48274, n48275, n48276, n48277, n48278,
         n48279, n48280, n48281, n48282, n48283, n48284, n48285, n48286,
         n48287, n48288, n48289, n48290, n48291, n48292, n48293, n48294,
         n48295, n48296, n48297, n48298, n48299, n48300, n48301, n48302,
         n48303, n48304, n48305, n48306, n48307, n48308, n48309, n48310,
         n48311, n48312, n48313, n48314, n48315, n48316, n48317, n48318,
         n48319, n48320, n48321, n48322, n48323, n48324, n48325, n48326,
         n48327, n48328, n48329, n48330, n48331, n48332, n48333, n48334,
         n48335, n48336, n48337, n48338, n48339, n48340, n48341, n48342,
         n48343, n48344, n48345, n48346, n48347, n48348, n48349, n48350,
         n48351, n48352, n48353, n48354, n48355, n48356, n48357, n48358,
         n48359, n48360, n48361, n48362, n48363, n48364, n48365, n48366,
         n48367, n48368, n48369, n48370, n48371, n48372, n48373, n48374,
         n48375, n48376, n48377, n48378, n48379, n48380, n48381, n48382,
         n48383, n48384, n48385, n48386, n48387, n48388, n48389, n48390,
         n48391, n48392, n48393, n48394, n48395, n48396, n48397, n48398,
         n48399, n48400, n48401, n48402, n48403, n48404, n48405, n48406,
         n48407, n48408, n48409, n48410, n48411, n48412, n48413, n48414,
         n48415, n48416, n48417, n48418, n48419, n48420, n48421, n48422,
         n48423, n48424, n48425, n48426, n48427, n48428, n48429, n48430,
         n48431, n48432, n48433, n48434, n48435, n48436, n48437, n48438,
         n48439, n48440, n48441, n48442, n48443, n48444, n48445, n48446,
         n48447, n48448, n48449, n48450, n48451, n48452, n48453, n48454,
         n48455, n48456, n48457, n48458, n48459, n48460, n48461, n48462,
         n48463, n48464, n48465, n48466, n48467, n48468, n48469, n48470,
         n48471, n48472, n48473, n48474, n48475, n48476, n48477, n48478,
         n48479, n48480, n48481, n48482, n48483, n48484, n48485, n48486,
         n48487, n48488, n48489, n48490, n48491, n48492, n48493, n48494,
         n48495, n48496, n48497, n48498, n48499, n48500, n48501, n48502,
         n48503, n48504, n48505, n48506, n48507, n48508, n48509, n48510,
         n48511, n48512, n48513, n48514, n48515, n48516, n48517, n48518,
         n48519, n48520, n48521, n48522, n48523, n48524, n48525, n48526,
         n48527, n48528, n48529, n48530, n48531, n48532, n48533, n48534,
         n48535, n48536, n48537, n48538, n48539, n48540, n48541, n48542,
         n48543, n48544, n48545, n48546, n48547, n48548, n48549, n48550,
         n48551, n48552, n48553, n48554, n48555, n48556, n48557, n48558,
         n48559, n48560, n48561, n48562, n48563, n48564, n48565, n48566,
         n48567, n48568, n48569, n48570, n48571, n48572, n48573, n48574,
         n48575, n48576, n48577, n48578, n48579, n48580, n48581, n48582,
         n48583, n48584, n48585, n48586, n48587, n48588, n48589, n48590,
         n48591, n48592, n48593, n48594, n48595, n48596, n48597, n48598,
         n48599, n48600, n48601, n48602, n48603, n48604, n48605, n48606,
         n48607, n48608, n48609, n48610, n48611, n48612, n48613, n48614,
         n48615, n48616, n48617, n48618, n48619, n48620, n48621, n48622,
         n48623, n48624, n48625, n48626, n48627, n48628, n48629, n48630,
         n48631, n48632, n48633, n48634, n48635, n48636, n48637, n48638,
         n48639, n48640, n48641, n48642, n48643, n48644, n48645, n48646,
         n48647, n48648, n48649, n48650, n48651, n48652, n48653, n48654,
         n48655, n48656, n48657, n48658, n48659, n48660, n48661, n48662,
         n48663, n48664, n48665, n48666, n48667, n48668, n48669, n48670,
         n48671, n48672, n48673, n48674, n48675, n48676, n48677, n48678,
         n48679, n48680, n48681, n48682, n48683, n48684, n48685, n48686,
         n48687, n48688, n48689, n48690, n48691, n48692, n48693, n48694,
         n48695, n48696, n48697, n48698, n48699, n48700, n48701, n48702,
         n48703, n48704, n48705, n48706, n48707, n48708, n48709, n48710,
         n48711, n48712, n48713, n48714, n48715, n48716, n48717, n48718,
         n48719, n48720, n48721, n48722, n48723, n48724, n48725, n48726,
         n48727, n48728, n48729, n48730, n48731, n48732, n48733, n48734,
         n48735, n48736, n48737, n48738, n48739, n48740, n48741, n48742,
         n48743, n48744, n48745, n48746, n48747, n48748, n48749, n48750,
         n48751, n48752, n48753, n48754, n48755, n48756, n48757, n48758,
         n48759, n48760, n48761, n48762, n48763, n48764, n48765, n48766,
         n48767, n48768, n48769, n48770, n48771, n48772, n48773, n48774,
         n48775, n48776, n48777, n48778, n48779, n48780, n48781, n48782,
         n48783, n48784, n48785, n48786, n48787, n48788, n48789, n48790,
         n48791, n48792, n48793, n48794, n48795, n48796, n48797, n48798,
         n48799, n48800, n48801, n48802, n48803, n48804, n48805, n48806,
         n48807, n48808, n48809, n48810, n48811, n48812, n48813, n48814,
         n48815, n48816, n48817, n48818, n48819, n48820, n48821, n48822,
         n48823, n48824, n48825, n48826, n48827, n48828, n48829, n48830,
         n48831, n48832, n48833, n48834, n48835, n48836, n48837, n48838,
         n48839, n48840, n48841, n48842, n48843, n48844, n48845, n48846,
         n48847, n48848, n48849, n48850, n48851, n48852, n48853, n48854,
         n48855, n48856, n48857, n48858, n48859, n48860, n48861, n48862,
         n48863, n48864, n48865, n48866, n48867, n48868, n48869, n48870,
         n48871, n48872, n48873, n48874, n48875, n48876, n48877, n48878,
         n48879, n48880, n48881, n48882, n48883, n48884, n48885, n48886,
         n48887, n48888, n48889, n48890, n48891, n48892, n48893, n48894,
         n48895, n48896, n48897, n48898, n48899, n48900, n48901, n48902,
         n48903, n48904, n48905, n48906, n48907, n48908, n48909, n48910,
         n48911, n48912, n48913, n48914, n48915, n48916, n48917, n48918,
         n48919, n48920, n48921, n48922, n48923, n48924, n48925, n48926,
         n48927, n48928, n48929, n48930, n48931, n48932, n48933, n48934,
         n48935, n48936, n48937, n48938, n48939, n48940, n48941, n48942,
         n48943, n48944, n48945, n48946, n48947, n48948, n48949, n48950,
         n48951, n48952, n48953, n48954, n48955, n48956, n48957, n48958,
         n48959, n48960, n48961, n48962, n48963, n48964, n48965, n48966,
         n48967, n48968, n48969, n48970, n48971, n48972, n48973, n48974,
         n48975, n48976, n48977, n48978, n48979, n48980, n48981, n48982,
         n48983, n48984, n48985, n48986, n48987, n48988, n48989, n48990,
         n48991, n48992, n48993, n48994, n48995, n48996, n48997, n48998,
         n48999, n49000, n49001, n49002, n49003, n49004, n49005, n49006,
         n49007, n49008, n49009, n49010, n49011, n49012, n49013, n49014,
         n49015, n49016, n49017, n49018, n49019, n49020, n49021, n49022,
         n49023, n49024, n49025, n49026, n49027, n49028, n49029, n49030,
         n49031, n49032, n49033, n49034, n49035, n49036, n49037, n49038,
         n49039, n49040, n49041, n49042, n49043, n49044, n49045, n49046,
         n49047, n49048, n49049, n49050, n49051, n49052, n49053, n49054,
         n49055, n49056, n49057, n49058, n49059, n49060, n49061, n49062,
         n49063, n49064, n49065, n49066, n49067, n49068, n49069, n49070,
         n49071, n49072, n49073, n49074, n49075, n49076, n49077, n49078,
         n49079, n49080, n49081, n49082, n49083, n49084, n49085, n49086,
         n49087, n49088, n49089, n49090, n49091, n49092, n49093, n49094,
         n49095, n49096, n49097, n49098, n49099, n49100, n49101, n49102,
         n49103, n49104, n49105, n49106, n49107, n49108, n49109, n49110,
         n49111, n49112, n49113, n49114, n49115, n49116, n49117, n49118,
         n49119, n49120, n49121, n49122, n49123, n49124, n49125, n49126,
         n49127, n49128, n49129, n49130, n49131, n49132, n49133, n49134,
         n49135, n49136, n49137, n49138, n49139, n49140, n49141, n49142,
         n49143, n49144, n49145, n49146, n49147, n49148, n49149, n49150,
         n49151, n49152, n49153, n49154, n49155, n49156, n49157, n49158,
         n49159, n49160, n49161, n49162, n49163, n49164, n49165, n49166,
         n49167, n49168, n49169, n49170, n49171, n49172, n49173, n49174,
         n49175, n49176, n49177, n49178, n49179, n49180, n49181, n49182,
         n49183, n49184, n49185, n49186, n49187, n49188, n49189, n49190,
         n49191, n49192, n49193, n49194, n49195, n49196, n49197, n49198,
         n49199, n49200, n49201, n49202, n49203, n49204, n49205, n49206,
         n49207, n49208, n49209, n49210, n49211, n49212, n49213, n49214,
         n49215, n49216, n49217, n49218, n49219, n49220, n49221, n49222,
         n49223, n49224, n49225, n49226, n49227, n49228, n49229, n49230,
         n49231, n49232, n49233, n49234, n49235, n49236, n49237, n49238,
         n49239, n49240, n49241, n49242, n49243, n49244, n49245, n49246,
         n49247, n49248, n49249, n49250, n49251, n49252, n49253, n49254,
         n49255, n49256, n49257, n49258, n49259, n49260, n49261, n49262,
         n49263, n49264, n49265, n49266, n49267, n49268, n49269, n49270,
         n49271, n49272, n49273, n49274, n49275, n49276, n49277, n49278,
         n49279, n49280, n49281, n49282, n49283, n49284, n49285, n49286,
         n49287, n49288, n49289, n49290, n49291, n49292, n49293, n49294,
         n49295, n49296, n49297, n49298, n49299, n49300, n49301, n49302,
         n49303, n49304, n49305, n49306, n49307, n49308, n49309, n49310,
         n49311, n49312, n49313, n49314, n49315, n49316, n49317, n49318,
         n49319, n49320, n49321, n49322, n49323, n49324, n49325, n49326,
         n49327, n49328, n49329, n49330, n49331, n49332, n49333, n49334,
         n49335, n49336, n49337, n49338, n49339, n49340, n49341, n49342,
         n49343, n49344, n49345, n49346, n49347, n49348, n49349, n49350,
         n49351, n49352, n49353, n49354, n49355, n49356, n49357, n49358,
         n49359, n49360, n49361, n49362, n49363, n49364, n49365, n49366,
         n49367, n49368, n49369, n49370, n49371, n49372, n49373, n49374,
         n49375, n49376, n49377, n49378, n49379, n49380, n49381, n49382,
         n49383, n49384, n49385, n49386, n49387, n49388, n49389, n49390,
         n49391, n49392, n49393, n49394, n49395, n49396, n49397, n49398,
         n49399, n49400, n49401, n49402, n49403, n49404, n49405, n49406,
         n49407, n49408, n49409, n49410, n49411, n49412, n49413, n49414,
         n49415, n49416, n49417, n49418, n49419, n49420, n49421, n49422,
         n49423, n49424, n49425, n49426, n49427, n49428, n49429, n49430,
         n49431, n49432, n49433, n49434, n49435, n49436, n49437, n49438,
         n49439, n49440, n49441, n49442, n49443, n49444, n49445, n49446,
         n49447, n49448, n49449, n49450, n49451, n49452, n49453, n49454,
         n49455, n49456, n49457, n49458, n49459, n49460, n49461, n49462,
         n49463, n49464, n49465, n49466, n49467, n49468, n49469, n49470,
         n49471, n49472, n49473, n49474, n49475, n49476, n49477, n49478,
         n49479, n49480, n49481, n49482, n49483, n49484, n49485, n49486,
         n49487, n49488, n49489, n49490, n49491, n49492, n49493, n49494,
         n49495, n49496, n49497, n49498, n49499, n49500, n49501, n49502,
         n49503, n49504, n49505, n49506, n49507, n49508, n49509, n49510,
         n49511, n49512, n49513, n49514, n49515, n49516, n49517, n49518,
         n49519, n49520, n49521, n49522, n49523, n49524, n49525, n49526,
         n49527, n49528, n49529, n49530, n49531, n49532, n49533, n49534,
         n49535, n49536, n49537, n49538, n49539, n49540, n49541, n49542,
         n49543, n49544, n49545, n49546, n49547, n49548, n49549, n49550,
         n49551, n49552, n49553, n49554, n49555, n49556, n49557, n49558,
         n49559, n49560, n49561, n49562, n49563, n49564, n49565, n49566,
         n49567, n49568, n49569, n49570, n49571, n49572, n49573, n49574,
         n49575, n49576, n49577, n49578, n49579, n49580, n49581, n49582,
         n49583, n49584, n49585, n49586, n49587, n49588, n49589, n49590,
         n49591, n49592, n49593, n49594, n49595, n49596, n49597, n49598,
         n49599, n49600, n49601, n49602, n49603, n49604, n49605, n49606,
         n49607, n49608, n49609, n49610, n49611, n49612, n49613, n49614,
         n49615, n49616, n49617, n49618, n49619, n49620, n49621, n49622,
         n49623, n49624, n49625, n49626, n49627, n49628, n49629, n49630,
         n49631, n49632, n49633, n49634, n49635, n49636, n49637, n49638,
         n49639, n49640, n49641, n49642, n49643, n49644, n49645, n49646,
         n49647, n49648, n49649, n49650, n49651, n49652, n49653, n49654,
         n49655, n49656, n49657, n49658, n49659, n49660, n49661, n49662,
         n49663, n49664, n49665, n49666, n49667, n49668, n49669, n49670,
         n49671, n49672, n49673, n49674, n49675, n49676, n49677, n49678,
         n49679, n49680, n49681, n49682, n49683, n49684, n49685, n49686,
         n49687, n49688, n49689, n49690, n49691, n49692, n49693, n49694,
         n49695, n49696, n49697, n49698, n49699, n49700, n49701, n49702,
         n49703, n49704, n49705, n49706, n49707, n49708, n49709, n49710,
         n49711, n49712, n49713, n49714, n49715, n49716, n49717, n49718,
         n49719, n49720, n49721, n49722, n49723, n49724, n49725, n49726,
         n49727, n49728, n49729, n49730, n49731, n49732, n49733, n49734,
         n49735, n49736, n49737, n49738, n49739, n49740, n49741, n49742,
         n49743, n49744, n49745, n49746, n49747, n49748, n49749, n49750,
         n49751, n49752, n49753, n49754, n49755, n49756, n49757, n49758,
         n49759, n49760, n49761, n49762, n49763, n49764, n49765, n49766,
         n49767, n49768, n49769, n49770, n49771, n49772, n49773, n49774,
         n49775, n49776, n49777, n49778, n49779, n49780, n49781, n49782,
         n49783, n49784, n49785, n49786, n49787, n49788, n49789, n49790,
         n49791, n49792, n49793, n49794, n49795, n49796, n49797, n49798,
         n49799, n49800, n49801, n49802, n49803, n49804, n49805, n49806,
         n49807, n49808, n49809, n49810, n49811, n49812, n49813, n49814,
         n49815, n49816, n49817, n49818, n49819, n49820, n49821, n49822,
         n49823, n49824, n49825, n49826, n49827, n49828, n49829, n49830,
         n49831, n49832, n49833, n49834, n49835, n49836, n49837, n49838,
         n49839, n49840, n49841, n49842, n49843, n49844, n49845, n49846,
         n49847, n49848, n49849, n49850, n49851, n49852, n49853, n49854,
         n49855, n49856, n49857, n49858, n49859, n49860, n49861, n49862,
         n49863, n49864, n49865, n49866, n49867, n49868, n49869, n49870,
         n49871, n49872, n49873, n49874, n49875, n49876, n49877, n49878,
         n49879, n49880, n49881, n49882, n49883, n49884, n49885, n49886,
         n49887, n49888, n49889, n49890, n49891, n49892, n49893, n49894,
         n49895, n49896, n49897, n49898, n49899, n49900, n49901, n49902,
         n49903, n49904, n49905, n49906, n49907, n49908, n49909, n49910,
         n49911, n49912, n49913, n49914, n49915, n49916, n49917, n49918,
         n49919, n49920, n49921, n49922, n49923, n49924, n49925, n49926,
         n49927, n49928, n49929, n49930, n49931, n49932, n49933, n49934,
         n49935, n49936, n49937, n49938, n49939, n49940, n49941, n49942,
         n49943, n49944, n49945, n49946, n49947, n49948, n49949, n49950,
         n49951, n49952, n49953, n49954, n49955, n49956, n49957, n49958,
         n49959, n49960, n49961, n49962, n49963, n49964, n49965, n49966,
         n49967, n49968, n49969, n49970, n49971, n49972, n49973, n49974,
         n49975, n49976, n49977, n49978, n49979, n49980, n49981, n49982,
         n49983, n49984, n49985, n49986, n49987, n49988, n49989, n49990,
         n49991, n49992, n49993, n49994, n49995, n49996, n49997, n49998,
         n49999, n50000, n50001, n50002, n50003, n50004, n50005, n50006,
         n50007, n50008, n50009, n50010, n50011, n50012, n50013, n50014,
         n50015, n50016, n50017, n50018, n50019, n50020, n50021, n50022,
         n50023, n50024, n50025, n50026, n50027, n50028, n50029, n50030,
         n50031, n50032, n50033, n50034, n50035, n50036, n50037, n50038,
         n50039, n50040, n50041, n50042, n50043, n50044, n50045, n50046,
         n50047, n50048, n50049, n50050, n50051, n50052, n50053, n50054,
         n50055, n50056, n50057, n50058, n50059, n50060, n50061, n50062,
         n50063, n50064, n50065, n50066, n50067, n50068, n50069, n50070,
         n50071, n50072, n50073, n50074, n50075, n50076, n50077, n50078,
         n50079, n50080, n50081, n50082, n50083, n50084, n50085, n50086,
         n50087, n50088, n50089, n50090, n50091, n50092, n50093, n50094,
         n50095, n50096, n50097, n50098, n50099, n50100, n50101, n50102,
         n50103, n50104, n50105, n50106, n50107, n50108, n50109, n50110,
         n50111, n50112, n50113, n50114, n50115, n50116, n50117, n50118,
         n50119, n50120, n50121, n50122, n50123, n50124, n50125, n50126,
         n50127, n50128, n50129, n50130, n50131, n50132, n50133, n50134,
         n50135, n50136, n50137, n50138, n50139, n50140, n50141, n50142,
         n50143, n50144, n50145, n50146, n50147, n50148, n50149, n50150,
         n50151, n50152, n50153, n50154, n50155, n50156, n50157, n50158,
         n50159, n50160, n50161, n50162, n50163, n50164, n50165, n50166,
         n50167, n50168, n50169, n50170, n50171, n50172, n50173, n50174,
         n50175, n50176, n50177, n50178, n50179, n50180, n50181, n50182,
         n50183, n50184, n50185, n50186, n50187, n50188, n50189, n50190,
         n50191, n50192, n50193, n50194, n50195, n50196, n50197, n50198,
         n50199, n50200, n50201, n50202, n50203, n50204, n50205, n50206,
         n50207, n50208, n50209, n50210, n50211, n50212, n50213, n50214,
         n50215, n50216, n50217, n50218, n50219, n50220, n50221, n50222,
         n50223, n50224, n50225, n50226, n50227, n50228, n50229, n50230,
         n50231, n50232, n50233, n50234, n50235, n50236, n50237, n50238,
         n50239, n50240, n50241, n50242, n50243, n50244, n50245, n50246,
         n50247, n50248, n50249, n50250, n50251, n50252, n50253, n50254,
         n50255, n50256, n50257, n50258, n50259, n50260, n50261, n50262,
         n50263, n50264, n50265, n50266, n50267, n50268, n50269, n50270,
         n50271, n50272, n50273, n50274, n50275, n50276, n50277, n50278,
         n50279, n50280, n50281, n50282, n50283, n50284, n50285, n50286,
         n50287, n50288, n50289, n50290, n50291, n50292, n50293, n50294,
         n50295, n50296, n50297, n50298, n50299, n50300, n50301, n50302,
         n50303, n50304, n50305, n50306, n50307, n50308, n50309, n50310,
         n50311, n50312, n50313, n50314, n50315, n50316, n50317, n50318,
         n50319, n50320, n50321, n50322, n50323, n50324, n50325, n50326,
         n50327, n50328, n50329, n50330, n50331, n50332, n50333, n50334,
         n50335, n50336, n50337, n50338, n50339, n50340, n50341, n50342,
         n50343, n50344, n50345, n50346, n50347, n50348, n50349, n50350,
         n50351, n50352, n50353, n50354, n50355, n50356, n50357, n50358,
         n50359, n50360, n50361, n50362, n50363, n50364, n50365, n50366,
         n50367, n50368, n50369, n50370, n50371, n50372, n50373, n50374,
         n50375, n50376, n50377, n50378, n50379, n50380, n50381, n50382,
         n50383, n50384, n50385, n50386, n50387, n50388, n50389, n50390,
         n50391, n50392, n50393, n50394, n50395, n50396, n50397, n50398,
         n50399, n50400, n50401, n50402, n50403, n50404, n50405, n50406,
         n50407, n50408, n50409, n50410, n50411, n50412, n50413, n50414,
         n50415, n50416, n50417, n50418, n50419, n50420, n50421, n50422,
         n50423, n50424, n50425, n50426, n50427, n50428, n50429, n50430,
         n50431, n50432, n50433, n50434, n50435, n50436, n50437, n50438,
         n50439, n50440, n50441, n50442, n50443, n50444, n50445, n50446,
         n50447, n50448, n50449, n50450, n50451, n50452, n50453, n50454,
         n50455, n50456, n50457, n50458, n50459, n50460, n50461, n50462,
         n50463, n50464, n50465, n50466, n50467, n50468, n50469, n50470,
         n50471, n50472, n50473, n50474, n50475, n50476, n50477, n50478,
         n50479, n50480, n50481, n50482, n50483, n50484, n50485, n50486,
         n50487, n50488, n50489, n50490, n50491, n50492, n50493, n50494,
         n50495, n50496, n50497, n50498, n50499, n50500, n50501, n50502,
         n50503, n50504, n50505, n50506, n50507, n50508, n50509, n50510,
         n50511, n50512, n50513, n50514, n50515, n50516, n50517, n50518,
         n50519, n50520, n50521, n50522, n50523, n50524, n50525, n50526,
         n50527, n50528, n50529, n50530, n50531, n50532, n50533, n50534,
         n50535, n50536, n50537, n50538, n50539, n50540, n50541, n50542,
         n50543, n50544, n50545, n50546, n50547, n50548, n50549, n50550,
         n50551, n50552, n50553, n50554, n50555, n50556, n50557, n50558,
         n50559, n50560, n50561, n50562, n50563, n50564, n50565, n50566,
         n50567, n50568, n50569, n50570, n50571, n50572, n50573, n50574,
         n50575, n50576, n50577, n50578, n50579, n50580, n50581, n50582,
         n50583, n50584, n50585, n50586, n50587, n50588, n50589, n50590,
         n50591, n50592, n50593, n50594, n50595, n50596, n50597, n50598,
         n50599, n50600, n50601, n50602, n50603, n50604, n50605, n50606,
         n50607, n50608, n50609, n50610, n50611, n50612, n50613, n50614,
         n50615, n50616, n50617, n50618, n50619, n50620, n50621, n50622,
         n50623, n50624, n50625, n50626, n50627, n50628, n50629, n50630,
         n50631, n50632, n50633, n50634, n50635, n50636, n50637, n50638,
         n50639, n50640, n50641, n50642, n50643, n50644, n50645, n50646,
         n50647, n50648, n50649, n50650, n50651, n50652, n50653, n50654,
         n50655, n50656, n50657, n50658, n50659, n50660, n50661, n50662,
         n50663, n50664, n50665, n50666, n50667, n50668, n50669, n50670,
         n50671, n50672, n50673, n50674, n50675, n50676, n50677, n50678,
         n50679, n50680, n50681, n50682, n50683, n50684, n50685, n50686,
         n50687, n50688, n50689, n50690, n50691, n50692, n50693, n50694,
         n50695, n50696, n50697, n50698, n50699, n50700, n50701, n50702,
         n50703, n50704, n50705, n50706, n50707, n50708, n50709, n50710,
         n50711, n50712, n50713, n50714, n50715, n50716, n50717, n50718,
         n50719, n50720, n50721, n50722, n50723, n50724, n50725, n50726,
         n50727, n50728, n50729, n50730, n50731, n50732, n50733, n50734,
         n50735, n50736, n50737, n50738, n50739, n50740, n50741, n50742,
         n50743, n50744, n50745, n50746, n50747, n50748, n50749, n50750,
         n50751, n50752, n50753, n50754, n50755, n50756, n50757, n50758,
         n50759, n50760, n50761, n50762, n50763, n50764, n50765, n50766,
         n50767, n50768, n50769, n50770, n50771, n50772, n50773, n50774,
         n50775, n50776, n50777, n50778, n50779, n50780, n50781, n50782,
         n50783, n50784, n50785, n50786, n50787, n50788, n50789, n50790,
         n50791, n50792, n50793, n50794, n50795, n50796, n50797, n50798,
         n50799, n50800, n50801, n50802, n50803, n50804, n50805, n50806,
         n50807, n50808, n50809, n50810, n50811, n50812, n50813, n50814,
         n50815, n50816, n50817, n50818, n50819, n50820, n50821, n50822,
         n50823, n50824, n50825, n50826, n50827, n50828, n50829, n50830,
         n50831, n50832, n50833, n50834, n50835, n50836, n50837, n50838,
         n50839, n50840, n50841, n50842, n50843, n50844, n50845, n50846,
         n50847, n50848, n50849, n50850, n50851, n50852, n50853, n50854,
         n50855, n50856, n50857, n50858, n50859, n50860, n50861, n50862,
         n50863, n50864, n50865, n50866, n50867, n50868, n50869, n50870,
         n50871, n50872, n50873, n50874, n50875, n50876, n50877, n50878,
         n50879, n50880, n50881, n50882, n50883, n50884, n50885, n50886,
         n50887, n50888, n50889, n50890, n50891, n50892, n50893, n50894,
         n50895, n50896, n50897, n50898, n50899, n50900, n50901, n50902,
         n50903, n50904, n50905, n50906, n50907, n50908, n50909, n50910,
         n50911, n50912, n50913, n50914, n50915, n50916, n50917, n50918,
         n50919, n50920, n50921, n50922, n50923, n50924, n50925, n50926,
         n50927, n50928, n50929, n50930, n50931, n50932, n50933, n50934,
         n50935, n50936, n50937, n50938, n50939, n50940, n50941, n50942,
         n50943, n50944, n50945, n50946, n50947, n50948, n50949, n50950,
         n50951, n50952, n50953, n50954, n50955, n50956, n50957, n50958,
         n50959, n50960, n50961, n50962, n50963, n50964, n50965, n50966,
         n50967, n50968, n50969, n50970, n50971, n50972, n50973, n50974,
         n50975, n50976, n50977, n50978, n50979, n50980, n50981, n50982,
         n50983, n50984, n50985, n50986, n50987, n50988, n50989, n50990,
         n50991, n50992, n50993, n50994, n50995, n50996, n50997, n50998,
         n50999, n51000, n51001, n51002, n51003, n51004, n51005, n51006,
         n51007, n51008, n51009, n51010, n51011, n51012, n51013, n51014,
         n51015, n51016, n51017, n51018, n51019, n51020, n51021, n51022,
         n51023, n51024, n51025, n51026, n51027, n51028, n51029, n51030,
         n51031, n51032, n51033, n51034, n51035, n51036, n51037, n51038,
         n51039, n51040, n51041, n51042, n51043, n51044, n51045, n51046,
         n51047, n51048, n51049, n51050, n51051, n51052, n51053, n51054,
         n51055, n51056, n51057, n51058, n51059, n51060, n51061, n51062,
         n51063, n51064, n51065, n51066, n51067, n51068, n51069, n51070,
         n51071, n51072, n51073, n51074, n51075, n51076, n51077, n51078,
         n51079, n51080, n51081, n51082, n51083, n51084, n51085, n51086,
         n51087, n51088, n51089, n51090, n51091, n51092, n51093, n51094,
         n51095, n51096, n51097, n51098, n51099, n51100, n51101, n51102,
         n51103, n51104, n51105, n51106, n51107, n51108, n51109, n51110,
         n51111, n51112, n51113, n51114, n51115, n51116, n51117, n51118,
         n51119, n51120, n51121, n51122, n51123, n51124, n51125, n51126,
         n51127, n51128, n51129, n51130, n51131, n51132, n51133, n51134,
         n51135, n51136, n51137, n51138, n51139, n51140, n51141, n51142,
         n51143, n51144, n51145, n51146, n51147, n51148, n51149, n51150,
         n51151, n51152, n51153, n51154, n51155, n51156, n51157, n51158,
         n51159, n51160, n51161, n51162, n51163, n51164, n51165, n51166,
         n51167, n51168, n51169, n51170, n51171, n51172, n51173, n51174,
         n51175, n51176, n51177, n51178, n51179, n51180, n51181, n51182,
         n51183, n51184, n51185, n51186, n51187, n51188, n51189, n51190,
         n51191, n51192, n51193, n51194, n51195, n51196, n51197, n51198,
         n51199, n51200, n51201, n51202, n51203, n51204, n51205, n51206,
         n51207, n51208, n51209, n51210, n51211, n51212, n51213, n51214,
         n51215, n51216, n51217, n51218, n51219, n51220, n51221, n51222,
         n51223, n51224, n51225, n51226, n51227, n51228, n51229, n51230,
         n51231, n51232, n51233, n51234, n51235, n51236, n51237, n51238,
         n51239, n51240, n51241, n51242, n51243, n51244, n51245, n51246,
         n51247, n51248, n51249, n51250, n51251, n51252, n51253, n51254,
         n51255, n51256, n51257, n51258, n51259, n51260, n51261, n51262,
         n51263, n51264, n51265, n51266, n51267, n51268, n51269, n51270,
         n51271, n51272, n51273, n51274, n51275, n51276, n51277, n51278,
         n51279, n51280, n51281, n51282, n51283, n51284, n51285, n51286,
         n51287, n51288, n51289, n51290, n51291, n51292, n51293, n51294,
         n51295, n51296, n51297, n51298, n51299, n51300, n51301, n51302,
         n51303, n51304, n51305, n51306, n51307, n51308, n51309, n51310,
         n51311, n51312, n51313, n51314, n51315, n51316, n51317, n51318,
         n51319, n51320, n51321, n51322, n51323, n51324, n51325, n51326,
         n51327, n51328, n51329, n51330, n51331, n51332, n51333, n51334,
         n51335, n51336, n51337, n51338, n51339, n51340, n51341, n51342,
         n51343, n51344, n51345, n51346, n51347, n51348, n51349, n51350,
         n51351, n51352, n51353, n51354, n51355, n51356, n51357, n51358,
         n51359, n51360, n51361, n51362, n51363, n51364, n51365, n51366,
         n51367, n51368, n51369, n51370, n51371, n51372, n51373, n51374,
         n51375, n51376, n51377, n51378, n51379, n51380, n51381, n51382,
         n51383, n51384, n51385, n51386, n51387, n51388, n51389, n51390,
         n51391, n51392, n51393, n51394, n51395, n51396, n51397, n51398,
         n51399, n51400, n51401, n51402, n51403, n51404, n51405, n51406,
         n51407, n51408, n51409, n51410, n51411, n51412, n51413, n51414,
         n51415, n51416, n51417, n51418, n51419, n51420, n51421, n51422,
         n51423, n51424, n51425, n51426, n51427, n51428, n51429, n51430,
         n51431, n51432, n51433, n51434, n51435, n51436, n51437, n51438,
         n51439, n51440, n51441, n51442, n51443, n51444, n51445, n51446,
         n51447, n51448, n51449, n51450, n51451, n51452, n51453, n51454,
         n51455, n51456, n51457, n51458, n51459, n51460, n51461, n51462,
         n51463, n51464, n51465, n51466, n51467, n51468, n51469, n51470,
         n51471, n51472, n51473, n51474, n51475, n51476, n51477, n51478,
         n51479, n51480, n51481, n51482, n51483, n51484, n51485, n51486,
         n51487, n51488, n51489, n51490, n51491, n51492, n51493, n51494,
         n51495, n51496, n51497, n51498, n51499, n51500, n51501, n51502,
         n51503, n51504, n51505, n51506, n51507, n51508, n51509, n51510,
         n51511, n51512, n51513, n51514, n51515, n51516, n51517, n51518,
         n51519, n51520, n51521, n51522, n51523, n51524, n51525, n51526,
         n51527, n51528, n51529, n51530, n51531, n51532, n51533, n51534,
         n51535, n51536, n51537, n51538, n51539, n51540, n51541, n51542,
         n51543, n51544, n51545, n51546, n51547, n51548, n51549, n51550,
         n51551, n51552, n51553, n51554, n51555, n51556, n51557, n51558,
         n51559, n51560, n51561, n51562, n51563, n51564, n51565, n51566,
         n51567, n51568, n51569, n51570, n51571, n51572, n51573, n51574,
         n51575, n51576, n51577, n51578, n51579, n51580, n51581, n51582,
         n51583, n51584, n51585, n51586, n51587, n51588, n51589, n51590,
         n51591, n51592, n51593, n51594, n51595, n51596, n51597, n51598,
         n51599, n51600, n51601, n51602, n51603, n51604, n51605, n51606,
         n51607, n51608, n51609, n51610, n51611, n51612, n51613, n51614,
         n51615, n51616, n51617, n51618, n51619, n51620, n51621, n51622,
         n51623, n51624, n51625, n51626, n51627, n51628, n51629, n51630,
         n51631, n51632, n51633, n51634, n51635, n51636, n51637, n51638,
         n51639, n51640, n51641, n51642, n51643, n51644, n51645, n51646,
         n51647, n51648, n51649, n51650, n51651, n51652, n51653, n51654,
         n51655, n51656, n51657, n51658, n51659, n51660, n51661, n51662,
         n51663, n51664, n51665, n51666, n51667, n51668, n51669, n51670,
         n51671, n51672, n51673, n51674, n51675, n51676, n51677, n51678,
         n51679, n51680, n51681, n51682, n51683, n51684, n51685, n51686,
         n51687, n51688, n51689, n51690, n51691, n51692, n51693, n51694,
         n51695, n51696, n51697, n51698, n51699, n51700, n51701, n51702,
         n51703, n51704, n51705, n51706, n51707, n51708, n51709, n51710,
         n51711, n51712, n51713, n51714, n51715, n51716, n51717, n51718,
         n51719, n51720, n51721, n51722, n51723, n51724, n51725, n51726,
         n51727, n51728, n51729, n51730, n51731, n51732, n51733, n51734,
         n51735, n51736, n51737, n51738, n51739, n51740, n51741, n51742,
         n51743, n51744, n51745, n51746, n51747, n51748, n51749, n51750,
         n51751, n51752, n51753, n51754, n51755, n51756, n51757, n51758,
         n51759, n51760, n51761, n51762, n51763, n51764, n51765, n51766,
         n51767, n51768, n51769, n51770, n51771, n51772, n51773, n51774,
         n51775, n51776, n51777, n51778, n51779, n51780, n51781, n51782,
         n51783, n51784, n51785, n51786, n51787, n51788, n51789, n51790,
         n51791, n51792, n51793, n51794, n51795, n51796, n51797, n51798,
         n51799, n51800, n51801, n51802, n51803, n51804, n51805, n51806,
         n51807, n51808, n51809, n51810, n51811, n51812, n51813, n51814,
         n51815, n51816, n51817, n51818, n51819, n51820, n51821, n51822,
         n51823, n51824, n51825, n51826, n51827, n51828, n51829, n51830,
         n51831, n51832, n51833, n51834, n51835, n51836, n51837, n51838,
         n51839, n51840, n51841, n51842, n51843, n51844, n51845, n51846,
         n51847, n51848, n51849, n51850, n51851, n51852, n51853, n51854,
         n51855, n51856, n51857, n51858, n51859, n51860, n51861, n51862,
         n51863, n51864, n51865, n51866, n51867, n51868, n51869, n51870,
         n51871, n51872, n51873, n51874, n51875, n51876, n51877, n51878,
         n51879, n51880, n51881, n51882, n51883, n51884, n51885, n51886,
         n51887, n51888, n51889, n51890, n51891, n51892, n51893, n51894,
         n51895, n51896, n51897, n51898, n51899, n51900, n51901, n51902,
         n51903, n51904, n51905, n51906, n51907, n51908, n51909, n51910,
         n51911, n51912, n51913, n51914, n51915, n51916, n51917, n51918,
         n51919, n51920, n51921, n51922, n51923, n51924, n51925, n51926,
         n51927, n51928, n51929, n51930, n51931, n51932, n51933, n51934,
         n51935, n51936, n51937, n51938, n51939, n51940, n51941, n51942,
         n51943, n51944, n51945, n51946, n51947, n51948, n51949, n51950,
         n51951, n51952, n51953, n51954, n51955, n51956, n51957, n51958,
         n51959, n51960, n51961, n51962, n51963, n51964, n51965, n51966,
         n51967, n51968, n51969, n51970, n51971, n51972, n51973, n51974,
         n51975, n51976, n51977, n51978, n51979, n51980, n51981, n51982,
         n51983, n51984, n51985, n51986, n51987, n51988, n51989, n51990,
         n51991, n51992, n51993, n51994, n51995, n51996, n51997, n51998,
         n51999, n52000, n52001, n52002, n52003, n52004, n52005, n52006,
         n52007, n52008, n52009, n52010, n52011, n52012, n52013, n52014,
         n52015, n52016, n52017, n52018, n52019, n52020, n52021, n52022,
         n52023, n52024, n52025, n52026, n52027, n52028, n52029, n52030,
         n52031, n52032, n52033, n52034, n52035, n52036, n52037, n52038,
         n52039, n52040, n52041, n52042, n52043, n52044, n52045, n52046,
         n52047, n52048, n52049, n52050, n52051, n52052, n52053, n52054,
         n52055, n52056, n52057, n52058, n52059, n52060, n52061, n52062,
         n52063, n52064, n52065, n52066, n52067, n52068, n52069, n52070,
         n52071, n52072, n52073, n52074, n52075, n52076, n52077, n52078,
         n52079, n52080, n52081, n52082, n52083, n52084, n52085, n52086,
         n52087, n52088, n52089, n52090, n52091, n52092, n52093, n52094,
         n52095, n52096, n52097, n52098, n52099, n52100, n52101, n52102,
         n52103, n52104, n52105, n52106, n52107, n52108, n52109, n52110,
         n52111, n52112, n52113, n52114, n52115, n52116, n52117, n52118,
         n52119, n52120, n52121, n52122, n52123, n52124, n52125, n52126,
         n52127, n52128, n52129, n52130, n52131, n52132, n52133, n52134,
         n52135, n52136, n52137, n52138, n52139, n52140, n52141, n52142,
         n52143, n52144, n52145, n52146, n52147, n52148, n52149, n52150,
         n52151, n52152, n52153, n52154, n52155, n52156, n52157, n52158,
         n52159, n52160, n52161, n52162, n52163, n52164, n52165, n52166,
         n52167, n52168, n52169, n52170, n52171, n52172, n52173, n52174,
         n52175, n52176, n52177, n52178, n52179, n52180, n52181, n52182,
         n52183, n52184, n52185, n52186, n52187, n52188, n52189, n52190,
         n52191, n52192, n52193, n52194, n52195, n52196, n52197, n52198,
         n52199, n52200, n52201, n52202, n52203, n52204, n52205, n52206,
         n52207, n52208, n52209, n52210, n52211, n52212, n52213, n52214,
         n52215, n52216, n52217, n52218, n52219, n52220, n52221, n52222,
         n52223, n52224, n52225, n52226, n52227, n52228, n52229, n52230,
         n52231, n52232, n52233, n52234, n52235, n52236, n52237, n52238,
         n52239, n52240, n52241, n52242, n52243, n52244, n52245, n52246,
         n52247, n52248, n52249, n52250, n52251, n52252, n52253, n52254,
         n52255, n52256, n52257, n52258, n52259, n52260, n52261, n52262,
         n52263, n52264, n52265, n52266, n52267, n52268, n52269, n52270,
         n52271, n52272, n52273, n52274, n52275, n52276, n52277, n52278,
         n52279, n52280, n52281, n52282, n52283, n52284, n52285, n52286,
         n52287, n52288, n52289, n52290, n52291, n52292, n52293, n52294,
         n52295, n52296, n52297, n52298, n52299, n52300, n52301, n52302,
         n52303, n52304, n52305, n52306, n52307, n52308, n52309, n52310,
         n52311, n52312, n52313, n52314, n52315, n52316, n52317, n52318,
         n52319, n52320, n52321, n52322, n52323, n52324, n52325, n52326,
         n52327, n52328, n52329, n52330, n52331, n52332, n52333, n52334,
         n52335, n52336, n52337, n52338, n52339, n52340, n52341, n52342,
         n52343, n52344, n52345, n52346, n52347, n52348, n52349, n52350,
         n52351, n52352, n52353, n52354, n52355, n52356, n52357, n52358,
         n52359, n52360, n52361, n52362, n52363, n52364, n52365, n52366,
         n52367, n52368, n52369, n52370, n52371, n52372, n52373, n52374,
         n52375, n52376, n52377, n52378, n52379, n52380, n52381, n52382,
         n52383, n52384, n52385, n52386, n52387, n52388, n52389, n52390,
         n52391, n52392, n52393, n52394, n52395, n52396, n52397, n52398,
         n52399, n52400, n52401, n52402, n52403, n52404, n52405, n52406,
         n52407, n52408, n52409, n52410, n52411, n52412, n52413, n52414,
         n52415, n52416, n52417, n52418, n52419, n52420, n52421, n52422,
         n52423, n52424, n52425, n52426, n52427, n52428, n52429, n52430,
         n52431, n52432, n52433, n52434, n52435, n52436, n52437, n52438,
         n52439, n52440, n52441, n52442, n52443, n52444, n52445, n52446,
         n52447, n52448, n52449, n52450, n52451, n52452, n52453, n52454,
         n52455, n52456, n52457, n52458, n52459, n52460, n52461, n52462,
         n52463, n52464, n52465, n52466, n52467, n52468, n52469, n52470,
         n52471, n52472, n52473, n52474, n52475, n52476, n52477, n52478,
         n52479, n52480, n52481, n52482, n52483, n52484, n52485, n52486,
         n52487, n52488, n52489, n52490, n52491, n52492, n52493, n52494,
         n52495, n52496, n52497, n52498, n52499, n52500, n52501, n52502,
         n52503, n52504, n52505, n52506, n52507, n52508, n52509, n52510,
         n52511, n52512, n52513, n52514, n52515, n52516, n52517, n52518,
         n52519, n52520, n52521, n52522, n52523, n52524, n52525, n52526,
         n52527, n52528, n52529, n52530, n52531, n52532, n52533, n52534,
         n52535, n52536, n52537, n52538, n52539, n52540, n52541, n52542,
         n52543, n52544, n52545, n52546, n52547, n52548, n52549, n52550,
         n52551, n52552, n52553, n52554, n52555, n52556, n52557, n52558,
         n52559, n52560, n52561, n52562, n52563, n52564, n52565, n52566,
         n52567, n52568, n52569, n52570, n52571, n52572, n52573, n52574,
         n52575, n52576, n52577, n52578, n52579, n52580, n52581, n52582,
         n52583, n52584, n52585, n52586, n52587, n52588, n52589, n52590,
         n52591, n52592, n52593, n52594, n52595, n52596, n52597, n52598,
         n52599, n52600, n52601, n52602, n52603, n52604, n52605, n52606,
         n52607, n52608, n52609, n52610, n52611, n52612, n52613, n52614,
         n52615, n52616, n52617, n52618, n52619, n52620, n52621, n52622,
         n52623, n52624, n52625, n52626, n52627, n52628, n52629, n52630,
         n52631, n52632, n52633, n52634, n52635, n52636, n52637, n52638,
         n52639, n52640, n52641, n52642, n52643, n52644, n52645, n52646,
         n52647, n52648, n52649, n52650, n52651, n52652, n52653, n52654,
         n52655, n52656, n52657, n52658, n52659, n52660, n52661, n52662,
         n52663, n52664, n52665, n52666, n52667, n52668, n52669, n52670,
         n52671, n52672, n52673, n52674, n52675, n52676, n52677, n52678,
         n52679, n52680, n52681, n52682, n52683, n52684, n52685, n52686,
         n52687, n52688, n52689, n52690, n52691, n52692, n52693, n52694,
         n52695, n52696, n52697, n52698, n52699, n52700, n52701, n52702,
         n52703, n52704, n52705, n52706, n52707, n52708, n52709, n52710,
         n52711, n52712, n52713, n52714, n52715, n52716, n52717, n52718,
         n52719, n52720, n52721, n52722, n52723, n52724, n52725, n52726,
         n52727, n52728, n52729, n52730, n52731, n52732, n52733, n52734,
         n52735, n52736, n52737, n52738, n52739, n52740, n52741, n52742,
         n52743, n52744, n52745, n52746, n52747, n52748, n52749, n52750,
         n52751, n52752, n52753, n52754, n52755, n52756, n52757, n52758,
         n52759, n52760, n52761, n52762, n52763, n52764, n52765, n52766,
         n52767, n52768, n52769, n52770, n52771, n52772, n52773, n52774,
         n52775, n52776, n52777, n52778, n52779, n52780, n52781, n52782,
         n52783, n52784, n52785, n52786, n52787, n52788, n52789, n52790,
         n52791, n52792, n52793, n52794, n52795, n52796, n52797, n52798,
         n52799, n52800, n52801, n52802, n52803, n52804, n52805, n52806,
         n52807, n52808, n52809, n52810, n52811, n52812, n52813, n52814,
         n52815, n52816, n52817, n52818, n52819, n52820, n52821, n52822,
         n52823, n52824, n52825, n52826, n52827, n52828, n52829, n52830,
         n52831, n52832, n52833, n52834, n52835, n52836, n52837, n52838,
         n52839, n52840, n52841, n52842, n52843, n52844, n52845, n52846,
         n52847, n52848, n52849, n52850, n52851, n52852, n52853, n52854,
         n52855, n52856, n52857, n52858, n52859, n52860, n52861, n52862,
         n52863, n52864, n52865, n52866, n52867, n52868, n52869, n52870,
         n52871, n52872, n52873, n52874, n52875, n52876, n52877, n52878,
         n52879, n52880, n52881, n52882, n52883, n52884, n52885, n52886,
         n52887, n52888, n52889, n52890, n52891, n52892, n52893, n52894,
         n52895, n52896, n52897, n52898, n52899, n52900, n52901, n52902,
         n52903, n52904, n52905, n52906, n52907, n52908, n52909, n52910,
         n52911, n52912, n52913, n52914, n52915, n52916, n52917, n52918,
         n52919, n52920, n52921, n52922, n52923, n52924, n52925, n52926,
         n52927, n52928, n52929, n52930, n52931, n52932, n52933, n52934,
         n52935, n52936, n52937, n52938, n52939, n52940, n52941, n52942,
         n52943, n52944, n52945, n52946, n52947, n52948, n52949, n52950,
         n52951, n52952, n52953, n52954, n52955, n52956, n52957, n52958,
         n52959, n52960, n52961, n52962, n52963, n52964, n52965, n52966,
         n52967, n52968, n52969, n52970, n52971, n52972, n52973, n52974,
         n52975, n52976, n52977, n52978, n52979, n52980, n52981, n52982,
         n52983, n52984, n52985, n52986, n52987, n52988, n52989, n52990,
         n52991, n52992, n52993, n52994, n52995, n52996, n52997, n52998,
         n52999, n53000, n53001, n53002, n53003, n53004, n53005, n53006,
         n53007, n53008, n53009, n53010, n53011, n53012, n53013, n53014,
         n53015, n53016, n53017, n53018, n53019, n53020, n53021, n53022,
         n53023, n53024, n53025, n53026, n53027, n53028, n53029, n53030,
         n53031, n53032, n53033, n53034, n53035, n53036, n53037, n53038,
         n53039, n53040, n53041, n53042, n53043, n53044, n53045, n53046,
         n53047, n53048, n53049, n53050, n53051, n53052, n53053, n53054,
         n53055, n53056, n53057, n53058, n53059, n53060, n53061, n53062,
         n53063, n53064, n53065, n53066, n53067, n53068, n53069, n53070,
         n53071, n53072, n53073, n53074, n53075, n53076, n53077, n53078,
         n53079, n53080, n53081, n53082, n53083, n53084, n53085, n53086,
         n53087, n53088, n53089, n53090, n53091, n53092, n53093, n53094,
         n53095, n53096, n53097, n53098, n53099, n53100, n53101, n53102,
         n53103, n53104, n53105, n53106, n53107, n53108, n53109, n53110,
         n53111, n53112, n53113, n53114, n53115, n53116, n53117, n53118,
         n53119, n53120, n53121, n53122, n53123, n53124, n53125, n53126,
         n53127, n53128, n53129, n53130, n53131, n53132, n53133, n53134,
         n53135, n53136, n53137, n53138, n53139, n53140, n53141, n53142,
         n53143, n53144, n53145, n53146, n53147, n53148, n53149, n53150,
         n53151, n53152, n53153, n53154, n53155, n53156, n53157, n53158,
         n53159, n53160, n53161, n53162, n53163, n53164, n53165, n53166,
         n53167, n53168, n53169, n53170, n53171, n53172, n53173, n53174,
         n53175, n53176, n53177, n53178, n53179, n53180, n53181, n53182,
         n53183, n53184, n53185, n53186, n53187, n53188, n53189, n53190,
         n53191, n53192, n53193, n53194, n53195, n53196, n53197, n53198,
         n53199, n53200, n53201, n53202, n53203, n53204, n53205, n53206,
         n53207, n53208, n53209, n53210, n53211, n53212, n53213, n53214,
         n53215, n53216, n53217, n53218, n53219, n53220, n53221, n53222,
         n53223, n53224, n53225, n53226, n53227, n53228, n53229, n53230,
         n53231, n53232, n53233, n53234, n53235, n53236, n53237, n53238,
         n53239, n53240, n53241, n53242, n53243, n53244, n53245, n53246,
         n53247, n53248, n53249, n53250, n53251, n53252, n53253, n53254,
         n53255, n53256, n53257, n53258, n53259, n53260, n53261, n53262,
         n53263, n53264, n53265, n53266, n53267, n53268, n53269, n53270,
         n53271, n53272, n53273, n53274, n53275, n53276, n53277, n53278,
         n53279, n53280, n53281, n53282, n53283, n53284, n53285, n53286,
         n53287, n53288, n53289, n53290, n53291, n53292, n53293, n53294,
         n53295, n53296, n53297, n53298, n53299, n53300, n53301, n53302,
         n53303, n53304, n53305, n53306, n53307, n53308, n53309, n53310,
         n53311, n53312, n53313, n53314, n53315, n53316, n53317, n53318,
         n53319, n53320, n53321, n53322, n53323, n53324, n53325, n53326,
         n53327, n53328, n53329, n53330, n53331, n53332, n53333, n53334,
         n53335, n53336, n53337, n53338, n53339, n53340, n53341, n53342,
         n53343, n53344, n53345, n53346, n53347, n53348, n53349, n53350,
         n53351, n53352, n53353, n53354, n53355, n53356, n53357, n53358,
         n53359, n53360, n53361, n53362, n53363, n53364, n53365, n53366,
         n53367, n53368, n53369, n53370, n53371, n53372, n53373, n53374,
         n53375, n53376, n53377, n53378, n53379, n53380, n53381, n53382,
         n53383, n53384, n53385, n53386, n53387, n53388, n53389, n53390,
         n53391, n53392, n53393, n53394, n53395, n53396, n53397, n53398,
         n53399, n53400, n53401, n53402, n53403, n53404, n53405, n53406,
         n53407, n53408, n53409, n53410, n53411, n53412, n53413, n53414,
         n53415, n53416, n53417, n53418, n53419, n53420, n53421, n53422,
         n53423, n53424, n53425, n53426, n53427, n53428, n53429, n53430,
         n53431, n53432, n53433, n53434, n53435, n53436, n53437, n53438,
         n53439, n53440, n53441, n53442, n53443, n53444, n53445, n53446,
         n53447, n53448, n53449, n53450, n53451, n53452, n53453, n53454,
         n53455, n53456, n53457, n53458, n53459, n53460, n53461, n53462,
         n53463, n53464, n53465, n53466, n53467, n53468, n53469, n53470,
         n53471, n53472, n53473, n53474, n53475, n53476, n53477, n53478,
         n53479, n53480, n53481, n53482, n53483, n53484, n53485, n53486,
         n53487, n53488, n53489, n53490, n53491, n53492, n53493, n53494,
         n53495, n53496, n53497, n53498, n53499, n53500, n53501, n53502,
         n53503, n53504, n53505, n53506, n53507, n53508, n53509, n53510,
         n53511, n53512, n53513, n53514, n53515, n53516, n53517, n53518,
         n53519, n53520, n53521, n53522, n53523, n53524, n53525, n53526,
         n53527, n53528, n53529, n53530, n53531, n53532, n53533, n53534,
         n53535, n53536, n53537, n53538, n53539, n53540, n53541, n53542,
         n53543, n53544, n53545, n53546, n53547, n53548, n53549, n53550,
         n53551, n53552, n53553, n53554, n53555, n53556, n53557, n53558,
         n53559, n53560, n53561, n53562, n53563, n53564, n53565, n53566,
         n53567, n53568, n53569, n53570, n53571, n53572, n53573, n53574,
         n53575, n53576, n53577, n53578, n53579, n53580, n53581, n53582,
         n53583, n53584, n53585, n53586, n53587, n53588, n53589, n53590,
         n53591, n53592, n53593, n53594, n53595, n53596, n53597, n53598,
         n53599, n53600, n53601, n53602, n53603, n53604, n53605, n53606,
         n53607, n53608, n53609, n53610, n53611, n53612, n53613, n53614,
         n53615, n53616, n53617, n53618, n53619, n53620, n53621, n53622,
         n53623, n53624, n53625, n53626, n53627, n53628, n53629, n53630,
         n53631, n53632, n53633, n53634, n53635, n53636, n53637, n53638,
         n53639, n53640, n53641, n53642, n53643, n53644, n53645, n53646,
         n53647, n53648, n53649, n53650, n53651, n53652, n53653, n53654,
         n53655, n53656, n53657, n53658, n53659, n53660, n53661, n53662,
         n53663, n53664, n53665, n53666, n53667, n53668, n53669, n53670,
         n53671, n53672, n53673, n53674, n53675, n53676, n53677, n53678,
         n53679, n53680, n53681, n53682, n53683, n53684, n53685, n53686,
         n53687, n53688, n53689, n53690, n53691, n53692, n53693, n53694,
         n53695, n53696, n53697, n53698, n53699, n53700, n53701, n53702,
         n53703, n53704, n53705, n53706, n53707, n53708, n53709, n53710,
         n53711, n53712, n53713, n53714, n53715, n53716, n53717, n53718,
         n53719, n53720, n53721, n53722, n53723, n53724, n53725, n53726,
         n53727, n53728, n53729, n53730, n53731, n53732, n53733, n53734,
         n53735, n53736, n53737, n53738, n53739, n53740, n53741, n53742,
         n53743, n53744, n53745, n53746, n53747, n53748, n53749, n53750,
         n53751, n53752, n53753, n53754, n53755, n53756, n53757, n53758,
         n53759, n53760, n53761, n53762, n53763, n53764, n53765, n53766,
         n53767, n53768, n53769, n53770;
  wire   [2:0] rc_i;
  wire   [1599:0] round_reg;

  DFF init_reg ( .D(1'b1), .CLK(clk), .RST(rst), .I(1'b0), .Q(init) );
  DFF \rc_i_reg[0]  ( .D(n1029), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[0])
         );
  DFF \rc_i_reg[1]  ( .D(rc_i[0]), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[1])
         );
  DFF \rc_i_reg[2]  ( .D(rc_i[1]), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[2])
         );
  DFF \round_reg_reg[0]  ( .D(out[0]), .CLK(clk), .RST(rst), .I(in[0]), .Q(
        round_reg[0]) );
  DFF \round_reg_reg[1]  ( .D(out[1]), .CLK(clk), .RST(rst), .I(in[1]), .Q(
        round_reg[1]) );
  DFF \round_reg_reg[2]  ( .D(out[2]), .CLK(clk), .RST(rst), .I(in[2]), .Q(
        round_reg[2]) );
  DFF \round_reg_reg[3]  ( .D(out[3]), .CLK(clk), .RST(rst), .I(in[3]), .Q(
        round_reg[3]) );
  DFF \round_reg_reg[4]  ( .D(out[4]), .CLK(clk), .RST(rst), .I(in[4]), .Q(
        round_reg[4]) );
  DFF \round_reg_reg[5]  ( .D(out[5]), .CLK(clk), .RST(rst), .I(in[5]), .Q(
        round_reg[5]) );
  DFF \round_reg_reg[6]  ( .D(out[6]), .CLK(clk), .RST(rst), .I(in[6]), .Q(
        round_reg[6]) );
  DFF \round_reg_reg[7]  ( .D(out[7]), .CLK(clk), .RST(rst), .I(in[7]), .Q(
        round_reg[7]) );
  DFF \round_reg_reg[8]  ( .D(out[8]), .CLK(clk), .RST(rst), .I(in[8]), .Q(
        round_reg[8]) );
  DFF \round_reg_reg[9]  ( .D(out[9]), .CLK(clk), .RST(rst), .I(in[9]), .Q(
        round_reg[9]) );
  DFF \round_reg_reg[10]  ( .D(out[10]), .CLK(clk), .RST(rst), .I(in[10]), .Q(
        round_reg[10]) );
  DFF \round_reg_reg[11]  ( .D(out[11]), .CLK(clk), .RST(rst), .I(in[11]), .Q(
        round_reg[11]) );
  DFF \round_reg_reg[12]  ( .D(out[12]), .CLK(clk), .RST(rst), .I(in[12]), .Q(
        round_reg[12]) );
  DFF \round_reg_reg[13]  ( .D(out[13]), .CLK(clk), .RST(rst), .I(in[13]), .Q(
        round_reg[13]) );
  DFF \round_reg_reg[14]  ( .D(out[14]), .CLK(clk), .RST(rst), .I(in[14]), .Q(
        round_reg[14]) );
  DFF \round_reg_reg[15]  ( .D(out[15]), .CLK(clk), .RST(rst), .I(in[15]), .Q(
        round_reg[15]) );
  DFF \round_reg_reg[16]  ( .D(out[16]), .CLK(clk), .RST(rst), .I(in[16]), .Q(
        round_reg[16]) );
  DFF \round_reg_reg[17]  ( .D(out[17]), .CLK(clk), .RST(rst), .I(in[17]), .Q(
        round_reg[17]) );
  DFF \round_reg_reg[18]  ( .D(out[18]), .CLK(clk), .RST(rst), .I(in[18]), .Q(
        round_reg[18]) );
  DFF \round_reg_reg[19]  ( .D(out[19]), .CLK(clk), .RST(rst), .I(in[19]), .Q(
        round_reg[19]) );
  DFF \round_reg_reg[20]  ( .D(out[20]), .CLK(clk), .RST(rst), .I(in[20]), .Q(
        round_reg[20]) );
  DFF \round_reg_reg[21]  ( .D(out[21]), .CLK(clk), .RST(rst), .I(in[21]), .Q(
        round_reg[21]) );
  DFF \round_reg_reg[22]  ( .D(out[22]), .CLK(clk), .RST(rst), .I(in[22]), .Q(
        round_reg[22]) );
  DFF \round_reg_reg[23]  ( .D(out[23]), .CLK(clk), .RST(rst), .I(in[23]), .Q(
        round_reg[23]) );
  DFF \round_reg_reg[24]  ( .D(out[24]), .CLK(clk), .RST(rst), .I(in[24]), .Q(
        round_reg[24]) );
  DFF \round_reg_reg[25]  ( .D(out[25]), .CLK(clk), .RST(rst), .I(in[25]), .Q(
        round_reg[25]) );
  DFF \round_reg_reg[26]  ( .D(out[26]), .CLK(clk), .RST(rst), .I(in[26]), .Q(
        round_reg[26]) );
  DFF \round_reg_reg[27]  ( .D(out[27]), .CLK(clk), .RST(rst), .I(in[27]), .Q(
        round_reg[27]) );
  DFF \round_reg_reg[28]  ( .D(out[28]), .CLK(clk), .RST(rst), .I(in[28]), .Q(
        round_reg[28]) );
  DFF \round_reg_reg[29]  ( .D(out[29]), .CLK(clk), .RST(rst), .I(in[29]), .Q(
        round_reg[29]) );
  DFF \round_reg_reg[30]  ( .D(out[30]), .CLK(clk), .RST(rst), .I(in[30]), .Q(
        round_reg[30]) );
  DFF \round_reg_reg[31]  ( .D(out[31]), .CLK(clk), .RST(rst), .I(in[31]), .Q(
        round_reg[31]) );
  DFF \round_reg_reg[32]  ( .D(out[32]), .CLK(clk), .RST(rst), .I(in[32]), .Q(
        round_reg[32]) );
  DFF \round_reg_reg[33]  ( .D(out[33]), .CLK(clk), .RST(rst), .I(in[33]), .Q(
        round_reg[33]) );
  DFF \round_reg_reg[34]  ( .D(out[34]), .CLK(clk), .RST(rst), .I(in[34]), .Q(
        round_reg[34]) );
  DFF \round_reg_reg[35]  ( .D(out[35]), .CLK(clk), .RST(rst), .I(in[35]), .Q(
        round_reg[35]) );
  DFF \round_reg_reg[36]  ( .D(out[36]), .CLK(clk), .RST(rst), .I(in[36]), .Q(
        round_reg[36]) );
  DFF \round_reg_reg[37]  ( .D(out[37]), .CLK(clk), .RST(rst), .I(in[37]), .Q(
        round_reg[37]) );
  DFF \round_reg_reg[38]  ( .D(out[38]), .CLK(clk), .RST(rst), .I(in[38]), .Q(
        round_reg[38]) );
  DFF \round_reg_reg[39]  ( .D(out[39]), .CLK(clk), .RST(rst), .I(in[39]), .Q(
        round_reg[39]) );
  DFF \round_reg_reg[40]  ( .D(out[40]), .CLK(clk), .RST(rst), .I(in[40]), .Q(
        round_reg[40]) );
  DFF \round_reg_reg[41]  ( .D(out[41]), .CLK(clk), .RST(rst), .I(in[41]), .Q(
        round_reg[41]) );
  DFF \round_reg_reg[42]  ( .D(out[42]), .CLK(clk), .RST(rst), .I(in[42]), .Q(
        round_reg[42]) );
  DFF \round_reg_reg[43]  ( .D(out[43]), .CLK(clk), .RST(rst), .I(in[43]), .Q(
        round_reg[43]) );
  DFF \round_reg_reg[44]  ( .D(out[44]), .CLK(clk), .RST(rst), .I(in[44]), .Q(
        round_reg[44]) );
  DFF \round_reg_reg[45]  ( .D(out[45]), .CLK(clk), .RST(rst), .I(in[45]), .Q(
        round_reg[45]) );
  DFF \round_reg_reg[46]  ( .D(out[46]), .CLK(clk), .RST(rst), .I(in[46]), .Q(
        round_reg[46]) );
  DFF \round_reg_reg[47]  ( .D(out[47]), .CLK(clk), .RST(rst), .I(in[47]), .Q(
        round_reg[47]) );
  DFF \round_reg_reg[48]  ( .D(out[48]), .CLK(clk), .RST(rst), .I(in[48]), .Q(
        round_reg[48]) );
  DFF \round_reg_reg[49]  ( .D(out[49]), .CLK(clk), .RST(rst), .I(in[49]), .Q(
        round_reg[49]) );
  DFF \round_reg_reg[50]  ( .D(out[50]), .CLK(clk), .RST(rst), .I(in[50]), .Q(
        round_reg[50]) );
  DFF \round_reg_reg[51]  ( .D(out[51]), .CLK(clk), .RST(rst), .I(in[51]), .Q(
        round_reg[51]) );
  DFF \round_reg_reg[52]  ( .D(out[52]), .CLK(clk), .RST(rst), .I(in[52]), .Q(
        round_reg[52]) );
  DFF \round_reg_reg[53]  ( .D(out[53]), .CLK(clk), .RST(rst), .I(in[53]), .Q(
        round_reg[53]) );
  DFF \round_reg_reg[54]  ( .D(out[54]), .CLK(clk), .RST(rst), .I(in[54]), .Q(
        round_reg[54]) );
  DFF \round_reg_reg[55]  ( .D(out[55]), .CLK(clk), .RST(rst), .I(in[55]), .Q(
        round_reg[55]) );
  DFF \round_reg_reg[56]  ( .D(out[56]), .CLK(clk), .RST(rst), .I(in[56]), .Q(
        round_reg[56]) );
  DFF \round_reg_reg[57]  ( .D(out[57]), .CLK(clk), .RST(rst), .I(in[57]), .Q(
        round_reg[57]) );
  DFF \round_reg_reg[58]  ( .D(out[58]), .CLK(clk), .RST(rst), .I(in[58]), .Q(
        round_reg[58]) );
  DFF \round_reg_reg[59]  ( .D(out[59]), .CLK(clk), .RST(rst), .I(in[59]), .Q(
        round_reg[59]) );
  DFF \round_reg_reg[60]  ( .D(out[60]), .CLK(clk), .RST(rst), .I(in[60]), .Q(
        round_reg[60]) );
  DFF \round_reg_reg[61]  ( .D(out[61]), .CLK(clk), .RST(rst), .I(in[61]), .Q(
        round_reg[61]) );
  DFF \round_reg_reg[62]  ( .D(out[62]), .CLK(clk), .RST(rst), .I(in[62]), .Q(
        round_reg[62]) );
  DFF \round_reg_reg[63]  ( .D(out[63]), .CLK(clk), .RST(rst), .I(in[63]), .Q(
        round_reg[63]) );
  DFF \round_reg_reg[64]  ( .D(out[64]), .CLK(clk), .RST(rst), .I(in[64]), .Q(
        round_reg[64]) );
  DFF \round_reg_reg[65]  ( .D(out[65]), .CLK(clk), .RST(rst), .I(in[65]), .Q(
        round_reg[65]) );
  DFF \round_reg_reg[66]  ( .D(out[66]), .CLK(clk), .RST(rst), .I(in[66]), .Q(
        round_reg[66]) );
  DFF \round_reg_reg[67]  ( .D(out[67]), .CLK(clk), .RST(rst), .I(in[67]), .Q(
        round_reg[67]) );
  DFF \round_reg_reg[68]  ( .D(out[68]), .CLK(clk), .RST(rst), .I(in[68]), .Q(
        round_reg[68]) );
  DFF \round_reg_reg[69]  ( .D(out[69]), .CLK(clk), .RST(rst), .I(in[69]), .Q(
        round_reg[69]) );
  DFF \round_reg_reg[70]  ( .D(out[70]), .CLK(clk), .RST(rst), .I(in[70]), .Q(
        round_reg[70]) );
  DFF \round_reg_reg[71]  ( .D(out[71]), .CLK(clk), .RST(rst), .I(in[71]), .Q(
        round_reg[71]) );
  DFF \round_reg_reg[72]  ( .D(out[72]), .CLK(clk), .RST(rst), .I(in[72]), .Q(
        round_reg[72]) );
  DFF \round_reg_reg[73]  ( .D(out[73]), .CLK(clk), .RST(rst), .I(in[73]), .Q(
        round_reg[73]) );
  DFF \round_reg_reg[74]  ( .D(out[74]), .CLK(clk), .RST(rst), .I(in[74]), .Q(
        round_reg[74]) );
  DFF \round_reg_reg[75]  ( .D(out[75]), .CLK(clk), .RST(rst), .I(in[75]), .Q(
        round_reg[75]) );
  DFF \round_reg_reg[76]  ( .D(out[76]), .CLK(clk), .RST(rst), .I(in[76]), .Q(
        round_reg[76]) );
  DFF \round_reg_reg[77]  ( .D(out[77]), .CLK(clk), .RST(rst), .I(in[77]), .Q(
        round_reg[77]) );
  DFF \round_reg_reg[78]  ( .D(out[78]), .CLK(clk), .RST(rst), .I(in[78]), .Q(
        round_reg[78]) );
  DFF \round_reg_reg[79]  ( .D(out[79]), .CLK(clk), .RST(rst), .I(in[79]), .Q(
        round_reg[79]) );
  DFF \round_reg_reg[80]  ( .D(out[80]), .CLK(clk), .RST(rst), .I(in[80]), .Q(
        round_reg[80]) );
  DFF \round_reg_reg[81]  ( .D(out[81]), .CLK(clk), .RST(rst), .I(in[81]), .Q(
        round_reg[81]) );
  DFF \round_reg_reg[82]  ( .D(out[82]), .CLK(clk), .RST(rst), .I(in[82]), .Q(
        round_reg[82]) );
  DFF \round_reg_reg[83]  ( .D(out[83]), .CLK(clk), .RST(rst), .I(in[83]), .Q(
        round_reg[83]) );
  DFF \round_reg_reg[84]  ( .D(out[84]), .CLK(clk), .RST(rst), .I(in[84]), .Q(
        round_reg[84]) );
  DFF \round_reg_reg[85]  ( .D(out[85]), .CLK(clk), .RST(rst), .I(in[85]), .Q(
        round_reg[85]) );
  DFF \round_reg_reg[86]  ( .D(out[86]), .CLK(clk), .RST(rst), .I(in[86]), .Q(
        round_reg[86]) );
  DFF \round_reg_reg[87]  ( .D(out[87]), .CLK(clk), .RST(rst), .I(in[87]), .Q(
        round_reg[87]) );
  DFF \round_reg_reg[88]  ( .D(out[88]), .CLK(clk), .RST(rst), .I(in[88]), .Q(
        round_reg[88]) );
  DFF \round_reg_reg[89]  ( .D(out[89]), .CLK(clk), .RST(rst), .I(in[89]), .Q(
        round_reg[89]) );
  DFF \round_reg_reg[90]  ( .D(out[90]), .CLK(clk), .RST(rst), .I(in[90]), .Q(
        round_reg[90]) );
  DFF \round_reg_reg[91]  ( .D(out[91]), .CLK(clk), .RST(rst), .I(in[91]), .Q(
        round_reg[91]) );
  DFF \round_reg_reg[92]  ( .D(out[92]), .CLK(clk), .RST(rst), .I(in[92]), .Q(
        round_reg[92]) );
  DFF \round_reg_reg[93]  ( .D(out[93]), .CLK(clk), .RST(rst), .I(in[93]), .Q(
        round_reg[93]) );
  DFF \round_reg_reg[94]  ( .D(out[94]), .CLK(clk), .RST(rst), .I(in[94]), .Q(
        round_reg[94]) );
  DFF \round_reg_reg[95]  ( .D(out[95]), .CLK(clk), .RST(rst), .I(in[95]), .Q(
        round_reg[95]) );
  DFF \round_reg_reg[96]  ( .D(out[96]), .CLK(clk), .RST(rst), .I(in[96]), .Q(
        round_reg[96]) );
  DFF \round_reg_reg[97]  ( .D(out[97]), .CLK(clk), .RST(rst), .I(in[97]), .Q(
        round_reg[97]) );
  DFF \round_reg_reg[98]  ( .D(out[98]), .CLK(clk), .RST(rst), .I(in[98]), .Q(
        round_reg[98]) );
  DFF \round_reg_reg[99]  ( .D(out[99]), .CLK(clk), .RST(rst), .I(in[99]), .Q(
        round_reg[99]) );
  DFF \round_reg_reg[100]  ( .D(out[100]), .CLK(clk), .RST(rst), .I(in[100]), 
        .Q(round_reg[100]) );
  DFF \round_reg_reg[101]  ( .D(out[101]), .CLK(clk), .RST(rst), .I(in[101]), 
        .Q(round_reg[101]) );
  DFF \round_reg_reg[102]  ( .D(out[102]), .CLK(clk), .RST(rst), .I(in[102]), 
        .Q(round_reg[102]) );
  DFF \round_reg_reg[103]  ( .D(out[103]), .CLK(clk), .RST(rst), .I(in[103]), 
        .Q(round_reg[103]) );
  DFF \round_reg_reg[104]  ( .D(out[104]), .CLK(clk), .RST(rst), .I(in[104]), 
        .Q(round_reg[104]) );
  DFF \round_reg_reg[105]  ( .D(out[105]), .CLK(clk), .RST(rst), .I(in[105]), 
        .Q(round_reg[105]) );
  DFF \round_reg_reg[106]  ( .D(out[106]), .CLK(clk), .RST(rst), .I(in[106]), 
        .Q(round_reg[106]) );
  DFF \round_reg_reg[107]  ( .D(out[107]), .CLK(clk), .RST(rst), .I(in[107]), 
        .Q(round_reg[107]) );
  DFF \round_reg_reg[108]  ( .D(out[108]), .CLK(clk), .RST(rst), .I(in[108]), 
        .Q(round_reg[108]) );
  DFF \round_reg_reg[109]  ( .D(out[109]), .CLK(clk), .RST(rst), .I(in[109]), 
        .Q(round_reg[109]) );
  DFF \round_reg_reg[110]  ( .D(out[110]), .CLK(clk), .RST(rst), .I(in[110]), 
        .Q(round_reg[110]) );
  DFF \round_reg_reg[111]  ( .D(out[111]), .CLK(clk), .RST(rst), .I(in[111]), 
        .Q(round_reg[111]) );
  DFF \round_reg_reg[112]  ( .D(out[112]), .CLK(clk), .RST(rst), .I(in[112]), 
        .Q(round_reg[112]) );
  DFF \round_reg_reg[113]  ( .D(out[113]), .CLK(clk), .RST(rst), .I(in[113]), 
        .Q(round_reg[113]) );
  DFF \round_reg_reg[114]  ( .D(out[114]), .CLK(clk), .RST(rst), .I(in[114]), 
        .Q(round_reg[114]) );
  DFF \round_reg_reg[115]  ( .D(out[115]), .CLK(clk), .RST(rst), .I(in[115]), 
        .Q(round_reg[115]) );
  DFF \round_reg_reg[116]  ( .D(out[116]), .CLK(clk), .RST(rst), .I(in[116]), 
        .Q(round_reg[116]) );
  DFF \round_reg_reg[117]  ( .D(out[117]), .CLK(clk), .RST(rst), .I(in[117]), 
        .Q(round_reg[117]) );
  DFF \round_reg_reg[118]  ( .D(out[118]), .CLK(clk), .RST(rst), .I(in[118]), 
        .Q(round_reg[118]) );
  DFF \round_reg_reg[119]  ( .D(out[119]), .CLK(clk), .RST(rst), .I(in[119]), 
        .Q(round_reg[119]) );
  DFF \round_reg_reg[120]  ( .D(out[120]), .CLK(clk), .RST(rst), .I(in[120]), 
        .Q(round_reg[120]) );
  DFF \round_reg_reg[121]  ( .D(out[121]), .CLK(clk), .RST(rst), .I(in[121]), 
        .Q(round_reg[121]) );
  DFF \round_reg_reg[122]  ( .D(out[122]), .CLK(clk), .RST(rst), .I(in[122]), 
        .Q(round_reg[122]) );
  DFF \round_reg_reg[123]  ( .D(out[123]), .CLK(clk), .RST(rst), .I(in[123]), 
        .Q(round_reg[123]) );
  DFF \round_reg_reg[124]  ( .D(out[124]), .CLK(clk), .RST(rst), .I(in[124]), 
        .Q(round_reg[124]) );
  DFF \round_reg_reg[125]  ( .D(out[125]), .CLK(clk), .RST(rst), .I(in[125]), 
        .Q(round_reg[125]) );
  DFF \round_reg_reg[126]  ( .D(out[126]), .CLK(clk), .RST(rst), .I(in[126]), 
        .Q(round_reg[126]) );
  DFF \round_reg_reg[127]  ( .D(out[127]), .CLK(clk), .RST(rst), .I(in[127]), 
        .Q(round_reg[127]) );
  DFF \round_reg_reg[128]  ( .D(out[128]), .CLK(clk), .RST(rst), .I(in[128]), 
        .Q(round_reg[128]) );
  DFF \round_reg_reg[129]  ( .D(out[129]), .CLK(clk), .RST(rst), .I(in[129]), 
        .Q(round_reg[129]) );
  DFF \round_reg_reg[130]  ( .D(out[130]), .CLK(clk), .RST(rst), .I(in[130]), 
        .Q(round_reg[130]) );
  DFF \round_reg_reg[131]  ( .D(out[131]), .CLK(clk), .RST(rst), .I(in[131]), 
        .Q(round_reg[131]) );
  DFF \round_reg_reg[132]  ( .D(out[132]), .CLK(clk), .RST(rst), .I(in[132]), 
        .Q(round_reg[132]) );
  DFF \round_reg_reg[133]  ( .D(out[133]), .CLK(clk), .RST(rst), .I(in[133]), 
        .Q(round_reg[133]) );
  DFF \round_reg_reg[134]  ( .D(out[134]), .CLK(clk), .RST(rst), .I(in[134]), 
        .Q(round_reg[134]) );
  DFF \round_reg_reg[135]  ( .D(out[135]), .CLK(clk), .RST(rst), .I(in[135]), 
        .Q(round_reg[135]) );
  DFF \round_reg_reg[136]  ( .D(out[136]), .CLK(clk), .RST(rst), .I(in[136]), 
        .Q(round_reg[136]) );
  DFF \round_reg_reg[137]  ( .D(out[137]), .CLK(clk), .RST(rst), .I(in[137]), 
        .Q(round_reg[137]) );
  DFF \round_reg_reg[138]  ( .D(out[138]), .CLK(clk), .RST(rst), .I(in[138]), 
        .Q(round_reg[138]) );
  DFF \round_reg_reg[139]  ( .D(out[139]), .CLK(clk), .RST(rst), .I(in[139]), 
        .Q(round_reg[139]) );
  DFF \round_reg_reg[140]  ( .D(out[140]), .CLK(clk), .RST(rst), .I(in[140]), 
        .Q(round_reg[140]) );
  DFF \round_reg_reg[141]  ( .D(out[141]), .CLK(clk), .RST(rst), .I(in[141]), 
        .Q(round_reg[141]) );
  DFF \round_reg_reg[142]  ( .D(out[142]), .CLK(clk), .RST(rst), .I(in[142]), 
        .Q(round_reg[142]) );
  DFF \round_reg_reg[143]  ( .D(out[143]), .CLK(clk), .RST(rst), .I(in[143]), 
        .Q(round_reg[143]) );
  DFF \round_reg_reg[144]  ( .D(out[144]), .CLK(clk), .RST(rst), .I(in[144]), 
        .Q(round_reg[144]) );
  DFF \round_reg_reg[145]  ( .D(out[145]), .CLK(clk), .RST(rst), .I(in[145]), 
        .Q(round_reg[145]) );
  DFF \round_reg_reg[146]  ( .D(out[146]), .CLK(clk), .RST(rst), .I(in[146]), 
        .Q(round_reg[146]) );
  DFF \round_reg_reg[147]  ( .D(out[147]), .CLK(clk), .RST(rst), .I(in[147]), 
        .Q(round_reg[147]) );
  DFF \round_reg_reg[148]  ( .D(out[148]), .CLK(clk), .RST(rst), .I(in[148]), 
        .Q(round_reg[148]) );
  DFF \round_reg_reg[149]  ( .D(out[149]), .CLK(clk), .RST(rst), .I(in[149]), 
        .Q(round_reg[149]) );
  DFF \round_reg_reg[150]  ( .D(out[150]), .CLK(clk), .RST(rst), .I(in[150]), 
        .Q(round_reg[150]) );
  DFF \round_reg_reg[151]  ( .D(out[151]), .CLK(clk), .RST(rst), .I(in[151]), 
        .Q(round_reg[151]) );
  DFF \round_reg_reg[152]  ( .D(out[152]), .CLK(clk), .RST(rst), .I(in[152]), 
        .Q(round_reg[152]) );
  DFF \round_reg_reg[153]  ( .D(out[153]), .CLK(clk), .RST(rst), .I(in[153]), 
        .Q(round_reg[153]) );
  DFF \round_reg_reg[154]  ( .D(out[154]), .CLK(clk), .RST(rst), .I(in[154]), 
        .Q(round_reg[154]) );
  DFF \round_reg_reg[155]  ( .D(out[155]), .CLK(clk), .RST(rst), .I(in[155]), 
        .Q(round_reg[155]) );
  DFF \round_reg_reg[156]  ( .D(out[156]), .CLK(clk), .RST(rst), .I(in[156]), 
        .Q(round_reg[156]) );
  DFF \round_reg_reg[157]  ( .D(out[157]), .CLK(clk), .RST(rst), .I(in[157]), 
        .Q(round_reg[157]) );
  DFF \round_reg_reg[158]  ( .D(out[158]), .CLK(clk), .RST(rst), .I(in[158]), 
        .Q(round_reg[158]) );
  DFF \round_reg_reg[159]  ( .D(out[159]), .CLK(clk), .RST(rst), .I(in[159]), 
        .Q(round_reg[159]) );
  DFF \round_reg_reg[160]  ( .D(out[160]), .CLK(clk), .RST(rst), .I(in[160]), 
        .Q(round_reg[160]) );
  DFF \round_reg_reg[161]  ( .D(out[161]), .CLK(clk), .RST(rst), .I(in[161]), 
        .Q(round_reg[161]) );
  DFF \round_reg_reg[162]  ( .D(out[162]), .CLK(clk), .RST(rst), .I(in[162]), 
        .Q(round_reg[162]) );
  DFF \round_reg_reg[163]  ( .D(out[163]), .CLK(clk), .RST(rst), .I(in[163]), 
        .Q(round_reg[163]) );
  DFF \round_reg_reg[164]  ( .D(out[164]), .CLK(clk), .RST(rst), .I(in[164]), 
        .Q(round_reg[164]) );
  DFF \round_reg_reg[165]  ( .D(out[165]), .CLK(clk), .RST(rst), .I(in[165]), 
        .Q(round_reg[165]) );
  DFF \round_reg_reg[166]  ( .D(out[166]), .CLK(clk), .RST(rst), .I(in[166]), 
        .Q(round_reg[166]) );
  DFF \round_reg_reg[167]  ( .D(out[167]), .CLK(clk), .RST(rst), .I(in[167]), 
        .Q(round_reg[167]) );
  DFF \round_reg_reg[168]  ( .D(out[168]), .CLK(clk), .RST(rst), .I(in[168]), 
        .Q(round_reg[168]) );
  DFF \round_reg_reg[169]  ( .D(out[169]), .CLK(clk), .RST(rst), .I(in[169]), 
        .Q(round_reg[169]) );
  DFF \round_reg_reg[170]  ( .D(out[170]), .CLK(clk), .RST(rst), .I(in[170]), 
        .Q(round_reg[170]) );
  DFF \round_reg_reg[171]  ( .D(out[171]), .CLK(clk), .RST(rst), .I(in[171]), 
        .Q(round_reg[171]) );
  DFF \round_reg_reg[172]  ( .D(out[172]), .CLK(clk), .RST(rst), .I(in[172]), 
        .Q(round_reg[172]) );
  DFF \round_reg_reg[173]  ( .D(out[173]), .CLK(clk), .RST(rst), .I(in[173]), 
        .Q(round_reg[173]) );
  DFF \round_reg_reg[174]  ( .D(out[174]), .CLK(clk), .RST(rst), .I(in[174]), 
        .Q(round_reg[174]) );
  DFF \round_reg_reg[175]  ( .D(out[175]), .CLK(clk), .RST(rst), .I(in[175]), 
        .Q(round_reg[175]) );
  DFF \round_reg_reg[176]  ( .D(out[176]), .CLK(clk), .RST(rst), .I(in[176]), 
        .Q(round_reg[176]) );
  DFF \round_reg_reg[177]  ( .D(out[177]), .CLK(clk), .RST(rst), .I(in[177]), 
        .Q(round_reg[177]) );
  DFF \round_reg_reg[178]  ( .D(out[178]), .CLK(clk), .RST(rst), .I(in[178]), 
        .Q(round_reg[178]) );
  DFF \round_reg_reg[179]  ( .D(out[179]), .CLK(clk), .RST(rst), .I(in[179]), 
        .Q(round_reg[179]) );
  DFF \round_reg_reg[180]  ( .D(out[180]), .CLK(clk), .RST(rst), .I(in[180]), 
        .Q(round_reg[180]) );
  DFF \round_reg_reg[181]  ( .D(out[181]), .CLK(clk), .RST(rst), .I(in[181]), 
        .Q(round_reg[181]) );
  DFF \round_reg_reg[182]  ( .D(out[182]), .CLK(clk), .RST(rst), .I(in[182]), 
        .Q(round_reg[182]) );
  DFF \round_reg_reg[183]  ( .D(out[183]), .CLK(clk), .RST(rst), .I(in[183]), 
        .Q(round_reg[183]) );
  DFF \round_reg_reg[184]  ( .D(out[184]), .CLK(clk), .RST(rst), .I(in[184]), 
        .Q(round_reg[184]) );
  DFF \round_reg_reg[185]  ( .D(out[185]), .CLK(clk), .RST(rst), .I(in[185]), 
        .Q(round_reg[185]) );
  DFF \round_reg_reg[186]  ( .D(out[186]), .CLK(clk), .RST(rst), .I(in[186]), 
        .Q(round_reg[186]) );
  DFF \round_reg_reg[187]  ( .D(out[187]), .CLK(clk), .RST(rst), .I(in[187]), 
        .Q(round_reg[187]) );
  DFF \round_reg_reg[188]  ( .D(out[188]), .CLK(clk), .RST(rst), .I(in[188]), 
        .Q(round_reg[188]) );
  DFF \round_reg_reg[189]  ( .D(out[189]), .CLK(clk), .RST(rst), .I(in[189]), 
        .Q(round_reg[189]) );
  DFF \round_reg_reg[190]  ( .D(out[190]), .CLK(clk), .RST(rst), .I(in[190]), 
        .Q(round_reg[190]) );
  DFF \round_reg_reg[191]  ( .D(out[191]), .CLK(clk), .RST(rst), .I(in[191]), 
        .Q(round_reg[191]) );
  DFF \round_reg_reg[192]  ( .D(out[192]), .CLK(clk), .RST(rst), .I(in[192]), 
        .Q(round_reg[192]) );
  DFF \round_reg_reg[193]  ( .D(out[193]), .CLK(clk), .RST(rst), .I(in[193]), 
        .Q(round_reg[193]) );
  DFF \round_reg_reg[194]  ( .D(out[194]), .CLK(clk), .RST(rst), .I(in[194]), 
        .Q(round_reg[194]) );
  DFF \round_reg_reg[195]  ( .D(out[195]), .CLK(clk), .RST(rst), .I(in[195]), 
        .Q(round_reg[195]) );
  DFF \round_reg_reg[196]  ( .D(out[196]), .CLK(clk), .RST(rst), .I(in[196]), 
        .Q(round_reg[196]) );
  DFF \round_reg_reg[197]  ( .D(out[197]), .CLK(clk), .RST(rst), .I(in[197]), 
        .Q(round_reg[197]) );
  DFF \round_reg_reg[198]  ( .D(out[198]), .CLK(clk), .RST(rst), .I(in[198]), 
        .Q(round_reg[198]) );
  DFF \round_reg_reg[199]  ( .D(out[199]), .CLK(clk), .RST(rst), .I(in[199]), 
        .Q(round_reg[199]) );
  DFF \round_reg_reg[200]  ( .D(out[200]), .CLK(clk), .RST(rst), .I(in[200]), 
        .Q(round_reg[200]) );
  DFF \round_reg_reg[201]  ( .D(out[201]), .CLK(clk), .RST(rst), .I(in[201]), 
        .Q(round_reg[201]) );
  DFF \round_reg_reg[202]  ( .D(out[202]), .CLK(clk), .RST(rst), .I(in[202]), 
        .Q(round_reg[202]) );
  DFF \round_reg_reg[203]  ( .D(out[203]), .CLK(clk), .RST(rst), .I(in[203]), 
        .Q(round_reg[203]) );
  DFF \round_reg_reg[204]  ( .D(out[204]), .CLK(clk), .RST(rst), .I(in[204]), 
        .Q(round_reg[204]) );
  DFF \round_reg_reg[205]  ( .D(out[205]), .CLK(clk), .RST(rst), .I(in[205]), 
        .Q(round_reg[205]) );
  DFF \round_reg_reg[206]  ( .D(out[206]), .CLK(clk), .RST(rst), .I(in[206]), 
        .Q(round_reg[206]) );
  DFF \round_reg_reg[207]  ( .D(out[207]), .CLK(clk), .RST(rst), .I(in[207]), 
        .Q(round_reg[207]) );
  DFF \round_reg_reg[208]  ( .D(out[208]), .CLK(clk), .RST(rst), .I(in[208]), 
        .Q(round_reg[208]) );
  DFF \round_reg_reg[209]  ( .D(out[209]), .CLK(clk), .RST(rst), .I(in[209]), 
        .Q(round_reg[209]) );
  DFF \round_reg_reg[210]  ( .D(out[210]), .CLK(clk), .RST(rst), .I(in[210]), 
        .Q(round_reg[210]) );
  DFF \round_reg_reg[211]  ( .D(out[211]), .CLK(clk), .RST(rst), .I(in[211]), 
        .Q(round_reg[211]) );
  DFF \round_reg_reg[212]  ( .D(out[212]), .CLK(clk), .RST(rst), .I(in[212]), 
        .Q(round_reg[212]) );
  DFF \round_reg_reg[213]  ( .D(out[213]), .CLK(clk), .RST(rst), .I(in[213]), 
        .Q(round_reg[213]) );
  DFF \round_reg_reg[214]  ( .D(out[214]), .CLK(clk), .RST(rst), .I(in[214]), 
        .Q(round_reg[214]) );
  DFF \round_reg_reg[215]  ( .D(out[215]), .CLK(clk), .RST(rst), .I(in[215]), 
        .Q(round_reg[215]) );
  DFF \round_reg_reg[216]  ( .D(out[216]), .CLK(clk), .RST(rst), .I(in[216]), 
        .Q(round_reg[216]) );
  DFF \round_reg_reg[217]  ( .D(out[217]), .CLK(clk), .RST(rst), .I(in[217]), 
        .Q(round_reg[217]) );
  DFF \round_reg_reg[218]  ( .D(out[218]), .CLK(clk), .RST(rst), .I(in[218]), 
        .Q(round_reg[218]) );
  DFF \round_reg_reg[219]  ( .D(out[219]), .CLK(clk), .RST(rst), .I(in[219]), 
        .Q(round_reg[219]) );
  DFF \round_reg_reg[220]  ( .D(out[220]), .CLK(clk), .RST(rst), .I(in[220]), 
        .Q(round_reg[220]) );
  DFF \round_reg_reg[221]  ( .D(out[221]), .CLK(clk), .RST(rst), .I(in[221]), 
        .Q(round_reg[221]) );
  DFF \round_reg_reg[222]  ( .D(out[222]), .CLK(clk), .RST(rst), .I(in[222]), 
        .Q(round_reg[222]) );
  DFF \round_reg_reg[223]  ( .D(out[223]), .CLK(clk), .RST(rst), .I(in[223]), 
        .Q(round_reg[223]) );
  DFF \round_reg_reg[224]  ( .D(out[224]), .CLK(clk), .RST(rst), .I(in[224]), 
        .Q(round_reg[224]) );
  DFF \round_reg_reg[225]  ( .D(out[225]), .CLK(clk), .RST(rst), .I(in[225]), 
        .Q(round_reg[225]) );
  DFF \round_reg_reg[226]  ( .D(out[226]), .CLK(clk), .RST(rst), .I(in[226]), 
        .Q(round_reg[226]) );
  DFF \round_reg_reg[227]  ( .D(out[227]), .CLK(clk), .RST(rst), .I(in[227]), 
        .Q(round_reg[227]) );
  DFF \round_reg_reg[228]  ( .D(out[228]), .CLK(clk), .RST(rst), .I(in[228]), 
        .Q(round_reg[228]) );
  DFF \round_reg_reg[229]  ( .D(out[229]), .CLK(clk), .RST(rst), .I(in[229]), 
        .Q(round_reg[229]) );
  DFF \round_reg_reg[230]  ( .D(out[230]), .CLK(clk), .RST(rst), .I(in[230]), 
        .Q(round_reg[230]) );
  DFF \round_reg_reg[231]  ( .D(out[231]), .CLK(clk), .RST(rst), .I(in[231]), 
        .Q(round_reg[231]) );
  DFF \round_reg_reg[232]  ( .D(out[232]), .CLK(clk), .RST(rst), .I(in[232]), 
        .Q(round_reg[232]) );
  DFF \round_reg_reg[233]  ( .D(out[233]), .CLK(clk), .RST(rst), .I(in[233]), 
        .Q(round_reg[233]) );
  DFF \round_reg_reg[234]  ( .D(out[234]), .CLK(clk), .RST(rst), .I(in[234]), 
        .Q(round_reg[234]) );
  DFF \round_reg_reg[235]  ( .D(out[235]), .CLK(clk), .RST(rst), .I(in[235]), 
        .Q(round_reg[235]) );
  DFF \round_reg_reg[236]  ( .D(out[236]), .CLK(clk), .RST(rst), .I(in[236]), 
        .Q(round_reg[236]) );
  DFF \round_reg_reg[237]  ( .D(out[237]), .CLK(clk), .RST(rst), .I(in[237]), 
        .Q(round_reg[237]) );
  DFF \round_reg_reg[238]  ( .D(out[238]), .CLK(clk), .RST(rst), .I(in[238]), 
        .Q(round_reg[238]) );
  DFF \round_reg_reg[239]  ( .D(out[239]), .CLK(clk), .RST(rst), .I(in[239]), 
        .Q(round_reg[239]) );
  DFF \round_reg_reg[240]  ( .D(out[240]), .CLK(clk), .RST(rst), .I(in[240]), 
        .Q(round_reg[240]) );
  DFF \round_reg_reg[241]  ( .D(out[241]), .CLK(clk), .RST(rst), .I(in[241]), 
        .Q(round_reg[241]) );
  DFF \round_reg_reg[242]  ( .D(out[242]), .CLK(clk), .RST(rst), .I(in[242]), 
        .Q(round_reg[242]) );
  DFF \round_reg_reg[243]  ( .D(out[243]), .CLK(clk), .RST(rst), .I(in[243]), 
        .Q(round_reg[243]) );
  DFF \round_reg_reg[244]  ( .D(out[244]), .CLK(clk), .RST(rst), .I(in[244]), 
        .Q(round_reg[244]) );
  DFF \round_reg_reg[245]  ( .D(out[245]), .CLK(clk), .RST(rst), .I(in[245]), 
        .Q(round_reg[245]) );
  DFF \round_reg_reg[246]  ( .D(out[246]), .CLK(clk), .RST(rst), .I(in[246]), 
        .Q(round_reg[246]) );
  DFF \round_reg_reg[247]  ( .D(out[247]), .CLK(clk), .RST(rst), .I(in[247]), 
        .Q(round_reg[247]) );
  DFF \round_reg_reg[248]  ( .D(out[248]), .CLK(clk), .RST(rst), .I(in[248]), 
        .Q(round_reg[248]) );
  DFF \round_reg_reg[249]  ( .D(out[249]), .CLK(clk), .RST(rst), .I(in[249]), 
        .Q(round_reg[249]) );
  DFF \round_reg_reg[250]  ( .D(out[250]), .CLK(clk), .RST(rst), .I(in[250]), 
        .Q(round_reg[250]) );
  DFF \round_reg_reg[251]  ( .D(out[251]), .CLK(clk), .RST(rst), .I(in[251]), 
        .Q(round_reg[251]) );
  DFF \round_reg_reg[252]  ( .D(out[252]), .CLK(clk), .RST(rst), .I(in[252]), 
        .Q(round_reg[252]) );
  DFF \round_reg_reg[253]  ( .D(out[253]), .CLK(clk), .RST(rst), .I(in[253]), 
        .Q(round_reg[253]) );
  DFF \round_reg_reg[254]  ( .D(out[254]), .CLK(clk), .RST(rst), .I(in[254]), 
        .Q(round_reg[254]) );
  DFF \round_reg_reg[255]  ( .D(out[255]), .CLK(clk), .RST(rst), .I(in[255]), 
        .Q(round_reg[255]) );
  DFF \round_reg_reg[256]  ( .D(out[256]), .CLK(clk), .RST(rst), .I(in[256]), 
        .Q(round_reg[256]) );
  DFF \round_reg_reg[257]  ( .D(out[257]), .CLK(clk), .RST(rst), .I(in[257]), 
        .Q(round_reg[257]) );
  DFF \round_reg_reg[258]  ( .D(out[258]), .CLK(clk), .RST(rst), .I(in[258]), 
        .Q(round_reg[258]) );
  DFF \round_reg_reg[259]  ( .D(out[259]), .CLK(clk), .RST(rst), .I(in[259]), 
        .Q(round_reg[259]) );
  DFF \round_reg_reg[260]  ( .D(out[260]), .CLK(clk), .RST(rst), .I(in[260]), 
        .Q(round_reg[260]) );
  DFF \round_reg_reg[261]  ( .D(out[261]), .CLK(clk), .RST(rst), .I(in[261]), 
        .Q(round_reg[261]) );
  DFF \round_reg_reg[262]  ( .D(out[262]), .CLK(clk), .RST(rst), .I(in[262]), 
        .Q(round_reg[262]) );
  DFF \round_reg_reg[263]  ( .D(out[263]), .CLK(clk), .RST(rst), .I(in[263]), 
        .Q(round_reg[263]) );
  DFF \round_reg_reg[264]  ( .D(out[264]), .CLK(clk), .RST(rst), .I(in[264]), 
        .Q(round_reg[264]) );
  DFF \round_reg_reg[265]  ( .D(out[265]), .CLK(clk), .RST(rst), .I(in[265]), 
        .Q(round_reg[265]) );
  DFF \round_reg_reg[266]  ( .D(out[266]), .CLK(clk), .RST(rst), .I(in[266]), 
        .Q(round_reg[266]) );
  DFF \round_reg_reg[267]  ( .D(out[267]), .CLK(clk), .RST(rst), .I(in[267]), 
        .Q(round_reg[267]) );
  DFF \round_reg_reg[268]  ( .D(out[268]), .CLK(clk), .RST(rst), .I(in[268]), 
        .Q(round_reg[268]) );
  DFF \round_reg_reg[269]  ( .D(out[269]), .CLK(clk), .RST(rst), .I(in[269]), 
        .Q(round_reg[269]) );
  DFF \round_reg_reg[270]  ( .D(out[270]), .CLK(clk), .RST(rst), .I(in[270]), 
        .Q(round_reg[270]) );
  DFF \round_reg_reg[271]  ( .D(out[271]), .CLK(clk), .RST(rst), .I(in[271]), 
        .Q(round_reg[271]) );
  DFF \round_reg_reg[272]  ( .D(out[272]), .CLK(clk), .RST(rst), .I(in[272]), 
        .Q(round_reg[272]) );
  DFF \round_reg_reg[273]  ( .D(out[273]), .CLK(clk), .RST(rst), .I(in[273]), 
        .Q(round_reg[273]) );
  DFF \round_reg_reg[274]  ( .D(out[274]), .CLK(clk), .RST(rst), .I(in[274]), 
        .Q(round_reg[274]) );
  DFF \round_reg_reg[275]  ( .D(out[275]), .CLK(clk), .RST(rst), .I(in[275]), 
        .Q(round_reg[275]) );
  DFF \round_reg_reg[276]  ( .D(out[276]), .CLK(clk), .RST(rst), .I(in[276]), 
        .Q(round_reg[276]) );
  DFF \round_reg_reg[277]  ( .D(out[277]), .CLK(clk), .RST(rst), .I(in[277]), 
        .Q(round_reg[277]) );
  DFF \round_reg_reg[278]  ( .D(out[278]), .CLK(clk), .RST(rst), .I(in[278]), 
        .Q(round_reg[278]) );
  DFF \round_reg_reg[279]  ( .D(out[279]), .CLK(clk), .RST(rst), .I(in[279]), 
        .Q(round_reg[279]) );
  DFF \round_reg_reg[280]  ( .D(out[280]), .CLK(clk), .RST(rst), .I(in[280]), 
        .Q(round_reg[280]) );
  DFF \round_reg_reg[281]  ( .D(out[281]), .CLK(clk), .RST(rst), .I(in[281]), 
        .Q(round_reg[281]) );
  DFF \round_reg_reg[282]  ( .D(out[282]), .CLK(clk), .RST(rst), .I(in[282]), 
        .Q(round_reg[282]) );
  DFF \round_reg_reg[283]  ( .D(out[283]), .CLK(clk), .RST(rst), .I(in[283]), 
        .Q(round_reg[283]) );
  DFF \round_reg_reg[284]  ( .D(out[284]), .CLK(clk), .RST(rst), .I(in[284]), 
        .Q(round_reg[284]) );
  DFF \round_reg_reg[285]  ( .D(out[285]), .CLK(clk), .RST(rst), .I(in[285]), 
        .Q(round_reg[285]) );
  DFF \round_reg_reg[286]  ( .D(out[286]), .CLK(clk), .RST(rst), .I(in[286]), 
        .Q(round_reg[286]) );
  DFF \round_reg_reg[287]  ( .D(out[287]), .CLK(clk), .RST(rst), .I(in[287]), 
        .Q(round_reg[287]) );
  DFF \round_reg_reg[288]  ( .D(out[288]), .CLK(clk), .RST(rst), .I(in[288]), 
        .Q(round_reg[288]) );
  DFF \round_reg_reg[289]  ( .D(out[289]), .CLK(clk), .RST(rst), .I(in[289]), 
        .Q(round_reg[289]) );
  DFF \round_reg_reg[290]  ( .D(out[290]), .CLK(clk), .RST(rst), .I(in[290]), 
        .Q(round_reg[290]) );
  DFF \round_reg_reg[291]  ( .D(out[291]), .CLK(clk), .RST(rst), .I(in[291]), 
        .Q(round_reg[291]) );
  DFF \round_reg_reg[292]  ( .D(out[292]), .CLK(clk), .RST(rst), .I(in[292]), 
        .Q(round_reg[292]) );
  DFF \round_reg_reg[293]  ( .D(out[293]), .CLK(clk), .RST(rst), .I(in[293]), 
        .Q(round_reg[293]) );
  DFF \round_reg_reg[294]  ( .D(out[294]), .CLK(clk), .RST(rst), .I(in[294]), 
        .Q(round_reg[294]) );
  DFF \round_reg_reg[295]  ( .D(out[295]), .CLK(clk), .RST(rst), .I(in[295]), 
        .Q(round_reg[295]) );
  DFF \round_reg_reg[296]  ( .D(out[296]), .CLK(clk), .RST(rst), .I(in[296]), 
        .Q(round_reg[296]) );
  DFF \round_reg_reg[297]  ( .D(out[297]), .CLK(clk), .RST(rst), .I(in[297]), 
        .Q(round_reg[297]) );
  DFF \round_reg_reg[298]  ( .D(out[298]), .CLK(clk), .RST(rst), .I(in[298]), 
        .Q(round_reg[298]) );
  DFF \round_reg_reg[299]  ( .D(out[299]), .CLK(clk), .RST(rst), .I(in[299]), 
        .Q(round_reg[299]) );
  DFF \round_reg_reg[300]  ( .D(out[300]), .CLK(clk), .RST(rst), .I(in[300]), 
        .Q(round_reg[300]) );
  DFF \round_reg_reg[301]  ( .D(out[301]), .CLK(clk), .RST(rst), .I(in[301]), 
        .Q(round_reg[301]) );
  DFF \round_reg_reg[302]  ( .D(out[302]), .CLK(clk), .RST(rst), .I(in[302]), 
        .Q(round_reg[302]) );
  DFF \round_reg_reg[303]  ( .D(out[303]), .CLK(clk), .RST(rst), .I(in[303]), 
        .Q(round_reg[303]) );
  DFF \round_reg_reg[304]  ( .D(out[304]), .CLK(clk), .RST(rst), .I(in[304]), 
        .Q(round_reg[304]) );
  DFF \round_reg_reg[305]  ( .D(out[305]), .CLK(clk), .RST(rst), .I(in[305]), 
        .Q(round_reg[305]) );
  DFF \round_reg_reg[306]  ( .D(out[306]), .CLK(clk), .RST(rst), .I(in[306]), 
        .Q(round_reg[306]) );
  DFF \round_reg_reg[307]  ( .D(out[307]), .CLK(clk), .RST(rst), .I(in[307]), 
        .Q(round_reg[307]) );
  DFF \round_reg_reg[308]  ( .D(out[308]), .CLK(clk), .RST(rst), .I(in[308]), 
        .Q(round_reg[308]) );
  DFF \round_reg_reg[309]  ( .D(out[309]), .CLK(clk), .RST(rst), .I(in[309]), 
        .Q(round_reg[309]) );
  DFF \round_reg_reg[310]  ( .D(out[310]), .CLK(clk), .RST(rst), .I(in[310]), 
        .Q(round_reg[310]) );
  DFF \round_reg_reg[311]  ( .D(out[311]), .CLK(clk), .RST(rst), .I(in[311]), 
        .Q(round_reg[311]) );
  DFF \round_reg_reg[312]  ( .D(out[312]), .CLK(clk), .RST(rst), .I(in[312]), 
        .Q(round_reg[312]) );
  DFF \round_reg_reg[313]  ( .D(out[313]), .CLK(clk), .RST(rst), .I(in[313]), 
        .Q(round_reg[313]) );
  DFF \round_reg_reg[314]  ( .D(out[314]), .CLK(clk), .RST(rst), .I(in[314]), 
        .Q(round_reg[314]) );
  DFF \round_reg_reg[315]  ( .D(out[315]), .CLK(clk), .RST(rst), .I(in[315]), 
        .Q(round_reg[315]) );
  DFF \round_reg_reg[316]  ( .D(out[316]), .CLK(clk), .RST(rst), .I(in[316]), 
        .Q(round_reg[316]) );
  DFF \round_reg_reg[317]  ( .D(out[317]), .CLK(clk), .RST(rst), .I(in[317]), 
        .Q(round_reg[317]) );
  DFF \round_reg_reg[318]  ( .D(out[318]), .CLK(clk), .RST(rst), .I(in[318]), 
        .Q(round_reg[318]) );
  DFF \round_reg_reg[319]  ( .D(out[319]), .CLK(clk), .RST(rst), .I(in[319]), 
        .Q(round_reg[319]) );
  DFF \round_reg_reg[320]  ( .D(out[320]), .CLK(clk), .RST(rst), .I(in[320]), 
        .Q(round_reg[320]) );
  DFF \round_reg_reg[321]  ( .D(out[321]), .CLK(clk), .RST(rst), .I(in[321]), 
        .Q(round_reg[321]) );
  DFF \round_reg_reg[322]  ( .D(out[322]), .CLK(clk), .RST(rst), .I(in[322]), 
        .Q(round_reg[322]) );
  DFF \round_reg_reg[323]  ( .D(out[323]), .CLK(clk), .RST(rst), .I(in[323]), 
        .Q(round_reg[323]) );
  DFF \round_reg_reg[324]  ( .D(out[324]), .CLK(clk), .RST(rst), .I(in[324]), 
        .Q(round_reg[324]) );
  DFF \round_reg_reg[325]  ( .D(out[325]), .CLK(clk), .RST(rst), .I(in[325]), 
        .Q(round_reg[325]) );
  DFF \round_reg_reg[326]  ( .D(out[326]), .CLK(clk), .RST(rst), .I(in[326]), 
        .Q(round_reg[326]) );
  DFF \round_reg_reg[327]  ( .D(out[327]), .CLK(clk), .RST(rst), .I(in[327]), 
        .Q(round_reg[327]) );
  DFF \round_reg_reg[328]  ( .D(out[328]), .CLK(clk), .RST(rst), .I(in[328]), 
        .Q(round_reg[328]) );
  DFF \round_reg_reg[329]  ( .D(out[329]), .CLK(clk), .RST(rst), .I(in[329]), 
        .Q(round_reg[329]) );
  DFF \round_reg_reg[330]  ( .D(out[330]), .CLK(clk), .RST(rst), .I(in[330]), 
        .Q(round_reg[330]) );
  DFF \round_reg_reg[331]  ( .D(out[331]), .CLK(clk), .RST(rst), .I(in[331]), 
        .Q(round_reg[331]) );
  DFF \round_reg_reg[332]  ( .D(out[332]), .CLK(clk), .RST(rst), .I(in[332]), 
        .Q(round_reg[332]) );
  DFF \round_reg_reg[333]  ( .D(out[333]), .CLK(clk), .RST(rst), .I(in[333]), 
        .Q(round_reg[333]) );
  DFF \round_reg_reg[334]  ( .D(out[334]), .CLK(clk), .RST(rst), .I(in[334]), 
        .Q(round_reg[334]) );
  DFF \round_reg_reg[335]  ( .D(out[335]), .CLK(clk), .RST(rst), .I(in[335]), 
        .Q(round_reg[335]) );
  DFF \round_reg_reg[336]  ( .D(out[336]), .CLK(clk), .RST(rst), .I(in[336]), 
        .Q(round_reg[336]) );
  DFF \round_reg_reg[337]  ( .D(out[337]), .CLK(clk), .RST(rst), .I(in[337]), 
        .Q(round_reg[337]) );
  DFF \round_reg_reg[338]  ( .D(out[338]), .CLK(clk), .RST(rst), .I(in[338]), 
        .Q(round_reg[338]) );
  DFF \round_reg_reg[339]  ( .D(out[339]), .CLK(clk), .RST(rst), .I(in[339]), 
        .Q(round_reg[339]) );
  DFF \round_reg_reg[340]  ( .D(out[340]), .CLK(clk), .RST(rst), .I(in[340]), 
        .Q(round_reg[340]) );
  DFF \round_reg_reg[341]  ( .D(out[341]), .CLK(clk), .RST(rst), .I(in[341]), 
        .Q(round_reg[341]) );
  DFF \round_reg_reg[342]  ( .D(out[342]), .CLK(clk), .RST(rst), .I(in[342]), 
        .Q(round_reg[342]) );
  DFF \round_reg_reg[343]  ( .D(out[343]), .CLK(clk), .RST(rst), .I(in[343]), 
        .Q(round_reg[343]) );
  DFF \round_reg_reg[344]  ( .D(out[344]), .CLK(clk), .RST(rst), .I(in[344]), 
        .Q(round_reg[344]) );
  DFF \round_reg_reg[345]  ( .D(out[345]), .CLK(clk), .RST(rst), .I(in[345]), 
        .Q(round_reg[345]) );
  DFF \round_reg_reg[346]  ( .D(out[346]), .CLK(clk), .RST(rst), .I(in[346]), 
        .Q(round_reg[346]) );
  DFF \round_reg_reg[347]  ( .D(out[347]), .CLK(clk), .RST(rst), .I(in[347]), 
        .Q(round_reg[347]) );
  DFF \round_reg_reg[348]  ( .D(out[348]), .CLK(clk), .RST(rst), .I(in[348]), 
        .Q(round_reg[348]) );
  DFF \round_reg_reg[349]  ( .D(out[349]), .CLK(clk), .RST(rst), .I(in[349]), 
        .Q(round_reg[349]) );
  DFF \round_reg_reg[350]  ( .D(out[350]), .CLK(clk), .RST(rst), .I(in[350]), 
        .Q(round_reg[350]) );
  DFF \round_reg_reg[351]  ( .D(out[351]), .CLK(clk), .RST(rst), .I(in[351]), 
        .Q(round_reg[351]) );
  DFF \round_reg_reg[352]  ( .D(out[352]), .CLK(clk), .RST(rst), .I(in[352]), 
        .Q(round_reg[352]) );
  DFF \round_reg_reg[353]  ( .D(out[353]), .CLK(clk), .RST(rst), .I(in[353]), 
        .Q(round_reg[353]) );
  DFF \round_reg_reg[354]  ( .D(out[354]), .CLK(clk), .RST(rst), .I(in[354]), 
        .Q(round_reg[354]) );
  DFF \round_reg_reg[355]  ( .D(out[355]), .CLK(clk), .RST(rst), .I(in[355]), 
        .Q(round_reg[355]) );
  DFF \round_reg_reg[356]  ( .D(out[356]), .CLK(clk), .RST(rst), .I(in[356]), 
        .Q(round_reg[356]) );
  DFF \round_reg_reg[357]  ( .D(out[357]), .CLK(clk), .RST(rst), .I(in[357]), 
        .Q(round_reg[357]) );
  DFF \round_reg_reg[358]  ( .D(out[358]), .CLK(clk), .RST(rst), .I(in[358]), 
        .Q(round_reg[358]) );
  DFF \round_reg_reg[359]  ( .D(out[359]), .CLK(clk), .RST(rst), .I(in[359]), 
        .Q(round_reg[359]) );
  DFF \round_reg_reg[360]  ( .D(out[360]), .CLK(clk), .RST(rst), .I(in[360]), 
        .Q(round_reg[360]) );
  DFF \round_reg_reg[361]  ( .D(out[361]), .CLK(clk), .RST(rst), .I(in[361]), 
        .Q(round_reg[361]) );
  DFF \round_reg_reg[362]  ( .D(out[362]), .CLK(clk), .RST(rst), .I(in[362]), 
        .Q(round_reg[362]) );
  DFF \round_reg_reg[363]  ( .D(out[363]), .CLK(clk), .RST(rst), .I(in[363]), 
        .Q(round_reg[363]) );
  DFF \round_reg_reg[364]  ( .D(out[364]), .CLK(clk), .RST(rst), .I(in[364]), 
        .Q(round_reg[364]) );
  DFF \round_reg_reg[365]  ( .D(out[365]), .CLK(clk), .RST(rst), .I(in[365]), 
        .Q(round_reg[365]) );
  DFF \round_reg_reg[366]  ( .D(out[366]), .CLK(clk), .RST(rst), .I(in[366]), 
        .Q(round_reg[366]) );
  DFF \round_reg_reg[367]  ( .D(out[367]), .CLK(clk), .RST(rst), .I(in[367]), 
        .Q(round_reg[367]) );
  DFF \round_reg_reg[368]  ( .D(out[368]), .CLK(clk), .RST(rst), .I(in[368]), 
        .Q(round_reg[368]) );
  DFF \round_reg_reg[369]  ( .D(out[369]), .CLK(clk), .RST(rst), .I(in[369]), 
        .Q(round_reg[369]) );
  DFF \round_reg_reg[370]  ( .D(out[370]), .CLK(clk), .RST(rst), .I(in[370]), 
        .Q(round_reg[370]) );
  DFF \round_reg_reg[371]  ( .D(out[371]), .CLK(clk), .RST(rst), .I(in[371]), 
        .Q(round_reg[371]) );
  DFF \round_reg_reg[372]  ( .D(out[372]), .CLK(clk), .RST(rst), .I(in[372]), 
        .Q(round_reg[372]) );
  DFF \round_reg_reg[373]  ( .D(out[373]), .CLK(clk), .RST(rst), .I(in[373]), 
        .Q(round_reg[373]) );
  DFF \round_reg_reg[374]  ( .D(out[374]), .CLK(clk), .RST(rst), .I(in[374]), 
        .Q(round_reg[374]) );
  DFF \round_reg_reg[375]  ( .D(out[375]), .CLK(clk), .RST(rst), .I(in[375]), 
        .Q(round_reg[375]) );
  DFF \round_reg_reg[376]  ( .D(out[376]), .CLK(clk), .RST(rst), .I(in[376]), 
        .Q(round_reg[376]) );
  DFF \round_reg_reg[377]  ( .D(out[377]), .CLK(clk), .RST(rst), .I(in[377]), 
        .Q(round_reg[377]) );
  DFF \round_reg_reg[378]  ( .D(out[378]), .CLK(clk), .RST(rst), .I(in[378]), 
        .Q(round_reg[378]) );
  DFF \round_reg_reg[379]  ( .D(out[379]), .CLK(clk), .RST(rst), .I(in[379]), 
        .Q(round_reg[379]) );
  DFF \round_reg_reg[380]  ( .D(out[380]), .CLK(clk), .RST(rst), .I(in[380]), 
        .Q(round_reg[380]) );
  DFF \round_reg_reg[381]  ( .D(out[381]), .CLK(clk), .RST(rst), .I(in[381]), 
        .Q(round_reg[381]) );
  DFF \round_reg_reg[382]  ( .D(out[382]), .CLK(clk), .RST(rst), .I(in[382]), 
        .Q(round_reg[382]) );
  DFF \round_reg_reg[383]  ( .D(out[383]), .CLK(clk), .RST(rst), .I(in[383]), 
        .Q(round_reg[383]) );
  DFF \round_reg_reg[384]  ( .D(out[384]), .CLK(clk), .RST(rst), .I(in[384]), 
        .Q(round_reg[384]) );
  DFF \round_reg_reg[385]  ( .D(out[385]), .CLK(clk), .RST(rst), .I(in[385]), 
        .Q(round_reg[385]) );
  DFF \round_reg_reg[386]  ( .D(out[386]), .CLK(clk), .RST(rst), .I(in[386]), 
        .Q(round_reg[386]) );
  DFF \round_reg_reg[387]  ( .D(out[387]), .CLK(clk), .RST(rst), .I(in[387]), 
        .Q(round_reg[387]) );
  DFF \round_reg_reg[388]  ( .D(out[388]), .CLK(clk), .RST(rst), .I(in[388]), 
        .Q(round_reg[388]) );
  DFF \round_reg_reg[389]  ( .D(out[389]), .CLK(clk), .RST(rst), .I(in[389]), 
        .Q(round_reg[389]) );
  DFF \round_reg_reg[390]  ( .D(out[390]), .CLK(clk), .RST(rst), .I(in[390]), 
        .Q(round_reg[390]) );
  DFF \round_reg_reg[391]  ( .D(out[391]), .CLK(clk), .RST(rst), .I(in[391]), 
        .Q(round_reg[391]) );
  DFF \round_reg_reg[392]  ( .D(out[392]), .CLK(clk), .RST(rst), .I(in[392]), 
        .Q(round_reg[392]) );
  DFF \round_reg_reg[393]  ( .D(out[393]), .CLK(clk), .RST(rst), .I(in[393]), 
        .Q(round_reg[393]) );
  DFF \round_reg_reg[394]  ( .D(out[394]), .CLK(clk), .RST(rst), .I(in[394]), 
        .Q(round_reg[394]) );
  DFF \round_reg_reg[395]  ( .D(out[395]), .CLK(clk), .RST(rst), .I(in[395]), 
        .Q(round_reg[395]) );
  DFF \round_reg_reg[396]  ( .D(out[396]), .CLK(clk), .RST(rst), .I(in[396]), 
        .Q(round_reg[396]) );
  DFF \round_reg_reg[397]  ( .D(out[397]), .CLK(clk), .RST(rst), .I(in[397]), 
        .Q(round_reg[397]) );
  DFF \round_reg_reg[398]  ( .D(out[398]), .CLK(clk), .RST(rst), .I(in[398]), 
        .Q(round_reg[398]) );
  DFF \round_reg_reg[399]  ( .D(out[399]), .CLK(clk), .RST(rst), .I(in[399]), 
        .Q(round_reg[399]) );
  DFF \round_reg_reg[400]  ( .D(out[400]), .CLK(clk), .RST(rst), .I(in[400]), 
        .Q(round_reg[400]) );
  DFF \round_reg_reg[401]  ( .D(out[401]), .CLK(clk), .RST(rst), .I(in[401]), 
        .Q(round_reg[401]) );
  DFF \round_reg_reg[402]  ( .D(out[402]), .CLK(clk), .RST(rst), .I(in[402]), 
        .Q(round_reg[402]) );
  DFF \round_reg_reg[403]  ( .D(out[403]), .CLK(clk), .RST(rst), .I(in[403]), 
        .Q(round_reg[403]) );
  DFF \round_reg_reg[404]  ( .D(out[404]), .CLK(clk), .RST(rst), .I(in[404]), 
        .Q(round_reg[404]) );
  DFF \round_reg_reg[405]  ( .D(out[405]), .CLK(clk), .RST(rst), .I(in[405]), 
        .Q(round_reg[405]) );
  DFF \round_reg_reg[406]  ( .D(out[406]), .CLK(clk), .RST(rst), .I(in[406]), 
        .Q(round_reg[406]) );
  DFF \round_reg_reg[407]  ( .D(out[407]), .CLK(clk), .RST(rst), .I(in[407]), 
        .Q(round_reg[407]) );
  DFF \round_reg_reg[408]  ( .D(out[408]), .CLK(clk), .RST(rst), .I(in[408]), 
        .Q(round_reg[408]) );
  DFF \round_reg_reg[409]  ( .D(out[409]), .CLK(clk), .RST(rst), .I(in[409]), 
        .Q(round_reg[409]) );
  DFF \round_reg_reg[410]  ( .D(out[410]), .CLK(clk), .RST(rst), .I(in[410]), 
        .Q(round_reg[410]) );
  DFF \round_reg_reg[411]  ( .D(out[411]), .CLK(clk), .RST(rst), .I(in[411]), 
        .Q(round_reg[411]) );
  DFF \round_reg_reg[412]  ( .D(out[412]), .CLK(clk), .RST(rst), .I(in[412]), 
        .Q(round_reg[412]) );
  DFF \round_reg_reg[413]  ( .D(out[413]), .CLK(clk), .RST(rst), .I(in[413]), 
        .Q(round_reg[413]) );
  DFF \round_reg_reg[414]  ( .D(out[414]), .CLK(clk), .RST(rst), .I(in[414]), 
        .Q(round_reg[414]) );
  DFF \round_reg_reg[415]  ( .D(out[415]), .CLK(clk), .RST(rst), .I(in[415]), 
        .Q(round_reg[415]) );
  DFF \round_reg_reg[416]  ( .D(out[416]), .CLK(clk), .RST(rst), .I(in[416]), 
        .Q(round_reg[416]) );
  DFF \round_reg_reg[417]  ( .D(out[417]), .CLK(clk), .RST(rst), .I(in[417]), 
        .Q(round_reg[417]) );
  DFF \round_reg_reg[418]  ( .D(out[418]), .CLK(clk), .RST(rst), .I(in[418]), 
        .Q(round_reg[418]) );
  DFF \round_reg_reg[419]  ( .D(out[419]), .CLK(clk), .RST(rst), .I(in[419]), 
        .Q(round_reg[419]) );
  DFF \round_reg_reg[420]  ( .D(out[420]), .CLK(clk), .RST(rst), .I(in[420]), 
        .Q(round_reg[420]) );
  DFF \round_reg_reg[421]  ( .D(out[421]), .CLK(clk), .RST(rst), .I(in[421]), 
        .Q(round_reg[421]) );
  DFF \round_reg_reg[422]  ( .D(out[422]), .CLK(clk), .RST(rst), .I(in[422]), 
        .Q(round_reg[422]) );
  DFF \round_reg_reg[423]  ( .D(out[423]), .CLK(clk), .RST(rst), .I(in[423]), 
        .Q(round_reg[423]) );
  DFF \round_reg_reg[424]  ( .D(out[424]), .CLK(clk), .RST(rst), .I(in[424]), 
        .Q(round_reg[424]) );
  DFF \round_reg_reg[425]  ( .D(out[425]), .CLK(clk), .RST(rst), .I(in[425]), 
        .Q(round_reg[425]) );
  DFF \round_reg_reg[426]  ( .D(out[426]), .CLK(clk), .RST(rst), .I(in[426]), 
        .Q(round_reg[426]) );
  DFF \round_reg_reg[427]  ( .D(out[427]), .CLK(clk), .RST(rst), .I(in[427]), 
        .Q(round_reg[427]) );
  DFF \round_reg_reg[428]  ( .D(out[428]), .CLK(clk), .RST(rst), .I(in[428]), 
        .Q(round_reg[428]) );
  DFF \round_reg_reg[429]  ( .D(out[429]), .CLK(clk), .RST(rst), .I(in[429]), 
        .Q(round_reg[429]) );
  DFF \round_reg_reg[430]  ( .D(out[430]), .CLK(clk), .RST(rst), .I(in[430]), 
        .Q(round_reg[430]) );
  DFF \round_reg_reg[431]  ( .D(out[431]), .CLK(clk), .RST(rst), .I(in[431]), 
        .Q(round_reg[431]) );
  DFF \round_reg_reg[432]  ( .D(out[432]), .CLK(clk), .RST(rst), .I(in[432]), 
        .Q(round_reg[432]) );
  DFF \round_reg_reg[433]  ( .D(out[433]), .CLK(clk), .RST(rst), .I(in[433]), 
        .Q(round_reg[433]) );
  DFF \round_reg_reg[434]  ( .D(out[434]), .CLK(clk), .RST(rst), .I(in[434]), 
        .Q(round_reg[434]) );
  DFF \round_reg_reg[435]  ( .D(out[435]), .CLK(clk), .RST(rst), .I(in[435]), 
        .Q(round_reg[435]) );
  DFF \round_reg_reg[436]  ( .D(out[436]), .CLK(clk), .RST(rst), .I(in[436]), 
        .Q(round_reg[436]) );
  DFF \round_reg_reg[437]  ( .D(out[437]), .CLK(clk), .RST(rst), .I(in[437]), 
        .Q(round_reg[437]) );
  DFF \round_reg_reg[438]  ( .D(out[438]), .CLK(clk), .RST(rst), .I(in[438]), 
        .Q(round_reg[438]) );
  DFF \round_reg_reg[439]  ( .D(out[439]), .CLK(clk), .RST(rst), .I(in[439]), 
        .Q(round_reg[439]) );
  DFF \round_reg_reg[440]  ( .D(out[440]), .CLK(clk), .RST(rst), .I(in[440]), 
        .Q(round_reg[440]) );
  DFF \round_reg_reg[441]  ( .D(out[441]), .CLK(clk), .RST(rst), .I(in[441]), 
        .Q(round_reg[441]) );
  DFF \round_reg_reg[442]  ( .D(out[442]), .CLK(clk), .RST(rst), .I(in[442]), 
        .Q(round_reg[442]) );
  DFF \round_reg_reg[443]  ( .D(out[443]), .CLK(clk), .RST(rst), .I(in[443]), 
        .Q(round_reg[443]) );
  DFF \round_reg_reg[444]  ( .D(out[444]), .CLK(clk), .RST(rst), .I(in[444]), 
        .Q(round_reg[444]) );
  DFF \round_reg_reg[445]  ( .D(out[445]), .CLK(clk), .RST(rst), .I(in[445]), 
        .Q(round_reg[445]) );
  DFF \round_reg_reg[446]  ( .D(out[446]), .CLK(clk), .RST(rst), .I(in[446]), 
        .Q(round_reg[446]) );
  DFF \round_reg_reg[447]  ( .D(out[447]), .CLK(clk), .RST(rst), .I(in[447]), 
        .Q(round_reg[447]) );
  DFF \round_reg_reg[448]  ( .D(out[448]), .CLK(clk), .RST(rst), .I(in[448]), 
        .Q(round_reg[448]) );
  DFF \round_reg_reg[449]  ( .D(out[449]), .CLK(clk), .RST(rst), .I(in[449]), 
        .Q(round_reg[449]) );
  DFF \round_reg_reg[450]  ( .D(out[450]), .CLK(clk), .RST(rst), .I(in[450]), 
        .Q(round_reg[450]) );
  DFF \round_reg_reg[451]  ( .D(out[451]), .CLK(clk), .RST(rst), .I(in[451]), 
        .Q(round_reg[451]) );
  DFF \round_reg_reg[452]  ( .D(out[452]), .CLK(clk), .RST(rst), .I(in[452]), 
        .Q(round_reg[452]) );
  DFF \round_reg_reg[453]  ( .D(out[453]), .CLK(clk), .RST(rst), .I(in[453]), 
        .Q(round_reg[453]) );
  DFF \round_reg_reg[454]  ( .D(out[454]), .CLK(clk), .RST(rst), .I(in[454]), 
        .Q(round_reg[454]) );
  DFF \round_reg_reg[455]  ( .D(out[455]), .CLK(clk), .RST(rst), .I(in[455]), 
        .Q(round_reg[455]) );
  DFF \round_reg_reg[456]  ( .D(out[456]), .CLK(clk), .RST(rst), .I(in[456]), 
        .Q(round_reg[456]) );
  DFF \round_reg_reg[457]  ( .D(out[457]), .CLK(clk), .RST(rst), .I(in[457]), 
        .Q(round_reg[457]) );
  DFF \round_reg_reg[458]  ( .D(out[458]), .CLK(clk), .RST(rst), .I(in[458]), 
        .Q(round_reg[458]) );
  DFF \round_reg_reg[459]  ( .D(out[459]), .CLK(clk), .RST(rst), .I(in[459]), 
        .Q(round_reg[459]) );
  DFF \round_reg_reg[460]  ( .D(out[460]), .CLK(clk), .RST(rst), .I(in[460]), 
        .Q(round_reg[460]) );
  DFF \round_reg_reg[461]  ( .D(out[461]), .CLK(clk), .RST(rst), .I(in[461]), 
        .Q(round_reg[461]) );
  DFF \round_reg_reg[462]  ( .D(out[462]), .CLK(clk), .RST(rst), .I(in[462]), 
        .Q(round_reg[462]) );
  DFF \round_reg_reg[463]  ( .D(out[463]), .CLK(clk), .RST(rst), .I(in[463]), 
        .Q(round_reg[463]) );
  DFF \round_reg_reg[464]  ( .D(out[464]), .CLK(clk), .RST(rst), .I(in[464]), 
        .Q(round_reg[464]) );
  DFF \round_reg_reg[465]  ( .D(out[465]), .CLK(clk), .RST(rst), .I(in[465]), 
        .Q(round_reg[465]) );
  DFF \round_reg_reg[466]  ( .D(out[466]), .CLK(clk), .RST(rst), .I(in[466]), 
        .Q(round_reg[466]) );
  DFF \round_reg_reg[467]  ( .D(out[467]), .CLK(clk), .RST(rst), .I(in[467]), 
        .Q(round_reg[467]) );
  DFF \round_reg_reg[468]  ( .D(out[468]), .CLK(clk), .RST(rst), .I(in[468]), 
        .Q(round_reg[468]) );
  DFF \round_reg_reg[469]  ( .D(out[469]), .CLK(clk), .RST(rst), .I(in[469]), 
        .Q(round_reg[469]) );
  DFF \round_reg_reg[470]  ( .D(out[470]), .CLK(clk), .RST(rst), .I(in[470]), 
        .Q(round_reg[470]) );
  DFF \round_reg_reg[471]  ( .D(out[471]), .CLK(clk), .RST(rst), .I(in[471]), 
        .Q(round_reg[471]) );
  DFF \round_reg_reg[472]  ( .D(out[472]), .CLK(clk), .RST(rst), .I(in[472]), 
        .Q(round_reg[472]) );
  DFF \round_reg_reg[473]  ( .D(out[473]), .CLK(clk), .RST(rst), .I(in[473]), 
        .Q(round_reg[473]) );
  DFF \round_reg_reg[474]  ( .D(out[474]), .CLK(clk), .RST(rst), .I(in[474]), 
        .Q(round_reg[474]) );
  DFF \round_reg_reg[475]  ( .D(out[475]), .CLK(clk), .RST(rst), .I(in[475]), 
        .Q(round_reg[475]) );
  DFF \round_reg_reg[476]  ( .D(out[476]), .CLK(clk), .RST(rst), .I(in[476]), 
        .Q(round_reg[476]) );
  DFF \round_reg_reg[477]  ( .D(out[477]), .CLK(clk), .RST(rst), .I(in[477]), 
        .Q(round_reg[477]) );
  DFF \round_reg_reg[478]  ( .D(out[478]), .CLK(clk), .RST(rst), .I(in[478]), 
        .Q(round_reg[478]) );
  DFF \round_reg_reg[479]  ( .D(out[479]), .CLK(clk), .RST(rst), .I(in[479]), 
        .Q(round_reg[479]) );
  DFF \round_reg_reg[480]  ( .D(out[480]), .CLK(clk), .RST(rst), .I(in[480]), 
        .Q(round_reg[480]) );
  DFF \round_reg_reg[481]  ( .D(out[481]), .CLK(clk), .RST(rst), .I(in[481]), 
        .Q(round_reg[481]) );
  DFF \round_reg_reg[482]  ( .D(out[482]), .CLK(clk), .RST(rst), .I(in[482]), 
        .Q(round_reg[482]) );
  DFF \round_reg_reg[483]  ( .D(out[483]), .CLK(clk), .RST(rst), .I(in[483]), 
        .Q(round_reg[483]) );
  DFF \round_reg_reg[484]  ( .D(out[484]), .CLK(clk), .RST(rst), .I(in[484]), 
        .Q(round_reg[484]) );
  DFF \round_reg_reg[485]  ( .D(out[485]), .CLK(clk), .RST(rst), .I(in[485]), 
        .Q(round_reg[485]) );
  DFF \round_reg_reg[486]  ( .D(out[486]), .CLK(clk), .RST(rst), .I(in[486]), 
        .Q(round_reg[486]) );
  DFF \round_reg_reg[487]  ( .D(out[487]), .CLK(clk), .RST(rst), .I(in[487]), 
        .Q(round_reg[487]) );
  DFF \round_reg_reg[488]  ( .D(out[488]), .CLK(clk), .RST(rst), .I(in[488]), 
        .Q(round_reg[488]) );
  DFF \round_reg_reg[489]  ( .D(out[489]), .CLK(clk), .RST(rst), .I(in[489]), 
        .Q(round_reg[489]) );
  DFF \round_reg_reg[490]  ( .D(out[490]), .CLK(clk), .RST(rst), .I(in[490]), 
        .Q(round_reg[490]) );
  DFF \round_reg_reg[491]  ( .D(out[491]), .CLK(clk), .RST(rst), .I(in[491]), 
        .Q(round_reg[491]) );
  DFF \round_reg_reg[492]  ( .D(out[492]), .CLK(clk), .RST(rst), .I(in[492]), 
        .Q(round_reg[492]) );
  DFF \round_reg_reg[493]  ( .D(out[493]), .CLK(clk), .RST(rst), .I(in[493]), 
        .Q(round_reg[493]) );
  DFF \round_reg_reg[494]  ( .D(out[494]), .CLK(clk), .RST(rst), .I(in[494]), 
        .Q(round_reg[494]) );
  DFF \round_reg_reg[495]  ( .D(out[495]), .CLK(clk), .RST(rst), .I(in[495]), 
        .Q(round_reg[495]) );
  DFF \round_reg_reg[496]  ( .D(out[496]), .CLK(clk), .RST(rst), .I(in[496]), 
        .Q(round_reg[496]) );
  DFF \round_reg_reg[497]  ( .D(out[497]), .CLK(clk), .RST(rst), .I(in[497]), 
        .Q(round_reg[497]) );
  DFF \round_reg_reg[498]  ( .D(out[498]), .CLK(clk), .RST(rst), .I(in[498]), 
        .Q(round_reg[498]) );
  DFF \round_reg_reg[499]  ( .D(out[499]), .CLK(clk), .RST(rst), .I(in[499]), 
        .Q(round_reg[499]) );
  DFF \round_reg_reg[500]  ( .D(out[500]), .CLK(clk), .RST(rst), .I(in[500]), 
        .Q(round_reg[500]) );
  DFF \round_reg_reg[501]  ( .D(out[501]), .CLK(clk), .RST(rst), .I(in[501]), 
        .Q(round_reg[501]) );
  DFF \round_reg_reg[502]  ( .D(out[502]), .CLK(clk), .RST(rst), .I(in[502]), 
        .Q(round_reg[502]) );
  DFF \round_reg_reg[503]  ( .D(out[503]), .CLK(clk), .RST(rst), .I(in[503]), 
        .Q(round_reg[503]) );
  DFF \round_reg_reg[504]  ( .D(out[504]), .CLK(clk), .RST(rst), .I(in[504]), 
        .Q(round_reg[504]) );
  DFF \round_reg_reg[505]  ( .D(out[505]), .CLK(clk), .RST(rst), .I(in[505]), 
        .Q(round_reg[505]) );
  DFF \round_reg_reg[506]  ( .D(out[506]), .CLK(clk), .RST(rst), .I(in[506]), 
        .Q(round_reg[506]) );
  DFF \round_reg_reg[507]  ( .D(out[507]), .CLK(clk), .RST(rst), .I(in[507]), 
        .Q(round_reg[507]) );
  DFF \round_reg_reg[508]  ( .D(out[508]), .CLK(clk), .RST(rst), .I(in[508]), 
        .Q(round_reg[508]) );
  DFF \round_reg_reg[509]  ( .D(out[509]), .CLK(clk), .RST(rst), .I(in[509]), 
        .Q(round_reg[509]) );
  DFF \round_reg_reg[510]  ( .D(out[510]), .CLK(clk), .RST(rst), .I(in[510]), 
        .Q(round_reg[510]) );
  DFF \round_reg_reg[511]  ( .D(out[511]), .CLK(clk), .RST(rst), .I(in[511]), 
        .Q(round_reg[511]) );
  DFF \round_reg_reg[512]  ( .D(out[512]), .CLK(clk), .RST(rst), .I(in[512]), 
        .Q(round_reg[512]) );
  DFF \round_reg_reg[513]  ( .D(out[513]), .CLK(clk), .RST(rst), .I(in[513]), 
        .Q(round_reg[513]) );
  DFF \round_reg_reg[514]  ( .D(out[514]), .CLK(clk), .RST(rst), .I(in[514]), 
        .Q(round_reg[514]) );
  DFF \round_reg_reg[515]  ( .D(out[515]), .CLK(clk), .RST(rst), .I(in[515]), 
        .Q(round_reg[515]) );
  DFF \round_reg_reg[516]  ( .D(out[516]), .CLK(clk), .RST(rst), .I(in[516]), 
        .Q(round_reg[516]) );
  DFF \round_reg_reg[517]  ( .D(out[517]), .CLK(clk), .RST(rst), .I(in[517]), 
        .Q(round_reg[517]) );
  DFF \round_reg_reg[518]  ( .D(out[518]), .CLK(clk), .RST(rst), .I(in[518]), 
        .Q(round_reg[518]) );
  DFF \round_reg_reg[519]  ( .D(out[519]), .CLK(clk), .RST(rst), .I(in[519]), 
        .Q(round_reg[519]) );
  DFF \round_reg_reg[520]  ( .D(out[520]), .CLK(clk), .RST(rst), .I(in[520]), 
        .Q(round_reg[520]) );
  DFF \round_reg_reg[521]  ( .D(out[521]), .CLK(clk), .RST(rst), .I(in[521]), 
        .Q(round_reg[521]) );
  DFF \round_reg_reg[522]  ( .D(out[522]), .CLK(clk), .RST(rst), .I(in[522]), 
        .Q(round_reg[522]) );
  DFF \round_reg_reg[523]  ( .D(out[523]), .CLK(clk), .RST(rst), .I(in[523]), 
        .Q(round_reg[523]) );
  DFF \round_reg_reg[524]  ( .D(out[524]), .CLK(clk), .RST(rst), .I(in[524]), 
        .Q(round_reg[524]) );
  DFF \round_reg_reg[525]  ( .D(out[525]), .CLK(clk), .RST(rst), .I(in[525]), 
        .Q(round_reg[525]) );
  DFF \round_reg_reg[526]  ( .D(out[526]), .CLK(clk), .RST(rst), .I(in[526]), 
        .Q(round_reg[526]) );
  DFF \round_reg_reg[527]  ( .D(out[527]), .CLK(clk), .RST(rst), .I(in[527]), 
        .Q(round_reg[527]) );
  DFF \round_reg_reg[528]  ( .D(out[528]), .CLK(clk), .RST(rst), .I(in[528]), 
        .Q(round_reg[528]) );
  DFF \round_reg_reg[529]  ( .D(out[529]), .CLK(clk), .RST(rst), .I(in[529]), 
        .Q(round_reg[529]) );
  DFF \round_reg_reg[530]  ( .D(out[530]), .CLK(clk), .RST(rst), .I(in[530]), 
        .Q(round_reg[530]) );
  DFF \round_reg_reg[531]  ( .D(out[531]), .CLK(clk), .RST(rst), .I(in[531]), 
        .Q(round_reg[531]) );
  DFF \round_reg_reg[532]  ( .D(out[532]), .CLK(clk), .RST(rst), .I(in[532]), 
        .Q(round_reg[532]) );
  DFF \round_reg_reg[533]  ( .D(out[533]), .CLK(clk), .RST(rst), .I(in[533]), 
        .Q(round_reg[533]) );
  DFF \round_reg_reg[534]  ( .D(out[534]), .CLK(clk), .RST(rst), .I(in[534]), 
        .Q(round_reg[534]) );
  DFF \round_reg_reg[535]  ( .D(out[535]), .CLK(clk), .RST(rst), .I(in[535]), 
        .Q(round_reg[535]) );
  DFF \round_reg_reg[536]  ( .D(out[536]), .CLK(clk), .RST(rst), .I(in[536]), 
        .Q(round_reg[536]) );
  DFF \round_reg_reg[537]  ( .D(out[537]), .CLK(clk), .RST(rst), .I(in[537]), 
        .Q(round_reg[537]) );
  DFF \round_reg_reg[538]  ( .D(out[538]), .CLK(clk), .RST(rst), .I(in[538]), 
        .Q(round_reg[538]) );
  DFF \round_reg_reg[539]  ( .D(out[539]), .CLK(clk), .RST(rst), .I(in[539]), 
        .Q(round_reg[539]) );
  DFF \round_reg_reg[540]  ( .D(out[540]), .CLK(clk), .RST(rst), .I(in[540]), 
        .Q(round_reg[540]) );
  DFF \round_reg_reg[541]  ( .D(out[541]), .CLK(clk), .RST(rst), .I(in[541]), 
        .Q(round_reg[541]) );
  DFF \round_reg_reg[542]  ( .D(out[542]), .CLK(clk), .RST(rst), .I(in[542]), 
        .Q(round_reg[542]) );
  DFF \round_reg_reg[543]  ( .D(out[543]), .CLK(clk), .RST(rst), .I(in[543]), 
        .Q(round_reg[543]) );
  DFF \round_reg_reg[544]  ( .D(out[544]), .CLK(clk), .RST(rst), .I(in[544]), 
        .Q(round_reg[544]) );
  DFF \round_reg_reg[545]  ( .D(out[545]), .CLK(clk), .RST(rst), .I(in[545]), 
        .Q(round_reg[545]) );
  DFF \round_reg_reg[546]  ( .D(out[546]), .CLK(clk), .RST(rst), .I(in[546]), 
        .Q(round_reg[546]) );
  DFF \round_reg_reg[547]  ( .D(out[547]), .CLK(clk), .RST(rst), .I(in[547]), 
        .Q(round_reg[547]) );
  DFF \round_reg_reg[548]  ( .D(out[548]), .CLK(clk), .RST(rst), .I(in[548]), 
        .Q(round_reg[548]) );
  DFF \round_reg_reg[549]  ( .D(out[549]), .CLK(clk), .RST(rst), .I(in[549]), 
        .Q(round_reg[549]) );
  DFF \round_reg_reg[550]  ( .D(out[550]), .CLK(clk), .RST(rst), .I(in[550]), 
        .Q(round_reg[550]) );
  DFF \round_reg_reg[551]  ( .D(out[551]), .CLK(clk), .RST(rst), .I(in[551]), 
        .Q(round_reg[551]) );
  DFF \round_reg_reg[552]  ( .D(out[552]), .CLK(clk), .RST(rst), .I(in[552]), 
        .Q(round_reg[552]) );
  DFF \round_reg_reg[553]  ( .D(out[553]), .CLK(clk), .RST(rst), .I(in[553]), 
        .Q(round_reg[553]) );
  DFF \round_reg_reg[554]  ( .D(out[554]), .CLK(clk), .RST(rst), .I(in[554]), 
        .Q(round_reg[554]) );
  DFF \round_reg_reg[555]  ( .D(out[555]), .CLK(clk), .RST(rst), .I(in[555]), 
        .Q(round_reg[555]) );
  DFF \round_reg_reg[556]  ( .D(out[556]), .CLK(clk), .RST(rst), .I(in[556]), 
        .Q(round_reg[556]) );
  DFF \round_reg_reg[557]  ( .D(out[557]), .CLK(clk), .RST(rst), .I(in[557]), 
        .Q(round_reg[557]) );
  DFF \round_reg_reg[558]  ( .D(out[558]), .CLK(clk), .RST(rst), .I(in[558]), 
        .Q(round_reg[558]) );
  DFF \round_reg_reg[559]  ( .D(out[559]), .CLK(clk), .RST(rst), .I(in[559]), 
        .Q(round_reg[559]) );
  DFF \round_reg_reg[560]  ( .D(out[560]), .CLK(clk), .RST(rst), .I(in[560]), 
        .Q(round_reg[560]) );
  DFF \round_reg_reg[561]  ( .D(out[561]), .CLK(clk), .RST(rst), .I(in[561]), 
        .Q(round_reg[561]) );
  DFF \round_reg_reg[562]  ( .D(out[562]), .CLK(clk), .RST(rst), .I(in[562]), 
        .Q(round_reg[562]) );
  DFF \round_reg_reg[563]  ( .D(out[563]), .CLK(clk), .RST(rst), .I(in[563]), 
        .Q(round_reg[563]) );
  DFF \round_reg_reg[564]  ( .D(out[564]), .CLK(clk), .RST(rst), .I(in[564]), 
        .Q(round_reg[564]) );
  DFF \round_reg_reg[565]  ( .D(out[565]), .CLK(clk), .RST(rst), .I(in[565]), 
        .Q(round_reg[565]) );
  DFF \round_reg_reg[566]  ( .D(out[566]), .CLK(clk), .RST(rst), .I(in[566]), 
        .Q(round_reg[566]) );
  DFF \round_reg_reg[567]  ( .D(out[567]), .CLK(clk), .RST(rst), .I(in[567]), 
        .Q(round_reg[567]) );
  DFF \round_reg_reg[568]  ( .D(out[568]), .CLK(clk), .RST(rst), .I(in[568]), 
        .Q(round_reg[568]) );
  DFF \round_reg_reg[569]  ( .D(out[569]), .CLK(clk), .RST(rst), .I(in[569]), 
        .Q(round_reg[569]) );
  DFF \round_reg_reg[570]  ( .D(out[570]), .CLK(clk), .RST(rst), .I(in[570]), 
        .Q(round_reg[570]) );
  DFF \round_reg_reg[571]  ( .D(out[571]), .CLK(clk), .RST(rst), .I(in[571]), 
        .Q(round_reg[571]) );
  DFF \round_reg_reg[572]  ( .D(out[572]), .CLK(clk), .RST(rst), .I(in[572]), 
        .Q(round_reg[572]) );
  DFF \round_reg_reg[573]  ( .D(out[573]), .CLK(clk), .RST(rst), .I(in[573]), 
        .Q(round_reg[573]) );
  DFF \round_reg_reg[574]  ( .D(out[574]), .CLK(clk), .RST(rst), .I(in[574]), 
        .Q(round_reg[574]) );
  DFF \round_reg_reg[575]  ( .D(out[575]), .CLK(clk), .RST(rst), .I(in[575]), 
        .Q(round_reg[575]) );
  DFF \round_reg_reg[576]  ( .D(out[576]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[576]) );
  DFF \round_reg_reg[577]  ( .D(out[577]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[577]) );
  DFF \round_reg_reg[578]  ( .D(out[578]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[578]) );
  DFF \round_reg_reg[579]  ( .D(out[579]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[579]) );
  DFF \round_reg_reg[580]  ( .D(out[580]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[580]) );
  DFF \round_reg_reg[581]  ( .D(out[581]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[581]) );
  DFF \round_reg_reg[582]  ( .D(out[582]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[582]) );
  DFF \round_reg_reg[583]  ( .D(out[583]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[583]) );
  DFF \round_reg_reg[584]  ( .D(out[584]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[584]) );
  DFF \round_reg_reg[585]  ( .D(out[585]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[585]) );
  DFF \round_reg_reg[586]  ( .D(out[586]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[586]) );
  DFF \round_reg_reg[587]  ( .D(out[587]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[587]) );
  DFF \round_reg_reg[588]  ( .D(out[588]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[588]) );
  DFF \round_reg_reg[589]  ( .D(out[589]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[589]) );
  DFF \round_reg_reg[590]  ( .D(out[590]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[590]) );
  DFF \round_reg_reg[591]  ( .D(out[591]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[591]) );
  DFF \round_reg_reg[592]  ( .D(out[592]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[592]) );
  DFF \round_reg_reg[593]  ( .D(out[593]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[593]) );
  DFF \round_reg_reg[594]  ( .D(out[594]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[594]) );
  DFF \round_reg_reg[595]  ( .D(out[595]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[595]) );
  DFF \round_reg_reg[596]  ( .D(out[596]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[596]) );
  DFF \round_reg_reg[597]  ( .D(out[597]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[597]) );
  DFF \round_reg_reg[598]  ( .D(out[598]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[598]) );
  DFF \round_reg_reg[599]  ( .D(out[599]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[599]) );
  DFF \round_reg_reg[600]  ( .D(out[600]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[600]) );
  DFF \round_reg_reg[601]  ( .D(out[601]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[601]) );
  DFF \round_reg_reg[602]  ( .D(out[602]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[602]) );
  DFF \round_reg_reg[603]  ( .D(out[603]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[603]) );
  DFF \round_reg_reg[604]  ( .D(out[604]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[604]) );
  DFF \round_reg_reg[605]  ( .D(out[605]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[605]) );
  DFF \round_reg_reg[606]  ( .D(out[606]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[606]) );
  DFF \round_reg_reg[607]  ( .D(out[607]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[607]) );
  DFF \round_reg_reg[608]  ( .D(out[608]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[608]) );
  DFF \round_reg_reg[609]  ( .D(out[609]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[609]) );
  DFF \round_reg_reg[610]  ( .D(out[610]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[610]) );
  DFF \round_reg_reg[611]  ( .D(out[611]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[611]) );
  DFF \round_reg_reg[612]  ( .D(out[612]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[612]) );
  DFF \round_reg_reg[613]  ( .D(out[613]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[613]) );
  DFF \round_reg_reg[614]  ( .D(out[614]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[614]) );
  DFF \round_reg_reg[615]  ( .D(out[615]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[615]) );
  DFF \round_reg_reg[616]  ( .D(out[616]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[616]) );
  DFF \round_reg_reg[617]  ( .D(out[617]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[617]) );
  DFF \round_reg_reg[618]  ( .D(out[618]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[618]) );
  DFF \round_reg_reg[619]  ( .D(out[619]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[619]) );
  DFF \round_reg_reg[620]  ( .D(out[620]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[620]) );
  DFF \round_reg_reg[621]  ( .D(out[621]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[621]) );
  DFF \round_reg_reg[622]  ( .D(out[622]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[622]) );
  DFF \round_reg_reg[623]  ( .D(out[623]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[623]) );
  DFF \round_reg_reg[624]  ( .D(out[624]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[624]) );
  DFF \round_reg_reg[625]  ( .D(out[625]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[625]) );
  DFF \round_reg_reg[626]  ( .D(out[626]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[626]) );
  DFF \round_reg_reg[627]  ( .D(out[627]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[627]) );
  DFF \round_reg_reg[628]  ( .D(out[628]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[628]) );
  DFF \round_reg_reg[629]  ( .D(out[629]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[629]) );
  DFF \round_reg_reg[630]  ( .D(out[630]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[630]) );
  DFF \round_reg_reg[631]  ( .D(out[631]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[631]) );
  DFF \round_reg_reg[632]  ( .D(out[632]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[632]) );
  DFF \round_reg_reg[633]  ( .D(out[633]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[633]) );
  DFF \round_reg_reg[634]  ( .D(out[634]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[634]) );
  DFF \round_reg_reg[635]  ( .D(out[635]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[635]) );
  DFF \round_reg_reg[636]  ( .D(out[636]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[636]) );
  DFF \round_reg_reg[637]  ( .D(out[637]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[637]) );
  DFF \round_reg_reg[638]  ( .D(out[638]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[638]) );
  DFF \round_reg_reg[639]  ( .D(out[639]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[639]) );
  DFF \round_reg_reg[640]  ( .D(out[640]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[640]) );
  DFF \round_reg_reg[641]  ( .D(out[641]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[641]) );
  DFF \round_reg_reg[642]  ( .D(out[642]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[642]) );
  DFF \round_reg_reg[643]  ( .D(out[643]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[643]) );
  DFF \round_reg_reg[644]  ( .D(out[644]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[644]) );
  DFF \round_reg_reg[645]  ( .D(out[645]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[645]) );
  DFF \round_reg_reg[646]  ( .D(out[646]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[646]) );
  DFF \round_reg_reg[647]  ( .D(out[647]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[647]) );
  DFF \round_reg_reg[648]  ( .D(out[648]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[648]) );
  DFF \round_reg_reg[649]  ( .D(out[649]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[649]) );
  DFF \round_reg_reg[650]  ( .D(out[650]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[650]) );
  DFF \round_reg_reg[651]  ( .D(out[651]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[651]) );
  DFF \round_reg_reg[652]  ( .D(out[652]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[652]) );
  DFF \round_reg_reg[653]  ( .D(out[653]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[653]) );
  DFF \round_reg_reg[654]  ( .D(out[654]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[654]) );
  DFF \round_reg_reg[655]  ( .D(out[655]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[655]) );
  DFF \round_reg_reg[656]  ( .D(out[656]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[656]) );
  DFF \round_reg_reg[657]  ( .D(out[657]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[657]) );
  DFF \round_reg_reg[658]  ( .D(out[658]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[658]) );
  DFF \round_reg_reg[659]  ( .D(out[659]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[659]) );
  DFF \round_reg_reg[660]  ( .D(out[660]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[660]) );
  DFF \round_reg_reg[661]  ( .D(out[661]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[661]) );
  DFF \round_reg_reg[662]  ( .D(out[662]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[662]) );
  DFF \round_reg_reg[663]  ( .D(out[663]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[663]) );
  DFF \round_reg_reg[664]  ( .D(out[664]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[664]) );
  DFF \round_reg_reg[665]  ( .D(out[665]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[665]) );
  DFF \round_reg_reg[666]  ( .D(out[666]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[666]) );
  DFF \round_reg_reg[667]  ( .D(out[667]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[667]) );
  DFF \round_reg_reg[668]  ( .D(out[668]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[668]) );
  DFF \round_reg_reg[669]  ( .D(out[669]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[669]) );
  DFF \round_reg_reg[670]  ( .D(out[670]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[670]) );
  DFF \round_reg_reg[671]  ( .D(out[671]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[671]) );
  DFF \round_reg_reg[672]  ( .D(out[672]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[672]) );
  DFF \round_reg_reg[673]  ( .D(out[673]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[673]) );
  DFF \round_reg_reg[674]  ( .D(out[674]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[674]) );
  DFF \round_reg_reg[675]  ( .D(out[675]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[675]) );
  DFF \round_reg_reg[676]  ( .D(out[676]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[676]) );
  DFF \round_reg_reg[677]  ( .D(out[677]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[677]) );
  DFF \round_reg_reg[678]  ( .D(out[678]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[678]) );
  DFF \round_reg_reg[679]  ( .D(out[679]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[679]) );
  DFF \round_reg_reg[680]  ( .D(out[680]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[680]) );
  DFF \round_reg_reg[681]  ( .D(out[681]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[681]) );
  DFF \round_reg_reg[682]  ( .D(out[682]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[682]) );
  DFF \round_reg_reg[683]  ( .D(out[683]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[683]) );
  DFF \round_reg_reg[684]  ( .D(out[684]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[684]) );
  DFF \round_reg_reg[685]  ( .D(out[685]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[685]) );
  DFF \round_reg_reg[686]  ( .D(out[686]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[686]) );
  DFF \round_reg_reg[687]  ( .D(out[687]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[687]) );
  DFF \round_reg_reg[688]  ( .D(out[688]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[688]) );
  DFF \round_reg_reg[689]  ( .D(out[689]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[689]) );
  DFF \round_reg_reg[690]  ( .D(out[690]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[690]) );
  DFF \round_reg_reg[691]  ( .D(out[691]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[691]) );
  DFF \round_reg_reg[692]  ( .D(out[692]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[692]) );
  DFF \round_reg_reg[693]  ( .D(out[693]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[693]) );
  DFF \round_reg_reg[694]  ( .D(out[694]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[694]) );
  DFF \round_reg_reg[695]  ( .D(out[695]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[695]) );
  DFF \round_reg_reg[696]  ( .D(out[696]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[696]) );
  DFF \round_reg_reg[697]  ( .D(out[697]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[697]) );
  DFF \round_reg_reg[698]  ( .D(out[698]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[698]) );
  DFF \round_reg_reg[699]  ( .D(out[699]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[699]) );
  DFF \round_reg_reg[700]  ( .D(out[700]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[700]) );
  DFF \round_reg_reg[701]  ( .D(out[701]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[701]) );
  DFF \round_reg_reg[702]  ( .D(out[702]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[702]) );
  DFF \round_reg_reg[703]  ( .D(out[703]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[703]) );
  DFF \round_reg_reg[704]  ( .D(out[704]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[704]) );
  DFF \round_reg_reg[705]  ( .D(out[705]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[705]) );
  DFF \round_reg_reg[706]  ( .D(out[706]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[706]) );
  DFF \round_reg_reg[707]  ( .D(out[707]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[707]) );
  DFF \round_reg_reg[708]  ( .D(out[708]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[708]) );
  DFF \round_reg_reg[709]  ( .D(out[709]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[709]) );
  DFF \round_reg_reg[710]  ( .D(out[710]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[710]) );
  DFF \round_reg_reg[711]  ( .D(out[711]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[711]) );
  DFF \round_reg_reg[712]  ( .D(out[712]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[712]) );
  DFF \round_reg_reg[713]  ( .D(out[713]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[713]) );
  DFF \round_reg_reg[714]  ( .D(out[714]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[714]) );
  DFF \round_reg_reg[715]  ( .D(out[715]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[715]) );
  DFF \round_reg_reg[716]  ( .D(out[716]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[716]) );
  DFF \round_reg_reg[717]  ( .D(out[717]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[717]) );
  DFF \round_reg_reg[718]  ( .D(out[718]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[718]) );
  DFF \round_reg_reg[719]  ( .D(out[719]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[719]) );
  DFF \round_reg_reg[720]  ( .D(out[720]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[720]) );
  DFF \round_reg_reg[721]  ( .D(out[721]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[721]) );
  DFF \round_reg_reg[722]  ( .D(out[722]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[722]) );
  DFF \round_reg_reg[723]  ( .D(out[723]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[723]) );
  DFF \round_reg_reg[724]  ( .D(out[724]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[724]) );
  DFF \round_reg_reg[725]  ( .D(out[725]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[725]) );
  DFF \round_reg_reg[726]  ( .D(out[726]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[726]) );
  DFF \round_reg_reg[727]  ( .D(out[727]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[727]) );
  DFF \round_reg_reg[728]  ( .D(out[728]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[728]) );
  DFF \round_reg_reg[729]  ( .D(out[729]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[729]) );
  DFF \round_reg_reg[730]  ( .D(out[730]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[730]) );
  DFF \round_reg_reg[731]  ( .D(out[731]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[731]) );
  DFF \round_reg_reg[732]  ( .D(out[732]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[732]) );
  DFF \round_reg_reg[733]  ( .D(out[733]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[733]) );
  DFF \round_reg_reg[734]  ( .D(out[734]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[734]) );
  DFF \round_reg_reg[735]  ( .D(out[735]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[735]) );
  DFF \round_reg_reg[736]  ( .D(out[736]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[736]) );
  DFF \round_reg_reg[737]  ( .D(out[737]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[737]) );
  DFF \round_reg_reg[738]  ( .D(out[738]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[738]) );
  DFF \round_reg_reg[739]  ( .D(out[739]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[739]) );
  DFF \round_reg_reg[740]  ( .D(out[740]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[740]) );
  DFF \round_reg_reg[741]  ( .D(out[741]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[741]) );
  DFF \round_reg_reg[742]  ( .D(out[742]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[742]) );
  DFF \round_reg_reg[743]  ( .D(out[743]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[743]) );
  DFF \round_reg_reg[744]  ( .D(out[744]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[744]) );
  DFF \round_reg_reg[745]  ( .D(out[745]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[745]) );
  DFF \round_reg_reg[746]  ( .D(out[746]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[746]) );
  DFF \round_reg_reg[747]  ( .D(out[747]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[747]) );
  DFF \round_reg_reg[748]  ( .D(out[748]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[748]) );
  DFF \round_reg_reg[749]  ( .D(out[749]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[749]) );
  DFF \round_reg_reg[750]  ( .D(out[750]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[750]) );
  DFF \round_reg_reg[751]  ( .D(out[751]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[751]) );
  DFF \round_reg_reg[752]  ( .D(out[752]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[752]) );
  DFF \round_reg_reg[753]  ( .D(out[753]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[753]) );
  DFF \round_reg_reg[754]  ( .D(out[754]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[754]) );
  DFF \round_reg_reg[755]  ( .D(out[755]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[755]) );
  DFF \round_reg_reg[756]  ( .D(out[756]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[756]) );
  DFF \round_reg_reg[757]  ( .D(out[757]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[757]) );
  DFF \round_reg_reg[758]  ( .D(out[758]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[758]) );
  DFF \round_reg_reg[759]  ( .D(out[759]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[759]) );
  DFF \round_reg_reg[760]  ( .D(out[760]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[760]) );
  DFF \round_reg_reg[761]  ( .D(out[761]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[761]) );
  DFF \round_reg_reg[762]  ( .D(out[762]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[762]) );
  DFF \round_reg_reg[763]  ( .D(out[763]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[763]) );
  DFF \round_reg_reg[764]  ( .D(out[764]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[764]) );
  DFF \round_reg_reg[765]  ( .D(out[765]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[765]) );
  DFF \round_reg_reg[766]  ( .D(out[766]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[766]) );
  DFF \round_reg_reg[767]  ( .D(out[767]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[767]) );
  DFF \round_reg_reg[768]  ( .D(out[768]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[768]) );
  DFF \round_reg_reg[769]  ( .D(out[769]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[769]) );
  DFF \round_reg_reg[770]  ( .D(out[770]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[770]) );
  DFF \round_reg_reg[771]  ( .D(out[771]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[771]) );
  DFF \round_reg_reg[772]  ( .D(out[772]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[772]) );
  DFF \round_reg_reg[773]  ( .D(out[773]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[773]) );
  DFF \round_reg_reg[774]  ( .D(out[774]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[774]) );
  DFF \round_reg_reg[775]  ( .D(out[775]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[775]) );
  DFF \round_reg_reg[776]  ( .D(out[776]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[776]) );
  DFF \round_reg_reg[777]  ( .D(out[777]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[777]) );
  DFF \round_reg_reg[778]  ( .D(out[778]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[778]) );
  DFF \round_reg_reg[779]  ( .D(out[779]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[779]) );
  DFF \round_reg_reg[780]  ( .D(out[780]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[780]) );
  DFF \round_reg_reg[781]  ( .D(out[781]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[781]) );
  DFF \round_reg_reg[782]  ( .D(out[782]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[782]) );
  DFF \round_reg_reg[783]  ( .D(out[783]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[783]) );
  DFF \round_reg_reg[784]  ( .D(out[784]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[784]) );
  DFF \round_reg_reg[785]  ( .D(out[785]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[785]) );
  DFF \round_reg_reg[786]  ( .D(out[786]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[786]) );
  DFF \round_reg_reg[787]  ( .D(out[787]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[787]) );
  DFF \round_reg_reg[788]  ( .D(out[788]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[788]) );
  DFF \round_reg_reg[789]  ( .D(out[789]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[789]) );
  DFF \round_reg_reg[790]  ( .D(out[790]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[790]) );
  DFF \round_reg_reg[791]  ( .D(out[791]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[791]) );
  DFF \round_reg_reg[792]  ( .D(out[792]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[792]) );
  DFF \round_reg_reg[793]  ( .D(out[793]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[793]) );
  DFF \round_reg_reg[794]  ( .D(out[794]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[794]) );
  DFF \round_reg_reg[795]  ( .D(out[795]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[795]) );
  DFF \round_reg_reg[796]  ( .D(out[796]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[796]) );
  DFF \round_reg_reg[797]  ( .D(out[797]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[797]) );
  DFF \round_reg_reg[798]  ( .D(out[798]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[798]) );
  DFF \round_reg_reg[799]  ( .D(out[799]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[799]) );
  DFF \round_reg_reg[800]  ( .D(out[800]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[800]) );
  DFF \round_reg_reg[801]  ( .D(out[801]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[801]) );
  DFF \round_reg_reg[802]  ( .D(out[802]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[802]) );
  DFF \round_reg_reg[803]  ( .D(out[803]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[803]) );
  DFF \round_reg_reg[804]  ( .D(out[804]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[804]) );
  DFF \round_reg_reg[805]  ( .D(out[805]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[805]) );
  DFF \round_reg_reg[806]  ( .D(out[806]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[806]) );
  DFF \round_reg_reg[807]  ( .D(out[807]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[807]) );
  DFF \round_reg_reg[808]  ( .D(out[808]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[808]) );
  DFF \round_reg_reg[809]  ( .D(out[809]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[809]) );
  DFF \round_reg_reg[810]  ( .D(out[810]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[810]) );
  DFF \round_reg_reg[811]  ( .D(out[811]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[811]) );
  DFF \round_reg_reg[812]  ( .D(out[812]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[812]) );
  DFF \round_reg_reg[813]  ( .D(out[813]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[813]) );
  DFF \round_reg_reg[814]  ( .D(out[814]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[814]) );
  DFF \round_reg_reg[815]  ( .D(out[815]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[815]) );
  DFF \round_reg_reg[816]  ( .D(out[816]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[816]) );
  DFF \round_reg_reg[817]  ( .D(out[817]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[817]) );
  DFF \round_reg_reg[818]  ( .D(out[818]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[818]) );
  DFF \round_reg_reg[819]  ( .D(out[819]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[819]) );
  DFF \round_reg_reg[820]  ( .D(out[820]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[820]) );
  DFF \round_reg_reg[821]  ( .D(out[821]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[821]) );
  DFF \round_reg_reg[822]  ( .D(out[822]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[822]) );
  DFF \round_reg_reg[823]  ( .D(out[823]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[823]) );
  DFF \round_reg_reg[824]  ( .D(out[824]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[824]) );
  DFF \round_reg_reg[825]  ( .D(out[825]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[825]) );
  DFF \round_reg_reg[826]  ( .D(out[826]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[826]) );
  DFF \round_reg_reg[827]  ( .D(out[827]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[827]) );
  DFF \round_reg_reg[828]  ( .D(out[828]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[828]) );
  DFF \round_reg_reg[829]  ( .D(out[829]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[829]) );
  DFF \round_reg_reg[830]  ( .D(out[830]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[830]) );
  DFF \round_reg_reg[831]  ( .D(out[831]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[831]) );
  DFF \round_reg_reg[832]  ( .D(out[832]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[832]) );
  DFF \round_reg_reg[833]  ( .D(out[833]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[833]) );
  DFF \round_reg_reg[834]  ( .D(out[834]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[834]) );
  DFF \round_reg_reg[835]  ( .D(out[835]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[835]) );
  DFF \round_reg_reg[836]  ( .D(out[836]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[836]) );
  DFF \round_reg_reg[837]  ( .D(out[837]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[837]) );
  DFF \round_reg_reg[838]  ( .D(out[838]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[838]) );
  DFF \round_reg_reg[839]  ( .D(out[839]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[839]) );
  DFF \round_reg_reg[840]  ( .D(out[840]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[840]) );
  DFF \round_reg_reg[841]  ( .D(out[841]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[841]) );
  DFF \round_reg_reg[842]  ( .D(out[842]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[842]) );
  DFF \round_reg_reg[843]  ( .D(out[843]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[843]) );
  DFF \round_reg_reg[844]  ( .D(out[844]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[844]) );
  DFF \round_reg_reg[845]  ( .D(out[845]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[845]) );
  DFF \round_reg_reg[846]  ( .D(out[846]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[846]) );
  DFF \round_reg_reg[847]  ( .D(out[847]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[847]) );
  DFF \round_reg_reg[848]  ( .D(out[848]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[848]) );
  DFF \round_reg_reg[849]  ( .D(out[849]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[849]) );
  DFF \round_reg_reg[850]  ( .D(out[850]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[850]) );
  DFF \round_reg_reg[851]  ( .D(out[851]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[851]) );
  DFF \round_reg_reg[852]  ( .D(out[852]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[852]) );
  DFF \round_reg_reg[853]  ( .D(out[853]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[853]) );
  DFF \round_reg_reg[854]  ( .D(out[854]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[854]) );
  DFF \round_reg_reg[855]  ( .D(out[855]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[855]) );
  DFF \round_reg_reg[856]  ( .D(out[856]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[856]) );
  DFF \round_reg_reg[857]  ( .D(out[857]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[857]) );
  DFF \round_reg_reg[858]  ( .D(out[858]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[858]) );
  DFF \round_reg_reg[859]  ( .D(out[859]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[859]) );
  DFF \round_reg_reg[860]  ( .D(out[860]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[860]) );
  DFF \round_reg_reg[861]  ( .D(out[861]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[861]) );
  DFF \round_reg_reg[862]  ( .D(out[862]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[862]) );
  DFF \round_reg_reg[863]  ( .D(out[863]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[863]) );
  DFF \round_reg_reg[864]  ( .D(out[864]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[864]) );
  DFF \round_reg_reg[865]  ( .D(out[865]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[865]) );
  DFF \round_reg_reg[866]  ( .D(out[866]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[866]) );
  DFF \round_reg_reg[867]  ( .D(out[867]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[867]) );
  DFF \round_reg_reg[868]  ( .D(out[868]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[868]) );
  DFF \round_reg_reg[869]  ( .D(out[869]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[869]) );
  DFF \round_reg_reg[870]  ( .D(out[870]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[870]) );
  DFF \round_reg_reg[871]  ( .D(out[871]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[871]) );
  DFF \round_reg_reg[872]  ( .D(out[872]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[872]) );
  DFF \round_reg_reg[873]  ( .D(out[873]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[873]) );
  DFF \round_reg_reg[874]  ( .D(out[874]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[874]) );
  DFF \round_reg_reg[875]  ( .D(out[875]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[875]) );
  DFF \round_reg_reg[876]  ( .D(out[876]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[876]) );
  DFF \round_reg_reg[877]  ( .D(out[877]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[877]) );
  DFF \round_reg_reg[878]  ( .D(out[878]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[878]) );
  DFF \round_reg_reg[879]  ( .D(out[879]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[879]) );
  DFF \round_reg_reg[880]  ( .D(out[880]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[880]) );
  DFF \round_reg_reg[881]  ( .D(out[881]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[881]) );
  DFF \round_reg_reg[882]  ( .D(out[882]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[882]) );
  DFF \round_reg_reg[883]  ( .D(out[883]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[883]) );
  DFF \round_reg_reg[884]  ( .D(out[884]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[884]) );
  DFF \round_reg_reg[885]  ( .D(out[885]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[885]) );
  DFF \round_reg_reg[886]  ( .D(out[886]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[886]) );
  DFF \round_reg_reg[887]  ( .D(out[887]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[887]) );
  DFF \round_reg_reg[888]  ( .D(out[888]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[888]) );
  DFF \round_reg_reg[889]  ( .D(out[889]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[889]) );
  DFF \round_reg_reg[890]  ( .D(out[890]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[890]) );
  DFF \round_reg_reg[891]  ( .D(out[891]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[891]) );
  DFF \round_reg_reg[892]  ( .D(out[892]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[892]) );
  DFF \round_reg_reg[893]  ( .D(out[893]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[893]) );
  DFF \round_reg_reg[894]  ( .D(out[894]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[894]) );
  DFF \round_reg_reg[895]  ( .D(out[895]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[895]) );
  DFF \round_reg_reg[896]  ( .D(out[896]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[896]) );
  DFF \round_reg_reg[897]  ( .D(out[897]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[897]) );
  DFF \round_reg_reg[898]  ( .D(out[898]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[898]) );
  DFF \round_reg_reg[899]  ( .D(out[899]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[899]) );
  DFF \round_reg_reg[900]  ( .D(out[900]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[900]) );
  DFF \round_reg_reg[901]  ( .D(out[901]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[901]) );
  DFF \round_reg_reg[902]  ( .D(out[902]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[902]) );
  DFF \round_reg_reg[903]  ( .D(out[903]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[903]) );
  DFF \round_reg_reg[904]  ( .D(out[904]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[904]) );
  DFF \round_reg_reg[905]  ( .D(out[905]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[905]) );
  DFF \round_reg_reg[906]  ( .D(out[906]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[906]) );
  DFF \round_reg_reg[907]  ( .D(out[907]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[907]) );
  DFF \round_reg_reg[908]  ( .D(out[908]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[908]) );
  DFF \round_reg_reg[909]  ( .D(out[909]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[909]) );
  DFF \round_reg_reg[910]  ( .D(out[910]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[910]) );
  DFF \round_reg_reg[911]  ( .D(out[911]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[911]) );
  DFF \round_reg_reg[912]  ( .D(out[912]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[912]) );
  DFF \round_reg_reg[913]  ( .D(out[913]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[913]) );
  DFF \round_reg_reg[914]  ( .D(out[914]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[914]) );
  DFF \round_reg_reg[915]  ( .D(out[915]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[915]) );
  DFF \round_reg_reg[916]  ( .D(out[916]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[916]) );
  DFF \round_reg_reg[917]  ( .D(out[917]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[917]) );
  DFF \round_reg_reg[918]  ( .D(out[918]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[918]) );
  DFF \round_reg_reg[919]  ( .D(out[919]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[919]) );
  DFF \round_reg_reg[920]  ( .D(out[920]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[920]) );
  DFF \round_reg_reg[921]  ( .D(out[921]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[921]) );
  DFF \round_reg_reg[922]  ( .D(out[922]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[922]) );
  DFF \round_reg_reg[923]  ( .D(out[923]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[923]) );
  DFF \round_reg_reg[924]  ( .D(out[924]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[924]) );
  DFF \round_reg_reg[925]  ( .D(out[925]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[925]) );
  DFF \round_reg_reg[926]  ( .D(out[926]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[926]) );
  DFF \round_reg_reg[927]  ( .D(out[927]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[927]) );
  DFF \round_reg_reg[928]  ( .D(out[928]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[928]) );
  DFF \round_reg_reg[929]  ( .D(out[929]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[929]) );
  DFF \round_reg_reg[930]  ( .D(out[930]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[930]) );
  DFF \round_reg_reg[931]  ( .D(out[931]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[931]) );
  DFF \round_reg_reg[932]  ( .D(out[932]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[932]) );
  DFF \round_reg_reg[933]  ( .D(out[933]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[933]) );
  DFF \round_reg_reg[934]  ( .D(out[934]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[934]) );
  DFF \round_reg_reg[935]  ( .D(out[935]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[935]) );
  DFF \round_reg_reg[936]  ( .D(out[936]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[936]) );
  DFF \round_reg_reg[937]  ( .D(out[937]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[937]) );
  DFF \round_reg_reg[938]  ( .D(out[938]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[938]) );
  DFF \round_reg_reg[939]  ( .D(out[939]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[939]) );
  DFF \round_reg_reg[940]  ( .D(out[940]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[940]) );
  DFF \round_reg_reg[941]  ( .D(out[941]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[941]) );
  DFF \round_reg_reg[942]  ( .D(out[942]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[942]) );
  DFF \round_reg_reg[943]  ( .D(out[943]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[943]) );
  DFF \round_reg_reg[944]  ( .D(out[944]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[944]) );
  DFF \round_reg_reg[945]  ( .D(out[945]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[945]) );
  DFF \round_reg_reg[946]  ( .D(out[946]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[946]) );
  DFF \round_reg_reg[947]  ( .D(out[947]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[947]) );
  DFF \round_reg_reg[948]  ( .D(out[948]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[948]) );
  DFF \round_reg_reg[949]  ( .D(out[949]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[949]) );
  DFF \round_reg_reg[950]  ( .D(out[950]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[950]) );
  DFF \round_reg_reg[951]  ( .D(out[951]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[951]) );
  DFF \round_reg_reg[952]  ( .D(out[952]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[952]) );
  DFF \round_reg_reg[953]  ( .D(out[953]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[953]) );
  DFF \round_reg_reg[954]  ( .D(out[954]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[954]) );
  DFF \round_reg_reg[955]  ( .D(out[955]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[955]) );
  DFF \round_reg_reg[956]  ( .D(out[956]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[956]) );
  DFF \round_reg_reg[957]  ( .D(out[957]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[957]) );
  DFF \round_reg_reg[958]  ( .D(out[958]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[958]) );
  DFF \round_reg_reg[959]  ( .D(out[959]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[959]) );
  DFF \round_reg_reg[960]  ( .D(out[960]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[960]) );
  DFF \round_reg_reg[961]  ( .D(out[961]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[961]) );
  DFF \round_reg_reg[962]  ( .D(out[962]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[962]) );
  DFF \round_reg_reg[963]  ( .D(out[963]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[963]) );
  DFF \round_reg_reg[964]  ( .D(out[964]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[964]) );
  DFF \round_reg_reg[965]  ( .D(out[965]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[965]) );
  DFF \round_reg_reg[966]  ( .D(out[966]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[966]) );
  DFF \round_reg_reg[967]  ( .D(out[967]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[967]) );
  DFF \round_reg_reg[968]  ( .D(out[968]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[968]) );
  DFF \round_reg_reg[969]  ( .D(out[969]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[969]) );
  DFF \round_reg_reg[970]  ( .D(out[970]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[970]) );
  DFF \round_reg_reg[971]  ( .D(out[971]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[971]) );
  DFF \round_reg_reg[972]  ( .D(out[972]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[972]) );
  DFF \round_reg_reg[973]  ( .D(out[973]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[973]) );
  DFF \round_reg_reg[974]  ( .D(out[974]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[974]) );
  DFF \round_reg_reg[975]  ( .D(out[975]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[975]) );
  DFF \round_reg_reg[976]  ( .D(out[976]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[976]) );
  DFF \round_reg_reg[977]  ( .D(out[977]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[977]) );
  DFF \round_reg_reg[978]  ( .D(out[978]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[978]) );
  DFF \round_reg_reg[979]  ( .D(out[979]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[979]) );
  DFF \round_reg_reg[980]  ( .D(out[980]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[980]) );
  DFF \round_reg_reg[981]  ( .D(out[981]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[981]) );
  DFF \round_reg_reg[982]  ( .D(out[982]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[982]) );
  DFF \round_reg_reg[983]  ( .D(out[983]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[983]) );
  DFF \round_reg_reg[984]  ( .D(out[984]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[984]) );
  DFF \round_reg_reg[985]  ( .D(out[985]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[985]) );
  DFF \round_reg_reg[986]  ( .D(out[986]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[986]) );
  DFF \round_reg_reg[987]  ( .D(out[987]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[987]) );
  DFF \round_reg_reg[988]  ( .D(out[988]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[988]) );
  DFF \round_reg_reg[989]  ( .D(out[989]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[989]) );
  DFF \round_reg_reg[990]  ( .D(out[990]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[990]) );
  DFF \round_reg_reg[991]  ( .D(out[991]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[991]) );
  DFF \round_reg_reg[992]  ( .D(out[992]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[992]) );
  DFF \round_reg_reg[993]  ( .D(out[993]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[993]) );
  DFF \round_reg_reg[994]  ( .D(out[994]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[994]) );
  DFF \round_reg_reg[995]  ( .D(out[995]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[995]) );
  DFF \round_reg_reg[996]  ( .D(out[996]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[996]) );
  DFF \round_reg_reg[997]  ( .D(out[997]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[997]) );
  DFF \round_reg_reg[998]  ( .D(out[998]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[998]) );
  DFF \round_reg_reg[999]  ( .D(out[999]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[999]) );
  DFF \round_reg_reg[1000]  ( .D(out[1000]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1000]) );
  DFF \round_reg_reg[1001]  ( .D(out[1001]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1001]) );
  DFF \round_reg_reg[1002]  ( .D(out[1002]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1002]) );
  DFF \round_reg_reg[1003]  ( .D(out[1003]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1003]) );
  DFF \round_reg_reg[1004]  ( .D(out[1004]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1004]) );
  DFF \round_reg_reg[1005]  ( .D(out[1005]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1005]) );
  DFF \round_reg_reg[1006]  ( .D(out[1006]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1006]) );
  DFF \round_reg_reg[1007]  ( .D(out[1007]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1007]) );
  DFF \round_reg_reg[1008]  ( .D(out[1008]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1008]) );
  DFF \round_reg_reg[1009]  ( .D(out[1009]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1009]) );
  DFF \round_reg_reg[1010]  ( .D(out[1010]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1010]) );
  DFF \round_reg_reg[1011]  ( .D(out[1011]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1011]) );
  DFF \round_reg_reg[1012]  ( .D(out[1012]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1012]) );
  DFF \round_reg_reg[1013]  ( .D(out[1013]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1013]) );
  DFF \round_reg_reg[1014]  ( .D(out[1014]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1014]) );
  DFF \round_reg_reg[1015]  ( .D(out[1015]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1015]) );
  DFF \round_reg_reg[1016]  ( .D(out[1016]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1016]) );
  DFF \round_reg_reg[1017]  ( .D(out[1017]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1017]) );
  DFF \round_reg_reg[1018]  ( .D(out[1018]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1018]) );
  DFF \round_reg_reg[1019]  ( .D(out[1019]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1019]) );
  DFF \round_reg_reg[1020]  ( .D(out[1020]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1020]) );
  DFF \round_reg_reg[1021]  ( .D(out[1021]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1021]) );
  DFF \round_reg_reg[1022]  ( .D(out[1022]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1022]) );
  DFF \round_reg_reg[1023]  ( .D(out[1023]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1023]) );
  DFF \round_reg_reg[1024]  ( .D(out[1024]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1024]) );
  DFF \round_reg_reg[1025]  ( .D(out[1025]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1025]) );
  DFF \round_reg_reg[1026]  ( .D(out[1026]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1026]) );
  DFF \round_reg_reg[1027]  ( .D(out[1027]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1027]) );
  DFF \round_reg_reg[1028]  ( .D(out[1028]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1028]) );
  DFF \round_reg_reg[1029]  ( .D(out[1029]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1029]) );
  DFF \round_reg_reg[1030]  ( .D(out[1030]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1030]) );
  DFF \round_reg_reg[1031]  ( .D(out[1031]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1031]) );
  DFF \round_reg_reg[1032]  ( .D(out[1032]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1032]) );
  DFF \round_reg_reg[1033]  ( .D(out[1033]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1033]) );
  DFF \round_reg_reg[1034]  ( .D(out[1034]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1034]) );
  DFF \round_reg_reg[1035]  ( .D(out[1035]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1035]) );
  DFF \round_reg_reg[1036]  ( .D(out[1036]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1036]) );
  DFF \round_reg_reg[1037]  ( .D(out[1037]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1037]) );
  DFF \round_reg_reg[1038]  ( .D(out[1038]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1038]) );
  DFF \round_reg_reg[1039]  ( .D(out[1039]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1039]) );
  DFF \round_reg_reg[1040]  ( .D(out[1040]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1040]) );
  DFF \round_reg_reg[1041]  ( .D(out[1041]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1041]) );
  DFF \round_reg_reg[1042]  ( .D(out[1042]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1042]) );
  DFF \round_reg_reg[1043]  ( .D(out[1043]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1043]) );
  DFF \round_reg_reg[1044]  ( .D(out[1044]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1044]) );
  DFF \round_reg_reg[1045]  ( .D(out[1045]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1045]) );
  DFF \round_reg_reg[1046]  ( .D(out[1046]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1046]) );
  DFF \round_reg_reg[1047]  ( .D(out[1047]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1047]) );
  DFF \round_reg_reg[1048]  ( .D(out[1048]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1048]) );
  DFF \round_reg_reg[1049]  ( .D(out[1049]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1049]) );
  DFF \round_reg_reg[1050]  ( .D(out[1050]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1050]) );
  DFF \round_reg_reg[1051]  ( .D(out[1051]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1051]) );
  DFF \round_reg_reg[1052]  ( .D(out[1052]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1052]) );
  DFF \round_reg_reg[1053]  ( .D(out[1053]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1053]) );
  DFF \round_reg_reg[1054]  ( .D(out[1054]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1054]) );
  DFF \round_reg_reg[1055]  ( .D(out[1055]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1055]) );
  DFF \round_reg_reg[1056]  ( .D(out[1056]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1056]) );
  DFF \round_reg_reg[1057]  ( .D(out[1057]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1057]) );
  DFF \round_reg_reg[1058]  ( .D(out[1058]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1058]) );
  DFF \round_reg_reg[1059]  ( .D(out[1059]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1059]) );
  DFF \round_reg_reg[1060]  ( .D(out[1060]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1060]) );
  DFF \round_reg_reg[1061]  ( .D(out[1061]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1061]) );
  DFF \round_reg_reg[1062]  ( .D(out[1062]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1062]) );
  DFF \round_reg_reg[1063]  ( .D(out[1063]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1063]) );
  DFF \round_reg_reg[1064]  ( .D(out[1064]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1064]) );
  DFF \round_reg_reg[1065]  ( .D(out[1065]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1065]) );
  DFF \round_reg_reg[1066]  ( .D(out[1066]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1066]) );
  DFF \round_reg_reg[1067]  ( .D(out[1067]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1067]) );
  DFF \round_reg_reg[1068]  ( .D(out[1068]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1068]) );
  DFF \round_reg_reg[1069]  ( .D(out[1069]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1069]) );
  DFF \round_reg_reg[1070]  ( .D(out[1070]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1070]) );
  DFF \round_reg_reg[1071]  ( .D(out[1071]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1071]) );
  DFF \round_reg_reg[1072]  ( .D(out[1072]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1072]) );
  DFF \round_reg_reg[1073]  ( .D(out[1073]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1073]) );
  DFF \round_reg_reg[1074]  ( .D(out[1074]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1074]) );
  DFF \round_reg_reg[1075]  ( .D(out[1075]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1075]) );
  DFF \round_reg_reg[1076]  ( .D(out[1076]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1076]) );
  DFF \round_reg_reg[1077]  ( .D(out[1077]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1077]) );
  DFF \round_reg_reg[1078]  ( .D(out[1078]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1078]) );
  DFF \round_reg_reg[1079]  ( .D(out[1079]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1079]) );
  DFF \round_reg_reg[1080]  ( .D(out[1080]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1080]) );
  DFF \round_reg_reg[1081]  ( .D(out[1081]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1081]) );
  DFF \round_reg_reg[1082]  ( .D(out[1082]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1082]) );
  DFF \round_reg_reg[1083]  ( .D(out[1083]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1083]) );
  DFF \round_reg_reg[1084]  ( .D(out[1084]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1084]) );
  DFF \round_reg_reg[1085]  ( .D(out[1085]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1085]) );
  DFF \round_reg_reg[1086]  ( .D(out[1086]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1086]) );
  DFF \round_reg_reg[1087]  ( .D(out[1087]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1087]) );
  DFF \round_reg_reg[1088]  ( .D(out[1088]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1088]) );
  DFF \round_reg_reg[1089]  ( .D(out[1089]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1089]) );
  DFF \round_reg_reg[1090]  ( .D(out[1090]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1090]) );
  DFF \round_reg_reg[1091]  ( .D(out[1091]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1091]) );
  DFF \round_reg_reg[1092]  ( .D(out[1092]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1092]) );
  DFF \round_reg_reg[1093]  ( .D(out[1093]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1093]) );
  DFF \round_reg_reg[1094]  ( .D(out[1094]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1094]) );
  DFF \round_reg_reg[1095]  ( .D(out[1095]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1095]) );
  DFF \round_reg_reg[1096]  ( .D(out[1096]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1096]) );
  DFF \round_reg_reg[1097]  ( .D(out[1097]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1097]) );
  DFF \round_reg_reg[1098]  ( .D(out[1098]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1098]) );
  DFF \round_reg_reg[1099]  ( .D(out[1099]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1099]) );
  DFF \round_reg_reg[1100]  ( .D(out[1100]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1100]) );
  DFF \round_reg_reg[1101]  ( .D(out[1101]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1101]) );
  DFF \round_reg_reg[1102]  ( .D(out[1102]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1102]) );
  DFF \round_reg_reg[1103]  ( .D(out[1103]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1103]) );
  DFF \round_reg_reg[1104]  ( .D(out[1104]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1104]) );
  DFF \round_reg_reg[1105]  ( .D(out[1105]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1105]) );
  DFF \round_reg_reg[1106]  ( .D(out[1106]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1106]) );
  DFF \round_reg_reg[1107]  ( .D(out[1107]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1107]) );
  DFF \round_reg_reg[1108]  ( .D(out[1108]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1108]) );
  DFF \round_reg_reg[1109]  ( .D(out[1109]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1109]) );
  DFF \round_reg_reg[1110]  ( .D(out[1110]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1110]) );
  DFF \round_reg_reg[1111]  ( .D(out[1111]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1111]) );
  DFF \round_reg_reg[1112]  ( .D(out[1112]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1112]) );
  DFF \round_reg_reg[1113]  ( .D(out[1113]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1113]) );
  DFF \round_reg_reg[1114]  ( .D(out[1114]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1114]) );
  DFF \round_reg_reg[1115]  ( .D(out[1115]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1115]) );
  DFF \round_reg_reg[1116]  ( .D(out[1116]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1116]) );
  DFF \round_reg_reg[1117]  ( .D(out[1117]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1117]) );
  DFF \round_reg_reg[1118]  ( .D(out[1118]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1118]) );
  DFF \round_reg_reg[1119]  ( .D(out[1119]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1119]) );
  DFF \round_reg_reg[1120]  ( .D(out[1120]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1120]) );
  DFF \round_reg_reg[1121]  ( .D(out[1121]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1121]) );
  DFF \round_reg_reg[1122]  ( .D(out[1122]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1122]) );
  DFF \round_reg_reg[1123]  ( .D(out[1123]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1123]) );
  DFF \round_reg_reg[1124]  ( .D(out[1124]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1124]) );
  DFF \round_reg_reg[1125]  ( .D(out[1125]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1125]) );
  DFF \round_reg_reg[1126]  ( .D(out[1126]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1126]) );
  DFF \round_reg_reg[1127]  ( .D(out[1127]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1127]) );
  DFF \round_reg_reg[1128]  ( .D(out[1128]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1128]) );
  DFF \round_reg_reg[1129]  ( .D(out[1129]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1129]) );
  DFF \round_reg_reg[1130]  ( .D(out[1130]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1130]) );
  DFF \round_reg_reg[1131]  ( .D(out[1131]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1131]) );
  DFF \round_reg_reg[1132]  ( .D(out[1132]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1132]) );
  DFF \round_reg_reg[1133]  ( .D(out[1133]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1133]) );
  DFF \round_reg_reg[1134]  ( .D(out[1134]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1134]) );
  DFF \round_reg_reg[1135]  ( .D(out[1135]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1135]) );
  DFF \round_reg_reg[1136]  ( .D(out[1136]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1136]) );
  DFF \round_reg_reg[1137]  ( .D(out[1137]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1137]) );
  DFF \round_reg_reg[1138]  ( .D(out[1138]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1138]) );
  DFF \round_reg_reg[1139]  ( .D(out[1139]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1139]) );
  DFF \round_reg_reg[1140]  ( .D(out[1140]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1140]) );
  DFF \round_reg_reg[1141]  ( .D(out[1141]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1141]) );
  DFF \round_reg_reg[1142]  ( .D(out[1142]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1142]) );
  DFF \round_reg_reg[1143]  ( .D(out[1143]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1143]) );
  DFF \round_reg_reg[1144]  ( .D(out[1144]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1144]) );
  DFF \round_reg_reg[1145]  ( .D(out[1145]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1145]) );
  DFF \round_reg_reg[1146]  ( .D(out[1146]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1146]) );
  DFF \round_reg_reg[1147]  ( .D(out[1147]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1147]) );
  DFF \round_reg_reg[1148]  ( .D(out[1148]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1148]) );
  DFF \round_reg_reg[1149]  ( .D(out[1149]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1149]) );
  DFF \round_reg_reg[1150]  ( .D(out[1150]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1150]) );
  DFF \round_reg_reg[1151]  ( .D(out[1151]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1151]) );
  DFF \round_reg_reg[1152]  ( .D(out[1152]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1152]) );
  DFF \round_reg_reg[1153]  ( .D(out[1153]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1153]) );
  DFF \round_reg_reg[1154]  ( .D(out[1154]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1154]) );
  DFF \round_reg_reg[1155]  ( .D(out[1155]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1155]) );
  DFF \round_reg_reg[1156]  ( .D(out[1156]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1156]) );
  DFF \round_reg_reg[1157]  ( .D(out[1157]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1157]) );
  DFF \round_reg_reg[1158]  ( .D(out[1158]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1158]) );
  DFF \round_reg_reg[1159]  ( .D(out[1159]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1159]) );
  DFF \round_reg_reg[1160]  ( .D(out[1160]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1160]) );
  DFF \round_reg_reg[1161]  ( .D(out[1161]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1161]) );
  DFF \round_reg_reg[1162]  ( .D(out[1162]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1162]) );
  DFF \round_reg_reg[1163]  ( .D(out[1163]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1163]) );
  DFF \round_reg_reg[1164]  ( .D(out[1164]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1164]) );
  DFF \round_reg_reg[1165]  ( .D(out[1165]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1165]) );
  DFF \round_reg_reg[1166]  ( .D(out[1166]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1166]) );
  DFF \round_reg_reg[1167]  ( .D(out[1167]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1167]) );
  DFF \round_reg_reg[1168]  ( .D(out[1168]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1168]) );
  DFF \round_reg_reg[1169]  ( .D(out[1169]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1169]) );
  DFF \round_reg_reg[1170]  ( .D(out[1170]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1170]) );
  DFF \round_reg_reg[1171]  ( .D(out[1171]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1171]) );
  DFF \round_reg_reg[1172]  ( .D(out[1172]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1172]) );
  DFF \round_reg_reg[1173]  ( .D(out[1173]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1173]) );
  DFF \round_reg_reg[1174]  ( .D(out[1174]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1174]) );
  DFF \round_reg_reg[1175]  ( .D(out[1175]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1175]) );
  DFF \round_reg_reg[1176]  ( .D(out[1176]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1176]) );
  DFF \round_reg_reg[1177]  ( .D(out[1177]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1177]) );
  DFF \round_reg_reg[1178]  ( .D(out[1178]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1178]) );
  DFF \round_reg_reg[1179]  ( .D(out[1179]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1179]) );
  DFF \round_reg_reg[1180]  ( .D(out[1180]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1180]) );
  DFF \round_reg_reg[1181]  ( .D(out[1181]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1181]) );
  DFF \round_reg_reg[1182]  ( .D(out[1182]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1182]) );
  DFF \round_reg_reg[1183]  ( .D(out[1183]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1183]) );
  DFF \round_reg_reg[1184]  ( .D(out[1184]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1184]) );
  DFF \round_reg_reg[1185]  ( .D(out[1185]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1185]) );
  DFF \round_reg_reg[1186]  ( .D(out[1186]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1186]) );
  DFF \round_reg_reg[1187]  ( .D(out[1187]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1187]) );
  DFF \round_reg_reg[1188]  ( .D(out[1188]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1188]) );
  DFF \round_reg_reg[1189]  ( .D(out[1189]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1189]) );
  DFF \round_reg_reg[1190]  ( .D(out[1190]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1190]) );
  DFF \round_reg_reg[1191]  ( .D(out[1191]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1191]) );
  DFF \round_reg_reg[1192]  ( .D(out[1192]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1192]) );
  DFF \round_reg_reg[1193]  ( .D(out[1193]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1193]) );
  DFF \round_reg_reg[1194]  ( .D(out[1194]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1194]) );
  DFF \round_reg_reg[1195]  ( .D(out[1195]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1195]) );
  DFF \round_reg_reg[1196]  ( .D(out[1196]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1196]) );
  DFF \round_reg_reg[1197]  ( .D(out[1197]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1197]) );
  DFF \round_reg_reg[1198]  ( .D(out[1198]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1198]) );
  DFF \round_reg_reg[1199]  ( .D(out[1199]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1199]) );
  DFF \round_reg_reg[1200]  ( .D(out[1200]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1200]) );
  DFF \round_reg_reg[1201]  ( .D(out[1201]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1201]) );
  DFF \round_reg_reg[1202]  ( .D(out[1202]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1202]) );
  DFF \round_reg_reg[1203]  ( .D(out[1203]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1203]) );
  DFF \round_reg_reg[1204]  ( .D(out[1204]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1204]) );
  DFF \round_reg_reg[1205]  ( .D(out[1205]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1205]) );
  DFF \round_reg_reg[1206]  ( .D(out[1206]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1206]) );
  DFF \round_reg_reg[1207]  ( .D(out[1207]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1207]) );
  DFF \round_reg_reg[1208]  ( .D(out[1208]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1208]) );
  DFF \round_reg_reg[1209]  ( .D(out[1209]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1209]) );
  DFF \round_reg_reg[1210]  ( .D(out[1210]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1210]) );
  DFF \round_reg_reg[1211]  ( .D(out[1211]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1211]) );
  DFF \round_reg_reg[1212]  ( .D(out[1212]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1212]) );
  DFF \round_reg_reg[1213]  ( .D(out[1213]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1213]) );
  DFF \round_reg_reg[1214]  ( .D(out[1214]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1214]) );
  DFF \round_reg_reg[1215]  ( .D(out[1215]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1215]) );
  DFF \round_reg_reg[1216]  ( .D(out[1216]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1216]) );
  DFF \round_reg_reg[1217]  ( .D(out[1217]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1217]) );
  DFF \round_reg_reg[1218]  ( .D(out[1218]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1218]) );
  DFF \round_reg_reg[1219]  ( .D(out[1219]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1219]) );
  DFF \round_reg_reg[1220]  ( .D(out[1220]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1220]) );
  DFF \round_reg_reg[1221]  ( .D(out[1221]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1221]) );
  DFF \round_reg_reg[1222]  ( .D(out[1222]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1222]) );
  DFF \round_reg_reg[1223]  ( .D(out[1223]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1223]) );
  DFF \round_reg_reg[1224]  ( .D(out[1224]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1224]) );
  DFF \round_reg_reg[1225]  ( .D(out[1225]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1225]) );
  DFF \round_reg_reg[1226]  ( .D(out[1226]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1226]) );
  DFF \round_reg_reg[1227]  ( .D(out[1227]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1227]) );
  DFF \round_reg_reg[1228]  ( .D(out[1228]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1228]) );
  DFF \round_reg_reg[1229]  ( .D(out[1229]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1229]) );
  DFF \round_reg_reg[1230]  ( .D(out[1230]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1230]) );
  DFF \round_reg_reg[1231]  ( .D(out[1231]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1231]) );
  DFF \round_reg_reg[1232]  ( .D(out[1232]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1232]) );
  DFF \round_reg_reg[1233]  ( .D(out[1233]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1233]) );
  DFF \round_reg_reg[1234]  ( .D(out[1234]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1234]) );
  DFF \round_reg_reg[1235]  ( .D(out[1235]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1235]) );
  DFF \round_reg_reg[1236]  ( .D(out[1236]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1236]) );
  DFF \round_reg_reg[1237]  ( .D(out[1237]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1237]) );
  DFF \round_reg_reg[1238]  ( .D(out[1238]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1238]) );
  DFF \round_reg_reg[1239]  ( .D(out[1239]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1239]) );
  DFF \round_reg_reg[1240]  ( .D(out[1240]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1240]) );
  DFF \round_reg_reg[1241]  ( .D(out[1241]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1241]) );
  DFF \round_reg_reg[1242]  ( .D(out[1242]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1242]) );
  DFF \round_reg_reg[1243]  ( .D(out[1243]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1243]) );
  DFF \round_reg_reg[1244]  ( .D(out[1244]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1244]) );
  DFF \round_reg_reg[1245]  ( .D(out[1245]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1245]) );
  DFF \round_reg_reg[1246]  ( .D(out[1246]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1246]) );
  DFF \round_reg_reg[1247]  ( .D(out[1247]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1247]) );
  DFF \round_reg_reg[1248]  ( .D(out[1248]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1248]) );
  DFF \round_reg_reg[1249]  ( .D(out[1249]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1249]) );
  DFF \round_reg_reg[1250]  ( .D(out[1250]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1250]) );
  DFF \round_reg_reg[1251]  ( .D(out[1251]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1251]) );
  DFF \round_reg_reg[1252]  ( .D(out[1252]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1252]) );
  DFF \round_reg_reg[1253]  ( .D(out[1253]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1253]) );
  DFF \round_reg_reg[1254]  ( .D(out[1254]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1254]) );
  DFF \round_reg_reg[1255]  ( .D(out[1255]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1255]) );
  DFF \round_reg_reg[1256]  ( .D(out[1256]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1256]) );
  DFF \round_reg_reg[1257]  ( .D(out[1257]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1257]) );
  DFF \round_reg_reg[1258]  ( .D(out[1258]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1258]) );
  DFF \round_reg_reg[1259]  ( .D(out[1259]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1259]) );
  DFF \round_reg_reg[1260]  ( .D(out[1260]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1260]) );
  DFF \round_reg_reg[1261]  ( .D(out[1261]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1261]) );
  DFF \round_reg_reg[1262]  ( .D(out[1262]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1262]) );
  DFF \round_reg_reg[1263]  ( .D(out[1263]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1263]) );
  DFF \round_reg_reg[1264]  ( .D(out[1264]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1264]) );
  DFF \round_reg_reg[1265]  ( .D(out[1265]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1265]) );
  DFF \round_reg_reg[1266]  ( .D(out[1266]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1266]) );
  DFF \round_reg_reg[1267]  ( .D(out[1267]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1267]) );
  DFF \round_reg_reg[1268]  ( .D(out[1268]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1268]) );
  DFF \round_reg_reg[1269]  ( .D(out[1269]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1269]) );
  DFF \round_reg_reg[1270]  ( .D(out[1270]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1270]) );
  DFF \round_reg_reg[1271]  ( .D(out[1271]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1271]) );
  DFF \round_reg_reg[1272]  ( .D(out[1272]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1272]) );
  DFF \round_reg_reg[1273]  ( .D(out[1273]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1273]) );
  DFF \round_reg_reg[1274]  ( .D(out[1274]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1274]) );
  DFF \round_reg_reg[1275]  ( .D(out[1275]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1275]) );
  DFF \round_reg_reg[1276]  ( .D(out[1276]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1276]) );
  DFF \round_reg_reg[1277]  ( .D(out[1277]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1277]) );
  DFF \round_reg_reg[1278]  ( .D(out[1278]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1278]) );
  DFF \round_reg_reg[1279]  ( .D(out[1279]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1279]) );
  DFF \round_reg_reg[1280]  ( .D(out[1280]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1280]) );
  DFF \round_reg_reg[1281]  ( .D(out[1281]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1281]) );
  DFF \round_reg_reg[1282]  ( .D(out[1282]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1282]) );
  DFF \round_reg_reg[1283]  ( .D(out[1283]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1283]) );
  DFF \round_reg_reg[1284]  ( .D(out[1284]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1284]) );
  DFF \round_reg_reg[1285]  ( .D(out[1285]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1285]) );
  DFF \round_reg_reg[1286]  ( .D(out[1286]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1286]) );
  DFF \round_reg_reg[1287]  ( .D(out[1287]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1287]) );
  DFF \round_reg_reg[1288]  ( .D(out[1288]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1288]) );
  DFF \round_reg_reg[1289]  ( .D(out[1289]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1289]) );
  DFF \round_reg_reg[1290]  ( .D(out[1290]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1290]) );
  DFF \round_reg_reg[1291]  ( .D(out[1291]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1291]) );
  DFF \round_reg_reg[1292]  ( .D(out[1292]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1292]) );
  DFF \round_reg_reg[1293]  ( .D(out[1293]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1293]) );
  DFF \round_reg_reg[1294]  ( .D(out[1294]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1294]) );
  DFF \round_reg_reg[1295]  ( .D(out[1295]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1295]) );
  DFF \round_reg_reg[1296]  ( .D(out[1296]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1296]) );
  DFF \round_reg_reg[1297]  ( .D(out[1297]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1297]) );
  DFF \round_reg_reg[1298]  ( .D(out[1298]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1298]) );
  DFF \round_reg_reg[1299]  ( .D(out[1299]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1299]) );
  DFF \round_reg_reg[1300]  ( .D(out[1300]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1300]) );
  DFF \round_reg_reg[1301]  ( .D(out[1301]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1301]) );
  DFF \round_reg_reg[1302]  ( .D(out[1302]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1302]) );
  DFF \round_reg_reg[1303]  ( .D(out[1303]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1303]) );
  DFF \round_reg_reg[1304]  ( .D(out[1304]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1304]) );
  DFF \round_reg_reg[1305]  ( .D(out[1305]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1305]) );
  DFF \round_reg_reg[1306]  ( .D(out[1306]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1306]) );
  DFF \round_reg_reg[1307]  ( .D(out[1307]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1307]) );
  DFF \round_reg_reg[1308]  ( .D(out[1308]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1308]) );
  DFF \round_reg_reg[1309]  ( .D(out[1309]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1309]) );
  DFF \round_reg_reg[1310]  ( .D(out[1310]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1310]) );
  DFF \round_reg_reg[1311]  ( .D(out[1311]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1311]) );
  DFF \round_reg_reg[1312]  ( .D(out[1312]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1312]) );
  DFF \round_reg_reg[1313]  ( .D(out[1313]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1313]) );
  DFF \round_reg_reg[1314]  ( .D(out[1314]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1314]) );
  DFF \round_reg_reg[1315]  ( .D(out[1315]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1315]) );
  DFF \round_reg_reg[1316]  ( .D(out[1316]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1316]) );
  DFF \round_reg_reg[1317]  ( .D(out[1317]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1317]) );
  DFF \round_reg_reg[1318]  ( .D(out[1318]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1318]) );
  DFF \round_reg_reg[1319]  ( .D(out[1319]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1319]) );
  DFF \round_reg_reg[1320]  ( .D(out[1320]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1320]) );
  DFF \round_reg_reg[1321]  ( .D(out[1321]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1321]) );
  DFF \round_reg_reg[1322]  ( .D(out[1322]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1322]) );
  DFF \round_reg_reg[1323]  ( .D(out[1323]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1323]) );
  DFF \round_reg_reg[1324]  ( .D(out[1324]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1324]) );
  DFF \round_reg_reg[1325]  ( .D(out[1325]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1325]) );
  DFF \round_reg_reg[1326]  ( .D(out[1326]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1326]) );
  DFF \round_reg_reg[1327]  ( .D(out[1327]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1327]) );
  DFF \round_reg_reg[1328]  ( .D(out[1328]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1328]) );
  DFF \round_reg_reg[1329]  ( .D(out[1329]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1329]) );
  DFF \round_reg_reg[1330]  ( .D(out[1330]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1330]) );
  DFF \round_reg_reg[1331]  ( .D(out[1331]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1331]) );
  DFF \round_reg_reg[1332]  ( .D(out[1332]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1332]) );
  DFF \round_reg_reg[1333]  ( .D(out[1333]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1333]) );
  DFF \round_reg_reg[1334]  ( .D(out[1334]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1334]) );
  DFF \round_reg_reg[1335]  ( .D(out[1335]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1335]) );
  DFF \round_reg_reg[1336]  ( .D(out[1336]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1336]) );
  DFF \round_reg_reg[1337]  ( .D(out[1337]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1337]) );
  DFF \round_reg_reg[1338]  ( .D(out[1338]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1338]) );
  DFF \round_reg_reg[1339]  ( .D(out[1339]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1339]) );
  DFF \round_reg_reg[1340]  ( .D(out[1340]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1340]) );
  DFF \round_reg_reg[1341]  ( .D(out[1341]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1341]) );
  DFF \round_reg_reg[1342]  ( .D(out[1342]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1342]) );
  DFF \round_reg_reg[1343]  ( .D(out[1343]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1343]) );
  DFF \round_reg_reg[1344]  ( .D(out[1344]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1344]) );
  DFF \round_reg_reg[1345]  ( .D(out[1345]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1345]) );
  DFF \round_reg_reg[1346]  ( .D(out[1346]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1346]) );
  DFF \round_reg_reg[1347]  ( .D(out[1347]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1347]) );
  DFF \round_reg_reg[1348]  ( .D(out[1348]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1348]) );
  DFF \round_reg_reg[1349]  ( .D(out[1349]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1349]) );
  DFF \round_reg_reg[1350]  ( .D(out[1350]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1350]) );
  DFF \round_reg_reg[1351]  ( .D(out[1351]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1351]) );
  DFF \round_reg_reg[1352]  ( .D(out[1352]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1352]) );
  DFF \round_reg_reg[1353]  ( .D(out[1353]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1353]) );
  DFF \round_reg_reg[1354]  ( .D(out[1354]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1354]) );
  DFF \round_reg_reg[1355]  ( .D(out[1355]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1355]) );
  DFF \round_reg_reg[1356]  ( .D(out[1356]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1356]) );
  DFF \round_reg_reg[1357]  ( .D(out[1357]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1357]) );
  DFF \round_reg_reg[1358]  ( .D(out[1358]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1358]) );
  DFF \round_reg_reg[1359]  ( .D(out[1359]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1359]) );
  DFF \round_reg_reg[1360]  ( .D(out[1360]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1360]) );
  DFF \round_reg_reg[1361]  ( .D(out[1361]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1361]) );
  DFF \round_reg_reg[1362]  ( .D(out[1362]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1362]) );
  DFF \round_reg_reg[1363]  ( .D(out[1363]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1363]) );
  DFF \round_reg_reg[1364]  ( .D(out[1364]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1364]) );
  DFF \round_reg_reg[1365]  ( .D(out[1365]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1365]) );
  DFF \round_reg_reg[1366]  ( .D(out[1366]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1366]) );
  DFF \round_reg_reg[1367]  ( .D(out[1367]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1367]) );
  DFF \round_reg_reg[1368]  ( .D(out[1368]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1368]) );
  DFF \round_reg_reg[1369]  ( .D(out[1369]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1369]) );
  DFF \round_reg_reg[1370]  ( .D(out[1370]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1370]) );
  DFF \round_reg_reg[1371]  ( .D(out[1371]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1371]) );
  DFF \round_reg_reg[1372]  ( .D(out[1372]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1372]) );
  DFF \round_reg_reg[1373]  ( .D(out[1373]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1373]) );
  DFF \round_reg_reg[1374]  ( .D(out[1374]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1374]) );
  DFF \round_reg_reg[1375]  ( .D(out[1375]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1375]) );
  DFF \round_reg_reg[1376]  ( .D(out[1376]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1376]) );
  DFF \round_reg_reg[1377]  ( .D(out[1377]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1377]) );
  DFF \round_reg_reg[1378]  ( .D(out[1378]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1378]) );
  DFF \round_reg_reg[1379]  ( .D(out[1379]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1379]) );
  DFF \round_reg_reg[1380]  ( .D(out[1380]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1380]) );
  DFF \round_reg_reg[1381]  ( .D(out[1381]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1381]) );
  DFF \round_reg_reg[1382]  ( .D(out[1382]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1382]) );
  DFF \round_reg_reg[1383]  ( .D(out[1383]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1383]) );
  DFF \round_reg_reg[1384]  ( .D(out[1384]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1384]) );
  DFF \round_reg_reg[1385]  ( .D(out[1385]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1385]) );
  DFF \round_reg_reg[1386]  ( .D(out[1386]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1386]) );
  DFF \round_reg_reg[1387]  ( .D(out[1387]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1387]) );
  DFF \round_reg_reg[1388]  ( .D(out[1388]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1388]) );
  DFF \round_reg_reg[1389]  ( .D(out[1389]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1389]) );
  DFF \round_reg_reg[1390]  ( .D(out[1390]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1390]) );
  DFF \round_reg_reg[1391]  ( .D(out[1391]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1391]) );
  DFF \round_reg_reg[1392]  ( .D(out[1392]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1392]) );
  DFF \round_reg_reg[1393]  ( .D(out[1393]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1393]) );
  DFF \round_reg_reg[1394]  ( .D(out[1394]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1394]) );
  DFF \round_reg_reg[1395]  ( .D(out[1395]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1395]) );
  DFF \round_reg_reg[1396]  ( .D(out[1396]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1396]) );
  DFF \round_reg_reg[1397]  ( .D(out[1397]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1397]) );
  DFF \round_reg_reg[1398]  ( .D(out[1398]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1398]) );
  DFF \round_reg_reg[1399]  ( .D(out[1399]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1399]) );
  DFF \round_reg_reg[1400]  ( .D(out[1400]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1400]) );
  DFF \round_reg_reg[1401]  ( .D(out[1401]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1401]) );
  DFF \round_reg_reg[1402]  ( .D(out[1402]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1402]) );
  DFF \round_reg_reg[1403]  ( .D(out[1403]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1403]) );
  DFF \round_reg_reg[1404]  ( .D(out[1404]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1404]) );
  DFF \round_reg_reg[1405]  ( .D(out[1405]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1405]) );
  DFF \round_reg_reg[1406]  ( .D(out[1406]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1406]) );
  DFF \round_reg_reg[1407]  ( .D(out[1407]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1407]) );
  DFF \round_reg_reg[1408]  ( .D(out[1408]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1408]) );
  DFF \round_reg_reg[1409]  ( .D(out[1409]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1409]) );
  DFF \round_reg_reg[1410]  ( .D(out[1410]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1410]) );
  DFF \round_reg_reg[1411]  ( .D(out[1411]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1411]) );
  DFF \round_reg_reg[1412]  ( .D(out[1412]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1412]) );
  DFF \round_reg_reg[1413]  ( .D(out[1413]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1413]) );
  DFF \round_reg_reg[1414]  ( .D(out[1414]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1414]) );
  DFF \round_reg_reg[1415]  ( .D(out[1415]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1415]) );
  DFF \round_reg_reg[1416]  ( .D(out[1416]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1416]) );
  DFF \round_reg_reg[1417]  ( .D(out[1417]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1417]) );
  DFF \round_reg_reg[1418]  ( .D(out[1418]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1418]) );
  DFF \round_reg_reg[1419]  ( .D(out[1419]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1419]) );
  DFF \round_reg_reg[1420]  ( .D(out[1420]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1420]) );
  DFF \round_reg_reg[1421]  ( .D(out[1421]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1421]) );
  DFF \round_reg_reg[1422]  ( .D(out[1422]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1422]) );
  DFF \round_reg_reg[1423]  ( .D(out[1423]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1423]) );
  DFF \round_reg_reg[1424]  ( .D(out[1424]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1424]) );
  DFF \round_reg_reg[1425]  ( .D(out[1425]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1425]) );
  DFF \round_reg_reg[1426]  ( .D(out[1426]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1426]) );
  DFF \round_reg_reg[1427]  ( .D(out[1427]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1427]) );
  DFF \round_reg_reg[1428]  ( .D(out[1428]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1428]) );
  DFF \round_reg_reg[1429]  ( .D(out[1429]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1429]) );
  DFF \round_reg_reg[1430]  ( .D(out[1430]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1430]) );
  DFF \round_reg_reg[1431]  ( .D(out[1431]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1431]) );
  DFF \round_reg_reg[1432]  ( .D(out[1432]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1432]) );
  DFF \round_reg_reg[1433]  ( .D(out[1433]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1433]) );
  DFF \round_reg_reg[1434]  ( .D(out[1434]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1434]) );
  DFF \round_reg_reg[1435]  ( .D(out[1435]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1435]) );
  DFF \round_reg_reg[1436]  ( .D(out[1436]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1436]) );
  DFF \round_reg_reg[1437]  ( .D(out[1437]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1437]) );
  DFF \round_reg_reg[1438]  ( .D(out[1438]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1438]) );
  DFF \round_reg_reg[1439]  ( .D(out[1439]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1439]) );
  DFF \round_reg_reg[1440]  ( .D(out[1440]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1440]) );
  DFF \round_reg_reg[1441]  ( .D(out[1441]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1441]) );
  DFF \round_reg_reg[1442]  ( .D(out[1442]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1442]) );
  DFF \round_reg_reg[1443]  ( .D(out[1443]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1443]) );
  DFF \round_reg_reg[1444]  ( .D(out[1444]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1444]) );
  DFF \round_reg_reg[1445]  ( .D(out[1445]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1445]) );
  DFF \round_reg_reg[1446]  ( .D(out[1446]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1446]) );
  DFF \round_reg_reg[1447]  ( .D(out[1447]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1447]) );
  DFF \round_reg_reg[1448]  ( .D(out[1448]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1448]) );
  DFF \round_reg_reg[1449]  ( .D(out[1449]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1449]) );
  DFF \round_reg_reg[1450]  ( .D(out[1450]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1450]) );
  DFF \round_reg_reg[1451]  ( .D(out[1451]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1451]) );
  DFF \round_reg_reg[1452]  ( .D(out[1452]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1452]) );
  DFF \round_reg_reg[1453]  ( .D(out[1453]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1453]) );
  DFF \round_reg_reg[1454]  ( .D(out[1454]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1454]) );
  DFF \round_reg_reg[1455]  ( .D(out[1455]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1455]) );
  DFF \round_reg_reg[1456]  ( .D(out[1456]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1456]) );
  DFF \round_reg_reg[1457]  ( .D(out[1457]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1457]) );
  DFF \round_reg_reg[1458]  ( .D(out[1458]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1458]) );
  DFF \round_reg_reg[1459]  ( .D(out[1459]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1459]) );
  DFF \round_reg_reg[1460]  ( .D(out[1460]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1460]) );
  DFF \round_reg_reg[1461]  ( .D(out[1461]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1461]) );
  DFF \round_reg_reg[1462]  ( .D(out[1462]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1462]) );
  DFF \round_reg_reg[1463]  ( .D(out[1463]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1463]) );
  DFF \round_reg_reg[1464]  ( .D(out[1464]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1464]) );
  DFF \round_reg_reg[1465]  ( .D(out[1465]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1465]) );
  DFF \round_reg_reg[1466]  ( .D(out[1466]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1466]) );
  DFF \round_reg_reg[1467]  ( .D(out[1467]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1467]) );
  DFF \round_reg_reg[1468]  ( .D(out[1468]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1468]) );
  DFF \round_reg_reg[1469]  ( .D(out[1469]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1469]) );
  DFF \round_reg_reg[1470]  ( .D(out[1470]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1470]) );
  DFF \round_reg_reg[1471]  ( .D(out[1471]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1471]) );
  DFF \round_reg_reg[1472]  ( .D(out[1472]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1472]) );
  DFF \round_reg_reg[1473]  ( .D(out[1473]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1473]) );
  DFF \round_reg_reg[1474]  ( .D(out[1474]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1474]) );
  DFF \round_reg_reg[1475]  ( .D(out[1475]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1475]) );
  DFF \round_reg_reg[1476]  ( .D(out[1476]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1476]) );
  DFF \round_reg_reg[1477]  ( .D(out[1477]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1477]) );
  DFF \round_reg_reg[1478]  ( .D(out[1478]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1478]) );
  DFF \round_reg_reg[1479]  ( .D(out[1479]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1479]) );
  DFF \round_reg_reg[1480]  ( .D(out[1480]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1480]) );
  DFF \round_reg_reg[1481]  ( .D(out[1481]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1481]) );
  DFF \round_reg_reg[1482]  ( .D(out[1482]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1482]) );
  DFF \round_reg_reg[1483]  ( .D(out[1483]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1483]) );
  DFF \round_reg_reg[1484]  ( .D(out[1484]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1484]) );
  DFF \round_reg_reg[1485]  ( .D(out[1485]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1485]) );
  DFF \round_reg_reg[1486]  ( .D(out[1486]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1486]) );
  DFF \round_reg_reg[1487]  ( .D(out[1487]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1487]) );
  DFF \round_reg_reg[1488]  ( .D(out[1488]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1488]) );
  DFF \round_reg_reg[1489]  ( .D(out[1489]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1489]) );
  DFF \round_reg_reg[1490]  ( .D(out[1490]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1490]) );
  DFF \round_reg_reg[1491]  ( .D(out[1491]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1491]) );
  DFF \round_reg_reg[1492]  ( .D(out[1492]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1492]) );
  DFF \round_reg_reg[1493]  ( .D(out[1493]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1493]) );
  DFF \round_reg_reg[1494]  ( .D(out[1494]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1494]) );
  DFF \round_reg_reg[1495]  ( .D(out[1495]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1495]) );
  DFF \round_reg_reg[1496]  ( .D(out[1496]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1496]) );
  DFF \round_reg_reg[1497]  ( .D(out[1497]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1497]) );
  DFF \round_reg_reg[1498]  ( .D(out[1498]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1498]) );
  DFF \round_reg_reg[1499]  ( .D(out[1499]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1499]) );
  DFF \round_reg_reg[1500]  ( .D(out[1500]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1500]) );
  DFF \round_reg_reg[1501]  ( .D(out[1501]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1501]) );
  DFF \round_reg_reg[1502]  ( .D(out[1502]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1502]) );
  DFF \round_reg_reg[1503]  ( .D(out[1503]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1503]) );
  DFF \round_reg_reg[1504]  ( .D(out[1504]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1504]) );
  DFF \round_reg_reg[1505]  ( .D(out[1505]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1505]) );
  DFF \round_reg_reg[1506]  ( .D(out[1506]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1506]) );
  DFF \round_reg_reg[1507]  ( .D(out[1507]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1507]) );
  DFF \round_reg_reg[1508]  ( .D(out[1508]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1508]) );
  DFF \round_reg_reg[1509]  ( .D(out[1509]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1509]) );
  DFF \round_reg_reg[1510]  ( .D(out[1510]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1510]) );
  DFF \round_reg_reg[1511]  ( .D(out[1511]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1511]) );
  DFF \round_reg_reg[1512]  ( .D(out[1512]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1512]) );
  DFF \round_reg_reg[1513]  ( .D(out[1513]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1513]) );
  DFF \round_reg_reg[1514]  ( .D(out[1514]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1514]) );
  DFF \round_reg_reg[1515]  ( .D(out[1515]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1515]) );
  DFF \round_reg_reg[1516]  ( .D(out[1516]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1516]) );
  DFF \round_reg_reg[1517]  ( .D(out[1517]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1517]) );
  DFF \round_reg_reg[1518]  ( .D(out[1518]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1518]) );
  DFF \round_reg_reg[1519]  ( .D(out[1519]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1519]) );
  DFF \round_reg_reg[1520]  ( .D(out[1520]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1520]) );
  DFF \round_reg_reg[1521]  ( .D(out[1521]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1521]) );
  DFF \round_reg_reg[1522]  ( .D(out[1522]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1522]) );
  DFF \round_reg_reg[1523]  ( .D(out[1523]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1523]) );
  DFF \round_reg_reg[1524]  ( .D(out[1524]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1524]) );
  DFF \round_reg_reg[1525]  ( .D(out[1525]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1525]) );
  DFF \round_reg_reg[1526]  ( .D(out[1526]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1526]) );
  DFF \round_reg_reg[1527]  ( .D(out[1527]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1527]) );
  DFF \round_reg_reg[1528]  ( .D(out[1528]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1528]) );
  DFF \round_reg_reg[1529]  ( .D(out[1529]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1529]) );
  DFF \round_reg_reg[1530]  ( .D(out[1530]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1530]) );
  DFF \round_reg_reg[1531]  ( .D(out[1531]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1531]) );
  DFF \round_reg_reg[1532]  ( .D(out[1532]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1532]) );
  DFF \round_reg_reg[1533]  ( .D(out[1533]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1533]) );
  DFF \round_reg_reg[1534]  ( .D(out[1534]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1534]) );
  DFF \round_reg_reg[1535]  ( .D(out[1535]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1535]) );
  DFF \round_reg_reg[1536]  ( .D(out[1536]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1536]) );
  DFF \round_reg_reg[1537]  ( .D(out[1537]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1537]) );
  DFF \round_reg_reg[1538]  ( .D(out[1538]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1538]) );
  DFF \round_reg_reg[1539]  ( .D(out[1539]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1539]) );
  DFF \round_reg_reg[1540]  ( .D(out[1540]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1540]) );
  DFF \round_reg_reg[1541]  ( .D(out[1541]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1541]) );
  DFF \round_reg_reg[1542]  ( .D(out[1542]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1542]) );
  DFF \round_reg_reg[1543]  ( .D(out[1543]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1543]) );
  DFF \round_reg_reg[1544]  ( .D(out[1544]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1544]) );
  DFF \round_reg_reg[1545]  ( .D(out[1545]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1545]) );
  DFF \round_reg_reg[1546]  ( .D(out[1546]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1546]) );
  DFF \round_reg_reg[1547]  ( .D(out[1547]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1547]) );
  DFF \round_reg_reg[1548]  ( .D(out[1548]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1548]) );
  DFF \round_reg_reg[1549]  ( .D(out[1549]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1549]) );
  DFF \round_reg_reg[1550]  ( .D(out[1550]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1550]) );
  DFF \round_reg_reg[1551]  ( .D(out[1551]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1551]) );
  DFF \round_reg_reg[1552]  ( .D(out[1552]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1552]) );
  DFF \round_reg_reg[1553]  ( .D(out[1553]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1553]) );
  DFF \round_reg_reg[1554]  ( .D(out[1554]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1554]) );
  DFF \round_reg_reg[1555]  ( .D(out[1555]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1555]) );
  DFF \round_reg_reg[1556]  ( .D(out[1556]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1556]) );
  DFF \round_reg_reg[1557]  ( .D(out[1557]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1557]) );
  DFF \round_reg_reg[1558]  ( .D(out[1558]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1558]) );
  DFF \round_reg_reg[1559]  ( .D(out[1559]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1559]) );
  DFF \round_reg_reg[1560]  ( .D(out[1560]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1560]) );
  DFF \round_reg_reg[1561]  ( .D(out[1561]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1561]) );
  DFF \round_reg_reg[1562]  ( .D(out[1562]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1562]) );
  DFF \round_reg_reg[1563]  ( .D(out[1563]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1563]) );
  DFF \round_reg_reg[1564]  ( .D(out[1564]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1564]) );
  DFF \round_reg_reg[1565]  ( .D(out[1565]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1565]) );
  DFF \round_reg_reg[1566]  ( .D(out[1566]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1566]) );
  DFF \round_reg_reg[1567]  ( .D(out[1567]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1567]) );
  DFF \round_reg_reg[1568]  ( .D(out[1568]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1568]) );
  DFF \round_reg_reg[1569]  ( .D(out[1569]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1569]) );
  DFF \round_reg_reg[1570]  ( .D(out[1570]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1570]) );
  DFF \round_reg_reg[1571]  ( .D(out[1571]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1571]) );
  DFF \round_reg_reg[1572]  ( .D(out[1572]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1572]) );
  DFF \round_reg_reg[1573]  ( .D(out[1573]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1573]) );
  DFF \round_reg_reg[1574]  ( .D(out[1574]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1574]) );
  DFF \round_reg_reg[1575]  ( .D(out[1575]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1575]) );
  DFF \round_reg_reg[1576]  ( .D(out[1576]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1576]) );
  DFF \round_reg_reg[1577]  ( .D(out[1577]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1577]) );
  DFF \round_reg_reg[1578]  ( .D(out[1578]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1578]) );
  DFF \round_reg_reg[1579]  ( .D(out[1579]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1579]) );
  DFF \round_reg_reg[1580]  ( .D(out[1580]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1580]) );
  DFF \round_reg_reg[1581]  ( .D(out[1581]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1581]) );
  DFF \round_reg_reg[1582]  ( .D(out[1582]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1582]) );
  DFF \round_reg_reg[1583]  ( .D(out[1583]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1583]) );
  DFF \round_reg_reg[1584]  ( .D(out[1584]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1584]) );
  DFF \round_reg_reg[1585]  ( .D(out[1585]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1585]) );
  DFF \round_reg_reg[1586]  ( .D(out[1586]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1586]) );
  DFF \round_reg_reg[1587]  ( .D(out[1587]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1587]) );
  DFF \round_reg_reg[1588]  ( .D(out[1588]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1588]) );
  DFF \round_reg_reg[1589]  ( .D(out[1589]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1589]) );
  DFF \round_reg_reg[1590]  ( .D(out[1590]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1590]) );
  DFF \round_reg_reg[1591]  ( .D(out[1591]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1591]) );
  DFF \round_reg_reg[1592]  ( .D(out[1592]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1592]) );
  DFF \round_reg_reg[1593]  ( .D(out[1593]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1593]) );
  DFF \round_reg_reg[1594]  ( .D(out[1594]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1594]) );
  DFF \round_reg_reg[1595]  ( .D(out[1595]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1595]) );
  DFF \round_reg_reg[1596]  ( .D(out[1596]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1596]) );
  DFF \round_reg_reg[1597]  ( .D(out[1597]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1597]) );
  DFF \round_reg_reg[1598]  ( .D(out[1598]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1598]) );
  DFF \round_reg_reg[1599]  ( .D(out[1599]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1599]) );
  XNOR U1032 ( .A(n40641), .B(n40640), .Z(n38766) );
  XNOR U1033 ( .A(n41717), .B(n41716), .Z(n37331) );
  XNOR U1034 ( .A(n35847), .B(n36797), .Z(n27933) );
  ANDN U1035 ( .B(n47651), .A(n47653), .Z(n49594) );
  AND U1036 ( .A(n50369), .B(n50403), .Z(n52817) );
  ANDN U1037 ( .B(n46623), .A(n46622), .Z(n46620) );
  AND U1038 ( .A(n50254), .B(n50255), .Z(n50252) );
  AND U1039 ( .A(n49102), .B(n49103), .Z(n49100) );
  ANDN U1040 ( .B(n47296), .A(n47297), .Z(n49794) );
  XNOR U1041 ( .A(n47245), .B(n45221), .Z(n40643) );
  XNOR U1042 ( .A(n45472), .B(n44280), .Z(n40967) );
  AND U1043 ( .A(n43943), .B(n43944), .Z(n45114) );
  XOR U1044 ( .A(n41860), .B(n39636), .Z(n37018) );
  AND U1045 ( .A(n33889), .B(n37895), .Z(n40901) );
  AND U1046 ( .A(n33844), .B(n33845), .Z(n39858) );
  NOR U1047 ( .A(n37131), .B(n37470), .Z(n38581) );
  ANDN U1048 ( .B(n36283), .A(n36285), .Z(n36284) );
  ANDN U1049 ( .B(n34564), .A(n34563), .Z(n34562) );
  XOR U1050 ( .A(n38510), .B(n35255), .Z(n34955) );
  XNOR U1051 ( .A(n32949), .B(n36268), .Z(n34320) );
  XOR U1052 ( .A(n34403), .B(n33062), .Z(n29324) );
  ANDN U1053 ( .B(n25529), .A(n25531), .Z(n28805) );
  XOR U1054 ( .A(n31109), .B(n26357), .Z(n24387) );
  AND U1055 ( .A(n28017), .B(n28019), .Z(n28410) );
  AND U1056 ( .A(n26937), .B(n27030), .Z(n27450) );
  AND U1057 ( .A(n29650), .B(n29651), .Z(n29649) );
  XOR U1058 ( .A(n26119), .B(n27060), .Z(n26280) );
  XNOR U1059 ( .A(n28358), .B(n23558), .Z(n21048) );
  XNOR U1060 ( .A(n23991), .B(n24791), .Z(n22040) );
  ANDN U1061 ( .B(n19911), .A(n19910), .Z(n19908) );
  ANDN U1062 ( .B(n13970), .A(n14379), .Z(n17120) );
  XNOR U1063 ( .A(n14488), .B(n11937), .Z(n13695) );
  NOR U1064 ( .A(n11542), .B(n11541), .Z(n13800) );
  AND U1065 ( .A(n8349), .B(n11533), .Z(n11658) );
  XNOR U1066 ( .A(n14473), .B(n9198), .Z(n9189) );
  XNOR U1067 ( .A(n52222), .B(n52099), .Z(n49080) );
  XNOR U1068 ( .A(n52342), .B(n52341), .Z(n50227) );
  XNOR U1069 ( .A(n52294), .B(n53133), .Z(n51547) );
  XNOR U1070 ( .A(round_reg[1511]), .B(n51947), .Z(n50689) );
  XNOR U1071 ( .A(round_reg[290]), .B(n50822), .Z(n50351) );
  ANDN U1072 ( .B(n48464), .A(n48463), .Z(n48461) );
  AND U1073 ( .A(n49504), .B(n49445), .Z(n50113) );
  ANDN U1074 ( .B(n47736), .A(n47738), .Z(n50953) );
  ANDN U1075 ( .B(n49349), .A(n49350), .Z(n50186) );
  ANDN U1076 ( .B(n49191), .A(n49190), .Z(n49188) );
  AND U1077 ( .A(n47208), .B(n47207), .Z(n52147) );
  XNOR U1078 ( .A(n50000), .B(n46914), .Z(n47388) );
  ANDN U1079 ( .B(n46136), .A(n46137), .Z(n52098) );
  AND U1080 ( .A(n49520), .B(n48782), .Z(n52280) );
  AND U1081 ( .A(n49725), .B(n49724), .Z(n49722) );
  ANDN U1082 ( .B(n47018), .A(n47019), .Z(n51008) );
  AND U1083 ( .A(n49744), .B(n50881), .Z(n51458) );
  ANDN U1084 ( .B(n51744), .A(n51745), .Z(n52060) );
  ANDN U1085 ( .B(n47830), .A(n47829), .Z(n47827) );
  ANDN U1086 ( .B(n49302), .A(n49301), .Z(n49299) );
  XOR U1087 ( .A(n49327), .B(n49326), .Z(n45734) );
  XNOR U1088 ( .A(n46824), .B(n46823), .Z(n41747) );
  XNOR U1089 ( .A(n51632), .B(n49682), .Z(n45928) );
  AND U1090 ( .A(n48172), .B(n48877), .Z(n48875) );
  XNOR U1091 ( .A(n49353), .B(n49352), .Z(n44837) );
  NAND U1092 ( .A(n47116), .B(n46958), .Z(n48448) );
  XOR U1093 ( .A(n47253), .B(n47252), .Z(n46120) );
  XOR U1094 ( .A(n48429), .B(n48428), .Z(n44173) );
  XNOR U1095 ( .A(n46409), .B(n46408), .Z(n42419) );
  XNOR U1096 ( .A(n50779), .B(n48437), .Z(n44523) );
  XNOR U1097 ( .A(n43589), .B(n42540), .Z(n42183) );
  XOR U1098 ( .A(n44474), .B(n44475), .Z(n37013) );
  ANDN U1099 ( .B(n41417), .A(n41416), .Z(n41414) );
  ANDN U1100 ( .B(n41823), .A(n42025), .Z(n43522) );
  XNOR U1101 ( .A(n41570), .B(n41569), .Z(n39692) );
  ANDN U1102 ( .B(n44296), .A(n44295), .Z(n44294) );
  AND U1103 ( .A(n42924), .B(n42925), .Z(n42923) );
  AND U1104 ( .A(n43012), .B(n43100), .Z(n44708) );
  XNOR U1105 ( .A(n42729), .B(n42730), .Z(n37963) );
  AND U1106 ( .A(n40163), .B(n40161), .Z(n45670) );
  ANDN U1107 ( .B(n40506), .A(n40505), .Z(n40503) );
  ANDN U1108 ( .B(n39721), .A(n45549), .Z(n46369) );
  XOR U1109 ( .A(n42118), .B(n42119), .Z(n36546) );
  ANDN U1110 ( .B(n42798), .A(n42800), .Z(n44427) );
  ANDN U1111 ( .B(n43242), .A(n45018), .Z(n45017) );
  ANDN U1112 ( .B(n44127), .A(n42998), .Z(n44126) );
  XNOR U1113 ( .A(n40096), .B(n40095), .Z(n36434) );
  XNOR U1114 ( .A(n41078), .B(n41077), .Z(n37517) );
  XNOR U1115 ( .A(n43569), .B(n39633), .Z(n34623) );
  XOR U1116 ( .A(n42963), .B(n42070), .Z(n37720) );
  AND U1117 ( .A(n37559), .B(n37560), .Z(n37558) );
  AND U1118 ( .A(n35971), .B(n36991), .Z(n36989) );
  AND U1119 ( .A(n36788), .B(n36337), .Z(n36786) );
  ANDN U1120 ( .B(n35123), .A(n35121), .Z(n41661) );
  ANDN U1121 ( .B(n37485), .A(n37135), .Z(n38576) );
  XNOR U1122 ( .A(n33910), .B(n33955), .Z(n34604) );
  AND U1123 ( .A(n33861), .B(n33862), .Z(n33859) );
  XOR U1124 ( .A(n37819), .B(n35727), .Z(n31705) );
  AND U1125 ( .A(n35706), .B(n34960), .Z(n37327) );
  ANDN U1126 ( .B(n34675), .A(n34674), .Z(n38763) );
  XNOR U1127 ( .A(n33450), .B(n33449), .Z(n31434) );
  XNOR U1128 ( .A(n33961), .B(n33960), .Z(n33359) );
  XNOR U1129 ( .A(n34160), .B(n34159), .Z(n31154) );
  XNOR U1130 ( .A(n38226), .B(n38225), .Z(n30743) );
  XOR U1131 ( .A(n31240), .B(n31329), .Z(n30155) );
  NOR U1132 ( .A(n29444), .B(n29443), .Z(n29442) );
  ANDN U1133 ( .B(n27547), .A(n27546), .Z(n27544) );
  NOR U1134 ( .A(n29140), .B(n29141), .Z(n31545) );
  ANDN U1135 ( .B(n27951), .A(n27813), .Z(n28563) );
  ANDN U1136 ( .B(n28209), .A(n27599), .Z(n36267) );
  NANDN U1137 ( .A(n30966), .B(n29625), .Z(n32137) );
  AND U1138 ( .A(n27483), .B(n27482), .Z(n29321) );
  NOR U1139 ( .A(n26946), .B(n27128), .Z(n27649) );
  AND U1140 ( .A(n29475), .B(n29476), .Z(n29473) );
  ANDN U1141 ( .B(n27461), .A(n27462), .Z(n28869) );
  AND U1142 ( .A(n31033), .B(n30925), .Z(n31789) );
  ANDN U1143 ( .B(n28581), .A(n28582), .Z(n30133) );
  AND U1144 ( .A(n27631), .B(n27632), .Z(n27629) );
  XOR U1145 ( .A(n29656), .B(n27579), .Z(n22982) );
  XNOR U1146 ( .A(n25214), .B(n23815), .Z(n19528) );
  XOR U1147 ( .A(n26950), .B(n21992), .Z(n19058) );
  AND U1148 ( .A(n22745), .B(n23657), .Z(n23656) );
  XNOR U1149 ( .A(n18852), .B(n18606), .Z(n18480) );
  XOR U1150 ( .A(n23719), .B(n22840), .Z(n17667) );
  AND U1151 ( .A(n20574), .B(n22326), .Z(n26478) );
  AND U1152 ( .A(n24653), .B(n24764), .Z(n24796) );
  AND U1153 ( .A(n22714), .B(n22712), .Z(n25407) );
  AND U1154 ( .A(n20578), .B(n20580), .Z(n24804) );
  ANDN U1155 ( .B(n20441), .A(n22900), .Z(n22897) );
  XNOR U1156 ( .A(n19311), .B(n20360), .Z(n18332) );
  AND U1157 ( .A(n20564), .B(n21969), .Z(n24513) );
  XNOR U1158 ( .A(n21201), .B(n20373), .Z(n17203) );
  XOR U1159 ( .A(n19015), .B(n20097), .Z(n17333) );
  XNOR U1160 ( .A(n21096), .B(n18100), .Z(n14941) );
  XNOR U1161 ( .A(n18037), .B(n18027), .Z(n13684) );
  XOR U1162 ( .A(n14944), .B(n14945), .Z(n12112) );
  AND U1163 ( .A(n15151), .B(n15149), .Z(n19473) );
  ANDN U1164 ( .B(n12462), .A(n16128), .Z(n17867) );
  AND U1165 ( .A(n17369), .B(n17370), .Z(n22664) );
  ANDN U1166 ( .B(n16549), .A(n14772), .Z(n19612) );
  XOR U1167 ( .A(n16466), .B(n15542), .Z(n14474) );
  XOR U1168 ( .A(n16776), .B(n16777), .Z(n13381) );
  XOR U1169 ( .A(n12741), .B(n11865), .Z(n9238) );
  AND U1170 ( .A(n7743), .B(n10248), .Z(n10431) );
  AND U1171 ( .A(n8626), .B(n9308), .Z(n9306) );
  ANDN U1172 ( .B(n9213), .A(n7979), .Z(n9211) );
  ANDN U1173 ( .B(n7388), .A(n7387), .Z(n7385) );
  AND U1174 ( .A(n7158), .B(n8338), .Z(n11236) );
  AND U1175 ( .A(n10573), .B(n10572), .Z(n10730) );
  AND U1176 ( .A(n11530), .B(n11531), .Z(n13845) );
  AND U1177 ( .A(n8162), .B(n11009), .Z(n11133) );
  XOR U1178 ( .A(n9908), .B(n6817), .Z(n7503) );
  ANDN U1179 ( .B(n8557), .A(n8458), .Z(n8556) );
  ANDN U1180 ( .B(n10556), .A(n8914), .Z(n10674) );
  XNOR U1181 ( .A(n6298), .B(n9183), .Z(n1732) );
  XNOR U1182 ( .A(n6244), .B(n8341), .Z(n1667) );
  XNOR U1183 ( .A(n52970), .B(n52969), .Z(n52081) );
  XNOR U1184 ( .A(n52010), .B(n52612), .Z(n50650) );
  XNOR U1185 ( .A(round_reg[963]), .B(n51985), .Z(n48334) );
  XNOR U1186 ( .A(round_reg[662]), .B(n48945), .Z(n47691) );
  XNOR U1187 ( .A(round_reg[196]), .B(n50505), .Z(n47274) );
  XNOR U1188 ( .A(round_reg[1495]), .B(n50995), .Z(n50602) );
  AND U1189 ( .A(n49645), .B(n49402), .Z(n51957) );
  AND U1190 ( .A(n47212), .B(n47211), .Z(n52151) );
  ANDN U1191 ( .B(n50088), .A(n50089), .Z(n51365) );
  ANDN U1192 ( .B(n46836), .A(n51282), .Z(n53469) );
  ANDN U1193 ( .B(n48215), .A(n48276), .Z(n50833) );
  XOR U1194 ( .A(n49521), .B(n48790), .Z(n44796) );
  AND U1195 ( .A(n47799), .B(n47800), .Z(n50776) );
  XNOR U1196 ( .A(n46794), .B(n47263), .Z(n44932) );
  AND U1197 ( .A(n48597), .B(n50393), .Z(n52765) );
  ANDN U1198 ( .B(n48157), .A(n51643), .Z(n51665) );
  AND U1199 ( .A(n50912), .B(n50913), .Z(n50910) );
  ANDN U1200 ( .B(n51884), .A(n50203), .Z(n52340) );
  ANDN U1201 ( .B(n47617), .A(n48880), .Z(n49831) );
  ANDN U1202 ( .B(n51044), .A(n49254), .Z(n52140) );
  ANDN U1203 ( .B(n47770), .A(n49120), .Z(n51142) );
  ANDN U1204 ( .B(n50605), .A(n50604), .Z(n50603) );
  XNOR U1205 ( .A(n46532), .B(n46531), .Z(n45403) );
  XNOR U1206 ( .A(n45727), .B(n45726), .Z(n41735) );
  AND U1207 ( .A(n49462), .B(n49500), .Z(n50105) );
  AND U1208 ( .A(n45878), .B(n45879), .Z(n50724) );
  AND U1209 ( .A(n47626), .B(n47627), .Z(n47624) );
  AND U1210 ( .A(n48926), .B(n48433), .Z(n48925) );
  XOR U1211 ( .A(n52047), .B(n51297), .Z(n50959) );
  ANDN U1212 ( .B(n49713), .A(n49712), .Z(n49711) );
  XNOR U1213 ( .A(n45451), .B(n48166), .Z(n44479) );
  ANDN U1214 ( .B(n49974), .A(n49975), .Z(n51858) );
  ANDN U1215 ( .B(n46960), .A(n46959), .Z(n46957) );
  XOR U1216 ( .A(n51394), .B(n49529), .Z(n44013) );
  AND U1217 ( .A(n48882), .B(n48181), .Z(n48881) );
  ANDN U1218 ( .B(n47366), .A(n48082), .Z(n49788) );
  XOR U1219 ( .A(n50102), .B(n50101), .Z(n43327) );
  XNOR U1220 ( .A(n47132), .B(n47131), .Z(n44686) );
  XNOR U1221 ( .A(n46498), .B(n48287), .Z(n46403) );
  XNOR U1222 ( .A(n47108), .B(n46798), .Z(n41874) );
  XNOR U1223 ( .A(n50144), .B(n50143), .Z(n43819) );
  XNOR U1224 ( .A(n49997), .B(n49996), .Z(n45415) );
  XNOR U1225 ( .A(n42519), .B(n42419), .Z(n40282) );
  XNOR U1226 ( .A(n45666), .B(n45135), .Z(n40311) );
  XNOR U1227 ( .A(n43346), .B(n43345), .Z(n41723) );
  XOR U1228 ( .A(n45370), .B(n45371), .Z(n40816) );
  XNOR U1229 ( .A(n43083), .B(n46034), .Z(n44104) );
  AND U1230 ( .A(n41277), .B(n41278), .Z(n41275) );
  AND U1231 ( .A(n40286), .B(n40285), .Z(n42197) );
  XNOR U1232 ( .A(n38708), .B(n38707), .Z(n35297) );
  AND U1233 ( .A(n43310), .B(n41478), .Z(n43963) );
  ANDN U1234 ( .B(n41955), .A(n41045), .Z(n45192) );
  AND U1235 ( .A(n41410), .B(n44090), .Z(n44457) );
  AND U1236 ( .A(n43359), .B(n43880), .Z(n43879) );
  AND U1237 ( .A(n43700), .B(n43701), .Z(n43699) );
  AND U1238 ( .A(n39506), .B(n46230), .Z(n46228) );
  ANDN U1239 ( .B(n45048), .A(n45049), .Z(n45923) );
  ANDN U1240 ( .B(n43473), .A(n42903), .Z(n43470) );
  AND U1241 ( .A(n42945), .B(n42946), .Z(n42943) );
  AND U1242 ( .A(n45003), .B(n43250), .Z(n45001) );
  AND U1243 ( .A(n40420), .B(n40838), .Z(n47062) );
  AND U1244 ( .A(n43216), .B(n42736), .Z(n43214) );
  XOR U1245 ( .A(n44945), .B(n42750), .Z(n43634) );
  AND U1246 ( .A(n42138), .B(n43128), .Z(n43126) );
  XOR U1247 ( .A(n41317), .B(n41318), .Z(n36389) );
  AND U1248 ( .A(n39914), .B(n41243), .Z(n45620) );
  AND U1249 ( .A(n39208), .B(n39206), .Z(n44760) );
  XOR U1250 ( .A(n44424), .B(n40807), .Z(n39516) );
  XOR U1251 ( .A(n42716), .B(n42717), .Z(n40669) );
  XNOR U1252 ( .A(n39156), .B(n39155), .Z(n36946) );
  AND U1253 ( .A(n42583), .B(n42582), .Z(n46006) );
  XOR U1254 ( .A(n42070), .B(n41490), .Z(n38438) );
  XNOR U1255 ( .A(n40465), .B(n40464), .Z(n38306) );
  ANDN U1256 ( .B(n43072), .A(n41271), .Z(n44171) );
  ANDN U1257 ( .B(n45532), .A(n43732), .Z(n46425) );
  XNOR U1258 ( .A(n45409), .B(n40710), .Z(n39825) );
  AND U1259 ( .A(n42990), .B(n42988), .Z(n45678) );
  ANDN U1260 ( .B(n43817), .A(n43407), .Z(n48796) );
  XOR U1261 ( .A(n39223), .B(n40348), .Z(n39312) );
  XNOR U1262 ( .A(n40215), .B(n40943), .Z(n38332) );
  XNOR U1263 ( .A(n43725), .B(n40920), .Z(n35376) );
  XNOR U1264 ( .A(n41513), .B(n41088), .Z(n37928) );
  XNOR U1265 ( .A(n39986), .B(n39985), .Z(n39982) );
  XOR U1266 ( .A(n39744), .B(n42804), .Z(n38419) );
  XNOR U1267 ( .A(n43498), .B(n43790), .Z(n36212) );
  XNOR U1268 ( .A(n42055), .B(n42054), .Z(n38843) );
  XOR U1269 ( .A(n37670), .B(n37044), .Z(n34849) );
  XNOR U1270 ( .A(n40186), .B(n34623), .Z(n33572) );
  XOR U1271 ( .A(n39242), .B(n38248), .Z(n34775) );
  XNOR U1272 ( .A(n38086), .B(n36308), .Z(n36712) );
  AND U1273 ( .A(n38289), .B(n35555), .Z(n39452) );
  AND U1274 ( .A(n36487), .B(n36060), .Z(n38356) );
  XNOR U1275 ( .A(n34179), .B(n34178), .Z(n30500) );
  AND U1276 ( .A(n35184), .B(n37249), .Z(n38926) );
  XNOR U1277 ( .A(n36471), .B(n36472), .Z(n31830) );
  XNOR U1278 ( .A(n39560), .B(n33480), .Z(n30532) );
  AND U1279 ( .A(n33403), .B(n33401), .Z(n38630) );
  AND U1280 ( .A(n33120), .B(n37611), .Z(n37608) );
  XOR U1281 ( .A(n36120), .B(n34681), .Z(n33541) );
  AND U1282 ( .A(n34917), .B(n34918), .Z(n36686) );
  AND U1283 ( .A(n36051), .B(n36049), .Z(n38022) );
  ANDN U1284 ( .B(n36328), .A(n36791), .Z(n36789) );
  XOR U1285 ( .A(n37487), .B(n37483), .Z(n37126) );
  ANDN U1286 ( .B(n34745), .A(n36373), .Z(n39836) );
  ANDN U1287 ( .B(n34725), .A(n34861), .Z(n39807) );
  ANDN U1288 ( .B(n36457), .A(n36296), .Z(n36456) );
  AND U1289 ( .A(n35987), .B(n36451), .Z(n36452) );
  AND U1290 ( .A(n33751), .B(n38841), .Z(n50070) );
  AND U1291 ( .A(n37131), .B(n37133), .Z(n37469) );
  XNOR U1292 ( .A(n33181), .B(n33180), .Z(n29946) );
  AND U1293 ( .A(n35908), .B(n35909), .Z(n35906) );
  ANDN U1294 ( .B(n34290), .A(n34291), .Z(n39532) );
  AND U1295 ( .A(n37233), .B(n37232), .Z(n39779) );
  XOR U1296 ( .A(n36216), .B(n35289), .Z(n27949) );
  ANDN U1297 ( .B(n37977), .A(n40070), .Z(n40299) );
  ANDN U1298 ( .B(n36758), .A(n38064), .Z(n40208) );
  AND U1299 ( .A(n37214), .B(n36256), .Z(n39760) );
  XOR U1300 ( .A(n35149), .B(n35396), .Z(n32142) );
  XNOR U1301 ( .A(n34790), .B(n36863), .Z(n32691) );
  AND U1302 ( .A(n33866), .B(n33867), .Z(n33864) );
  AND U1303 ( .A(n35174), .B(n35175), .Z(n35172) );
  AND U1304 ( .A(n34517), .B(n35678), .Z(n35676) );
  XNOR U1305 ( .A(n33675), .B(n35751), .Z(n33942) );
  ANDN U1306 ( .B(n33895), .A(n33896), .Z(n41756) );
  XNOR U1307 ( .A(n36582), .B(n36249), .Z(n32689) );
  XOR U1308 ( .A(n34432), .B(n38527), .Z(n30260) );
  XNOR U1309 ( .A(n33329), .B(n33328), .Z(n28995) );
  AND U1310 ( .A(n37961), .B(n33595), .Z(n40346) );
  XNOR U1311 ( .A(n36174), .B(n34949), .Z(n29071) );
  XNOR U1312 ( .A(n33490), .B(n33489), .Z(n31068) );
  AND U1313 ( .A(n36573), .B(n36574), .Z(n36572) );
  XNOR U1314 ( .A(n34020), .B(n33717), .Z(n31542) );
  XOR U1315 ( .A(n31261), .B(n30258), .Z(n28531) );
  XNOR U1316 ( .A(n33412), .B(n30743), .Z(n30096) );
  XNOR U1317 ( .A(n31212), .B(n29067), .Z(n29029) );
  XOR U1318 ( .A(n31177), .B(n31178), .Z(n29806) );
  ANDN U1319 ( .B(n26592), .A(n26593), .Z(n28369) );
  AND U1320 ( .A(n30410), .B(n29198), .Z(n30408) );
  ANDN U1321 ( .B(n29012), .A(n29011), .Z(n32374) );
  AND U1322 ( .A(n26802), .B(n28143), .Z(n34954) );
  ANDN U1323 ( .B(n32642), .A(n28307), .Z(n34536) );
  AND U1324 ( .A(n28413), .B(n28822), .Z(n28819) );
  AND U1325 ( .A(n27086), .B(n28606), .Z(n28605) );
  AND U1326 ( .A(n28525), .B(n28526), .Z(n28523) );
  ANDN U1327 ( .B(n28691), .A(n28689), .Z(n29868) );
  AND U1328 ( .A(n28667), .B(n29404), .Z(n34269) );
  AND U1329 ( .A(n27531), .B(n27533), .Z(n37729) );
  ANDN U1330 ( .B(n26355), .A(n27660), .Z(n36761) );
  ANDN U1331 ( .B(n32075), .A(n27208), .Z(n33601) );
  XOR U1332 ( .A(n29920), .B(n26854), .Z(n24694) );
  ANDN U1333 ( .B(n27869), .A(n27766), .Z(n38231) );
  ANDN U1334 ( .B(n27523), .A(n27522), .Z(n27520) );
  ANDN U1335 ( .B(n26363), .A(n27132), .Z(n27131) );
  NOR U1336 ( .A(n29478), .B(n30392), .Z(n31431) );
  XOR U1337 ( .A(n31023), .B(n31024), .Z(n26640) );
  AND U1338 ( .A(n27551), .B(n27552), .Z(n27549) );
  AND U1339 ( .A(n27554), .B(n27555), .Z(n28967) );
  XNOR U1340 ( .A(n29883), .B(n31713), .Z(n22354) );
  ANDN U1341 ( .B(n30801), .A(n30599), .Z(n34064) );
  XOR U1342 ( .A(n28159), .B(n30725), .Z(n25109) );
  AND U1343 ( .A(n30103), .B(n28286), .Z(n31125) );
  AND U1344 ( .A(n28907), .B(n29259), .Z(n29256) );
  ANDN U1345 ( .B(n28376), .A(n26606), .Z(n35354) );
  ANDN U1346 ( .B(n31616), .A(n30841), .Z(n32764) );
  ANDN U1347 ( .B(n31442), .A(n30396), .Z(n38952) );
  XNOR U1348 ( .A(n26015), .B(n29279), .Z(n24402) );
  XNOR U1349 ( .A(n28417), .B(n28416), .Z(n22495) );
  AND U1350 ( .A(n28055), .B(n27382), .Z(n28054) );
  AND U1351 ( .A(n27444), .B(n27004), .Z(n27442) );
  XNOR U1352 ( .A(n28061), .B(n29311), .Z(n22534) );
  XNOR U1353 ( .A(n29705), .B(n27900), .Z(n23839) );
  XNOR U1354 ( .A(n31799), .B(n29650), .Z(n29373) );
  XNOR U1355 ( .A(n25199), .B(n25198), .Z(n22223) );
  XNOR U1356 ( .A(n29911), .B(n30726), .Z(n25152) );
  XNOR U1357 ( .A(n30225), .B(n30130), .Z(n23065) );
  XNOR U1358 ( .A(n27637), .B(n26763), .Z(n24926) );
  XNOR U1359 ( .A(n26199), .B(n27408), .Z(n23978) );
  XNOR U1360 ( .A(n27577), .B(n28870), .Z(n23442) );
  XNOR U1361 ( .A(n26246), .B(n26245), .Z(n25382) );
  XNOR U1362 ( .A(n27583), .B(n26795), .Z(n23964) );
  XOR U1363 ( .A(n24034), .B(n24035), .Z(n21450) );
  XNOR U1364 ( .A(n27873), .B(n24379), .Z(n21810) );
  XOR U1365 ( .A(n27795), .B(n27796), .Z(n21803) );
  ANDN U1366 ( .B(n20000), .A(n19861), .Z(n21582) );
  ANDN U1367 ( .B(n21555), .A(n21554), .Z(n21552) );
  XOR U1368 ( .A(n23073), .B(n20220), .Z(n22416) );
  ANDN U1369 ( .B(n23456), .A(n23457), .Z(n26277) );
  ANDN U1370 ( .B(n23679), .A(n23467), .Z(n32442) );
  AND U1371 ( .A(n23926), .B(n24475), .Z(n24717) );
  AND U1372 ( .A(n19572), .B(n19573), .Z(n19570) );
  AND U1373 ( .A(n24046), .B(n22073), .Z(n24754) );
  AND U1374 ( .A(n20749), .B(n20186), .Z(n20747) );
  ANDN U1375 ( .B(n21416), .A(n22018), .Z(n25497) );
  NOR U1376 ( .A(n22057), .B(n22056), .Z(n22054) );
  XNOR U1377 ( .A(n25191), .B(n24058), .Z(n24042) );
  XOR U1378 ( .A(n26459), .B(n21868), .Z(n21856) );
  XOR U1379 ( .A(n24352), .B(n24326), .Z(n21865) );
  AND U1380 ( .A(n23453), .B(n23454), .Z(n23451) );
  AND U1381 ( .A(n20949), .B(n20950), .Z(n20947) );
  AND U1382 ( .A(n20898), .B(n22137), .Z(n22136) );
  XOR U1383 ( .A(n19747), .B(n19746), .Z(n14158) );
  XNOR U1384 ( .A(n19557), .B(n18393), .Z(n16331) );
  XOR U1385 ( .A(n24952), .B(n22696), .Z(n17608) );
  XNOR U1386 ( .A(n19136), .B(n19135), .Z(n17994) );
  XNOR U1387 ( .A(n19677), .B(n19676), .Z(n19444) );
  ANDN U1388 ( .B(n24322), .A(n25386), .Z(n25385) );
  AND U1389 ( .A(n23163), .B(n23161), .Z(n30153) );
  XOR U1390 ( .A(n21458), .B(n21666), .Z(n16998) );
  XNOR U1391 ( .A(n20704), .B(n20703), .Z(n17646) );
  XOR U1392 ( .A(n19595), .B(n20672), .Z(n16868) );
  XOR U1393 ( .A(n22185), .B(n19956), .Z(n15256) );
  XNOR U1394 ( .A(n16031), .B(n16032), .Z(n13435) );
  XOR U1395 ( .A(n19669), .B(n16502), .Z(n13324) );
  XNOR U1396 ( .A(n18277), .B(n18276), .Z(n17314) );
  XNOR U1397 ( .A(n18369), .B(n16674), .Z(n17711) );
  XNOR U1398 ( .A(n20594), .B(n15635), .Z(n15801) );
  AND U1399 ( .A(n14698), .B(n15137), .Z(n15136) );
  ANDN U1400 ( .B(n19638), .A(n19645), .Z(n19643) );
  AND U1401 ( .A(n15168), .B(n15169), .Z(n15166) );
  ANDN U1402 ( .B(n17682), .A(n16135), .Z(n16132) );
  AND U1403 ( .A(n18115), .B(n17151), .Z(n19188) );
  AND U1404 ( .A(n12859), .B(n12860), .Z(n12857) );
  AND U1405 ( .A(n15224), .B(n14052), .Z(n18826) );
  AND U1406 ( .A(n13584), .B(n13585), .Z(n13582) );
  NOR U1407 ( .A(n16142), .B(n17694), .Z(n17692) );
  AND U1408 ( .A(n14405), .B(n14407), .Z(n19277) );
  XOR U1409 ( .A(n13504), .B(n13505), .Z(n12339) );
  XNOR U1410 ( .A(n14103), .B(n14104), .Z(n12607) );
  AND U1411 ( .A(n14782), .B(n14783), .Z(n14780) );
  AND U1412 ( .A(n15112), .B(n16652), .Z(n17996) );
  AND U1413 ( .A(n13255), .B(n14169), .Z(n14166) );
  ANDN U1414 ( .B(n15141), .A(n17256), .Z(n21687) );
  AND U1415 ( .A(n12823), .B(n12824), .Z(n12821) );
  XOR U1416 ( .A(n16018), .B(n16019), .Z(n12219) );
  AND U1417 ( .A(n16337), .B(n16880), .Z(n18491) );
  XOR U1418 ( .A(n22489), .B(n17766), .Z(n11831) );
  AND U1419 ( .A(n13109), .B(n13110), .Z(n19377) );
  AND U1420 ( .A(n15811), .B(n15812), .Z(n15809) );
  XNOR U1421 ( .A(n12817), .B(n12816), .Z(n10604) );
  XNOR U1422 ( .A(n16177), .B(n16176), .Z(n10741) );
  AND U1423 ( .A(n17156), .B(n17157), .Z(n17154) );
  XNOR U1424 ( .A(n15078), .B(n16263), .Z(n9524) );
  XNOR U1425 ( .A(n11122), .B(n12468), .Z(n9142) );
  XOR U1426 ( .A(n11820), .B(n10182), .Z(n9734) );
  XNOR U1427 ( .A(n10561), .B(n7794), .Z(n5064) );
  XOR U1428 ( .A(n7499), .B(n6821), .Z(n4928) );
  XOR U1429 ( .A(n8100), .B(n7008), .Z(n4958) );
  ANDN U1430 ( .B(n8419), .A(n8418), .Z(n8416) );
  ANDN U1431 ( .B(n8072), .A(n8071), .Z(n8069) );
  AND U1432 ( .A(n9286), .B(n9287), .Z(n9284) );
  AND U1433 ( .A(n8929), .B(n6574), .Z(n9014) );
  AND U1434 ( .A(n12131), .B(n8695), .Z(n12262) );
  AND U1435 ( .A(n8826), .B(n12434), .Z(n12666) );
  XNOR U1436 ( .A(n6335), .B(n6424), .Z(n5173) );
  XNOR U1437 ( .A(n6343), .B(n6477), .Z(n5179) );
  ANDN U1438 ( .B(n12900), .A(n8308), .Z(n13353) );
  AND U1439 ( .A(n7943), .B(n10661), .Z(n10808) );
  ANDN U1440 ( .B(n7043), .A(n8150), .Z(n10876) );
  ANDN U1441 ( .B(n6994), .A(n6993), .Z(n10453) );
  XOR U1442 ( .A(n13163), .B(n9062), .Z(n9040) );
  AND U1443 ( .A(n9083), .B(n9082), .Z(n9096) );
  ANDN U1444 ( .B(n10037), .A(n10036), .Z(n11162) );
  XOR U1445 ( .A(n11309), .B(n7638), .Z(n1688) );
  XOR U1446 ( .A(n7557), .B(n7558), .Z(n2168) );
  ANDN U1447 ( .B(n6545), .A(n8922), .Z(n8921) );
  AND U1448 ( .A(n7734), .B(n7659), .Z(n7733) );
  XOR U1449 ( .A(n6470), .B(n6471), .Z(n3656) );
  XOR U1450 ( .A(n9172), .B(n9173), .Z(n3890) );
  XNOR U1451 ( .A(n6043), .B(n6042), .Z(n2203) );
  XNOR U1452 ( .A(n8844), .B(n8843), .Z(n2440) );
  XNOR U1453 ( .A(n6294), .B(n9090), .Z(n1727) );
  XNOR U1454 ( .A(n6310), .B(n9497), .Z(n1745) );
  XOR U1455 ( .A(n5408), .B(n2248), .Z(n4508) );
  XNOR U1456 ( .A(n2332), .B(n7120), .Z(n1043) );
  XNOR U1457 ( .A(n3137), .B(n2280), .Z(n2685) );
  XNOR U1458 ( .A(n4872), .B(n2241), .Z(n1670) );
  AND U1459 ( .A(n4461), .B(n4462), .Z(n4459) );
  AND U1460 ( .A(n4517), .B(n4518), .Z(n4515) );
  AND U1461 ( .A(n4607), .B(n4608), .Z(n4605) );
  ANDN U1462 ( .B(n4679), .A(n4680), .Z(n4678) );
  ANDN U1463 ( .B(n4933), .A(n4741), .Z(n4931) );
  AND U1464 ( .A(n4965), .B(n4764), .Z(n4963) );
  NOR U1465 ( .A(n5753), .B(n1104), .Z(n5752) );
  AND U1466 ( .A(n1502), .B(n1221), .Z(n1501) );
  XNOR U1467 ( .A(n52225), .B(n52224), .Z(n51696) );
  XNOR U1468 ( .A(n52516), .B(n52271), .Z(n50110) );
  XOR U1469 ( .A(n52456), .B(n52227), .Z(n50739) );
  XOR U1470 ( .A(n53313), .B(n53620), .Z(n51199) );
  XNOR U1471 ( .A(n52586), .B(n52585), .Z(n50735) );
  XOR U1472 ( .A(n52338), .B(n52907), .Z(n51468) );
  XNOR U1473 ( .A(n53093), .B(n53092), .Z(n50984) );
  XNOR U1474 ( .A(n52301), .B(n52300), .Z(n51564) );
  XOR U1475 ( .A(round_reg[837]), .B(n48453), .Z(n46972) );
  XNOR U1476 ( .A(round_reg[157]), .B(n48517), .Z(n49007) );
  XNOR U1477 ( .A(round_reg[880]), .B(n48938), .Z(n47043) );
  XOR U1478 ( .A(round_reg[1136]), .B(n51818), .Z(n51251) );
  XNOR U1479 ( .A(round_reg[1146]), .B(n51620), .Z(n50035) );
  XNOR U1480 ( .A(round_reg[287]), .B(n50453), .Z(n48431) );
  XNOR U1481 ( .A(round_reg[78]), .B(n48957), .Z(n50492) );
  XNOR U1482 ( .A(round_reg[769]), .B(n50127), .Z(n46333) );
  AND U1483 ( .A(n49003), .B(n49002), .Z(n49000) );
  ANDN U1484 ( .B(n47426), .A(n48614), .Z(n52548) );
  AND U1485 ( .A(n46329), .B(n46327), .Z(n51546) );
  AND U1486 ( .A(n51294), .B(n49060), .Z(n53529) );
  ANDN U1487 ( .B(n48587), .A(n48588), .Z(n48764) );
  ANDN U1488 ( .B(n47768), .A(n47769), .Z(n49611) );
  ANDN U1489 ( .B(n50810), .A(n50809), .Z(n50807) );
  ANDN U1490 ( .B(n50178), .A(n48849), .Z(n51152) );
  AND U1491 ( .A(n48515), .B(n46325), .Z(n48513) );
  ANDN U1492 ( .B(n50584), .A(n48704), .Z(n52146) );
  ANDN U1493 ( .B(n48063), .A(n48064), .Z(n52364) );
  ANDN U1494 ( .B(n46050), .A(n46051), .Z(n51012) );
  ANDN U1495 ( .B(n49721), .A(n49720), .Z(n49718) );
  AND U1496 ( .A(n47507), .B(n47508), .Z(n47505) );
  ANDN U1497 ( .B(n47008), .A(n46854), .Z(n52401) );
  ANDN U1498 ( .B(n48692), .A(n48655), .Z(n51596) );
  ANDN U1499 ( .B(n49971), .A(n49972), .Z(n51852) );
  AND U1500 ( .A(n51319), .B(n50303), .Z(n51704) );
  ANDN U1501 ( .B(n48536), .A(n48535), .Z(n48533) );
  AND U1502 ( .A(n48897), .B(n48898), .Z(n48895) );
  ANDN U1503 ( .B(n50313), .A(n47230), .Z(n51802) );
  AND U1504 ( .A(n47865), .B(n49781), .Z(n52406) );
  ANDN U1505 ( .B(n46964), .A(n46963), .Z(n46961) );
  AND U1506 ( .A(n49305), .B(n49941), .Z(n51000) );
  XOR U1507 ( .A(n52048), .B(n51291), .Z(n47567) );
  AND U1508 ( .A(n46143), .B(n46144), .Z(n46141) );
  ANDN U1509 ( .B(n49389), .A(n49390), .Z(n52323) );
  ANDN U1510 ( .B(n48330), .A(n46777), .Z(n51986) );
  ANDN U1511 ( .B(n49198), .A(n49197), .Z(n49195) );
  XNOR U1512 ( .A(n47995), .B(n47972), .Z(n45828) );
  ANDN U1513 ( .B(n46477), .A(n46476), .Z(n46474) );
  AND U1514 ( .A(n48233), .B(n48234), .Z(n48231) );
  XNOR U1515 ( .A(n46428), .B(n46427), .Z(n44469) );
  XNOR U1516 ( .A(n49885), .B(n46583), .Z(n43671) );
  XNOR U1517 ( .A(n46706), .B(n46913), .Z(n46166) );
  AND U1518 ( .A(n50165), .B(n50166), .Z(n50164) );
  XNOR U1519 ( .A(n48349), .B(n48107), .Z(n45371) );
  XNOR U1520 ( .A(n46584), .B(n49395), .Z(n45519) );
  AND U1521 ( .A(n49460), .B(n49458), .Z(n49816) );
  ANDN U1522 ( .B(n48992), .A(n50802), .Z(n51791) );
  AND U1523 ( .A(n51277), .B(n51278), .Z(n51276) );
  XNOR U1524 ( .A(n46127), .B(n45937), .Z(n42219) );
  XOR U1525 ( .A(n51387), .B(n51388), .Z(n46496) );
  XOR U1526 ( .A(n47237), .B(n47236), .Z(n45664) );
  XNOR U1527 ( .A(n46349), .B(n46348), .Z(n42309) );
  XOR U1528 ( .A(n45093), .B(n43665), .Z(n41135) );
  XNOR U1529 ( .A(n47099), .B(n43680), .Z(n40858) );
  XOR U1530 ( .A(n43559), .B(n46007), .Z(n40261) );
  XNOR U1531 ( .A(n44947), .B(n41649), .Z(n43638) );
  XNOR U1532 ( .A(n45785), .B(n44220), .Z(n41020) );
  XNOR U1533 ( .A(n43597), .B(n43598), .Z(n41463) );
  ANDN U1534 ( .B(n41186), .A(n41185), .Z(n41183) );
  AND U1535 ( .A(n43082), .B(n43028), .Z(n44684) );
  XOR U1536 ( .A(n44261), .B(n43905), .Z(n39890) );
  AND U1537 ( .A(n40769), .B(n40770), .Z(n40767) );
  XNOR U1538 ( .A(n47399), .B(n43853), .Z(n41568) );
  AND U1539 ( .A(n42989), .B(n44137), .Z(n44136) );
  ANDN U1540 ( .B(n42765), .A(n42766), .Z(n44735) );
  XOR U1541 ( .A(n43065), .B(n43066), .Z(n41413) );
  AND U1542 ( .A(n40460), .B(n40459), .Z(n44542) );
  AND U1543 ( .A(n40156), .B(n42399), .Z(n42398) );
  AND U1544 ( .A(n45207), .B(n43842), .Z(n45205) );
  AND U1545 ( .A(n43172), .B(n43174), .Z(n43697) );
  AND U1546 ( .A(n41007), .B(n41005), .Z(n46173) );
  AND U1547 ( .A(n42940), .B(n43363), .Z(n43886) );
  AND U1548 ( .A(n40409), .B(n40594), .Z(n40593) );
  XNOR U1549 ( .A(n43994), .B(n40360), .Z(n34617) );
  XNOR U1550 ( .A(n41142), .B(n41141), .Z(n40827) );
  XOR U1551 ( .A(n41481), .B(n41482), .Z(n38128) );
  AND U1552 ( .A(n43518), .B(n43519), .Z(n43516) );
  AND U1553 ( .A(n40488), .B(n40489), .Z(n40486) );
  AND U1554 ( .A(n42289), .B(n42290), .Z(n45108) );
  AND U1555 ( .A(n43353), .B(n44228), .Z(n45706) );
  AND U1556 ( .A(n40602), .B(n40636), .Z(n40634) );
  NOR U1557 ( .A(n40682), .B(n40914), .Z(n40912) );
  XNOR U1558 ( .A(n44656), .B(n40223), .Z(n42711) );
  AND U1559 ( .A(n41999), .B(n43923), .Z(n45150) );
  NOR U1560 ( .A(n43233), .B(n44818), .Z(n44817) );
  ANDN U1561 ( .B(n43469), .A(n41693), .Z(n47323) );
  ANDN U1562 ( .B(n42260), .A(n42259), .Z(n42257) );
  XNOR U1563 ( .A(n40905), .B(n41024), .Z(n37008) );
  ANDN U1564 ( .B(n42865), .A(n45552), .Z(n46727) );
  XNOR U1565 ( .A(n49696), .B(n44651), .Z(n38586) );
  ANDN U1566 ( .B(n44235), .A(n40951), .Z(n44234) );
  XNOR U1567 ( .A(n40429), .B(n40428), .Z(n39596) );
  XNOR U1568 ( .A(n39759), .B(n39758), .Z(n38801) );
  ANDN U1569 ( .B(n42096), .A(n42095), .Z(n42093) );
  AND U1570 ( .A(n41812), .B(n41811), .Z(n46592) );
  AND U1571 ( .A(n43669), .B(n41859), .Z(n45174) );
  ANDN U1572 ( .B(n41291), .A(n41290), .Z(n41288) );
  XOR U1573 ( .A(n45609), .B(n43794), .Z(n39271) );
  AND U1574 ( .A(n42622), .B(n43806), .Z(n46202) );
  ANDN U1575 ( .B(n41285), .A(n41286), .Z(n41873) );
  XNOR U1576 ( .A(n41685), .B(n42758), .Z(n37420) );
  XNOR U1577 ( .A(n40674), .B(n39949), .Z(n34638) );
  XOR U1578 ( .A(n45398), .B(n40723), .Z(n39296) );
  XOR U1579 ( .A(n45851), .B(n41319), .Z(n39493) );
  AND U1580 ( .A(n39910), .B(n41237), .Z(n45633) );
  XOR U1581 ( .A(n39652), .B(n39651), .Z(n35938) );
  XNOR U1582 ( .A(n42122), .B(n40830), .Z(n39468) );
  AND U1583 ( .A(n43205), .B(n42740), .Z(n43203) );
  ANDN U1584 ( .B(n44965), .A(n41018), .Z(n44964) );
  ANDN U1585 ( .B(n41949), .A(n45194), .Z(n45193) );
  XOR U1586 ( .A(n40216), .B(n40215), .Z(n37714) );
  XNOR U1587 ( .A(n42226), .B(n42693), .Z(n35301) );
  XNOR U1588 ( .A(n41398), .B(n41397), .Z(n35944) );
  NAND U1589 ( .A(n40847), .B(n40411), .Z(n47105) );
  XNOR U1590 ( .A(n43274), .B(n45977), .Z(n35940) );
  ANDN U1591 ( .B(n43246), .A(n45016), .Z(n45013) );
  XOR U1592 ( .A(n39180), .B(n39179), .Z(n36359) );
  XNOR U1593 ( .A(n43619), .B(n40616), .Z(n36308) );
  XOR U1594 ( .A(n40469), .B(n40468), .Z(n38096) );
  XNOR U1595 ( .A(n39834), .B(n40378), .Z(n36794) );
  XNOR U1596 ( .A(n39793), .B(n36779), .Z(n36559) );
  XNOR U1597 ( .A(n43494), .B(n37011), .Z(n36105) );
  XNOR U1598 ( .A(n37766), .B(n36356), .Z(n36261) );
  XOR U1599 ( .A(n38684), .B(n38683), .Z(n36020) );
  XNOR U1600 ( .A(n37720), .B(n37933), .Z(n36193) );
  XNOR U1601 ( .A(n39923), .B(n35861), .Z(n31926) );
  AND U1602 ( .A(n33938), .B(n33939), .Z(n33936) );
  XOR U1603 ( .A(n38946), .B(n34472), .Z(n34424) );
  AND U1604 ( .A(n33979), .B(n33980), .Z(n33977) );
  XOR U1605 ( .A(n37142), .B(n34813), .Z(n29318) );
  AND U1606 ( .A(n34893), .B(n34892), .Z(n37944) );
  AND U1607 ( .A(n32856), .B(n33253), .Z(n38112) );
  NOR U1608 ( .A(n33989), .B(n33988), .Z(n33986) );
  AND U1609 ( .A(n33086), .B(n37093), .Z(n39553) );
  AND U1610 ( .A(n37298), .B(n37297), .Z(n37295) );
  ANDN U1611 ( .B(n35836), .A(n36017), .Z(n36403) );
  AND U1612 ( .A(n34479), .B(n34478), .Z(n38483) );
  ANDN U1613 ( .B(n34662), .A(n34661), .Z(n34659) );
  AND U1614 ( .A(n37762), .B(n38512), .Z(n38528) );
  AND U1615 ( .A(n34260), .B(n33627), .Z(n36365) );
  AND U1616 ( .A(n36463), .B(n36879), .Z(n36877) );
  XOR U1617 ( .A(n38296), .B(n38289), .Z(n35806) );
  XOR U1618 ( .A(n46186), .B(n35423), .Z(n32830) );
  ANDN U1619 ( .B(n35531), .A(n35101), .Z(n35530) );
  XNOR U1620 ( .A(n34250), .B(n34748), .Z(n32415) );
  AND U1621 ( .A(n36151), .B(n36150), .Z(n37739) );
  AND U1622 ( .A(n36266), .B(n36590), .Z(n36589) );
  AND U1623 ( .A(n34330), .B(n36774), .Z(n36772) );
  ANDN U1624 ( .B(n34943), .A(n34942), .Z(n34940) );
  ANDN U1625 ( .B(n35459), .A(n35458), .Z(n35457) );
  XNOR U1626 ( .A(n37174), .B(n35019), .Z(n33381) );
  XOR U1627 ( .A(n37544), .B(n35228), .Z(n31584) );
  AND U1628 ( .A(n38062), .B(n36747), .Z(n42387) );
  AND U1629 ( .A(n36745), .B(n38073), .Z(n40213) );
  ANDN U1630 ( .B(n37386), .A(n37387), .Z(n39614) );
  AND U1631 ( .A(n38015), .B(n38014), .Z(n38468) );
  AND U1632 ( .A(n35537), .B(n33437), .Z(n35925) );
  ANDN U1633 ( .B(n36062), .A(n36063), .Z(n38035) );
  AND U1634 ( .A(n33080), .B(n34739), .Z(n39829) );
  XNOR U1635 ( .A(n32618), .B(n34503), .Z(n31148) );
  AND U1636 ( .A(n36802), .B(n36801), .Z(n37415) );
  ANDN U1637 ( .B(n37281), .A(n37280), .Z(n37279) );
  AND U1638 ( .A(n36784), .B(n36335), .Z(n36781) );
  AND U1639 ( .A(n37483), .B(n37482), .Z(n38583) );
  XNOR U1640 ( .A(n35893), .B(n34666), .Z(n30524) );
  XOR U1641 ( .A(n39983), .B(n37649), .Z(n37353) );
  XOR U1642 ( .A(n35768), .B(n34832), .Z(n32547) );
  AND U1643 ( .A(n34468), .B(n34469), .Z(n34466) );
  XNOR U1644 ( .A(n35396), .B(n35395), .Z(n32402) );
  AND U1645 ( .A(n36723), .B(n36724), .Z(n36721) );
  ANDN U1646 ( .B(n35262), .A(n36577), .Z(n38994) );
  ANDN U1647 ( .B(n34762), .A(n34763), .Z(n38921) );
  XNOR U1648 ( .A(n34211), .B(n33880), .Z(n29922) );
  AND U1649 ( .A(n33322), .B(n34149), .Z(n34148) );
  XNOR U1650 ( .A(n34227), .B(n32211), .Z(n31772) );
  XOR U1651 ( .A(n33539), .B(n33538), .Z(n30507) );
  ANDN U1652 ( .B(n35266), .A(n35267), .Z(n37763) );
  XNOR U1653 ( .A(n38527), .B(n36243), .Z(n29943) );
  XNOR U1654 ( .A(n33368), .B(n33367), .Z(n30248) );
  XNOR U1655 ( .A(n34575), .B(n32961), .Z(n33303) );
  AND U1656 ( .A(n35727), .B(n35728), .Z(n35725) );
  XNOR U1657 ( .A(n32386), .B(n33852), .Z(n28836) );
  XOR U1658 ( .A(n33823), .B(n34020), .Z(n29734) );
  XNOR U1659 ( .A(n35289), .B(n32924), .Z(n31116) );
  XOR U1660 ( .A(n29045), .B(n35190), .Z(n28394) );
  XNOR U1661 ( .A(n27932), .B(n27933), .Z(n27632) );
  XNOR U1662 ( .A(n33946), .B(n30583), .Z(n30685) );
  XNOR U1663 ( .A(n33044), .B(n32511), .Z(n26324) );
  XNOR U1664 ( .A(n32694), .B(n31340), .Z(n30773) );
  XNOR U1665 ( .A(n36751), .B(n31539), .Z(n28207) );
  XNOR U1666 ( .A(n27936), .B(n27937), .Z(n27621) );
  AND U1667 ( .A(n29815), .B(n30680), .Z(n31134) );
  XOR U1668 ( .A(n31816), .B(n28942), .Z(n23587) );
  AND U1669 ( .A(n26808), .B(n26807), .Z(n32417) );
  XNOR U1670 ( .A(n32156), .B(n29664), .Z(n23149) );
  AND U1671 ( .A(n27745), .B(n26430), .Z(n30498) );
  AND U1672 ( .A(n27447), .B(n27022), .Z(n27446) );
  ANDN U1673 ( .B(n27713), .A(n28329), .Z(n31933) );
  XNOR U1674 ( .A(n27729), .B(n28271), .Z(n28725) );
  AND U1675 ( .A(n29092), .B(n27976), .Z(n32033) );
  AND U1676 ( .A(n28487), .B(n29177), .Z(n31151) );
  XNOR U1677 ( .A(n27901), .B(n27900), .Z(n22517) );
  AND U1678 ( .A(n29088), .B(n28647), .Z(n32876) );
  AND U1679 ( .A(n26737), .B(n26736), .Z(n26734) );
  ANDN U1680 ( .B(n30409), .A(n30410), .Z(n32615) );
  ANDN U1681 ( .B(n27297), .A(n27298), .Z(n28546) );
  AND U1682 ( .A(n27822), .B(n27821), .Z(n32566) );
  AND U1683 ( .A(n29550), .B(n30114), .Z(n34248) );
  XNOR U1684 ( .A(n27898), .B(n27897), .Z(n25551) );
  XOR U1685 ( .A(n31198), .B(n31199), .Z(n30021) );
  AND U1686 ( .A(n27626), .B(n27627), .Z(n27926) );
  XNOR U1687 ( .A(n30383), .B(n28342), .Z(n29450) );
  AND U1688 ( .A(n28629), .B(n28630), .Z(n28627) );
  XNOR U1689 ( .A(n26980), .B(n29502), .Z(n26904) );
  XNOR U1690 ( .A(n28270), .B(n25968), .Z(n25865) );
  ANDN U1691 ( .B(n29829), .A(n29828), .Z(n29827) );
  AND U1692 ( .A(n30832), .B(n30833), .Z(n30830) );
  AND U1693 ( .A(n28233), .B(n28234), .Z(n28231) );
  AND U1694 ( .A(n30052), .B(n29898), .Z(n30051) );
  ANDN U1695 ( .B(n28120), .A(n28119), .Z(n28117) );
  AND U1696 ( .A(n29001), .B(n29000), .Z(n30815) );
  XNOR U1697 ( .A(n30965), .B(n29627), .Z(n24006) );
  AND U1698 ( .A(n31090), .B(n30844), .Z(n31619) );
  AND U1699 ( .A(n30335), .B(n30859), .Z(n31639) );
  AND U1700 ( .A(n29011), .B(n26159), .Z(n32358) );
  AND U1701 ( .A(n27245), .B(n27246), .Z(n30195) );
  AND U1702 ( .A(n29702), .B(n28312), .Z(n34531) );
  ANDN U1703 ( .B(n28221), .A(n29160), .Z(n30669) );
  ANDN U1704 ( .B(n25846), .A(n25847), .Z(n29914) );
  ANDN U1705 ( .B(n27474), .A(n27475), .Z(n29314) );
  XOR U1706 ( .A(n27994), .B(n27995), .Z(n26284) );
  AND U1707 ( .A(n29513), .B(n28285), .Z(n30102) );
  ANDN U1708 ( .B(n28046), .A(n27371), .Z(n28044) );
  ANDN U1709 ( .B(n29723), .A(n27079), .Z(n30065) );
  ANDN U1710 ( .B(n27231), .A(n27232), .Z(n27229) );
  XOR U1711 ( .A(n30985), .B(n28109), .Z(n24518) );
  AND U1712 ( .A(n28106), .B(n30994), .Z(n30992) );
  XNOR U1713 ( .A(n28714), .B(n28713), .Z(n23250) );
  XOR U1714 ( .A(n25513), .B(n28291), .Z(n25356) );
  AND U1715 ( .A(n27536), .B(n27537), .Z(n27534) );
  AND U1716 ( .A(n28922), .B(n29276), .Z(n29274) );
  XNOR U1717 ( .A(n26258), .B(n26257), .Z(n26053) );
  AND U1718 ( .A(n26946), .B(n27650), .Z(n36859) );
  XNOR U1719 ( .A(n26409), .B(n26408), .Z(n23253) );
  XNOR U1720 ( .A(n26880), .B(n26879), .Z(n24943) );
  XNOR U1721 ( .A(n26792), .B(n26791), .Z(n23015) );
  AND U1722 ( .A(n30588), .B(n30585), .Z(n31040) );
  XNOR U1723 ( .A(n26764), .B(n26763), .Z(n23864) );
  XNOR U1724 ( .A(n25710), .B(n26484), .Z(n24154) );
  XOR U1725 ( .A(n26712), .B(n26711), .Z(n22809) );
  XNOR U1726 ( .A(n26507), .B(n26506), .Z(n21221) );
  XOR U1727 ( .A(n26769), .B(n29013), .Z(n24930) );
  XNOR U1728 ( .A(n27202), .B(n27778), .Z(n25170) );
  XOR U1729 ( .A(n26056), .B(n29705), .Z(n24899) );
  XNOR U1730 ( .A(n25727), .B(n25726), .Z(n22342) );
  XNOR U1731 ( .A(n32316), .B(n29134), .Z(n25706) );
  XNOR U1732 ( .A(n27580), .B(n27579), .Z(n23024) );
  XNOR U1733 ( .A(n25581), .B(n25580), .Z(n21593) );
  XNOR U1734 ( .A(n27031), .B(n26377), .Z(n24745) );
  XNOR U1735 ( .A(n25476), .B(n25475), .Z(n21983) );
  XNOR U1736 ( .A(n28289), .B(n25361), .Z(n22450) );
  XOR U1737 ( .A(n26521), .B(n23978), .Z(n22301) );
  XNOR U1738 ( .A(n25168), .B(n23602), .Z(n24155) );
  XNOR U1739 ( .A(n23592), .B(n24805), .Z(n20580) );
  XNOR U1740 ( .A(n22223), .B(n22222), .Z(n20689) );
  XOR U1741 ( .A(n23505), .B(n23850), .Z(n21285) );
  AND U1742 ( .A(n20437), .B(n22896), .Z(n22894) );
  ANDN U1743 ( .B(n20590), .A(n21612), .Z(n21611) );
  AND U1744 ( .A(n20023), .B(n20024), .Z(n20021) );
  ANDN U1745 ( .B(n23173), .A(n23171), .Z(n30284) );
  NOR U1746 ( .A(n21655), .B(n21654), .Z(n24456) );
  AND U1747 ( .A(n20617), .B(n21810), .Z(n24495) );
  AND U1748 ( .A(n20410), .B(n19160), .Z(n21379) );
  AND U1749 ( .A(n23921), .B(n21403), .Z(n24168) );
  AND U1750 ( .A(n20351), .B(n21412), .Z(n25508) );
  AND U1751 ( .A(n22083), .B(n19571), .Z(n25097) );
  AND U1752 ( .A(n20541), .B(n21360), .Z(n21359) );
  ANDN U1753 ( .B(n22291), .A(n24113), .Z(n24111) );
  XOR U1754 ( .A(n20370), .B(n20163), .Z(n16464) );
  AND U1755 ( .A(n22908), .B(n22909), .Z(n22907) );
  AND U1756 ( .A(n23471), .B(n23668), .Z(n32831) );
  AND U1757 ( .A(n21542), .B(n21540), .Z(n23939) );
  XOR U1758 ( .A(n24790), .B(n22040), .Z(n18632) );
  XOR U1759 ( .A(n22814), .B(n20119), .Z(n16663) );
  ANDN U1760 ( .B(n18912), .A(n18911), .Z(n18909) );
  AND U1761 ( .A(n27903), .B(n19627), .Z(n31756) );
  AND U1762 ( .A(n21569), .B(n21570), .Z(n21567) );
  XNOR U1763 ( .A(n25285), .B(n24664), .Z(n20130) );
  AND U1764 ( .A(n23532), .B(n23530), .Z(n27304) );
  AND U1765 ( .A(n20232), .B(n20230), .Z(n23496) );
  AND U1766 ( .A(n23225), .B(n25135), .Z(n33465) );
  AND U1767 ( .A(n22055), .B(n22056), .Z(n23487) );
  AND U1768 ( .A(n19567), .B(n19569), .Z(n19686) );
  XNOR U1769 ( .A(n23520), .B(n18977), .Z(n15879) );
  AND U1770 ( .A(n24876), .B(n24878), .Z(n30508) );
  AND U1771 ( .A(n21677), .B(n22109), .Z(n29657) );
  AND U1772 ( .A(n20945), .B(n20944), .Z(n25945) );
  AND U1773 ( .A(n19165), .B(n26345), .Z(n26343) );
  AND U1774 ( .A(n21699), .B(n21418), .Z(n21698) );
  XOR U1775 ( .A(n25667), .B(n20457), .Z(n19297) );
  AND U1776 ( .A(n21761), .B(n21762), .Z(n21759) );
  ANDN U1777 ( .B(n22844), .A(n22843), .Z(n22841) );
  XOR U1778 ( .A(n19419), .B(n18264), .Z(n14970) );
  ANDN U1779 ( .B(n19933), .A(n19932), .Z(n19930) );
  XNOR U1780 ( .A(n20481), .B(n20480), .Z(n17589) );
  AND U1781 ( .A(n19939), .B(n19941), .Z(n20834) );
  XOR U1782 ( .A(n18461), .B(n18460), .Z(n16154) );
  AND U1783 ( .A(n21924), .B(n21923), .Z(n29252) );
  AND U1784 ( .A(n23167), .B(n23297), .Z(n24872) );
  XOR U1785 ( .A(n20414), .B(n20415), .Z(n19370) );
  XNOR U1786 ( .A(n20664), .B(n20663), .Z(n16757) );
  XNOR U1787 ( .A(n18926), .B(n18925), .Z(n16892) );
  XNOR U1788 ( .A(n19653), .B(n20277), .Z(n17009) );
  XOR U1789 ( .A(n20989), .B(n20988), .Z(n16813) );
  XNOR U1790 ( .A(n21256), .B(n20884), .Z(n15694) );
  XNOR U1791 ( .A(n19712), .B(n19711), .Z(n16068) );
  XNOR U1792 ( .A(n19336), .B(n20910), .Z(n18090) );
  XNOR U1793 ( .A(n20153), .B(n20703), .Z(n17140) );
  XNOR U1794 ( .A(n16036), .B(n19791), .Z(n13817) );
  XNOR U1795 ( .A(n17228), .B(n17229), .Z(n13564) );
  XNOR U1796 ( .A(n16877), .B(n16878), .Z(n14791) );
  XOR U1797 ( .A(n17940), .B(n16930), .Z(n12293) );
  XOR U1798 ( .A(n16322), .B(n15555), .Z(n10286) );
  XOR U1799 ( .A(n15696), .B(n14973), .Z(n12914) );
  ANDN U1800 ( .B(n17424), .A(n16435), .Z(n16432) );
  AND U1801 ( .A(n15003), .B(n15005), .Z(n16354) );
  AND U1802 ( .A(n16351), .B(n17353), .Z(n17352) );
  ANDN U1803 ( .B(n14484), .A(n14485), .Z(n15035) );
  ANDN U1804 ( .B(n15065), .A(n15064), .Z(n15062) );
  AND U1805 ( .A(n12835), .B(n12833), .Z(n14940) );
  AND U1806 ( .A(n14339), .B(n13606), .Z(n14337) );
  AND U1807 ( .A(n15398), .B(n19008), .Z(n19006) );
  XOR U1808 ( .A(n18689), .B(n18690), .Z(n13928) );
  AND U1809 ( .A(n15214), .B(n15216), .Z(n18443) );
  XOR U1810 ( .A(n13952), .B(n13142), .Z(n12284) );
  AND U1811 ( .A(n13365), .B(n15297), .Z(n17201) );
  AND U1812 ( .A(n15576), .B(n15577), .Z(n15574) );
  ANDN U1813 ( .B(n15515), .A(n15514), .Z(n15512) );
  ANDN U1814 ( .B(n14375), .A(n13105), .Z(n14373) );
  XOR U1815 ( .A(n15450), .B(n14242), .Z(n15280) );
  XNOR U1816 ( .A(n12836), .B(n11949), .Z(n11711) );
  ANDN U1817 ( .B(n14969), .A(n13179), .Z(n21346) );
  XOR U1818 ( .A(n17761), .B(n17384), .Z(n14651) );
  ANDN U1819 ( .B(n14087), .A(n14085), .Z(n19385) );
  ANDN U1820 ( .B(n13860), .A(n13859), .Z(n13857) );
  ANDN U1821 ( .B(n13775), .A(n14578), .Z(n14576) );
  ANDN U1822 ( .B(n14425), .A(n14424), .Z(n14422) );
  AND U1823 ( .A(n13900), .B(n13901), .Z(n15433) );
  XOR U1824 ( .A(n18142), .B(n15014), .Z(n12437) );
  XOR U1825 ( .A(n19206), .B(n12474), .Z(n15204) );
  XNOR U1826 ( .A(n17727), .B(n14692), .Z(n9450) );
  XOR U1827 ( .A(n17697), .B(n14548), .Z(n11819) );
  XNOR U1828 ( .A(n18484), .B(n16969), .Z(n10690) );
  AND U1829 ( .A(n16142), .B(n14557), .Z(n16141) );
  XNOR U1830 ( .A(n13296), .B(n13295), .Z(n12299) );
  AND U1831 ( .A(n16686), .B(n16687), .Z(n16685) );
  XOR U1832 ( .A(n18372), .B(n13255), .Z(n14153) );
  XNOR U1833 ( .A(n15730), .B(n11568), .Z(n9028) );
  XNOR U1834 ( .A(n12559), .B(n9142), .Z(n8948) );
  XNOR U1835 ( .A(n11810), .B(n11733), .Z(n9742) );
  XOR U1836 ( .A(n12310), .B(n11340), .Z(n8574) );
  XOR U1837 ( .A(n7294), .B(n6729), .Z(n4918) );
  XOR U1838 ( .A(n7919), .B(n7920), .Z(n4952) );
  ANDN U1839 ( .B(n9059), .A(n8984), .Z(n9058) );
  XOR U1840 ( .A(n8825), .B(n8826), .Z(n5300) );
  AND U1841 ( .A(n9998), .B(n9997), .Z(n11035) );
  AND U1842 ( .A(n8583), .B(n6441), .Z(n8581) );
  AND U1843 ( .A(n8008), .B(n8007), .Z(n8005) );
  AND U1844 ( .A(n6929), .B(n6930), .Z(n7718) );
  ANDN U1845 ( .B(n6703), .A(n6702), .Z(n6700) );
  AND U1846 ( .A(n7629), .B(n7630), .Z(n7627) );
  ANDN U1847 ( .B(n10046), .A(n7993), .Z(n10170) );
  ANDN U1848 ( .B(n10227), .A(n7969), .Z(n10355) );
  ANDN U1849 ( .B(n10881), .A(n8152), .Z(n10999) );
  XNOR U1850 ( .A(n6352), .B(n6530), .Z(n4293) );
  AND U1851 ( .A(n7790), .B(n10416), .Z(n10560) );
  AND U1852 ( .A(n8489), .B(n11995), .Z(n12148) );
  XOR U1853 ( .A(n11636), .B(n8554), .Z(n8530) );
  ANDN U1854 ( .B(n7903), .A(n7904), .Z(n8981) );
  AND U1855 ( .A(n11542), .B(n9606), .Z(n11540) );
  ANDN U1856 ( .B(n11152), .A(n9285), .Z(n11150) );
  ANDN U1857 ( .B(n6897), .A(n6896), .Z(n6894) );
  AND U1858 ( .A(n8907), .B(n8828), .Z(n8906) );
  AND U1859 ( .A(n9005), .B(n8957), .Z(n9004) );
  AND U1860 ( .A(n6817), .B(n6818), .Z(n6815) );
  AND U1861 ( .A(n8755), .B(n6465), .Z(n8754) );
  AND U1862 ( .A(n8113), .B(n8114), .Z(n8112) );
  XNOR U1863 ( .A(n7527), .B(n6243), .Z(n3444) );
  AND U1864 ( .A(n7083), .B(n7084), .Z(n7081) );
  ANDN U1865 ( .B(n10028), .A(n7598), .Z(n10026) );
  XNOR U1866 ( .A(n6224), .B(n8179), .Z(n1969) );
  XOR U1867 ( .A(n10960), .B(n9400), .Z(n3778) );
  AND U1868 ( .A(n7253), .B(n7254), .Z(n7251) );
  ANDN U1869 ( .B(n7896), .A(n7895), .Z(n7893) );
  XNOR U1870 ( .A(n6059), .B(n6058), .Z(n3843) );
  AND U1871 ( .A(n7615), .B(n7617), .Z(n8727) );
  XOR U1872 ( .A(n11681), .B(n11682), .Z(n3911) );
  AND U1873 ( .A(n8071), .B(n8070), .Z(n9180) );
  AND U1874 ( .A(n7544), .B(n7545), .Z(n7542) );
  ANDN U1875 ( .B(n8912), .A(n8913), .Z(n11553) );
  XNOR U1876 ( .A(n6239), .B(n8287), .Z(n1662) );
  XNOR U1877 ( .A(n3668), .B(n2438), .Z(n2742) );
  XNOR U1878 ( .A(n2339), .B(n9371), .Z(n3587) );
  AND U1879 ( .A(n4509), .B(n4510), .Z(n4507) );
  AND U1880 ( .A(n4513), .B(n4514), .Z(n4511) );
  ANDN U1881 ( .B(n4633), .A(n4634), .Z(n4631) );
  AND U1882 ( .A(n4669), .B(n4670), .Z(n4667) );
  ANDN U1883 ( .B(n4727), .A(n4461), .Z(n4726) );
  AND U1884 ( .A(n4486), .B(n4743), .Z(n4742) );
  AND U1885 ( .A(n4541), .B(n4773), .Z(n4772) );
  AND U1886 ( .A(n4731), .B(n4922), .Z(n4920) );
  ANDN U1887 ( .B(n5009), .A(n4799), .Z(n5007) );
  AND U1888 ( .A(n5026), .B(n4807), .Z(n5024) );
  AND U1889 ( .A(n4813), .B(n5035), .Z(n5033) );
  AND U1890 ( .A(n4929), .B(n4476), .Z(n5148) );
  AND U1891 ( .A(n5622), .B(n5621), .Z(n5619) );
  AND U1892 ( .A(n5714), .B(n5893), .Z(n5889) );
  ANDN U1893 ( .B(n5989), .A(n1111), .Z(n6315) );
  ANDN U1894 ( .B(n1155), .A(n6044), .Z(n6363) );
  XOR U1895 ( .A(n1282), .B(n1283), .Z(out[943]) );
  AND U1896 ( .A(n1336), .B(n1337), .Z(n1334) );
  NOR U1897 ( .A(n1361), .B(n1360), .Z(n1358) );
  AND U1898 ( .A(n1532), .B(n1273), .Z(n1531) );
  AND U1899 ( .A(n1609), .B(n1405), .Z(n1608) );
  AND U1900 ( .A(n1659), .B(n1497), .Z(n1658) );
  NOR U1901 ( .A(n1668), .B(n1502), .Z(n1665) );
  AND U1902 ( .A(n1768), .B(n1554), .Z(n1765) );
  AND U1903 ( .A(n1852), .B(n1597), .Z(n1849) );
  ANDN U1904 ( .B(n2758), .A(n2757), .Z(n2755) );
  ANDN U1905 ( .B(n2790), .A(n2789), .Z(n2787) );
  ANDN U1906 ( .B(n3183), .A(n2732), .Z(n3437) );
  XNOR U1907 ( .A(n52278), .B(n52277), .Z(n51448) );
  XNOR U1908 ( .A(n51916), .B(n52606), .Z(n51595) );
  XNOR U1909 ( .A(n52286), .B(n52285), .Z(n51462) );
  XNOR U1910 ( .A(n51952), .B(n51951), .Z(n51710) );
  XNOR U1911 ( .A(n51692), .B(n52105), .Z(n51243) );
  XNOR U1912 ( .A(n51922), .B(n51921), .Z(n49427) );
  XOR U1913 ( .A(n51925), .B(n51924), .Z(n51141) );
  XNOR U1914 ( .A(n51681), .B(n51680), .Z(n48566) );
  XNOR U1915 ( .A(n52535), .B(n52458), .Z(n52176) );
  XNOR U1916 ( .A(n51938), .B(n52519), .Z(n50741) );
  XNOR U1917 ( .A(n52423), .B(n52450), .Z(n48879) );
  XNOR U1918 ( .A(n53262), .B(n51659), .Z(n48445) );
  XNOR U1919 ( .A(n51764), .B(n51763), .Z(n49901) );
  XNOR U1920 ( .A(n52430), .B(n52429), .Z(n51464) );
  XNOR U1921 ( .A(n52825), .B(n52363), .Z(n50745) );
  XNOR U1922 ( .A(n52133), .B(n52132), .Z(n50744) );
  XNOR U1923 ( .A(n53104), .B(n52422), .Z(n49857) );
  XNOR U1924 ( .A(n52766), .B(n52603), .Z(n51579) );
  XNOR U1925 ( .A(n52729), .B(n53298), .Z(n48365) );
  XNOR U1926 ( .A(n51830), .B(n52676), .Z(n52313) );
  XNOR U1927 ( .A(n52662), .B(n52627), .Z(n50136) );
  XNOR U1928 ( .A(n52650), .B(n52810), .Z(n51567) );
  XOR U1929 ( .A(n52126), .B(n51945), .Z(n50738) );
  XNOR U1930 ( .A(round_reg[481]), .B(n49175), .Z(n49407) );
  XOR U1931 ( .A(round_reg[251]), .B(n49080), .Z(n46869) );
  XNOR U1932 ( .A(round_reg[1164]), .B(n51140), .Z(n50279) );
  XNOR U1933 ( .A(round_reg[478]), .B(n50650), .Z(n48543) );
  XOR U1934 ( .A(round_reg[804]), .B(n48449), .Z(n46958) );
  XNOR U1935 ( .A(round_reg[50]), .B(n50404), .Z(n48753) );
  XNOR U1936 ( .A(round_reg[125]), .B(n50949), .Z(n48149) );
  XNOR U1937 ( .A(round_reg[763]), .B(n50984), .Z(n47430) );
  XNOR U1938 ( .A(round_reg[159]), .B(n52025), .Z(n51376) );
  AND U1939 ( .A(n48025), .B(n47155), .Z(n50477) );
  AND U1940 ( .A(n47349), .B(n48562), .Z(n48567) );
  ANDN U1941 ( .B(n48161), .A(n51370), .Z(n51657) );
  ANDN U1942 ( .B(n46613), .A(n46612), .Z(n46610) );
  AND U1943 ( .A(n47497), .B(n47498), .Z(n47495) );
  AND U1944 ( .A(n48904), .B(n48905), .Z(n51382) );
  ANDN U1945 ( .B(n48240), .A(n48241), .Z(n51360) );
  ANDN U1946 ( .B(n47421), .A(n48620), .Z(n52537) );
  ANDN U1947 ( .B(n48937), .A(n48431), .Z(n51173) );
  XNOR U1948 ( .A(n47526), .B(n50245), .Z(n46940) );
  ANDN U1949 ( .B(n50679), .A(n50678), .Z(n50676) );
  ANDN U1950 ( .B(n47947), .A(n47946), .Z(n47944) );
  AND U1951 ( .A(n49909), .B(n49910), .Z(n52320) );
  AND U1952 ( .A(n49755), .B(n49754), .Z(n50893) );
  ANDN U1953 ( .B(n47088), .A(n47089), .Z(n47346) );
  AND U1954 ( .A(n50799), .B(n50800), .Z(n50797) );
  XNOR U1955 ( .A(n46884), .B(n46883), .Z(n45514) );
  AND U1956 ( .A(n47727), .B(n47728), .Z(n47725) );
  ANDN U1957 ( .B(n50205), .A(n50204), .Z(n50202) );
  AND U1958 ( .A(n49481), .B(n48731), .Z(n50242) );
  XOR U1959 ( .A(n48243), .B(n47126), .Z(n46176) );
  ANDN U1960 ( .B(n48300), .A(n48298), .Z(n49244) );
  XNOR U1961 ( .A(n47580), .B(n48107), .Z(n45247) );
  XNOR U1962 ( .A(n47244), .B(n47243), .Z(n43765) );
  ANDN U1963 ( .B(n48497), .A(n48498), .Z(n51015) );
  XNOR U1964 ( .A(n49326), .B(n50197), .Z(n46877) );
  AND U1965 ( .A(n48293), .B(n48294), .Z(n48291) );
  XNOR U1966 ( .A(n47683), .B(n47682), .Z(n43102) );
  AND U1967 ( .A(n50069), .B(n50063), .Z(n50068) );
  XNOR U1968 ( .A(n46273), .B(n47694), .Z(n43767) );
  XNOR U1969 ( .A(n46684), .B(n48987), .Z(n48548) );
  AND U1970 ( .A(n49842), .B(n49933), .Z(n49932) );
  AND U1971 ( .A(n50601), .B(n50602), .Z(n50600) );
  ANDN U1972 ( .B(n47289), .A(n47290), .Z(n49799) );
  ANDN U1973 ( .B(n47824), .A(n47823), .Z(n47821) );
  XNOR U1974 ( .A(n48194), .B(n48193), .Z(n43088) );
  XNOR U1975 ( .A(n47476), .B(n47475), .Z(n45080) );
  XNOR U1976 ( .A(n49783), .B(n46850), .Z(n44410) );
  XNOR U1977 ( .A(n49536), .B(n49535), .Z(n45861) );
  ANDN U1978 ( .B(n48531), .A(n48530), .Z(n48528) );
  ANDN U1979 ( .B(n51581), .A(n50464), .Z(n52695) );
  AND U1980 ( .A(n49710), .B(n49709), .Z(n49708) );
  ANDN U1981 ( .B(n47776), .A(n47777), .Z(n49613) );
  XOR U1982 ( .A(n49438), .B(n47454), .Z(n41883) );
  ANDN U1983 ( .B(n46490), .A(n46489), .Z(n46487) );
  ANDN U1984 ( .B(n50094), .A(n50223), .Z(n52295) );
  AND U1985 ( .A(n46972), .B(n47967), .Z(n48451) );
  XOR U1986 ( .A(n49441), .B(n49352), .Z(n43925) );
  XNOR U1987 ( .A(n45428), .B(n45427), .Z(n40853) );
  XNOR U1988 ( .A(n47094), .B(n46191), .Z(n45279) );
  AND U1989 ( .A(n48097), .B(n48919), .Z(n48918) );
  XNOR U1990 ( .A(n51746), .B(n50588), .Z(n45953) );
  ANDN U1991 ( .B(n47364), .A(n47365), .Z(n50496) );
  XNOR U1992 ( .A(n48245), .B(n50570), .Z(n42301) );
  XOR U1993 ( .A(n47414), .B(n48320), .Z(n44743) );
  XNOR U1994 ( .A(n50763), .B(n48265), .Z(n45085) );
  XOR U1995 ( .A(n46595), .B(n48494), .Z(n43916) );
  ANDN U1996 ( .B(n49965), .A(n49966), .Z(n51856) );
  XNOR U1997 ( .A(n48773), .B(n48311), .Z(n44191) );
  XNOR U1998 ( .A(n49624), .B(n46328), .Z(n46936) );
  AND U1999 ( .A(n48873), .B(n48178), .Z(n48871) );
  AND U2000 ( .A(n49282), .B(n49150), .Z(n52562) );
  ANDN U2001 ( .B(n48671), .A(n49660), .Z(n49659) );
  XNOR U2002 ( .A(n50491), .B(n48005), .Z(n47266) );
  XNOR U2003 ( .A(n46641), .B(n42498), .Z(n42836) );
  XNOR U2004 ( .A(n45663), .B(n45664), .Z(n40154) );
  XNOR U2005 ( .A(n43573), .B(n43574), .Z(n41620) );
  XNOR U2006 ( .A(n42395), .B(n47331), .Z(n42263) );
  XNOR U2007 ( .A(n46341), .B(n42513), .Z(n42136) );
  XOR U2008 ( .A(n42510), .B(n45131), .Z(n43435) );
  XNOR U2009 ( .A(n44549), .B(n44550), .Z(n43982) );
  XNOR U2010 ( .A(n45145), .B(n49726), .Z(n41340) );
  XNOR U2011 ( .A(n45849), .B(n45453), .Z(n41334) );
  XOR U2012 ( .A(n47063), .B(n44523), .Z(n40587) );
  AND U2013 ( .A(n43265), .B(n43266), .Z(n43264) );
  ANDN U2014 ( .B(n40702), .A(n40701), .Z(n40699) );
  NOR U2015 ( .A(n43180), .B(n45207), .Z(n47384) );
  XNOR U2016 ( .A(n43367), .B(n42937), .Z(n41917) );
  ANDN U2017 ( .B(n41869), .A(n41868), .Z(n41866) );
  AND U2018 ( .A(n41545), .B(n41544), .Z(n45650) );
  ANDN U2019 ( .B(n40644), .A(n46397), .Z(n46396) );
  AND U2020 ( .A(n40748), .B(n40749), .Z(n40746) );
  AND U2021 ( .A(n40121), .B(n40122), .Z(n40119) );
  AND U2022 ( .A(n43158), .B(n43159), .Z(n43157) );
  ANDN U2023 ( .B(n44059), .A(n44060), .Z(n44891) );
  ANDN U2024 ( .B(n42410), .A(n40722), .Z(n44900) );
  AND U2025 ( .A(n40456), .B(n40457), .Z(n40454) );
  XOR U2026 ( .A(n41242), .B(n39915), .Z(n38458) );
  XNOR U2027 ( .A(n40534), .B(n39799), .Z(n39454) );
  XOR U2028 ( .A(n44977), .B(n42994), .Z(n37173) );
  AND U2029 ( .A(n41177), .B(n43927), .Z(n45139) );
  AND U2030 ( .A(n42439), .B(n42438), .Z(n42436) );
  XNOR U2031 ( .A(n44080), .B(n42005), .Z(n39219) );
  XNOR U2032 ( .A(n42551), .B(n41077), .Z(n36413) );
  ANDN U2033 ( .B(n42479), .A(n42478), .Z(n42477) );
  XNOR U2034 ( .A(n40419), .B(n40420), .Z(n38963) );
  XOR U2035 ( .A(n43668), .B(n43669), .Z(n39266) );
  XNOR U2036 ( .A(n40086), .B(n39841), .Z(n37071) );
  AND U2037 ( .A(n41497), .B(n41498), .Z(n41495) );
  ANDN U2038 ( .B(n44097), .A(n41404), .Z(n44249) );
  ANDN U2039 ( .B(n41144), .A(n43727), .Z(n43726) );
  XOR U2040 ( .A(n40127), .B(n40301), .Z(n37219) );
  XNOR U2041 ( .A(n40374), .B(n40373), .Z(n35632) );
  AND U2042 ( .A(n42941), .B(n42942), .Z(n42939) );
  ANDN U2043 ( .B(n40751), .A(n40752), .Z(n43558) );
  ANDN U2044 ( .B(n41647), .A(n41028), .Z(n42657) );
  AND U2045 ( .A(n43660), .B(n42705), .Z(n46667) );
  AND U2046 ( .A(n43696), .B(n43850), .Z(n45201) );
  AND U2047 ( .A(n41349), .B(n41351), .Z(n45043) );
  AND U2048 ( .A(n42274), .B(n42273), .Z(n45088) );
  XOR U2049 ( .A(n46751), .B(n41192), .Z(n40347) );
  ANDN U2050 ( .B(n39512), .A(n39513), .Z(n43993) );
  XOR U2051 ( .A(n40906), .B(n40905), .Z(n38912) );
  AND U2052 ( .A(n45136), .B(n44394), .Z(n45133) );
  ANDN U2053 ( .B(n39568), .A(n41787), .Z(n41786) );
  XNOR U2054 ( .A(n41490), .B(n39362), .Z(n37707) );
  XOR U2055 ( .A(n38690), .B(n38689), .Z(n36423) );
  ANDN U2056 ( .B(n40242), .A(n40241), .Z(n40239) );
  ANDN U2057 ( .B(n41828), .A(n43526), .Z(n43525) );
  AND U2058 ( .A(n41434), .B(n40169), .Z(n41433) );
  AND U2059 ( .A(n39955), .B(n45918), .Z(n47582) );
  XOR U2060 ( .A(n45607), .B(n43805), .Z(n39282) );
  XNOR U2061 ( .A(n41984), .B(n41213), .Z(n39242) );
  XNOR U2062 ( .A(n41997), .B(n41996), .Z(n37051) );
  AND U2063 ( .A(n41258), .B(n44170), .Z(n44168) );
  XOR U2064 ( .A(n44944), .B(n41141), .Z(n39389) );
  XNOR U2065 ( .A(n42886), .B(n42693), .Z(n38486) );
  AND U2066 ( .A(n40599), .B(n40600), .Z(n40597) );
  XOR U2067 ( .A(n38449), .B(n42055), .Z(n35929) );
  ANDN U2068 ( .B(n41781), .A(n41780), .Z(n41778) );
  XOR U2069 ( .A(n44446), .B(n44447), .Z(n39849) );
  AND U2070 ( .A(n41247), .B(n39897), .Z(n45638) );
  XOR U2071 ( .A(n43626), .B(n40661), .Z(n38113) );
  AND U2072 ( .A(n39196), .B(n39197), .Z(n39194) );
  XNOR U2073 ( .A(n39818), .B(n42575), .Z(n39011) );
  XOR U2074 ( .A(n46306), .B(n43741), .Z(n42947) );
  XNOR U2075 ( .A(n45837), .B(n41323), .Z(n38620) );
  AND U2076 ( .A(n40185), .B(n40183), .Z(n43317) );
  ANDN U2077 ( .B(n41012), .A(n42980), .Z(n42979) );
  ANDN U2078 ( .B(n41124), .A(n42271), .Z(n42269) );
  XOR U2079 ( .A(n38624), .B(n40542), .Z(n35630) );
  XNOR U2080 ( .A(n39356), .B(n39355), .Z(n35619) );
  AND U2081 ( .A(n42782), .B(n44006), .Z(n45411) );
  XOR U2082 ( .A(n36211), .B(n36212), .Z(n33661) );
  XNOR U2083 ( .A(n45675), .B(n35611), .Z(n37989) );
  XNOR U2084 ( .A(n39324), .B(n37328), .Z(n35357) );
  XNOR U2085 ( .A(n34618), .B(n35591), .Z(n33314) );
  XOR U2086 ( .A(n34638), .B(n39010), .Z(n36565) );
  XOR U2087 ( .A(n34628), .B(n39239), .Z(n33694) );
  XNOR U2088 ( .A(n40996), .B(n37890), .Z(n37207) );
  XOR U2089 ( .A(n37330), .B(n37331), .Z(n35706) );
  AND U2090 ( .A(n34556), .B(n34557), .Z(n39148) );
  AND U2091 ( .A(n34385), .B(n34416), .Z(n34414) );
  NOR U2092 ( .A(n33681), .B(n33680), .Z(n37004) );
  AND U2093 ( .A(n37456), .B(n37360), .Z(n37638) );
  AND U2094 ( .A(n33391), .B(n33392), .Z(n38638) );
  ANDN U2095 ( .B(n33248), .A(n37594), .Z(n39065) );
  AND U2096 ( .A(n35912), .B(n35913), .Z(n35910) );
  AND U2097 ( .A(n34923), .B(n34921), .Z(n36684) );
  AND U2098 ( .A(n36986), .B(n35961), .Z(n37628) );
  AND U2099 ( .A(n36883), .B(n36881), .Z(n42813) );
  AND U2100 ( .A(n35063), .B(n35064), .Z(n35061) );
  XNOR U2101 ( .A(n34591), .B(n34592), .Z(n32378) );
  AND U2102 ( .A(n34653), .B(n34654), .Z(n34651) );
  AND U2103 ( .A(n34947), .B(n37442), .Z(n37441) );
  ANDN U2104 ( .B(n36385), .A(n34876), .Z(n39792) );
  XNOR U2105 ( .A(n33477), .B(n33476), .Z(n32064) );
  NOR U2106 ( .A(n34917), .B(n36687), .Z(n42002) );
  XNOR U2107 ( .A(n38752), .B(n36845), .Z(n36138) );
  XNOR U2108 ( .A(n37119), .B(n34734), .Z(n32836) );
  XNOR U2109 ( .A(n39581), .B(n33082), .Z(n30266) );
  ANDN U2110 ( .B(n37571), .A(n35726), .Z(n37569) );
  XOR U2111 ( .A(n38778), .B(n34962), .Z(n33238) );
  AND U2112 ( .A(n37280), .B(n36072), .Z(n39293) );
  AND U2113 ( .A(n33652), .B(n33653), .Z(n33650) );
  XNOR U2114 ( .A(n38386), .B(n38387), .Z(n30038) );
  XNOR U2115 ( .A(n33487), .B(n33486), .Z(n30125) );
  AND U2116 ( .A(n33111), .B(n33112), .Z(n33109) );
  XOR U2117 ( .A(n33718), .B(n33717), .Z(n30215) );
  XNOR U2118 ( .A(n38251), .B(n34589), .Z(n30519) );
  XNOR U2119 ( .A(n32970), .B(n33493), .Z(n28825) );
  AND U2120 ( .A(n33989), .B(n34266), .Z(n36360) );
  AND U2121 ( .A(n36472), .B(n36871), .Z(n36869) );
  AND U2122 ( .A(n35153), .B(n34694), .Z(n37507) );
  ANDN U2123 ( .B(n35839), .A(n36007), .Z(n36418) );
  XNOR U2124 ( .A(n37829), .B(n37828), .Z(n31001) );
  XNOR U2125 ( .A(n32636), .B(n32637), .Z(n32427) );
  XNOR U2126 ( .A(n35871), .B(n37771), .Z(n31539) );
  ANDN U2127 ( .B(n38414), .A(n36753), .Z(n42465) );
  ANDN U2128 ( .B(n34239), .A(n34238), .Z(n34236) );
  AND U2129 ( .A(n35135), .B(n35134), .Z(n37539) );
  ANDN U2130 ( .B(n38709), .A(n38390), .Z(n40048) );
  AND U2131 ( .A(n33970), .B(n33971), .Z(n33968) );
  XNOR U2132 ( .A(n33365), .B(n33364), .Z(n29736) );
  AND U2133 ( .A(n35438), .B(n34982), .Z(n35436) );
  ANDN U2134 ( .B(n37556), .A(n37555), .Z(n37553) );
  ANDN U2135 ( .B(n36102), .A(n36101), .Z(n36099) );
  XNOR U2136 ( .A(n33244), .B(n34213), .Z(n31579) );
  XNOR U2137 ( .A(n32257), .B(n32256), .Z(n28887) );
  XNOR U2138 ( .A(n36500), .B(n33049), .Z(n31159) );
  AND U2139 ( .A(n40062), .B(n37985), .Z(n40275) );
  AND U2140 ( .A(n34780), .B(n34779), .Z(n35496) );
  ANDN U2141 ( .B(n37286), .A(n37285), .Z(n37283) );
  AND U2142 ( .A(n37915), .B(n35291), .Z(n40341) );
  AND U2143 ( .A(n36066), .B(n36484), .Z(n36482) );
  ANDN U2144 ( .B(n36064), .A(n36494), .Z(n38346) );
  AND U2145 ( .A(n34757), .B(n34756), .Z(n38905) );
  XNOR U2146 ( .A(n35353), .B(n33960), .Z(n29166) );
  AND U2147 ( .A(n34173), .B(n34172), .Z(n35100) );
  ANDN U2148 ( .B(n36021), .A(n34513), .Z(n36019) );
  XNOR U2149 ( .A(n35949), .B(n34138), .Z(n31440) );
  XOR U2150 ( .A(n32373), .B(n33604), .Z(n32053) );
  XNOR U2151 ( .A(n33742), .B(n32754), .Z(n32101) );
  XOR U2152 ( .A(n35501), .B(n36216), .Z(n31834) );
  ANDN U2153 ( .B(n34245), .A(n34246), .Z(n36271) );
  AND U2154 ( .A(n34208), .B(n35432), .Z(n46363) );
  XOR U2155 ( .A(n32742), .B(n33386), .Z(n30784) );
  XOR U2156 ( .A(n38323), .B(n34179), .Z(n30959) );
  AND U2157 ( .A(n35219), .B(n35220), .Z(n35218) );
  ANDN U2158 ( .B(n35186), .A(n37251), .Z(n38931) );
  XNOR U2159 ( .A(n37212), .B(n27947), .Z(n27531) );
  XNOR U2160 ( .A(n31137), .B(n31913), .Z(n31898) );
  XNOR U2161 ( .A(n35394), .B(n32402), .Z(n28475) );
  XNOR U2162 ( .A(n32922), .B(n32585), .Z(n28645) );
  XNOR U2163 ( .A(n32762), .B(n30491), .Z(n31086) );
  XNOR U2164 ( .A(n30066), .B(n33445), .Z(n30088) );
  XNOR U2165 ( .A(n30207), .B(n30208), .Z(n27330) );
  XOR U2166 ( .A(n30781), .B(n31832), .Z(n29233) );
  XNOR U2167 ( .A(n30864), .B(n30865), .Z(n30328) );
  XNOR U2168 ( .A(n31824), .B(n31068), .Z(n29878) );
  ANDN U2169 ( .B(n27866), .A(n27865), .Z(n27864) );
  XNOR U2170 ( .A(n32013), .B(n28690), .Z(n29129) );
  AND U2171 ( .A(n27089), .B(n27090), .Z(n27087) );
  AND U2172 ( .A(n28942), .B(n28943), .Z(n28940) );
  AND U2173 ( .A(n28165), .B(n28167), .Z(n28448) );
  XNOR U2174 ( .A(n26264), .B(n26263), .Z(n25252) );
  ANDN U2175 ( .B(n26604), .A(n28737), .Z(n28734) );
  XOR U2176 ( .A(n29580), .B(n29581), .Z(n28901) );
  XOR U2177 ( .A(n32542), .B(n27622), .Z(n26757) );
  AND U2178 ( .A(n28586), .B(n28587), .Z(n30135) );
  ANDN U2179 ( .B(n29617), .A(n29615), .Z(n34708) );
  NOR U2180 ( .A(n26747), .B(n26746), .Z(n26744) );
  XNOR U2181 ( .A(n25873), .B(n26727), .Z(n24262) );
  XOR U2182 ( .A(n31966), .B(n28682), .Z(n24293) );
  AND U2183 ( .A(n28776), .B(n27833), .Z(n30533) );
  ANDN U2184 ( .B(n27183), .A(n27892), .Z(n29069) );
  ANDN U2185 ( .B(n28193), .A(n28191), .Z(n36341) );
  AND U2186 ( .A(n28335), .B(n27230), .Z(n28334) );
  AND U2187 ( .A(n27591), .B(n28212), .Z(n36322) );
  XNOR U2188 ( .A(n26342), .B(n26378), .Z(n25079) );
  AND U2189 ( .A(n26993), .B(n26994), .Z(n33058) );
  XOR U2190 ( .A(n31282), .B(n28206), .Z(n29953) );
  AND U2191 ( .A(n27546), .B(n27545), .Z(n28964) );
  AND U2192 ( .A(n28147), .B(n28149), .Z(n29445) );
  AND U2193 ( .A(n28492), .B(n30667), .Z(n31167) );
  AND U2194 ( .A(n26492), .B(n29419), .Z(n29418) );
  XNOR U2195 ( .A(n28543), .B(n27264), .Z(n28900) );
  ANDN U2196 ( .B(n28850), .A(n29219), .Z(n29762) );
  XNOR U2197 ( .A(n30622), .B(n29812), .Z(n23071) );
  ANDN U2198 ( .B(n30611), .A(n30694), .Z(n30692) );
  XOR U2199 ( .A(n31540), .B(n27689), .Z(n31182) );
  AND U2200 ( .A(n27999), .B(n31483), .Z(n31481) );
  AND U2201 ( .A(n28674), .B(n29411), .Z(n29999) );
  ANDN U2202 ( .B(n28244), .A(n28154), .Z(n34998) );
  AND U2203 ( .A(n30841), .B(n30842), .Z(n30839) );
  NOR U2204 ( .A(n28203), .B(n28202), .Z(n28200) );
  XOR U2205 ( .A(n32508), .B(n28072), .Z(n25025) );
  AND U2206 ( .A(n31342), .B(n28975), .Z(n32290) );
  AND U2207 ( .A(n28660), .B(n29399), .Z(n34318) );
  XNOR U2208 ( .A(n30725), .B(n30724), .Z(n22793) );
  XNOR U2209 ( .A(n26252), .B(n30319), .Z(n23810) );
  AND U2210 ( .A(n26677), .B(n26678), .Z(n26675) );
  ANDN U2211 ( .B(n32772), .A(n30837), .Z(n32770) );
  ANDN U2212 ( .B(n29388), .A(n29387), .Z(n34132) );
  XNOR U2213 ( .A(n27071), .B(n27070), .Z(n24661) );
  AND U2214 ( .A(n26902), .B(n26903), .Z(n26900) );
  XNOR U2215 ( .A(n28291), .B(n28290), .Z(n23019) );
  XOR U2216 ( .A(n27354), .B(n25581), .Z(n24783) );
  XNOR U2217 ( .A(n27888), .B(n27887), .Z(n23422) );
  AND U2218 ( .A(n27599), .B(n27600), .Z(n27597) );
  AND U2219 ( .A(n27917), .B(n29381), .Z(n30602) );
  AND U2220 ( .A(n31859), .B(n31197), .Z(n32482) );
  ANDN U2221 ( .B(n27743), .A(n26437), .Z(n27741) );
  AND U2222 ( .A(n29478), .B(n29480), .Z(n30391) );
  ANDN U2223 ( .B(n29029), .A(n29033), .Z(n29030) );
  AND U2224 ( .A(n26174), .B(n26175), .Z(n30028) );
  ANDN U2225 ( .B(n30192), .A(n27855), .Z(n30190) );
  XOR U2226 ( .A(n26867), .B(n26866), .Z(n23914) );
  AND U2227 ( .A(n25850), .B(n25852), .Z(n29942) );
  ANDN U2228 ( .B(n28524), .A(n28525), .Z(n29570) );
  AND U2229 ( .A(n28409), .B(n28022), .Z(n32676) );
  AND U2230 ( .A(n29336), .B(n29335), .Z(n31814) );
  AND U2231 ( .A(n30417), .B(n30418), .Z(n30415) );
  XNOR U2232 ( .A(n26518), .B(n27923), .Z(n21725) );
  XOR U2233 ( .A(n30154), .B(n26971), .Z(n27038) );
  XNOR U2234 ( .A(n24315), .B(n26153), .Z(n25405) );
  XNOR U2235 ( .A(n26350), .B(n28271), .Z(n25182) );
  XNOR U2236 ( .A(n26082), .B(n30479), .Z(n22325) );
  XOR U2237 ( .A(n28780), .B(n25262), .Z(n24146) );
  XOR U2238 ( .A(n31665), .B(n27276), .Z(n25401) );
  XNOR U2239 ( .A(n29041), .B(n26081), .Z(n23592) );
  XNOR U2240 ( .A(n26530), .B(n26782), .Z(n25227) );
  ANDN U2241 ( .B(n28706), .A(n28806), .Z(n30202) );
  AND U2242 ( .A(n29801), .B(n30689), .Z(n31140) );
  XOR U2243 ( .A(n27398), .B(n27399), .Z(n22994) );
  XNOR U2244 ( .A(n26694), .B(n26693), .Z(n23436) );
  AND U2245 ( .A(n28391), .B(n27503), .Z(n28389) );
  NOR U2246 ( .A(n28279), .B(n27109), .Z(n29516) );
  ANDN U2247 ( .B(n31205), .A(n30348), .Z(n31524) );
  XNOR U2248 ( .A(n29843), .B(n29954), .Z(n21819) );
  XNOR U2249 ( .A(n29277), .B(n26768), .Z(n25362) );
  ANDN U2250 ( .B(n27476), .A(n28515), .Z(n29025) );
  XNOR U2251 ( .A(n26244), .B(n25382), .Z(n22926) );
  XOR U2252 ( .A(n26018), .B(n23015), .Z(n21252) );
  XNOR U2253 ( .A(n24445), .B(n22624), .Z(n21741) );
  XNOR U2254 ( .A(n21583), .B(n21584), .Z(n19861) );
  XNOR U2255 ( .A(n27669), .B(n24798), .Z(n21524) );
  AND U2256 ( .A(n21793), .B(n21794), .Z(n21791) );
  AND U2257 ( .A(n20881), .B(n20882), .Z(n20879) );
  AND U2258 ( .A(n24130), .B(n24129), .Z(n24679) );
  ANDN U2259 ( .B(n20164), .A(n19891), .Z(n21217) );
  AND U2260 ( .A(n19156), .B(n21370), .Z(n26375) );
  XNOR U2261 ( .A(n19042), .B(n22585), .Z(n19740) );
  AND U2262 ( .A(n23543), .B(n22722), .Z(n23542) );
  AND U2263 ( .A(n20557), .B(n20558), .Z(n20555) );
  XOR U2264 ( .A(n27451), .B(n23660), .Z(n19720) );
  AND U2265 ( .A(n22203), .B(n22205), .Z(n22966) );
  ANDN U2266 ( .B(n19745), .A(n19744), .Z(n19742) );
  ANDN U2267 ( .B(n20513), .A(n20512), .Z(n20510) );
  AND U2268 ( .A(n22292), .B(n24687), .Z(n26514) );
  AND U2269 ( .A(n23650), .B(n22737), .Z(n23649) );
  AND U2270 ( .A(n21855), .B(n21854), .Z(n24914) );
  AND U2271 ( .A(n23215), .B(n22455), .Z(n23214) );
  AND U2272 ( .A(n22444), .B(n20931), .Z(n22442) );
  ANDN U2273 ( .B(n20960), .A(n20959), .Z(n20957) );
  XOR U2274 ( .A(n24188), .B(n22780), .Z(n16397) );
  AND U2275 ( .A(n21798), .B(n23803), .Z(n24502) );
  ANDN U2276 ( .B(n25138), .A(n23238), .Z(n35866) );
  AND U2277 ( .A(n20863), .B(n20861), .Z(n27261) );
  AND U2278 ( .A(n22048), .B(n22049), .Z(n22046) );
  ANDN U2279 ( .B(n18851), .A(n18850), .Z(n18848) );
  AND U2280 ( .A(n20725), .B(n20726), .Z(n20723) );
  XNOR U2281 ( .A(n21253), .B(n20017), .Z(n19069) );
  ANDN U2282 ( .B(n23452), .A(n23453), .Z(n26273) );
  ANDN U2283 ( .B(n20584), .A(n20585), .Z(n24809) );
  XOR U2284 ( .A(n21933), .B(n20264), .Z(n16766) );
  NOR U2285 ( .A(n23292), .B(n23172), .Z(n24882) );
  AND U2286 ( .A(n19972), .B(n19973), .Z(n22989) );
  ANDN U2287 ( .B(n21656), .A(n21743), .Z(n23514) );
  AND U2288 ( .A(n21808), .B(n20625), .Z(n21806) );
  AND U2289 ( .A(n19340), .B(n20313), .Z(n20311) );
  AND U2290 ( .A(n23672), .B(n23671), .Z(n25904) );
  ANDN U2291 ( .B(n21641), .A(n20231), .Z(n24425) );
  XOR U2292 ( .A(n21769), .B(n21770), .Z(n18369) );
  XNOR U2293 ( .A(n19983), .B(n24726), .Z(n16727) );
  AND U2294 ( .A(n19786), .B(n19527), .Z(n19784) );
  ANDN U2295 ( .B(n20691), .A(n20690), .Z(n20688) );
  AND U2296 ( .A(n21047), .B(n21049), .Z(n24201) );
  ANDN U2297 ( .B(n22848), .A(n22847), .Z(n22846) );
  XNOR U2298 ( .A(n18460), .B(n20480), .Z(n20074) );
  AND U2299 ( .A(n21354), .B(n21345), .Z(n21353) );
  ANDN U2300 ( .B(n22693), .A(n22691), .Z(n23399) );
  AND U2301 ( .A(n21018), .B(n21980), .Z(n25463) );
  AND U2302 ( .A(n20888), .B(n22142), .Z(n22141) );
  ANDN U2303 ( .B(n22773), .A(n22772), .Z(n22771) );
  XOR U2304 ( .A(n23174), .B(n23175), .Z(n18860) );
  AND U2305 ( .A(n21868), .B(n21869), .Z(n21866) );
  XNOR U2306 ( .A(n18819), .B(n18818), .Z(n15671) );
  XOR U2307 ( .A(n20006), .B(n18926), .Z(n18283) );
  XNOR U2308 ( .A(n21341), .B(n21813), .Z(n15635) );
  AND U2309 ( .A(n22125), .B(n22124), .Z(n22122) );
  XNOR U2310 ( .A(n20013), .B(n20252), .Z(n17177) );
  XNOR U2311 ( .A(n21383), .B(n20374), .Z(n18683) );
  NOR U2312 ( .A(n20492), .B(n22399), .Z(n22807) );
  XOR U2313 ( .A(n25737), .B(n21920), .Z(n22184) );
  ANDN U2314 ( .B(n24140), .A(n21526), .Z(n25160) );
  XNOR U2315 ( .A(n21461), .B(n22904), .Z(n15962) );
  ANDN U2316 ( .B(n22424), .A(n20764), .Z(n22423) );
  AND U2317 ( .A(n20929), .B(n22435), .Z(n25450) );
  XOR U2318 ( .A(n22797), .B(n22798), .Z(n18738) );
  AND U2319 ( .A(n24049), .B(n22077), .Z(n24743) );
  XNOR U2320 ( .A(n18264), .B(n18263), .Z(n17055) );
  XNOR U2321 ( .A(n19193), .B(n20277), .Z(n18828) );
  AND U2322 ( .A(n22057), .B(n22151), .Z(n24773) );
  XNOR U2323 ( .A(n20086), .B(n20226), .Z(n18442) );
  XOR U2324 ( .A(n19427), .B(n20570), .Z(n17440) );
  XNOR U2325 ( .A(n19839), .B(n19838), .Z(n16737) );
  XOR U2326 ( .A(n19823), .B(n19746), .Z(n15265) );
  AND U2327 ( .A(n22969), .B(n23119), .Z(n23118) );
  XNOR U2328 ( .A(n17395), .B(n17394), .Z(n14007) );
  XNOR U2329 ( .A(n17143), .B(n19556), .Z(n15611) );
  XNOR U2330 ( .A(n18038), .B(n17601), .Z(n13683) );
  XNOR U2331 ( .A(n17139), .B(n17140), .Z(n15788) );
  XNOR U2332 ( .A(n20838), .B(n16531), .Z(n14865) );
  XNOR U2333 ( .A(n13869), .B(n12366), .Z(n12090) );
  AND U2334 ( .A(n17163), .B(n17161), .Z(n18107) );
  ANDN U2335 ( .B(n14622), .A(n15178), .Z(n25208) );
  ANDN U2336 ( .B(n15301), .A(n12799), .Z(n15298) );
  ANDN U2337 ( .B(n13785), .A(n13783), .Z(n14991) );
  AND U2338 ( .A(n14586), .B(n14588), .Z(n19449) );
  AND U2339 ( .A(n15712), .B(n15711), .Z(n15709) );
  AND U2340 ( .A(n17404), .B(n14598), .Z(n19943) );
  ANDN U2341 ( .B(n14708), .A(n14706), .Z(n17255) );
  AND U2342 ( .A(n16288), .B(n15992), .Z(n16287) );
  ANDN U2343 ( .B(n13679), .A(n13678), .Z(n13676) );
  AND U2344 ( .A(n14433), .B(n14434), .Z(n14431) );
  ANDN U2345 ( .B(n13060), .A(n13059), .Z(n13057) );
  XOR U2346 ( .A(n15090), .B(n15091), .Z(n11777) );
  AND U2347 ( .A(n13113), .B(n13114), .Z(n19381) );
  XOR U2348 ( .A(n16030), .B(n13435), .Z(n10401) );
  ANDN U2349 ( .B(n15677), .A(n14868), .Z(n16965) );
  AND U2350 ( .A(n13266), .B(n13268), .Z(n14148) );
  AND U2351 ( .A(n15310), .B(n15311), .Z(n15308) );
  AND U2352 ( .A(n14035), .B(n14036), .Z(n14033) );
  AND U2353 ( .A(n15369), .B(n14421), .Z(n16260) );
  AND U2354 ( .A(n15820), .B(n18624), .Z(n19079) );
  ANDN U2355 ( .B(n19110), .A(n16711), .Z(n19113) );
  AND U2356 ( .A(n14050), .B(n15227), .Z(n18431) );
  XNOR U2357 ( .A(n12068), .B(n12963), .Z(n9118) );
  AND U2358 ( .A(n16777), .B(n15987), .Z(n17103) );
  AND U2359 ( .A(n16435), .B(n16433), .Z(n17948) );
  ANDN U2360 ( .B(n17675), .A(n12449), .Z(n17673) );
  ANDN U2361 ( .B(n15161), .A(n15160), .Z(n15158) );
  AND U2362 ( .A(n14658), .B(n13225), .Z(n16463) );
  NOR U2363 ( .A(n14495), .B(n13713), .Z(n14493) );
  ANDN U2364 ( .B(n13452), .A(n13450), .Z(n18873) );
  AND U2365 ( .A(n15575), .B(n16329), .Z(n16831) );
  AND U2366 ( .A(n16137), .B(n16138), .Z(n16136) );
  ANDN U2367 ( .B(n14939), .A(n14938), .Z(n14936) );
  XNOR U2368 ( .A(n11848), .B(n11847), .Z(n9939) );
  XOR U2369 ( .A(n11323), .B(n14592), .Z(n10878) );
  XNOR U2370 ( .A(n17492), .B(n12895), .Z(n9783) );
  AND U2371 ( .A(n14275), .B(n14225), .Z(n18927) );
  ANDN U2372 ( .B(n16849), .A(n14027), .Z(n18449) );
  XNOR U2373 ( .A(n14732), .B(n14183), .Z(n10396) );
  AND U2374 ( .A(n13324), .B(n13325), .Z(n13322) );
  AND U2375 ( .A(n16315), .B(n15063), .Z(n17662) );
  ANDN U2376 ( .B(n14875), .A(n16675), .Z(n16672) );
  AND U2377 ( .A(n14630), .B(n14631), .Z(n15475) );
  XNOR U2378 ( .A(n12205), .B(n12793), .Z(n11325) );
  XNOR U2379 ( .A(n12125), .B(n12124), .Z(n9872) );
  ANDN U2380 ( .B(n16231), .A(n16278), .Z(n17040) );
  AND U2381 ( .A(n14285), .B(n14284), .Z(n14282) );
  AND U2382 ( .A(n14458), .B(n14459), .Z(n14456) );
  ANDN U2383 ( .B(n16694), .A(n16693), .Z(n16692) );
  XOR U2384 ( .A(n17446), .B(n14069), .Z(n11909) );
  XNOR U2385 ( .A(n13306), .B(n13305), .Z(n10868) );
  XOR U2386 ( .A(n22810), .B(n14782), .Z(n14188) );
  XNOR U2387 ( .A(n11898), .B(n11897), .Z(n9790) );
  XNOR U2388 ( .A(n11976), .B(n14154), .Z(n9623) );
  ANDN U2389 ( .B(n16017), .A(n16155), .Z(n17695) );
  XNOR U2390 ( .A(n15046), .B(n12768), .Z(n9107) );
  XNOR U2391 ( .A(n9112), .B(n9113), .Z(n6649) );
  XOR U2392 ( .A(n9527), .B(n9526), .Z(n6726) );
  AND U2393 ( .A(n7813), .B(n7717), .Z(n7812) );
  AND U2394 ( .A(n8384), .B(n8317), .Z(n8383) );
  XOR U2395 ( .A(n12187), .B(n9038), .Z(n5145) );
  ANDN U2396 ( .B(n9021), .A(n6595), .Z(n9019) );
  ANDN U2397 ( .B(n8578), .A(n8522), .Z(n8576) );
  AND U2398 ( .A(n7840), .B(n7842), .Z(n8954) );
  AND U2399 ( .A(n7539), .B(n7540), .Z(n7537) );
  XNOR U2400 ( .A(n6054), .B(n6053), .Z(n5584) );
  ANDN U2401 ( .B(n6901), .A(n6900), .Z(n6898) );
  AND U2402 ( .A(n11470), .B(n8432), .Z(n11644) );
  AND U2403 ( .A(n12154), .B(n12155), .Z(n12309) );
  XNOR U2404 ( .A(n6347), .B(n6503), .Z(n5187) );
  XOR U2405 ( .A(n9451), .B(n7292), .Z(n7273) );
  AND U2406 ( .A(n10003), .B(n10004), .Z(n11051) );
  XOR U2407 ( .A(n11449), .B(n7743), .Z(n1692) );
  AND U2408 ( .A(n9406), .B(n11274), .Z(n11272) );
  AND U2409 ( .A(n9742), .B(n8395), .Z(n9740) );
  AND U2410 ( .A(n6482), .B(n6483), .Z(n6480) );
  AND U2411 ( .A(n8894), .B(n8970), .Z(n8969) );
  AND U2412 ( .A(n7804), .B(n10568), .Z(n10566) );
  AND U2413 ( .A(n7599), .B(n7600), .Z(n7597) );
  AND U2414 ( .A(n6508), .B(n6509), .Z(n6506) );
  AND U2415 ( .A(n6535), .B(n6536), .Z(n6533) );
  XOR U2416 ( .A(n8789), .B(n6491), .Z(n2552) );
  ANDN U2417 ( .B(n6571), .A(n9013), .Z(n9012) );
  ANDN U2418 ( .B(n7050), .A(n7049), .Z(n7047) );
  AND U2419 ( .A(n7876), .B(n7877), .Z(n7874) );
  ANDN U2420 ( .B(n6540), .A(n8873), .Z(n8919) );
  AND U2421 ( .A(n6604), .B(n9028), .Z(n9072) );
  XNOR U2422 ( .A(n12503), .B(n8162), .Z(n3831) );
  XOR U2423 ( .A(n11529), .B(n11530), .Z(n3677) );
  AND U2424 ( .A(n6804), .B(n6805), .Z(n6802) );
  XOR U2425 ( .A(n16937), .B(n8619), .Z(n3751) );
  XNOR U2426 ( .A(n10600), .B(n9689), .Z(n3764) );
  XNOR U2427 ( .A(n6248), .B(n8646), .Z(n1675) );
  AND U2428 ( .A(n10032), .B(n10030), .Z(n11169) );
  XNOR U2429 ( .A(n11709), .B(n7872), .Z(n3808) );
  ANDN U2430 ( .B(n7687), .A(n7686), .Z(n7684) );
  XNOR U2431 ( .A(n6048), .B(n6047), .Z(n3834) );
  NOR U2432 ( .A(n11996), .B(n11995), .Z(n16617) );
  AND U2433 ( .A(n7092), .B(n7093), .Z(n7090) );
  NOR U2434 ( .A(n7912), .B(n7911), .Z(n8983) );
  NOR U2435 ( .A(n6689), .B(n6688), .Z(n7124) );
  XOR U2436 ( .A(n7566), .B(n7567), .Z(n4365) );
  ANDN U2437 ( .B(n9219), .A(n7983), .Z(n9217) );
  XOR U2438 ( .A(n9313), .B(n9314), .Z(n4948) );
  XOR U2439 ( .A(n6705), .B(n6706), .Z(n6173) );
  AND U2440 ( .A(n7904), .B(n7905), .Z(n7902) );
  XOR U2441 ( .A(n11217), .B(n7168), .Z(n5785) );
  XOR U2442 ( .A(n18743), .B(n7734), .Z(n4134) );
  XNOR U2443 ( .A(n6204), .B(n7890), .Z(n1946) );
  AND U2444 ( .A(n7522), .B(n9994), .Z(n10018) );
  XNOR U2445 ( .A(n8973), .B(n8972), .Z(n3238) );
  AND U2446 ( .A(n7883), .B(n10542), .Z(n10681) );
  XNOR U2447 ( .A(n6302), .B(n9282), .Z(n1736) );
  ANDN U2448 ( .B(n11986), .A(n13728), .Z(n14755) );
  XNOR U2449 ( .A(n6326), .B(n9819), .Z(n1758) );
  XNOR U2450 ( .A(n6041), .B(n2203), .Z(n5791) );
  XNOR U2451 ( .A(n3893), .B(n2297), .Z(n2941) );
  XNOR U2452 ( .A(n4226), .B(n1662), .Z(n3967) );
  AND U2453 ( .A(n4444), .B(n4445), .Z(n4442) );
  AND U2454 ( .A(n4505), .B(n4506), .Z(n4503) );
  NANDN U2455 ( .A(n4551), .B(n4552), .Z(n4550) );
  ANDN U2456 ( .B(n4568), .A(n4567), .Z(n4565) );
  AND U2457 ( .A(n4587), .B(n4588), .Z(n4585) );
  NOR U2458 ( .A(n4626), .B(n4625), .Z(n4623) );
  AND U2459 ( .A(n4637), .B(n4638), .Z(n4635) );
  AND U2460 ( .A(n4696), .B(n4695), .Z(n4693) );
  ANDN U2461 ( .B(n4959), .A(n4755), .Z(n4957) );
  AND U2462 ( .A(n4435), .B(n4894), .Z(n5118) );
  AND U2463 ( .A(n4472), .B(n4925), .Z(n5146) );
  AND U2464 ( .A(n4554), .B(n4994), .Z(n5200) );
  ANDN U2465 ( .B(n4997), .A(n4558), .Z(n5203) );
  AND U2466 ( .A(n5000), .B(n4562), .Z(n5205) );
  AND U2467 ( .A(n5617), .B(n5618), .Z(n5615) );
  ANDN U2468 ( .B(n5713), .A(n5714), .Z(n5712) );
  AND U2469 ( .A(n5716), .B(n1044), .Z(n5715) );
  AND U2470 ( .A(n5777), .B(n1141), .Z(n5776) );
  AND U2471 ( .A(n5797), .B(n1173), .Z(n5796) );
  AND U2472 ( .A(n5725), .B(n5923), .Z(n5919) );
  AND U2473 ( .A(n5838), .B(n6140), .Z(n6136) );
  ANDN U2474 ( .B(n5908), .A(n1047), .Z(n6250) );
  ANDN U2475 ( .B(n5918), .A(n1055), .Z(n6258) );
  XOR U2476 ( .A(n1290), .B(n1291), .Z(out[941]) );
  NOR U2477 ( .A(n1357), .B(n1356), .Z(n1354) );
  AND U2478 ( .A(n1380), .B(n1381), .Z(n1378) );
  XOR U2479 ( .A(n1446), .B(n1447), .Z(out[906]) );
  AND U2480 ( .A(n1269), .B(n1530), .Z(n1529) );
  AND U2481 ( .A(n1536), .B(n1280), .Z(n1535) );
  AND U2482 ( .A(n1542), .B(n1284), .Z(n1541) );
  AND U2483 ( .A(n1565), .B(n1325), .Z(n1564) );
  AND U2484 ( .A(n1601), .B(n1384), .Z(n1600) );
  AND U2485 ( .A(n1611), .B(n1408), .Z(n1610) );
  AND U2486 ( .A(n1657), .B(n1493), .Z(n1656) );
  AND U2487 ( .A(n1848), .B(n1595), .Z(n1845) );
  AND U2488 ( .A(n1319), .B(n1786), .Z(n2061) );
  ANDN U2489 ( .B(n2714), .A(n2713), .Z(n2711) );
  XOR U2490 ( .A(n2910), .B(n2911), .Z(out[588]) );
  AND U2491 ( .A(n3020), .B(n2766), .Z(n3019) );
  AND U2492 ( .A(n3032), .B(n2793), .Z(n3031) );
  AND U2493 ( .A(n3081), .B(n2872), .Z(n3080) );
  AND U2494 ( .A(n3098), .B(n2896), .Z(n3097) );
  NOR U2495 ( .A(n3327), .B(n3326), .Z(n3324) );
  NOR U2496 ( .A(n3361), .B(n3360), .Z(n3358) );
  ANDN U2497 ( .B(n3151), .A(n2692), .Z(n3408) );
  AND U2498 ( .A(n2756), .B(n3211), .Z(n3455) );
  AND U2499 ( .A(n3239), .B(n2788), .Z(n3479) );
  ANDN U2500 ( .B(n3278), .A(n2832), .Z(n3511) );
  ANDN U2501 ( .B(n2875), .A(n3316), .Z(n3541) );
  ANDN U2502 ( .B(n3365), .A(n2927), .Z(n3578) );
  ANDN U2503 ( .B(n3369), .A(n2931), .Z(n3580) );
  AND U2504 ( .A(n4079), .B(n1821), .Z(n4077) );
  ANDN U2505 ( .B(n3946), .A(n4150), .Z(n4148) );
  ANDN U2506 ( .B(n4178), .A(n3426), .Z(n4357) );
  XNOR U2507 ( .A(n52476), .B(n52475), .Z(n52332) );
  XNOR U2508 ( .A(n52708), .B(n51921), .Z(n51434) );
  XOR U2509 ( .A(n52669), .B(n52222), .Z(n51094) );
  XNOR U2510 ( .A(n53167), .B(n52707), .Z(n51721) );
  XNOR U2511 ( .A(n52871), .B(n52802), .Z(n52113) );
  XNOR U2512 ( .A(n53261), .B(n53385), .Z(n52523) );
  XNOR U2513 ( .A(n51455), .B(n52491), .Z(n51349) );
  XNOR U2514 ( .A(n52578), .B(n52577), .Z(n49608) );
  XNOR U2515 ( .A(n52641), .B(n52640), .Z(n49795) );
  XNOR U2516 ( .A(n52715), .B(n52191), .Z(n52028) );
  XNOR U2517 ( .A(n53373), .B(n52362), .Z(n51397) );
  XNOR U2518 ( .A(n53030), .B(n52178), .Z(n51582) );
  XNOR U2519 ( .A(n52395), .B(n52654), .Z(n52089) );
  XNOR U2520 ( .A(n52697), .B(n52696), .Z(n50507) );
  XNOR U2521 ( .A(n52400), .B(n52399), .Z(n51332) );
  XNOR U2522 ( .A(n52569), .B(n52568), .Z(n50835) );
  XOR U2523 ( .A(n52682), .B(n52345), .Z(n51624) );
  XOR U2524 ( .A(n51924), .B(n52417), .Z(n51708) );
  XOR U2525 ( .A(n53054), .B(n53212), .Z(n51789) );
  XOR U2526 ( .A(n51917), .B(n51916), .Z(n48701) );
  XOR U2527 ( .A(n52581), .B(n52907), .Z(n50434) );
  XNOR U2528 ( .A(n52350), .B(n52780), .Z(n51399) );
  XNOR U2529 ( .A(n52773), .B(n52887), .Z(n49955) );
  XOR U2530 ( .A(n52933), .B(n52772), .Z(n50520) );
  XNOR U2531 ( .A(n52202), .B(n52589), .Z(n50834) );
  XNOR U2532 ( .A(n53243), .B(n53242), .Z(n51205) );
  XNOR U2533 ( .A(n52917), .B(n52542), .Z(n50815) );
  XNOR U2534 ( .A(n52122), .B(n52121), .Z(n51539) );
  XOR U2535 ( .A(n52774), .B(n52450), .Z(n50448) );
  XNOR U2536 ( .A(n52855), .B(n52854), .Z(n52303) );
  XNOR U2537 ( .A(round_reg[1400]), .B(n49977), .Z(n47424) );
  XOR U2538 ( .A(round_reg[758]), .B(n48445), .Z(n46962) );
  XNOR U2539 ( .A(round_reg[418]), .B(n50745), .Z(n49725) );
  XOR U2540 ( .A(round_reg[165]), .B(n48566), .Z(n51472) );
  XNOR U2541 ( .A(round_reg[861]), .B(n51032), .Z(n47558) );
  XNOR U2542 ( .A(round_reg[1337]), .B(n50828), .Z(n47432) );
  XOR U2543 ( .A(round_reg[882]), .B(n51466), .Z(n45884) );
  ANDN U2544 ( .B(n51806), .A(n50685), .Z(n51805) );
  ANDN U2545 ( .B(n47666), .A(n47665), .Z(n47663) );
  ANDN U2546 ( .B(n48489), .A(n48491), .Z(n51356) );
  ANDN U2547 ( .B(n48675), .A(n49662), .Z(n49661) );
  ANDN U2548 ( .B(n49735), .A(n49736), .Z(n50889) );
  ANDN U2549 ( .B(n49765), .A(n49764), .Z(n50898) );
  ANDN U2550 ( .B(n50781), .A(n50783), .Z(n51562) );
  AND U2551 ( .A(n50004), .B(n50005), .Z(n50003) );
  ANDN U2552 ( .B(n50037), .A(n50036), .Z(n50034) );
  ANDN U2553 ( .B(n48642), .A(n48233), .Z(n52465) );
  AND U2554 ( .A(n49411), .B(n49655), .Z(n51950) );
  AND U2555 ( .A(n48855), .B(n48853), .Z(n49281) );
  XOR U2556 ( .A(n48012), .B(n49536), .Z(n44461) );
  XNOR U2557 ( .A(n47056), .B(n45751), .Z(n43457) );
  XNOR U2558 ( .A(n47151), .B(n47150), .Z(n43581) );
  ANDN U2559 ( .B(n46952), .A(n46951), .Z(n46949) );
  XNOR U2560 ( .A(n45437), .B(n51022), .Z(n45723) );
  ANDN U2561 ( .B(n51210), .A(n50580), .Z(n51673) );
  ANDN U2562 ( .B(n47774), .A(n49125), .Z(n51139) );
  ANDN U2563 ( .B(n48591), .A(n48592), .Z(n48771) );
  ANDN U2564 ( .B(n47353), .A(n48521), .Z(n48519) );
  ANDN U2565 ( .B(n49887), .A(n49889), .Z(n50209) );
  ANDN U2566 ( .B(n46973), .A(n46972), .Z(n47966) );
  ANDN U2567 ( .B(n49101), .A(n49102), .Z(n50469) );
  ANDN U2568 ( .B(n45876), .A(n45875), .Z(n45873) );
  AND U2569 ( .A(n50878), .B(n50879), .Z(n51460) );
  AND U2570 ( .A(n48092), .B(n48922), .Z(n48921) );
  AND U2571 ( .A(n45882), .B(n45883), .Z(n50713) );
  ANDN U2572 ( .B(n48159), .A(n48160), .Z(n50193) );
  AND U2573 ( .A(n48819), .B(n51638), .Z(n53302) );
  ANDN U2574 ( .B(n50576), .A(n47191), .Z(n51473) );
  ANDN U2575 ( .B(n48544), .A(n48543), .Z(n48541) );
  XOR U2576 ( .A(n49439), .B(n49438), .Z(n41649) );
  ANDN U2577 ( .B(n46984), .A(n46983), .Z(n46981) );
  XNOR U2578 ( .A(n48039), .B(n50570), .Z(n44673) );
  AND U2579 ( .A(n49222), .B(n48347), .Z(n49796) );
  ANDN U2580 ( .B(n47091), .A(n47092), .Z(n47348) );
  XOR U2581 ( .A(n51799), .B(n50325), .Z(n45958) );
  ANDN U2582 ( .B(n46323), .A(n46324), .Z(n47338) );
  XOR U2583 ( .A(n47115), .B(n48447), .Z(n47110) );
  XNOR U2584 ( .A(n48883), .B(n47248), .Z(n44488) );
  XNOR U2585 ( .A(n47259), .B(n47258), .Z(n44774) );
  ANDN U2586 ( .B(n50387), .A(n50388), .Z(n53023) );
  ANDN U2587 ( .B(n47834), .A(n47833), .Z(n47831) );
  XNOR U2588 ( .A(n47126), .B(n46531), .Z(n46601) );
  AND U2589 ( .A(n49930), .B(n49931), .Z(n49929) );
  AND U2590 ( .A(n49006), .B(n49007), .Z(n49004) );
  AND U2591 ( .A(n48755), .B(n48753), .Z(n52305) );
  AND U2592 ( .A(n48861), .B(n49284), .Z(n51105) );
  ANDN U2593 ( .B(n48980), .A(n46621), .Z(n53681) );
  XNOR U2594 ( .A(n47236), .B(n48320), .Z(n44223) );
  XNOR U2595 ( .A(n46544), .B(n46543), .Z(n45443) );
  AND U2596 ( .A(n50620), .B(n49528), .Z(n50914) );
  XNOR U2597 ( .A(n46921), .B(n46920), .Z(n42210) );
  ANDN U2598 ( .B(n50085), .A(n50086), .Z(n51832) );
  ANDN U2599 ( .B(n47553), .A(n47941), .Z(n47940) );
  AND U2600 ( .A(n47647), .B(n47649), .Z(n52064) );
  ANDN U2601 ( .B(n46970), .A(n46969), .Z(n46967) );
  XOR U2602 ( .A(n47356), .B(n47355), .Z(n42329) );
  XNOR U2603 ( .A(n48694), .B(n49823), .Z(n42513) );
  AND U2604 ( .A(n46858), .B(n47014), .Z(n52381) );
  ANDN U2605 ( .B(n46486), .A(n46485), .Z(n46483) );
  XOR U2606 ( .A(n50569), .B(n46532), .Z(n43319) );
  AND U2607 ( .A(n48033), .B(n46240), .Z(n50481) );
  XNOR U2608 ( .A(n50589), .B(n50588), .Z(n42855) );
  ANDN U2609 ( .B(n50321), .A(n50320), .Z(n50319) );
  XNOR U2610 ( .A(n46100), .B(n50787), .Z(n48401) );
  ANDN U2611 ( .B(n50251), .A(n50250), .Z(n50248) );
  XNOR U2612 ( .A(n47520), .B(n47519), .Z(n43719) );
  XNOR U2613 ( .A(n47307), .B(n44837), .Z(n39504) );
  XNOR U2614 ( .A(n45080), .B(n45079), .Z(n41131) );
  XNOR U2615 ( .A(n43670), .B(n43671), .Z(n41857) );
  XNOR U2616 ( .A(n46553), .B(n45203), .Z(n40107) );
  XNOR U2617 ( .A(n44618), .B(n44619), .Z(n41100) );
  XNOR U2618 ( .A(n48379), .B(n45569), .Z(n42608) );
  XNOR U2619 ( .A(n45504), .B(n49969), .Z(n45018) );
  XNOR U2620 ( .A(n44680), .B(n44679), .Z(n41258) );
  XNOR U2621 ( .A(n46589), .B(n44859), .Z(n40739) );
  XNOR U2622 ( .A(n44535), .B(n44534), .Z(n40770) );
  XNOR U2623 ( .A(n46513), .B(n42219), .Z(n42620) );
  XOR U2624 ( .A(n43073), .B(n45925), .Z(n45049) );
  XNOR U2625 ( .A(n45657), .B(n43562), .Z(n40398) );
  XNOR U2626 ( .A(n43463), .B(n44017), .Z(n40711) );
  XNOR U2627 ( .A(n45719), .B(n43303), .Z(n43880) );
  XNOR U2628 ( .A(n43643), .B(n43644), .Z(n43526) );
  XOR U2629 ( .A(n47584), .B(n39965), .Z(n39245) );
  AND U2630 ( .A(n43365), .B(n43366), .Z(n43364) );
  AND U2631 ( .A(n41312), .B(n44383), .Z(n48191) );
  AND U2632 ( .A(n42245), .B(n42244), .Z(n46298) );
  ANDN U2633 ( .B(n44293), .A(n42289), .Z(n46243) );
  AND U2634 ( .A(n43289), .B(n40236), .Z(n45337) );
  ANDN U2635 ( .B(n40391), .A(n40390), .Z(n40388) );
  AND U2636 ( .A(n43176), .B(n43178), .Z(n43689) );
  AND U2637 ( .A(n43229), .B(n43228), .Z(n46096) );
  AND U2638 ( .A(n42173), .B(n41621), .Z(n43572) );
  ANDN U2639 ( .B(n41225), .A(n42955), .Z(n42954) );
  ANDN U2640 ( .B(n42808), .A(n42809), .Z(n43531) );
  ANDN U2641 ( .B(n41934), .A(n41932), .Z(n44259) );
  AND U2642 ( .A(n42869), .B(n41772), .Z(n42866) );
  ANDN U2643 ( .B(n42117), .A(n42116), .Z(n42114) );
  ANDN U2644 ( .B(n43387), .A(n40947), .Z(n43385) );
  AND U2645 ( .A(n43693), .B(n43694), .Z(n47394) );
  XNOR U2646 ( .A(n41579), .B(n41578), .Z(n38961) );
  ANDN U2647 ( .B(n45055), .A(n39957), .Z(n45926) );
  AND U2648 ( .A(n41983), .B(n42962), .Z(n44594) );
  XNOR U2649 ( .A(n42721), .B(n42722), .Z(n40207) );
  AND U2650 ( .A(n41909), .B(n41910), .Z(n41907) );
  AND U2651 ( .A(n43938), .B(n43427), .Z(n44388) );
  XNOR U2652 ( .A(n44958), .B(n42973), .Z(n37001) );
  AND U2653 ( .A(n40807), .B(n40808), .Z(n40805) );
  AND U2654 ( .A(n42815), .B(n40257), .Z(n43058) );
  AND U2655 ( .A(n43233), .B(n43234), .Z(n43231) );
  AND U2656 ( .A(n41549), .B(n40938), .Z(n49286) );
  AND U2657 ( .A(n40645), .B(n40643), .Z(n46452) );
  XOR U2658 ( .A(n44919), .B(n42741), .Z(n39010) );
  AND U2659 ( .A(n43809), .B(n43808), .Z(n46206) );
  ANDN U2660 ( .B(n40743), .A(n40744), .Z(n43553) );
  XOR U2661 ( .A(n41557), .B(n40488), .Z(n38294) );
  AND U2662 ( .A(n42762), .B(n42763), .Z(n42761) );
  AND U2663 ( .A(n44103), .B(n41542), .Z(n45700) );
  AND U2664 ( .A(n42374), .B(n42375), .Z(n45475) );
  AND U2665 ( .A(n39510), .B(n43505), .Z(n46217) );
  XNOR U2666 ( .A(n42351), .B(n42352), .Z(n39144) );
  XNOR U2667 ( .A(n41491), .B(n41479), .Z(n40766) );
  AND U2668 ( .A(n42986), .B(n42984), .Z(n45689) );
  XOR U2669 ( .A(n39675), .B(n42050), .Z(n37472) );
  AND U2670 ( .A(n40726), .B(n40727), .Z(n42781) );
  AND U2671 ( .A(n44475), .B(n44248), .Z(n53114) );
  ANDN U2672 ( .B(n41464), .A(n41463), .Z(n41461) );
  XNOR U2673 ( .A(n39970), .B(n41091), .Z(n38298) );
  AND U2674 ( .A(n41468), .B(n41632), .Z(n42678) );
  XNOR U2675 ( .A(n40301), .B(n40705), .Z(n38124) );
  XOR U2676 ( .A(n43136), .B(n42236), .Z(n36393) );
  XNOR U2677 ( .A(n39110), .B(n39109), .Z(n38878) );
  AND U2678 ( .A(n40418), .B(n40416), .Z(n40850) );
  XNOR U2679 ( .A(n42785), .B(n42784), .Z(n36364) );
  XNOR U2680 ( .A(n40507), .B(n39155), .Z(n37710) );
  AND U2681 ( .A(n42994), .B(n42995), .Z(n42992) );
  XNOR U2682 ( .A(n38982), .B(n43452), .Z(n37258) );
  AND U2683 ( .A(n43698), .B(n43847), .Z(n45210) );
  AND U2684 ( .A(n45910), .B(n45905), .Z(n46069) );
  XOR U2685 ( .A(n39704), .B(n39703), .Z(n33922) );
  AND U2686 ( .A(n41824), .B(n41822), .Z(n46574) );
  AND U2687 ( .A(n40424), .B(n40842), .Z(n47066) );
  XNOR U2688 ( .A(n43476), .B(n43475), .Z(n37868) );
  XNOR U2689 ( .A(n38810), .B(n38809), .Z(n36209) );
  XNOR U2690 ( .A(n39236), .B(n40542), .Z(n36347) );
  AND U2691 ( .A(n41293), .B(n41442), .Z(n41440) );
  XNOR U2692 ( .A(n39576), .B(n38448), .Z(n35598) );
  AND U2693 ( .A(n43936), .B(n43935), .Z(n45130) );
  XNOR U2694 ( .A(n42804), .B(n41891), .Z(n38972) );
  ANDN U2695 ( .B(n39727), .A(n39726), .Z(n39724) );
  XOR U2696 ( .A(n40530), .B(n40529), .Z(n37802) );
  AND U2697 ( .A(n42751), .B(n42749), .Z(n43708) );
  AND U2698 ( .A(n41359), .B(n41357), .Z(n45042) );
  ANDN U2699 ( .B(n44068), .A(n44069), .Z(n44894) );
  AND U2700 ( .A(n41318), .B(n42910), .Z(n49541) );
  XOR U2701 ( .A(n41148), .B(n41147), .Z(n36976) );
  XOR U2702 ( .A(n41488), .B(n41489), .Z(n37840) );
  XOR U2703 ( .A(n45446), .B(n44018), .Z(n44904) );
  AND U2704 ( .A(n43248), .B(n45012), .Z(n45009) );
  AND U2705 ( .A(n42241), .B(n42242), .Z(n42239) );
  XNOR U2706 ( .A(n35943), .B(n35942), .Z(n35104) );
  XNOR U2707 ( .A(n38896), .B(n39740), .Z(n36529) );
  XNOR U2708 ( .A(n35604), .B(n35603), .Z(n34100) );
  XNOR U2709 ( .A(n37479), .B(n40992), .Z(n37203) );
  XOR U2710 ( .A(n45168), .B(n35929), .Z(n37973) );
  XNOR U2711 ( .A(n39397), .B(n37517), .Z(n34266) );
  XNOR U2712 ( .A(n42778), .B(n39454), .Z(n38054) );
  XOR U2713 ( .A(n35787), .B(n37845), .Z(n33505) );
  XNOR U2714 ( .A(n38954), .B(n36420), .Z(n34142) );
  XOR U2715 ( .A(n39158), .B(n39533), .Z(n37104) );
  XNOR U2716 ( .A(n40157), .B(n38163), .Z(n36651) );
  XOR U2717 ( .A(n38250), .B(n37427), .Z(n35449) );
  XNOR U2718 ( .A(n39497), .B(n35792), .Z(n37952) );
  XNOR U2719 ( .A(n38670), .B(n38401), .Z(n34245) );
  XOR U2720 ( .A(n38154), .B(n36908), .Z(n37158) );
  ANDN U2721 ( .B(n33695), .A(n33694), .Z(n33692) );
  AND U2722 ( .A(n36260), .B(n36261), .Z(n37764) );
  ANDN U2723 ( .B(n34343), .A(n34344), .Z(n37028) );
  AND U2724 ( .A(n37991), .B(n37989), .Z(n38389) );
  AND U2725 ( .A(n33680), .B(n34776), .Z(n34774) );
  ANDN U2726 ( .B(n35044), .A(n35043), .Z(n35041) );
  AND U2727 ( .A(n36035), .B(n36036), .Z(n36034) );
  AND U2728 ( .A(n33792), .B(n35357), .Z(n35355) );
  AND U2729 ( .A(n34420), .B(n34418), .Z(n40922) );
  ANDN U2730 ( .B(n33663), .A(n33662), .Z(n33660) );
  AND U2731 ( .A(n34096), .B(n34076), .Z(n34094) );
  ANDN U2732 ( .B(n38240), .A(n34596), .Z(n38259) );
  XNOR U2733 ( .A(n37342), .B(n35657), .Z(n32972) );
  ANDN U2734 ( .B(n34696), .A(n35163), .Z(n37495) );
  AND U2735 ( .A(n35195), .B(n35196), .Z(n37744) );
  XOR U2736 ( .A(n35694), .B(n34259), .Z(n32343) );
  ANDN U2737 ( .B(n37474), .A(n37128), .Z(n38578) );
  AND U2738 ( .A(n36188), .B(n36189), .Z(n36187) );
  XOR U2739 ( .A(n35069), .B(n35070), .Z(n31635) );
  ANDN U2740 ( .B(n36795), .A(n33160), .Z(n37047) );
  XNOR U2741 ( .A(n32842), .B(n37299), .Z(n32411) );
  XNOR U2742 ( .A(n35506), .B(n35335), .Z(n29286) );
  XNOR U2743 ( .A(n34364), .B(n34363), .Z(n30517) );
  AND U2744 ( .A(n34844), .B(n33984), .Z(n35318) );
  ANDN U2745 ( .B(n33580), .A(n33581), .Z(n40194) );
  AND U2746 ( .A(n33314), .B(n33315), .Z(n33312) );
  AND U2747 ( .A(n34753), .B(n34754), .Z(n34751) );
  AND U2748 ( .A(n34131), .B(n34549), .Z(n39151) );
  XOR U2749 ( .A(n34587), .B(n34588), .Z(n31842) );
  AND U2750 ( .A(n34196), .B(n34197), .Z(n34194) );
  ANDN U2751 ( .B(n35286), .A(n37915), .Z(n37955) );
  AND U2752 ( .A(n34969), .B(n34970), .Z(n36121) );
  XOR U2753 ( .A(n33736), .B(n38226), .Z(n28982) );
  ANDN U2754 ( .B(n33348), .A(n36715), .Z(n37147) );
  XNOR U2755 ( .A(n32931), .B(n33421), .Z(n32806) );
  XNOR U2756 ( .A(n36116), .B(n35732), .Z(n32571) );
  ANDN U2757 ( .B(n35126), .A(n34051), .Z(n41687) );
  AND U2758 ( .A(n35816), .B(n35559), .Z(n39457) );
  AND U2759 ( .A(n34242), .B(n34243), .Z(n34240) );
  AND U2760 ( .A(n35840), .B(n35838), .Z(n40075) );
  ANDN U2761 ( .B(n36050), .A(n36491), .Z(n38354) );
  XNOR U2762 ( .A(n32502), .B(n32501), .Z(n31030) );
  AND U2763 ( .A(n35809), .B(n35808), .Z(n38290) );
  XOR U2764 ( .A(n45765), .B(n38716), .Z(n31660) );
  XNOR U2765 ( .A(n34225), .B(n34224), .Z(n30493) );
  AND U2766 ( .A(n36309), .B(n35342), .Z(n36306) );
  ANDN U2767 ( .B(n34309), .A(n35759), .Z(n38303) );
  AND U2768 ( .A(n33115), .B(n33116), .Z(n33113) );
  XOR U2769 ( .A(n37123), .B(n37092), .Z(n31474) );
  AND U2770 ( .A(n34284), .B(n34282), .Z(n39526) );
  XNOR U2771 ( .A(n34526), .B(n37810), .Z(n32191) );
  AND U2772 ( .A(n33790), .B(n33402), .Z(n39339) );
  AND U2773 ( .A(n34733), .B(n34735), .Z(n39578) );
  XNOR U2774 ( .A(n34326), .B(n37771), .Z(n33226) );
  AND U2775 ( .A(n36014), .B(n35842), .Z(n40123) );
  XNOR U2776 ( .A(n33147), .B(n38225), .Z(n31632) );
  AND U2777 ( .A(n34014), .B(n35391), .Z(n35390) );
  XNOR U2778 ( .A(n33447), .B(n34956), .Z(n31547) );
  AND U2779 ( .A(n37225), .B(n37224), .Z(n39784) );
  ANDN U2780 ( .B(n35253), .A(n37762), .Z(n39005) );
  XOR U2781 ( .A(n38699), .B(n38396), .Z(n30371) );
  XNOR U2782 ( .A(n35957), .B(n33270), .Z(n32018) );
  ANDN U2783 ( .B(n36588), .A(n37207), .Z(n40994) );
  XNOR U2784 ( .A(n33642), .B(n38757), .Z(n31968) );
  ANDN U2785 ( .B(n35462), .A(n35461), .Z(n35460) );
  AND U2786 ( .A(n35009), .B(n35010), .Z(n36668) );
  XNOR U2787 ( .A(n37294), .B(n33376), .Z(n30129) );
  XNOR U2788 ( .A(n34529), .B(n32534), .Z(n31127) );
  XNOR U2789 ( .A(n34398), .B(n34397), .Z(n29528) );
  XNOR U2790 ( .A(n34113), .B(n34112), .Z(n29747) );
  ANDN U2791 ( .B(n33429), .A(n33430), .Z(n35105) );
  AND U2792 ( .A(n35146), .B(n35144), .Z(n38860) );
  XNOR U2793 ( .A(n33513), .B(n33512), .Z(n30764) );
  AND U2794 ( .A(n36805), .B(n36804), .Z(n37410) );
  XOR U2795 ( .A(n32877), .B(n32878), .Z(n32464) );
  XNOR U2796 ( .A(n34015), .B(n33493), .Z(n31348) );
  XNOR U2797 ( .A(n38517), .B(n35263), .Z(n31106) );
  AND U2798 ( .A(n35437), .B(n34984), .Z(n40904) );
  XOR U2799 ( .A(n33063), .B(n33062), .Z(n31598) );
  AND U2800 ( .A(n34152), .B(n33460), .Z(n34150) );
  AND U2801 ( .A(n33975), .B(n33976), .Z(n33973) );
  XOR U2802 ( .A(n34214), .B(n34213), .Z(n30247) );
  AND U2803 ( .A(n36780), .B(n36330), .Z(n36777) );
  ANDN U2804 ( .B(n36515), .A(n35851), .Z(n38391) );
  AND U2805 ( .A(n36867), .B(n36868), .Z(n42927) );
  XNOR U2806 ( .A(n34359), .B(n36499), .Z(n30483) );
  AND U2807 ( .A(n34806), .B(n36698), .Z(n38094) );
  AND U2808 ( .A(n35142), .B(n35141), .Z(n35139) );
  XNOR U2809 ( .A(n40051), .B(n38007), .Z(n32579) );
  ANDN U2810 ( .B(n34581), .A(n35446), .Z(n35664) );
  XNOR U2811 ( .A(n35187), .B(n34690), .Z(n31322) );
  XNOR U2812 ( .A(n29926), .B(n29927), .Z(n25862) );
  XNOR U2813 ( .A(n31854), .B(n31855), .Z(n30349) );
  XNOR U2814 ( .A(n29736), .B(n33363), .Z(n30457) );
  XNOR U2815 ( .A(n33851), .B(n28836), .Z(n29824) );
  XNOR U2816 ( .A(n36560), .B(n29166), .Z(n28181) );
  XOR U2817 ( .A(n28421), .B(n35675), .Z(n26435) );
  XNOR U2818 ( .A(n30903), .B(n31862), .Z(n30357) );
  AND U2819 ( .A(n31921), .B(n33225), .Z(n33325) );
  ANDN U2820 ( .B(n30976), .A(n29635), .Z(n32133) );
  XNOR U2821 ( .A(n32042), .B(n27970), .Z(n29086) );
  ANDN U2822 ( .B(n30405), .A(n30406), .Z(n32608) );
  AND U2823 ( .A(n26204), .B(n29240), .Z(n29777) );
  AND U2824 ( .A(n29683), .B(n29704), .Z(n29703) );
  ANDN U2825 ( .B(n28252), .A(n30565), .Z(n31575) );
  AND U2826 ( .A(n28454), .B(n28444), .Z(n28453) );
  NOR U2827 ( .A(n28001), .B(n28000), .Z(n27998) );
  XOR U2828 ( .A(n31694), .B(n29718), .Z(n23917) );
  ANDN U2829 ( .B(n27353), .A(n26549), .Z(n27352) );
  AND U2830 ( .A(n27824), .B(n27825), .Z(n32563) );
  AND U2831 ( .A(n29688), .B(n29689), .Z(n29686) );
  AND U2832 ( .A(n27604), .B(n28207), .Z(n36181) );
  AND U2833 ( .A(n30576), .B(n28532), .Z(n31260) );
  AND U2834 ( .A(n27276), .B(n27275), .Z(n29739) );
  AND U2835 ( .A(n26745), .B(n26746), .Z(n30522) );
  AND U2836 ( .A(n28350), .B(n28351), .Z(n28348) );
  XOR U2837 ( .A(n32022), .B(n29205), .Z(n22945) );
  AND U2838 ( .A(n28933), .B(n28934), .Z(n30900) );
  ANDN U2839 ( .B(n28645), .A(n31007), .Z(n31004) );
  ANDN U2840 ( .B(n30638), .A(n30637), .Z(n33483) );
  AND U2841 ( .A(n26888), .B(n27194), .Z(n29044) );
  XNOR U2842 ( .A(n25117), .B(n25116), .Z(n23690) );
  AND U2843 ( .A(n30373), .B(n27684), .Z(n34157) );
  AND U2844 ( .A(n31491), .B(n27991), .Z(n31489) );
  ANDN U2845 ( .B(n27480), .A(n28507), .Z(n29018) );
  XNOR U2846 ( .A(n27955), .B(n27240), .Z(n21606) );
  XOR U2847 ( .A(n27851), .B(n27704), .Z(n23513) );
  XNOR U2848 ( .A(n27700), .B(n26702), .Z(n22521) );
  AND U2849 ( .A(n29470), .B(n29471), .Z(n29468) );
  AND U2850 ( .A(n27865), .B(n27772), .Z(n35922) );
  AND U2851 ( .A(n27330), .B(n27329), .Z(n27328) );
  AND U2852 ( .A(n26602), .B(n28475), .Z(n31753) );
  AND U2853 ( .A(n31624), .B(n31092), .Z(n32761) );
  AND U2854 ( .A(n30970), .B(n30971), .Z(n30969) );
  XNOR U2855 ( .A(n27663), .B(n26245), .Z(n26944) );
  AND U2856 ( .A(n27222), .B(n27224), .Z(n31722) );
  XOR U2857 ( .A(n28332), .B(n27708), .Z(n26134) );
  AND U2858 ( .A(n29372), .B(n28843), .Z(n30791) );
  AND U2859 ( .A(n29357), .B(n29643), .Z(n30915) );
  AND U2860 ( .A(n29607), .B(n29609), .Z(n34787) );
  XOR U2861 ( .A(n33379), .B(n30447), .Z(n24824) );
  XNOR U2862 ( .A(n27846), .B(n27728), .Z(n21368) );
  AND U2863 ( .A(n26594), .B(n28467), .Z(n28742) );
  XOR U2864 ( .A(n27204), .B(n25937), .Z(n25757) );
  ANDN U2865 ( .B(n29902), .A(n29901), .Z(n29899) );
  XNOR U2866 ( .A(n27199), .B(n29390), .Z(n23139) );
  XNOR U2867 ( .A(n26779), .B(n25521), .Z(n25839) );
  XNOR U2868 ( .A(n27849), .B(n30806), .Z(n25045) );
  AND U2869 ( .A(n26171), .B(n26172), .Z(n26169) );
  XOR U2870 ( .A(n26541), .B(n26540), .Z(n24904) );
  ANDN U2871 ( .B(n30088), .A(n30087), .Z(n30085) );
  XNOR U2872 ( .A(n26588), .B(n29156), .Z(n22820) );
  ANDN U2873 ( .B(n28140), .A(n32408), .Z(n32406) );
  AND U2874 ( .A(n28854), .B(n29226), .Z(n29760) );
  AND U2875 ( .A(n27623), .B(n27621), .Z(n27935) );
  AND U2876 ( .A(n27040), .B(n26957), .Z(n31336) );
  AND U2877 ( .A(n28484), .B(n28483), .Z(n29154) );
  ANDN U2878 ( .B(n28680), .A(n29126), .Z(n30272) );
  ANDN U2879 ( .B(n27564), .A(n29836), .Z(n30626) );
  ANDN U2880 ( .B(n30398), .A(n31773), .Z(n38697) );
  XNOR U2881 ( .A(n25263), .B(n25262), .Z(n23812) );
  AND U2882 ( .A(n29327), .B(n29017), .Z(n31265) );
  ANDN U2883 ( .B(n28774), .A(n28833), .Z(n30769) );
  XNOR U2884 ( .A(n28009), .B(n30106), .Z(n24442) );
  AND U2885 ( .A(n28189), .B(n26313), .Z(n28187) );
  XNOR U2886 ( .A(n28652), .B(n26703), .Z(n25490) );
  XOR U2887 ( .A(n26730), .B(n31008), .Z(n22790) );
  ANDN U2888 ( .B(n26330), .A(n26329), .Z(n26327) );
  XOR U2889 ( .A(n25103), .B(n25102), .Z(n24399) );
  XOR U2890 ( .A(n30720), .B(n29091), .Z(n29208) );
  XNOR U2891 ( .A(n26863), .B(n28109), .Z(n25032) );
  ANDN U2892 ( .B(n26847), .A(n26846), .Z(n26845) );
  XNOR U2893 ( .A(n27101), .B(n26257), .Z(n23869) );
  AND U2894 ( .A(n30845), .B(n30846), .Z(n30843) );
  AND U2895 ( .A(n29891), .B(n31740), .Z(n32051) );
  AND U2896 ( .A(n32077), .B(n31725), .Z(n32076) );
  XNOR U2897 ( .A(n25825), .B(n26577), .Z(n23505) );
  AND U2898 ( .A(n29223), .B(n29224), .Z(n29222) );
  XNOR U2899 ( .A(n27060), .B(n27059), .Z(n24849) );
  XNOR U2900 ( .A(n26911), .B(n27283), .Z(n23573) );
  AND U2901 ( .A(n27916), .B(n27915), .Z(n31014) );
  XNOR U2902 ( .A(n24312), .B(n23566), .Z(n23880) );
  XNOR U2903 ( .A(n24351), .B(n23065), .Z(n21880) );
  XNOR U2904 ( .A(n24902), .B(n23436), .Z(n22702) );
  XNOR U2905 ( .A(n24600), .B(n22495), .Z(n22734) );
  XNOR U2906 ( .A(n26508), .B(n25008), .Z(n20578) );
  XNOR U2907 ( .A(n25215), .B(n23253), .Z(n19786) );
  XNOR U2908 ( .A(n25205), .B(n25206), .Z(n21262) );
  XOR U2909 ( .A(n24850), .B(n22504), .Z(n21615) );
  XNOR U2910 ( .A(n29808), .B(n23964), .Z(n23213) );
  XNOR U2911 ( .A(n25096), .B(n21221), .Z(n19576) );
  AND U2912 ( .A(n21037), .B(n21177), .Z(n26818) );
  AND U2913 ( .A(n22162), .B(n22044), .Z(n24780) );
  AND U2914 ( .A(n23652), .B(n22741), .Z(n23651) );
  AND U2915 ( .A(n21564), .B(n21565), .Z(n21562) );
  AND U2916 ( .A(n21012), .B(n21983), .Z(n22791) );
  AND U2917 ( .A(n20925), .B(n22431), .Z(n25459) );
  AND U2918 ( .A(n22237), .B(n22470), .Z(n28132) );
  AND U2919 ( .A(n23267), .B(n24082), .Z(n24081) );
  AND U2920 ( .A(n22770), .B(n21051), .Z(n27922) );
  AND U2921 ( .A(n22483), .B(n22484), .Z(n22482) );
  XNOR U2922 ( .A(n19735), .B(n19734), .Z(n18203) );
  ANDN U2923 ( .B(n23388), .A(n23389), .Z(n23409) );
  AND U2924 ( .A(n25647), .B(n23202), .Z(n30872) );
  AND U2925 ( .A(n21902), .B(n21903), .Z(n21901) );
  ANDN U2926 ( .B(n23375), .A(n22596), .Z(n26637) );
  AND U2927 ( .A(n21080), .B(n21128), .Z(n21126) );
  AND U2928 ( .A(n22592), .B(n22591), .Z(n22589) );
  NOR U2929 ( .A(n20574), .B(n20576), .Z(n24802) );
  ANDN U2930 ( .B(n22739), .A(n22738), .Z(n22736) );
  AND U2931 ( .A(n22802), .B(n23344), .Z(n26917) );
  AND U2932 ( .A(n20613), .B(n21802), .Z(n24508) );
  ANDN U2933 ( .B(n20055), .A(n20054), .Z(n24023) );
  ANDN U2934 ( .B(n21941), .A(n21940), .Z(n21938) );
  AND U2935 ( .A(n22927), .B(n23187), .Z(n26243) );
  XNOR U2936 ( .A(n21093), .B(n21092), .Z(n15299) );
  XNOR U2937 ( .A(n20045), .B(n22258), .Z(n16664) );
  AND U2938 ( .A(n20805), .B(n25126), .Z(n25923) );
  XOR U2939 ( .A(n24357), .B(n21972), .Z(n20707) );
  NOR U2940 ( .A(n21312), .B(n21311), .Z(n21309) );
  AND U2941 ( .A(n23207), .B(n23208), .Z(n23205) );
  XNOR U2942 ( .A(n19466), .B(n19465), .Z(n18517) );
  NOR U2943 ( .A(n20648), .B(n20647), .Z(n20645) );
  AND U2944 ( .A(n22696), .B(n22695), .Z(n23397) );
  AND U2945 ( .A(n21200), .B(n20426), .Z(n26061) );
  AND U2946 ( .A(n20586), .B(n21610), .Z(n21609) );
  AND U2947 ( .A(n20492), .B(n20494), .Z(n22398) );
  ANDN U2948 ( .B(n19894), .A(n19895), .Z(n20368) );
  AND U2949 ( .A(n23622), .B(n20262), .Z(n25863) );
  AND U2950 ( .A(n23899), .B(n24155), .Z(n24152) );
  AND U2951 ( .A(n22156), .B(n22038), .Z(n22154) );
  AND U2952 ( .A(n19620), .B(n21102), .Z(n31516) );
  AND U2953 ( .A(n23953), .B(n23949), .Z(n23950) );
  AND U2954 ( .A(n23382), .B(n23383), .Z(n23380) );
  XNOR U2955 ( .A(n23155), .B(n23154), .Z(n19551) );
  XNOR U2956 ( .A(n20380), .B(n20379), .Z(n18154) );
  AND U2957 ( .A(n20001), .B(n19860), .Z(n19999) );
  XNOR U2958 ( .A(n20902), .B(n20602), .Z(n17750) );
  NOR U2959 ( .A(n20946), .B(n20945), .Z(n20943) );
  XOR U2960 ( .A(n20476), .B(n19852), .Z(n17186) );
  AND U2961 ( .A(n21850), .B(n21852), .Z(n23830) );
  XNOR U2962 ( .A(n18552), .B(n18551), .Z(n15196) );
  AND U2963 ( .A(n22052), .B(n22053), .Z(n22050) );
  XNOR U2964 ( .A(n19459), .B(n19877), .Z(n18563) );
  XOR U2965 ( .A(n20324), .B(n20325), .Z(n18591) );
  AND U2966 ( .A(n21031), .B(n21170), .Z(n21168) );
  ANDN U2967 ( .B(n21130), .A(n21132), .Z(n22756) );
  ANDN U2968 ( .B(n21405), .A(n20345), .Z(n25504) );
  XNOR U2969 ( .A(n19516), .B(n18757), .Z(n18266) );
  XOR U2970 ( .A(n22659), .B(n22658), .Z(n15339) );
  AND U2971 ( .A(n19744), .B(n19743), .Z(n20417) );
  XNOR U2972 ( .A(n23179), .B(n21507), .Z(n18557) );
  XNOR U2973 ( .A(n19139), .B(n21281), .Z(n17479) );
  ANDN U2974 ( .B(n19805), .A(n20888), .Z(n25575) );
  XNOR U2975 ( .A(n25034), .B(n23341), .Z(n17338) );
  NOR U2976 ( .A(n23548), .B(n23644), .Z(n24611) );
  AND U2977 ( .A(n20588), .B(n22315), .Z(n26473) );
  AND U2978 ( .A(n24333), .B(n25393), .Z(n25392) );
  AND U2979 ( .A(n18850), .B(n22933), .Z(n22952) );
  ANDN U2980 ( .B(n20730), .A(n20729), .Z(n20727) );
  XNOR U2981 ( .A(n19702), .B(n19701), .Z(n15644) );
  ANDN U2982 ( .B(n20452), .A(n22698), .Z(n25657) );
  XOR U2983 ( .A(n24962), .B(n22692), .Z(n20448) );
  AND U2984 ( .A(n23302), .B(n23303), .Z(n23301) );
  XOR U2985 ( .A(n19167), .B(n19095), .Z(n16529) );
  XNOR U2986 ( .A(n20141), .B(n23385), .Z(n16616) );
  ANDN U2987 ( .B(n22239), .A(n22480), .Z(n24215) );
  XOR U2988 ( .A(n23477), .B(n20988), .Z(n18234) );
  ANDN U2989 ( .B(n20213), .A(n20212), .Z(n20210) );
  XNOR U2990 ( .A(n18343), .B(n20097), .Z(n17795) );
  AND U2991 ( .A(n19858), .B(n19857), .Z(n19855) );
  ANDN U2992 ( .B(n21925), .A(n21924), .Z(n21922) );
  AND U2993 ( .A(n22563), .B(n23362), .Z(n25961) );
  XOR U2994 ( .A(n20488), .B(n20487), .Z(n16613) );
  AND U2995 ( .A(n20927), .B(n20928), .Z(n22523) );
  XOR U2996 ( .A(n24665), .B(n24664), .Z(n17744) );
  XOR U2997 ( .A(n19558), .B(n19557), .Z(n17143) );
  AND U2998 ( .A(n19626), .B(n21465), .Z(n27902) );
  ANDN U2999 ( .B(n19928), .A(n19926), .Z(n19975) );
  AND U3000 ( .A(n21568), .B(n23931), .Z(n24486) );
  XNOR U3001 ( .A(n20305), .B(n18502), .Z(n18072) );
  XOR U3002 ( .A(n18220), .B(n18221), .Z(n12953) );
  XNOR U3003 ( .A(n17937), .B(n17203), .Z(n16429) );
  XNOR U3004 ( .A(n15639), .B(n22537), .Z(n17375) );
  XNOR U3005 ( .A(n19309), .B(n15875), .Z(n14425) );
  XNOR U3006 ( .A(n19710), .B(n16068), .Z(n14710) );
  XNOR U3007 ( .A(n18367), .B(n17853), .Z(n17707) );
  XOR U3008 ( .A(n19680), .B(n16108), .Z(n13883) );
  XOR U3009 ( .A(n18090), .B(n21975), .Z(n17827) );
  XNOR U3010 ( .A(n15955), .B(n15956), .Z(n12938) );
  XNOR U3011 ( .A(n19438), .B(n16088), .Z(n13827) );
  ANDN U3012 ( .B(n15982), .A(n17078), .Z(n17609) );
  AND U3013 ( .A(n12806), .B(n12804), .Z(n13366) );
  XOR U3014 ( .A(n13540), .B(n13079), .Z(n12236) );
  AND U3015 ( .A(n14232), .B(n17242), .Z(n18939) );
  AND U3016 ( .A(n14947), .B(n12826), .Z(n21143) );
  NOR U3017 ( .A(n15109), .B(n15110), .Z(n16646) );
  ANDN U3018 ( .B(n14577), .A(n13776), .Z(n20146) );
  XOR U3019 ( .A(n15940), .B(n13185), .Z(n12193) );
  ANDN U3020 ( .B(n18654), .A(n15513), .Z(n18989) );
  XOR U3021 ( .A(n14248), .B(n13753), .Z(n12407) );
  XNOR U3022 ( .A(n17362), .B(n17361), .Z(n11722) );
  AND U3023 ( .A(n15868), .B(n15084), .Z(n15878) );
  AND U3024 ( .A(n14945), .B(n15187), .Z(n15686) );
  ANDN U3025 ( .B(n14550), .A(n14551), .Z(n16012) );
  AND U3026 ( .A(n15572), .B(n15573), .Z(n15570) );
  AND U3027 ( .A(n14077), .B(n14079), .Z(n15763) );
  AND U3028 ( .A(n17155), .B(n18117), .Z(n19190) );
  AND U3029 ( .A(n17709), .B(n15715), .Z(n18720) );
  AND U3030 ( .A(n15091), .B(n13414), .Z(n17286) );
  NOR U3031 ( .A(n14505), .B(n13735), .Z(n14503) );
  AND U3032 ( .A(n15979), .B(n15980), .Z(n15977) );
  ANDN U3033 ( .B(n13037), .A(n13905), .Z(n16054) );
  AND U3034 ( .A(n12564), .B(n12565), .Z(n12562) );
  ANDN U3035 ( .B(n13688), .A(n14648), .Z(n18047) );
  AND U3036 ( .A(n16768), .B(n17437), .Z(n17434) );
  ANDN U3037 ( .B(n13501), .A(n13502), .Z(n27877) );
  XOR U3038 ( .A(n19081), .B(n15824), .Z(n9890) );
  ANDN U3039 ( .B(n17382), .A(n17383), .Z(n22580) );
  XOR U3040 ( .A(n16824), .B(n16315), .Z(n10981) );
  XOR U3041 ( .A(n14174), .B(n13251), .Z(n11346) );
  ANDN U3042 ( .B(n15448), .A(n15447), .Z(n15446) );
  AND U3043 ( .A(n12354), .B(n15793), .Z(n16949) );
  ANDN U3044 ( .B(n14295), .A(n15122), .Z(n17999) );
  ANDN U3045 ( .B(n13562), .A(n13561), .Z(n13559) );
  ANDN U3046 ( .B(n13968), .A(n13969), .Z(n19366) );
  AND U3047 ( .A(n14864), .B(n15666), .Z(n15664) );
  XNOR U3048 ( .A(n13289), .B(n12661), .Z(n10057) );
  AND U3049 ( .A(n17778), .B(n17779), .Z(n17808) );
  AND U3050 ( .A(n14700), .B(n14702), .Z(n17263) );
  XNOR U3051 ( .A(n12970), .B(n12969), .Z(n9859) );
  XNOR U3052 ( .A(n12721), .B(n12720), .Z(n10738) );
  ANDN U3053 ( .B(n16237), .A(n16235), .Z(n22131) );
  XNOR U3054 ( .A(n12597), .B(n12596), .Z(n10116) );
  XOR U3055 ( .A(n14204), .B(n13584), .Z(n13556) );
  AND U3056 ( .A(n13684), .B(n13682), .Z(n14477) );
  ANDN U3057 ( .B(n13456), .A(n13457), .Z(n18882) );
  ANDN U3058 ( .B(n16421), .A(n16422), .Z(n16419) );
  AND U3059 ( .A(n14685), .B(n14684), .Z(n18663) );
  AND U3060 ( .A(n14494), .B(n13715), .Z(n17021) );
  XNOR U3061 ( .A(n11862), .B(n12022), .Z(n9119) );
  ANDN U3062 ( .B(n12039), .A(n12040), .Z(n16348) );
  XOR U3063 ( .A(n15365), .B(n15366), .Z(n10942) );
  ANDN U3064 ( .B(n14723), .A(n13506), .Z(n16723) );
  AND U3065 ( .A(n17170), .B(n14353), .Z(n20036) );
  AND U3066 ( .A(n13258), .B(n13260), .Z(n14144) );
  ANDN U3067 ( .B(n14573), .A(n13779), .Z(n14571) );
  ANDN U3068 ( .B(n14873), .A(n14874), .Z(n15033) );
  ANDN U3069 ( .B(n16145), .A(n14560), .Z(n16143) );
  ANDN U3070 ( .B(n14754), .A(n14752), .Z(n18899) );
  AND U3071 ( .A(n14628), .B(n14626), .Z(n16489) );
  XNOR U3072 ( .A(n12625), .B(n12624), .Z(n11196) );
  AND U3073 ( .A(n18689), .B(n15801), .Z(n20592) );
  XNOR U3074 ( .A(n14186), .B(n13442), .Z(n11301) );
  XNOR U3075 ( .A(n11571), .B(n13422), .Z(n9242) );
  NOR U3076 ( .A(n15276), .B(n15788), .Z(n17137) );
  AND U3077 ( .A(n17452), .B(n14074), .Z(n17449) );
  AND U3078 ( .A(n14316), .B(n15673), .Z(n20850) );
  AND U3079 ( .A(n12869), .B(n12870), .Z(n12867) );
  AND U3080 ( .A(n16569), .B(n14779), .Z(n22784) );
  ANDN U3081 ( .B(n18085), .A(n18739), .Z(n18737) );
  AND U3082 ( .A(n19267), .B(n14846), .Z(n19281) );
  AND U3083 ( .A(n14961), .B(n13173), .Z(n21278) );
  ANDN U3084 ( .B(n13660), .A(n13194), .Z(n19736) );
  XOR U3085 ( .A(n9530), .B(n11050), .Z(n9995) );
  XNOR U3086 ( .A(n11969), .B(n9872), .Z(n7473) );
  XOR U3087 ( .A(n9101), .B(n9923), .Z(n6832) );
  XNOR U3088 ( .A(n10052), .B(n9426), .Z(n7989) );
  XNOR U3089 ( .A(n10399), .B(n10607), .Z(n9686) );
  XNOR U3090 ( .A(n9652), .B(n9651), .Z(n6794) );
  XNOR U3091 ( .A(n9630), .B(n10291), .Z(n8644) );
  AND U3092 ( .A(n9841), .B(n9842), .Z(n10955) );
  ANDN U3093 ( .B(n7644), .A(n7643), .Z(n7641) );
  AND U3094 ( .A(n7328), .B(n7327), .Z(n7325) );
  ANDN U3095 ( .B(n6716), .A(n6715), .Z(n6713) );
  XNOR U3096 ( .A(n6727), .B(n6728), .Z(n6380) );
  AND U3097 ( .A(n6769), .B(n6770), .Z(n6767) );
  AND U3098 ( .A(n8730), .B(n12260), .Z(n12436) );
  XOR U3099 ( .A(n9405), .B(n9406), .Z(n8248) );
  AND U3100 ( .A(n13004), .B(n6515), .Z(n13508) );
  ANDN U3101 ( .B(n14128), .A(n6569), .Z(n15043) );
  AND U3102 ( .A(n6471), .B(n6472), .Z(n12570) );
  AND U3103 ( .A(n6744), .B(n6742), .Z(n7211) );
  ANDN U3104 ( .B(n7100), .A(n7101), .Z(n8229) );
  ANDN U3105 ( .B(n6603), .A(n9029), .Z(n9027) );
  XOR U3106 ( .A(n12642), .B(n8962), .Z(n1933) );
  ANDN U3107 ( .B(n6456), .A(n6455), .Z(n6453) );
  AND U3108 ( .A(n6845), .B(n6846), .Z(n6843) );
  ANDN U3109 ( .B(n8575), .A(n8574), .Z(n8572) );
  ANDN U3110 ( .B(n9721), .A(n9722), .Z(n11822) );
  ANDN U3111 ( .B(n6487), .A(n8772), .Z(n8795) );
  XNOR U3112 ( .A(n8910), .B(n8909), .Z(n3234) );
  ANDN U3113 ( .B(n8033), .A(n8032), .Z(n8030) );
  AND U3114 ( .A(n8165), .B(n8166), .Z(n8163) );
  XOR U3115 ( .A(n9134), .B(n6631), .Z(n3311) );
  AND U3116 ( .A(n9038), .B(n10798), .Z(n10910) );
  XNOR U3117 ( .A(n6219), .B(n8116), .Z(n1961) );
  ANDN U3118 ( .B(n6500), .A(n6499), .Z(n6497) );
  AND U3119 ( .A(n6859), .B(n6860), .Z(n6857) );
  AND U3120 ( .A(n6651), .B(n7071), .Z(n7069) );
  AND U3121 ( .A(n6886), .B(n6887), .Z(n6884) );
  XNOR U3122 ( .A(n7134), .B(n7135), .Z(n3743) );
  ANDN U3123 ( .B(n6920), .A(n6919), .Z(n6917) );
  AND U3124 ( .A(n6944), .B(n6945), .Z(n6942) );
  XNOR U3125 ( .A(n6234), .B(n8233), .Z(n1973) );
  XNOR U3126 ( .A(n6003), .B(n6002), .Z(n3791) );
  AND U3127 ( .A(n7612), .B(n7613), .Z(n7610) );
  AND U3128 ( .A(n10895), .B(n10896), .Z(n12357) );
  AND U3129 ( .A(n7256), .B(n7257), .Z(n8374) );
  AND U3130 ( .A(n7314), .B(n7313), .Z(n8429) );
  ANDN U3131 ( .B(n8004), .A(n8003), .Z(n8001) );
  AND U3132 ( .A(n7689), .B(n7690), .Z(n8822) );
  AND U3133 ( .A(n7898), .B(n7899), .Z(n8986) );
  AND U3134 ( .A(n9739), .B(n7341), .Z(n9737) );
  XOR U3135 ( .A(n10002), .B(n10003), .Z(n5153) );
  AND U3136 ( .A(n8519), .B(n8567), .Z(n12163) );
  ANDN U3137 ( .B(n6597), .A(n6596), .Z(n6594) );
  ANDN U3138 ( .B(n8609), .A(n8608), .Z(n8606) );
  AND U3139 ( .A(n7009), .B(n7007), .Z(n10447) );
  AND U3140 ( .A(n7845), .B(n7844), .Z(n8949) );
  AND U3141 ( .A(n11149), .B(n8190), .Z(n11147) );
  ANDN U3142 ( .B(n6443), .A(n6442), .Z(n6440) );
  XOR U3143 ( .A(n6620), .B(n6621), .Z(n6011) );
  AND U3144 ( .A(n10445), .B(n8109), .Z(n10454) );
  ANDN U3145 ( .B(n7393), .A(n7392), .Z(n7390) );
  ANDN U3146 ( .B(n8975), .A(n8976), .Z(n11690) );
  ANDN U3147 ( .B(n11199), .A(n7199), .Z(n11343) );
  AND U3148 ( .A(n8320), .B(n8387), .Z(n8386) );
  XNOR U3149 ( .A(n8784), .B(n8783), .Z(n2432) );
  XNOR U3150 ( .A(n6209), .B(n7998), .Z(n1951) );
  XNOR U3151 ( .A(n6214), .B(n8049), .Z(n1955) );
  XOR U3152 ( .A(n8185), .B(n8186), .Z(n4583) );
  XNOR U3153 ( .A(n6253), .B(n9396), .Z(n4237) );
  AND U3154 ( .A(n11546), .B(n10678), .Z(n11727) );
  ANDN U3155 ( .B(n8665), .A(n12290), .Z(n12599) );
  AND U3156 ( .A(n6561), .B(n8933), .Z(n9009) );
  XNOR U3157 ( .A(n6306), .B(n9403), .Z(n1741) );
  XNOR U3158 ( .A(n6314), .B(n9603), .Z(n1749) );
  XNOR U3159 ( .A(n2220), .B(n2221), .Z(n1676) );
  XNOR U3160 ( .A(n3150), .B(n2294), .Z(n2693) );
  XNOR U3161 ( .A(n3652), .B(n2410), .Z(n2722) );
  XNOR U3162 ( .A(n3678), .B(n2445), .Z(n2746) );
  XNOR U3163 ( .A(n2434), .B(n4092), .Z(n1480) );
  AND U3164 ( .A(n4412), .B(n4413), .Z(n4410) );
  AND U3165 ( .A(n4615), .B(n4616), .Z(n4613) );
  AND U3166 ( .A(n4626), .B(n4825), .Z(n4824) );
  ANDN U3167 ( .B(n4969), .A(n4767), .Z(n4966) );
  ANDN U3168 ( .B(n4976), .A(n4771), .Z(n4974) );
  AND U3169 ( .A(n4827), .B(n5052), .Z(n5050) );
  AND U3170 ( .A(n5076), .B(n4845), .Z(n5074) );
  AND U3171 ( .A(n4849), .B(n5082), .Z(n5080) );
  AND U3172 ( .A(n5088), .B(n4853), .Z(n5086) );
  AND U3173 ( .A(n4452), .B(n4904), .Z(n5134) );
  AND U3174 ( .A(n4660), .B(n5079), .Z(n5275) );
  AND U3175 ( .A(n4668), .B(n5085), .Z(n5284) );
  AND U3176 ( .A(n5689), .B(n5690), .Z(n5687) );
  ANDN U3177 ( .B(n5724), .A(n5725), .Z(n5723) );
  ANDN U3178 ( .B(n5944), .A(n5740), .Z(n5940) );
  AND U3179 ( .A(n6185), .B(n5859), .Z(n6181) );
  AND U3180 ( .A(n6240), .B(n5888), .Z(n6236) );
  AND U3181 ( .A(n1043), .B(n5898), .Z(n6245) );
  ANDN U3182 ( .B(n5913), .A(n1051), .Z(n6254) );
  ANDN U3183 ( .B(n6009), .A(n1131), .Z(n6336) );
  XOR U3184 ( .A(n1318), .B(n1319), .Z(out[935]) );
  XOR U3185 ( .A(n1414), .B(n1415), .Z(out[913]) );
  AND U3186 ( .A(n1623), .B(n1901), .Z(n1898) );
  AND U3187 ( .A(n1629), .B(n1913), .Z(n1910) );
  ANDN U3188 ( .B(n1243), .A(n1699), .Z(n1996) );
  AND U3189 ( .A(n1742), .B(n1279), .Z(n2026) );
  AND U3190 ( .A(n1283), .B(n1746), .Z(n2029) );
  ANDN U3191 ( .B(n1351), .A(n1817), .Z(n2087) );
  ANDN U3192 ( .B(n1953), .A(n1471), .Z(n2189) );
  XOR U3193 ( .A(n2851), .B(n2852), .Z(out[600]) );
  AND U3194 ( .A(n3013), .B(n2754), .Z(n3012) );
  AND U3195 ( .A(n2821), .B(n3050), .Z(n3049) );
  AND U3196 ( .A(n3331), .B(n3096), .Z(n3328) );
  AND U3197 ( .A(n3100), .B(n3339), .Z(n3336) );
  ANDN U3198 ( .B(n2836), .A(n3282), .Z(n3513) );
  ANDN U3199 ( .B(n2863), .A(n3301), .Z(n3533) );
  AND U3200 ( .A(n2911), .B(n3346), .Z(n3568) );
  AND U3201 ( .A(n3932), .B(n2949), .Z(n3931) );
  AND U3202 ( .A(n3934), .B(n2983), .Z(n3933) );
  AND U3203 ( .A(n3938), .B(n3036), .Z(n3937) );
  AND U3204 ( .A(n3948), .B(n3148), .Z(n3947) );
  AND U3205 ( .A(n3967), .B(n4007), .Z(n4005) );
  AND U3206 ( .A(n4012), .B(n4013), .Z(n4011) );
  AND U3207 ( .A(n4073), .B(n1033), .Z(n4071) );
  AND U3208 ( .A(n4090), .B(n3185), .Z(n4088) );
  AND U3209 ( .A(n4095), .B(n3556), .Z(n4093) );
  ANDN U3210 ( .B(n4112), .A(n3922), .Z(n4110) );
  AND U3211 ( .A(n4042), .B(n1670), .Z(n4256) );
  AND U3212 ( .A(n1722), .B(n4045), .Z(n4260) );
  ANDN U3213 ( .B(n1770), .A(n4048), .Z(n4261) );
  ANDN U3214 ( .B(n2111), .A(n4076), .Z(n4276) );
  AND U3215 ( .A(n2236), .B(n4087), .Z(n4288) );
  AND U3216 ( .A(n4150), .B(n3117), .Z(n4341) );
  ANDN U3217 ( .B(n2001), .A(n2000), .Z(n5124) );
  ANDN U3218 ( .B(n1433), .A(n1432), .Z(n1430) );
  AND U3219 ( .A(n1539), .B(n1540), .Z(n1537) );
  AND U3220 ( .A(n1568), .B(n1569), .Z(n1566) );
  ANDN U3221 ( .B(n1593), .A(n1592), .Z(n1590) );
  AND U3222 ( .A(n1916), .B(n1917), .Z(n1914) );
  AND U3223 ( .A(n1822), .B(n1820), .Z(n2148) );
  AND U3224 ( .A(n2813), .B(n2814), .Z(n2811) );
  AND U3225 ( .A(n2904), .B(n2905), .Z(n2902) );
  AND U3226 ( .A(n3010), .B(n3011), .Z(n3008) );
  AND U3227 ( .A(n3427), .B(n3428), .Z(n3425) );
  AND U3228 ( .A(n3459), .B(n3460), .Z(n3457) );
  AND U3229 ( .A(n3586), .B(n3587), .Z(n3584) );
  AND U3230 ( .A(n3672), .B(n3673), .Z(n3670) );
  AND U3231 ( .A(n3724), .B(n1037), .Z(n3723) );
  ANDN U3232 ( .B(n3918), .A(n1212), .Z(n3917) );
  AND U3233 ( .A(n3991), .B(n1345), .Z(n3990) );
  XNOR U3234 ( .A(n1030), .B(n1031), .Z(out[9]) );
  ANDN U3235 ( .B(n1032), .A(n1033), .Z(n1030) );
  XNOR U3236 ( .A(n1034), .B(n1035), .Z(out[99]) );
  ANDN U3237 ( .B(n1036), .A(n1037), .Z(n1034) );
  XNOR U3238 ( .A(n1038), .B(n1039), .Z(out[999]) );
  ANDN U3239 ( .B(n1040), .A(n1041), .Z(n1038) );
  XOR U3240 ( .A(n1042), .B(n1043), .Z(out[998]) );
  NOR U3241 ( .A(n1044), .B(n1045), .Z(n1042) );
  XNOR U3242 ( .A(n1046), .B(n1047), .Z(out[997]) );
  NOR U3243 ( .A(n1048), .B(n1049), .Z(n1046) );
  XNOR U3244 ( .A(n1050), .B(n1051), .Z(out[996]) );
  ANDN U3245 ( .B(n1052), .A(n1053), .Z(n1050) );
  XNOR U3246 ( .A(n1054), .B(n1055), .Z(out[995]) );
  ANDN U3247 ( .B(n1056), .A(n1057), .Z(n1054) );
  XNOR U3248 ( .A(n1058), .B(n1059), .Z(out[994]) );
  ANDN U3249 ( .B(n1060), .A(n1061), .Z(n1058) );
  XNOR U3250 ( .A(n1062), .B(n1063), .Z(out[993]) );
  ANDN U3251 ( .B(n1064), .A(n1065), .Z(n1062) );
  XNOR U3252 ( .A(n1066), .B(n1067), .Z(out[992]) );
  AND U3253 ( .A(n1068), .B(n1069), .Z(n1066) );
  XNOR U3254 ( .A(n1070), .B(n1071), .Z(out[991]) );
  ANDN U3255 ( .B(n1072), .A(n1073), .Z(n1070) );
  XNOR U3256 ( .A(n1074), .B(n1075), .Z(out[990]) );
  NOR U3257 ( .A(n1076), .B(n1077), .Z(n1074) );
  XNOR U3258 ( .A(n1078), .B(n1079), .Z(out[98]) );
  AND U3259 ( .A(n1080), .B(n1081), .Z(n1078) );
  XNOR U3260 ( .A(n1082), .B(n1083), .Z(out[989]) );
  AND U3261 ( .A(n1084), .B(n1085), .Z(n1082) );
  XOR U3262 ( .A(n1086), .B(n1087), .Z(out[988]) );
  AND U3263 ( .A(n1088), .B(n1089), .Z(n1086) );
  XNOR U3264 ( .A(n1090), .B(n1091), .Z(out[987]) );
  AND U3265 ( .A(n1092), .B(n1093), .Z(n1090) );
  XNOR U3266 ( .A(n1094), .B(n1095), .Z(out[986]) );
  ANDN U3267 ( .B(n1096), .A(n1097), .Z(n1094) );
  XNOR U3268 ( .A(n1098), .B(n1099), .Z(out[985]) );
  NOR U3269 ( .A(n1100), .B(n1101), .Z(n1098) );
  XNOR U3270 ( .A(n1102), .B(n1103), .Z(out[984]) );
  ANDN U3271 ( .B(n1104), .A(n1105), .Z(n1102) );
  XNOR U3272 ( .A(n1106), .B(n1107), .Z(out[983]) );
  ANDN U3273 ( .B(n1108), .A(n1109), .Z(n1106) );
  XNOR U3274 ( .A(n1110), .B(n1111), .Z(out[982]) );
  NOR U3275 ( .A(n1112), .B(n1113), .Z(n1110) );
  XNOR U3276 ( .A(n1114), .B(n1115), .Z(out[981]) );
  ANDN U3277 ( .B(n1116), .A(n1117), .Z(n1114) );
  XNOR U3278 ( .A(n1118), .B(n1119), .Z(out[980]) );
  NOR U3279 ( .A(n1120), .B(n1121), .Z(n1118) );
  XNOR U3280 ( .A(n1122), .B(n1123), .Z(out[97]) );
  AND U3281 ( .A(n1124), .B(n1125), .Z(n1122) );
  XNOR U3282 ( .A(n1126), .B(n1127), .Z(out[979]) );
  ANDN U3283 ( .B(n1128), .A(n1129), .Z(n1126) );
  XNOR U3284 ( .A(n1130), .B(n1131), .Z(out[978]) );
  NOR U3285 ( .A(n1132), .B(n1133), .Z(n1130) );
  XNOR U3286 ( .A(n1134), .B(n1135), .Z(out[977]) );
  ANDN U3287 ( .B(n1136), .A(n1137), .Z(n1134) );
  XNOR U3288 ( .A(n1138), .B(n1139), .Z(out[976]) );
  ANDN U3289 ( .B(n1140), .A(n1141), .Z(n1138) );
  XNOR U3290 ( .A(n1142), .B(n1143), .Z(out[975]) );
  NOR U3291 ( .A(n1144), .B(n1145), .Z(n1142) );
  XNOR U3292 ( .A(n1146), .B(n1147), .Z(out[974]) );
  ANDN U3293 ( .B(n1148), .A(n1149), .Z(n1146) );
  XNOR U3294 ( .A(n1150), .B(n1151), .Z(out[973]) );
  ANDN U3295 ( .B(n1152), .A(n1153), .Z(n1150) );
  XOR U3296 ( .A(n1154), .B(n1155), .Z(out[972]) );
  NOR U3297 ( .A(n1156), .B(n1157), .Z(n1154) );
  XOR U3298 ( .A(n1158), .B(n1159), .Z(out[971]) );
  NOR U3299 ( .A(n1160), .B(n1161), .Z(n1158) );
  XNOR U3300 ( .A(n1162), .B(n1163), .Z(out[970]) );
  AND U3301 ( .A(n1164), .B(n1165), .Z(n1162) );
  XOR U3302 ( .A(n1166), .B(n1167), .Z(out[96]) );
  NOR U3303 ( .A(n1168), .B(n1169), .Z(n1166) );
  XNOR U3304 ( .A(n1170), .B(n1171), .Z(out[969]) );
  ANDN U3305 ( .B(n1172), .A(n1173), .Z(n1170) );
  XOR U3306 ( .A(n1174), .B(n1175), .Z(out[968]) );
  ANDN U3307 ( .B(n1176), .A(n1177), .Z(n1174) );
  XNOR U3308 ( .A(n1178), .B(n1179), .Z(out[967]) );
  ANDN U3309 ( .B(n1180), .A(n1181), .Z(n1178) );
  XNOR U3310 ( .A(n1182), .B(n1183), .Z(out[966]) );
  ANDN U3311 ( .B(n1184), .A(n1185), .Z(n1182) );
  XOR U3312 ( .A(n1186), .B(n1187), .Z(out[965]) );
  NOR U3313 ( .A(n1188), .B(n1189), .Z(n1186) );
  XNOR U3314 ( .A(n1190), .B(n1191), .Z(out[964]) );
  NOR U3315 ( .A(n1192), .B(n1193), .Z(n1190) );
  XOR U3316 ( .A(n1194), .B(n1195), .Z(out[963]) );
  NOR U3317 ( .A(n1196), .B(n1197), .Z(n1194) );
  XNOR U3318 ( .A(n1198), .B(n1199), .Z(out[962]) );
  AND U3319 ( .A(n1200), .B(n1201), .Z(n1198) );
  XNOR U3320 ( .A(n1202), .B(n1203), .Z(out[961]) );
  AND U3321 ( .A(n1204), .B(n1205), .Z(n1202) );
  XNOR U3322 ( .A(n1206), .B(n1207), .Z(out[960]) );
  NOR U3323 ( .A(n1208), .B(n1209), .Z(n1206) );
  XNOR U3324 ( .A(n1210), .B(n1211), .Z(out[95]) );
  AND U3325 ( .A(n1212), .B(n1213), .Z(n1210) );
  XNOR U3326 ( .A(n1214), .B(n1215), .Z(out[959]) );
  ANDN U3327 ( .B(n1216), .A(n1217), .Z(n1214) );
  XNOR U3328 ( .A(n1218), .B(n1219), .Z(out[958]) );
  ANDN U3329 ( .B(n1220), .A(n1221), .Z(n1218) );
  XNOR U3330 ( .A(n1222), .B(n1223), .Z(out[957]) );
  ANDN U3331 ( .B(n1224), .A(n1225), .Z(n1222) );
  XNOR U3332 ( .A(n1226), .B(n1227), .Z(out[956]) );
  ANDN U3333 ( .B(n1228), .A(n1229), .Z(n1226) );
  XNOR U3334 ( .A(n1230), .B(n1231), .Z(out[955]) );
  ANDN U3335 ( .B(n1232), .A(n1233), .Z(n1230) );
  XNOR U3336 ( .A(n1234), .B(n1235), .Z(out[954]) );
  ANDN U3337 ( .B(n1236), .A(n1237), .Z(n1234) );
  XNOR U3338 ( .A(n1238), .B(n1239), .Z(out[953]) );
  AND U3339 ( .A(n1240), .B(n1241), .Z(n1238) );
  XOR U3340 ( .A(n1242), .B(n1243), .Z(out[952]) );
  NOR U3341 ( .A(n1244), .B(n1245), .Z(n1242) );
  XNOR U3342 ( .A(n1246), .B(n1247), .Z(out[951]) );
  AND U3343 ( .A(n1248), .B(n1249), .Z(n1246) );
  XNOR U3344 ( .A(n1250), .B(n1251), .Z(out[950]) );
  ANDN U3345 ( .B(n1252), .A(n1253), .Z(n1250) );
  XOR U3346 ( .A(n1254), .B(n1255), .Z(out[94]) );
  NOR U3347 ( .A(n1256), .B(n1257), .Z(n1254) );
  XNOR U3348 ( .A(n1258), .B(n1259), .Z(out[949]) );
  AND U3349 ( .A(n1260), .B(n1261), .Z(n1258) );
  XNOR U3350 ( .A(n1262), .B(n1263), .Z(out[948]) );
  ANDN U3351 ( .B(n1264), .A(n1265), .Z(n1262) );
  XNOR U3352 ( .A(n1266), .B(n1267), .Z(out[947]) );
  ANDN U3353 ( .B(n1268), .A(n1269), .Z(n1266) );
  XNOR U3354 ( .A(n1270), .B(n1271), .Z(out[946]) );
  ANDN U3355 ( .B(n1272), .A(n1273), .Z(n1270) );
  XNOR U3356 ( .A(n1274), .B(n1275), .Z(out[945]) );
  AND U3357 ( .A(n1276), .B(n1277), .Z(n1274) );
  XOR U3358 ( .A(n1278), .B(n1279), .Z(out[944]) );
  NOR U3359 ( .A(n1280), .B(n1281), .Z(n1278) );
  NOR U3360 ( .A(n1284), .B(n1285), .Z(n1282) );
  XOR U3361 ( .A(n1286), .B(n1287), .Z(out[942]) );
  NOR U3362 ( .A(n1288), .B(n1289), .Z(n1286) );
  NOR U3363 ( .A(n1292), .B(n1293), .Z(n1290) );
  XOR U3364 ( .A(n1294), .B(n1295), .Z(out[940]) );
  NOR U3365 ( .A(n1296), .B(n1297), .Z(n1294) );
  XNOR U3366 ( .A(n1298), .B(n1299), .Z(out[93]) );
  AND U3367 ( .A(n1300), .B(n1301), .Z(n1298) );
  XOR U3368 ( .A(n1302), .B(n1303), .Z(out[939]) );
  ANDN U3369 ( .B(n1304), .A(n1305), .Z(n1302) );
  XOR U3370 ( .A(n1306), .B(n1307), .Z(out[938]) );
  NOR U3371 ( .A(n1308), .B(n1309), .Z(n1306) );
  XNOR U3372 ( .A(n1310), .B(n1311), .Z(out[937]) );
  ANDN U3373 ( .B(n1312), .A(n1313), .Z(n1310) );
  XOR U3374 ( .A(n1314), .B(n1315), .Z(out[936]) );
  NOR U3375 ( .A(n1316), .B(n1317), .Z(n1314) );
  NOR U3376 ( .A(n1320), .B(n1321), .Z(n1318) );
  XNOR U3377 ( .A(n1322), .B(n1323), .Z(out[934]) );
  ANDN U3378 ( .B(n1324), .A(n1325), .Z(n1322) );
  XNOR U3379 ( .A(n1326), .B(n1327), .Z(out[933]) );
  ANDN U3380 ( .B(n1328), .A(n1329), .Z(n1326) );
  XOR U3381 ( .A(n1330), .B(n1331), .Z(out[932]) );
  ANDN U3382 ( .B(n1332), .A(n1333), .Z(n1330) );
  XNOR U3383 ( .A(n1334), .B(n1335), .Z(out[931]) );
  XOR U3384 ( .A(n1338), .B(n1339), .Z(out[930]) );
  ANDN U3385 ( .B(n1340), .A(n1341), .Z(n1338) );
  XNOR U3386 ( .A(n1342), .B(n1343), .Z(out[92]) );
  ANDN U3387 ( .B(n1344), .A(n1345), .Z(n1342) );
  XOR U3388 ( .A(n1346), .B(n1347), .Z(out[929]) );
  ANDN U3389 ( .B(n1348), .A(n1349), .Z(n1346) );
  XOR U3390 ( .A(n1350), .B(n1351), .Z(out[928]) );
  ANDN U3391 ( .B(n1352), .A(n1353), .Z(n1350) );
  XNOR U3392 ( .A(n1354), .B(n1355), .Z(out[927]) );
  XNOR U3393 ( .A(n1358), .B(n1359), .Z(out[926]) );
  XNOR U3394 ( .A(n1362), .B(n1363), .Z(out[925]) );
  ANDN U3395 ( .B(n1364), .A(n1365), .Z(n1362) );
  XOR U3396 ( .A(n1366), .B(n1367), .Z(out[924]) );
  ANDN U3397 ( .B(n1368), .A(n1369), .Z(n1366) );
  XOR U3398 ( .A(n1370), .B(n1371), .Z(out[923]) );
  ANDN U3399 ( .B(n1372), .A(n1373), .Z(n1370) );
  XNOR U3400 ( .A(n1374), .B(n1375), .Z(out[922]) );
  ANDN U3401 ( .B(n1376), .A(n1377), .Z(n1374) );
  XNOR U3402 ( .A(n1378), .B(n1379), .Z(out[921]) );
  XOR U3403 ( .A(n1382), .B(n1383), .Z(out[920]) );
  NOR U3404 ( .A(n1384), .B(n1385), .Z(n1382) );
  XNOR U3405 ( .A(n1386), .B(n1387), .Z(out[91]) );
  ANDN U3406 ( .B(n1388), .A(n1389), .Z(n1386) );
  XNOR U3407 ( .A(n1390), .B(n1391), .Z(out[919]) );
  AND U3408 ( .A(n1392), .B(n1393), .Z(n1390) );
  XNOR U3409 ( .A(n1394), .B(n1395), .Z(out[918]) );
  AND U3410 ( .A(n1396), .B(n1397), .Z(n1394) );
  XNOR U3411 ( .A(n1398), .B(n1399), .Z(out[917]) );
  AND U3412 ( .A(n1400), .B(n1401), .Z(n1398) );
  XNOR U3413 ( .A(n1402), .B(n1403), .Z(out[916]) );
  ANDN U3414 ( .B(n1404), .A(n1405), .Z(n1402) );
  XOR U3415 ( .A(n1406), .B(n1407), .Z(out[915]) );
  NOR U3416 ( .A(n1408), .B(n1409), .Z(n1406) );
  XNOR U3417 ( .A(n1410), .B(n1411), .Z(out[914]) );
  ANDN U3418 ( .B(n1412), .A(n1413), .Z(n1410) );
  ANDN U3419 ( .B(n1416), .A(n1417), .Z(n1414) );
  XNOR U3420 ( .A(n1418), .B(n1419), .Z(out[912]) );
  AND U3421 ( .A(n1420), .B(n1421), .Z(n1418) );
  XNOR U3422 ( .A(n1422), .B(n1423), .Z(out[911]) );
  AND U3423 ( .A(n1424), .B(n1425), .Z(n1422) );
  XNOR U3424 ( .A(n1426), .B(n1427), .Z(out[910]) );
  AND U3425 ( .A(n1428), .B(n1429), .Z(n1426) );
  XOR U3426 ( .A(n1430), .B(n1431), .Z(out[90]) );
  XNOR U3427 ( .A(n1434), .B(n1435), .Z(out[909]) );
  ANDN U3428 ( .B(n1436), .A(n1437), .Z(n1434) );
  XNOR U3429 ( .A(n1438), .B(n1439), .Z(out[908]) );
  AND U3430 ( .A(n1440), .B(n1441), .Z(n1438) );
  XOR U3431 ( .A(n1442), .B(n1443), .Z(out[907]) );
  NOR U3432 ( .A(n1444), .B(n1445), .Z(n1442) );
  ANDN U3433 ( .B(n1448), .A(n1449), .Z(n1446) );
  XNOR U3434 ( .A(n1450), .B(n1451), .Z(out[905]) );
  AND U3435 ( .A(n1452), .B(n1453), .Z(n1450) );
  XOR U3436 ( .A(n1454), .B(n1455), .Z(out[904]) );
  AND U3437 ( .A(n1456), .B(n1457), .Z(n1454) );
  XNOR U3438 ( .A(n1458), .B(n1459), .Z(out[903]) );
  AND U3439 ( .A(n1460), .B(n1461), .Z(n1458) );
  XNOR U3440 ( .A(n1462), .B(n1463), .Z(out[902]) );
  ANDN U3441 ( .B(n1464), .A(n1465), .Z(n1462) );
  XNOR U3442 ( .A(n1466), .B(n1467), .Z(out[901]) );
  AND U3443 ( .A(n1468), .B(n1469), .Z(n1466) );
  XNOR U3444 ( .A(n1470), .B(n1471), .Z(out[900]) );
  ANDN U3445 ( .B(n1472), .A(n1473), .Z(n1470) );
  XOR U3446 ( .A(n1474), .B(n1475), .Z(out[8]) );
  ANDN U3447 ( .B(n1476), .A(n1477), .Z(n1474) );
  XNOR U3448 ( .A(n1478), .B(n1479), .Z(out[89]) );
  AND U3449 ( .A(n1480), .B(n1481), .Z(n1478) );
  XNOR U3450 ( .A(n1482), .B(n1483), .Z(out[899]) );
  AND U3451 ( .A(n1484), .B(n1485), .Z(n1482) );
  XNOR U3452 ( .A(n1486), .B(n1487), .Z(out[898]) );
  ANDN U3453 ( .B(n1488), .A(n1489), .Z(n1486) );
  XNOR U3454 ( .A(n1490), .B(n1491), .Z(out[897]) );
  ANDN U3455 ( .B(n1492), .A(n1493), .Z(n1490) );
  XNOR U3456 ( .A(n1494), .B(n1495), .Z(out[896]) );
  ANDN U3457 ( .B(n1496), .A(n1497), .Z(n1494) );
  XNOR U3458 ( .A(n1498), .B(n1216), .Z(out[895]) );
  ANDN U3459 ( .B(n1499), .A(n1500), .Z(n1498) );
  XNOR U3460 ( .A(n1501), .B(n1220), .Z(out[894]) );
  XOR U3461 ( .A(n1503), .B(n1225), .Z(out[893]) );
  ANDN U3462 ( .B(n1504), .A(n1224), .Z(n1503) );
  XNOR U3463 ( .A(n1505), .B(n1228), .Z(out[892]) );
  ANDN U3464 ( .B(n1229), .A(n1506), .Z(n1505) );
  XNOR U3465 ( .A(n1507), .B(n1232), .Z(out[891]) );
  ANDN U3466 ( .B(n1508), .A(n1509), .Z(n1507) );
  XNOR U3467 ( .A(n1510), .B(n1236), .Z(out[890]) );
  ANDN U3468 ( .B(n1511), .A(n1512), .Z(n1510) );
  XNOR U3469 ( .A(n1513), .B(n1514), .Z(out[88]) );
  AND U3470 ( .A(n1515), .B(n1516), .Z(n1513) );
  XNOR U3471 ( .A(n1517), .B(n1241), .Z(out[889]) );
  NOR U3472 ( .A(n1518), .B(n1240), .Z(n1517) );
  XOR U3473 ( .A(n1519), .B(n1245), .Z(out[888]) );
  ANDN U3474 ( .B(n1244), .A(n1520), .Z(n1519) );
  XNOR U3475 ( .A(n1521), .B(n1249), .Z(out[887]) );
  NOR U3476 ( .A(n1522), .B(n1248), .Z(n1521) );
  XNOR U3477 ( .A(n1523), .B(n1252), .Z(out[886]) );
  ANDN U3478 ( .B(n1253), .A(n1524), .Z(n1523) );
  XNOR U3479 ( .A(n1525), .B(n1261), .Z(out[885]) );
  NOR U3480 ( .A(n1526), .B(n1260), .Z(n1525) );
  XNOR U3481 ( .A(n1527), .B(n1264), .Z(out[884]) );
  ANDN U3482 ( .B(n1265), .A(n1528), .Z(n1527) );
  XNOR U3483 ( .A(n1529), .B(n1268), .Z(out[883]) );
  XNOR U3484 ( .A(n1531), .B(n1272), .Z(out[882]) );
  XNOR U3485 ( .A(n1533), .B(n1277), .Z(out[881]) );
  NOR U3486 ( .A(n1534), .B(n1276), .Z(n1533) );
  XOR U3487 ( .A(n1535), .B(n1281), .Z(out[880]) );
  XNOR U3488 ( .A(n1537), .B(n1538), .Z(out[87]) );
  XOR U3489 ( .A(n1541), .B(n1285), .Z(out[879]) );
  XOR U3490 ( .A(n1543), .B(n1289), .Z(out[878]) );
  ANDN U3491 ( .B(n1288), .A(n1544), .Z(n1543) );
  IV U3492 ( .A(n1545), .Z(n1288) );
  XOR U3493 ( .A(n1546), .B(n1293), .Z(out[877]) );
  ANDN U3494 ( .B(n1292), .A(n1547), .Z(n1546) );
  XOR U3495 ( .A(n1548), .B(n1297), .Z(out[876]) );
  ANDN U3496 ( .B(n1296), .A(n1549), .Z(n1548) );
  IV U3497 ( .A(n1550), .Z(n1296) );
  XOR U3498 ( .A(n1551), .B(n1305), .Z(out[875]) );
  NOR U3499 ( .A(n1552), .B(n1304), .Z(n1551) );
  XOR U3500 ( .A(n1553), .B(n1309), .Z(out[874]) );
  ANDN U3501 ( .B(n1308), .A(n1554), .Z(n1553) );
  IV U3502 ( .A(n1555), .Z(n1308) );
  XOR U3503 ( .A(n1556), .B(n1313), .Z(out[873]) );
  NOR U3504 ( .A(n1557), .B(n1312), .Z(n1556) );
  XOR U3505 ( .A(n1558), .B(n1317), .Z(out[872]) );
  ANDN U3506 ( .B(n1316), .A(n1559), .Z(n1558) );
  IV U3507 ( .A(n1560), .Z(n1316) );
  XOR U3508 ( .A(n1561), .B(n1321), .Z(out[871]) );
  ANDN U3509 ( .B(n1320), .A(n1562), .Z(n1561) );
  IV U3510 ( .A(n1563), .Z(n1320) );
  XNOR U3511 ( .A(n1564), .B(n1324), .Z(out[870]) );
  XNOR U3512 ( .A(n1566), .B(n1567), .Z(out[86]) );
  XNOR U3513 ( .A(n1570), .B(n1328), .Z(out[869]) );
  ANDN U3514 ( .B(n1329), .A(n1571), .Z(n1570) );
  XOR U3515 ( .A(n1572), .B(n1333), .Z(out[868]) );
  NOR U3516 ( .A(n1573), .B(n1332), .Z(n1572) );
  XNOR U3517 ( .A(n1574), .B(n1337), .Z(out[867]) );
  NOR U3518 ( .A(n1336), .B(n1575), .Z(n1574) );
  XOR U3519 ( .A(n1576), .B(n1341), .Z(out[866]) );
  NOR U3520 ( .A(n1577), .B(n1340), .Z(n1576) );
  XOR U3521 ( .A(n1578), .B(n1349), .Z(out[865]) );
  NOR U3522 ( .A(n1579), .B(n1348), .Z(n1578) );
  XOR U3523 ( .A(n1580), .B(n1353), .Z(out[864]) );
  NOR U3524 ( .A(n1581), .B(n1352), .Z(n1580) );
  XOR U3525 ( .A(n1582), .B(n1356), .Z(out[863]) );
  ANDN U3526 ( .B(n1357), .A(n1583), .Z(n1582) );
  XOR U3527 ( .A(n1584), .B(n1360), .Z(out[862]) );
  ANDN U3528 ( .B(n1361), .A(n1585), .Z(n1584) );
  XOR U3529 ( .A(n1586), .B(n1365), .Z(out[861]) );
  ANDN U3530 ( .B(n1587), .A(n1364), .Z(n1586) );
  XOR U3531 ( .A(n1588), .B(n1369), .Z(out[860]) );
  NOR U3532 ( .A(n1589), .B(n1368), .Z(n1588) );
  XOR U3533 ( .A(n1590), .B(n1591), .Z(out[85]) );
  XOR U3534 ( .A(n1594), .B(n1373), .Z(out[859]) );
  NOR U3535 ( .A(n1595), .B(n1372), .Z(n1594) );
  XOR U3536 ( .A(n1596), .B(n1377), .Z(out[858]) );
  NOR U3537 ( .A(n1597), .B(n1376), .Z(n1596) );
  XNOR U3538 ( .A(n1598), .B(n1381), .Z(out[857]) );
  ANDN U3539 ( .B(n1599), .A(n1380), .Z(n1598) );
  XOR U3540 ( .A(n1600), .B(n1385), .Z(out[856]) );
  XNOR U3541 ( .A(n1602), .B(n1393), .Z(out[855]) );
  ANDN U3542 ( .B(n1603), .A(n1392), .Z(n1602) );
  XNOR U3543 ( .A(n1604), .B(n1397), .Z(out[854]) );
  ANDN U3544 ( .B(n1605), .A(n1396), .Z(n1604) );
  XNOR U3545 ( .A(n1606), .B(n1401), .Z(out[853]) );
  ANDN U3546 ( .B(n1607), .A(n1400), .Z(n1606) );
  XNOR U3547 ( .A(n1608), .B(n1404), .Z(out[852]) );
  XOR U3548 ( .A(n1610), .B(n1409), .Z(out[851]) );
  XNOR U3549 ( .A(n1612), .B(n1412), .Z(out[850]) );
  ANDN U3550 ( .B(n1413), .A(n1613), .Z(n1612) );
  XNOR U3551 ( .A(n1614), .B(n1615), .Z(out[84]) );
  AND U3552 ( .A(n1616), .B(n1617), .Z(n1614) );
  XOR U3553 ( .A(n1618), .B(n1417), .Z(out[849]) );
  NOR U3554 ( .A(n1619), .B(n1416), .Z(n1618) );
  XNOR U3555 ( .A(n1620), .B(n1421), .Z(out[848]) );
  NOR U3556 ( .A(n1621), .B(n1420), .Z(n1620) );
  XNOR U3557 ( .A(n1622), .B(n1425), .Z(out[847]) );
  NOR U3558 ( .A(n1623), .B(n1424), .Z(n1622) );
  XNOR U3559 ( .A(n1624), .B(n1429), .Z(out[846]) );
  ANDN U3560 ( .B(n1625), .A(n1428), .Z(n1624) );
  XNOR U3561 ( .A(n1626), .B(n1436), .Z(out[845]) );
  ANDN U3562 ( .B(n1437), .A(n1627), .Z(n1626) );
  XNOR U3563 ( .A(n1628), .B(n1441), .Z(out[844]) );
  NOR U3564 ( .A(n1629), .B(n1440), .Z(n1628) );
  XOR U3565 ( .A(n1630), .B(n1445), .Z(out[843]) );
  ANDN U3566 ( .B(n1444), .A(n1631), .Z(n1630) );
  XNOR U3567 ( .A(n1632), .B(n1448), .Z(out[842]) );
  ANDN U3568 ( .B(n1449), .A(n1633), .Z(n1632) );
  XNOR U3569 ( .A(n1634), .B(n1453), .Z(out[841]) );
  ANDN U3570 ( .B(n1635), .A(n1452), .Z(n1634) );
  XNOR U3571 ( .A(n1636), .B(n1457), .Z(out[840]) );
  NOR U3572 ( .A(n1637), .B(n1456), .Z(n1636) );
  XNOR U3573 ( .A(n1638), .B(n1639), .Z(out[83]) );
  AND U3574 ( .A(n1640), .B(n1641), .Z(n1638) );
  XNOR U3575 ( .A(n1642), .B(n1461), .Z(out[839]) );
  ANDN U3576 ( .B(n1643), .A(n1460), .Z(n1642) );
  XNOR U3577 ( .A(n1644), .B(n1464), .Z(out[838]) );
  ANDN U3578 ( .B(n1465), .A(n1645), .Z(n1644) );
  XNOR U3579 ( .A(n1646), .B(n1469), .Z(out[837]) );
  NOR U3580 ( .A(n1647), .B(n1468), .Z(n1646) );
  XNOR U3581 ( .A(n1648), .B(n1472), .Z(out[836]) );
  ANDN U3582 ( .B(n1649), .A(n1650), .Z(n1648) );
  XNOR U3583 ( .A(n1651), .B(n1485), .Z(out[835]) );
  NOR U3584 ( .A(n1652), .B(n1484), .Z(n1651) );
  XNOR U3585 ( .A(n1653), .B(n1488), .Z(out[834]) );
  ANDN U3586 ( .B(n1654), .A(n1655), .Z(n1653) );
  XNOR U3587 ( .A(n1656), .B(n1492), .Z(out[833]) );
  XNOR U3588 ( .A(n1658), .B(n1496), .Z(out[832]) );
  XNOR U3589 ( .A(n1660), .B(n1217), .Z(out[831]) );
  IV U3590 ( .A(n1500), .Z(n1217) );
  XOR U3591 ( .A(n1661), .B(n1662), .Z(n1500) );
  ANDN U3592 ( .B(n1663), .A(n1499), .Z(n1660) );
  IV U3593 ( .A(n1664), .Z(n1499) );
  XNOR U3594 ( .A(n1665), .B(n1221), .Z(out[830]) );
  XOR U3595 ( .A(n1666), .B(n1667), .Z(n1221) );
  XOR U3596 ( .A(n1669), .B(n1670), .Z(out[82]) );
  ANDN U3597 ( .B(n1671), .A(n1672), .Z(n1669) );
  XOR U3598 ( .A(n1673), .B(n1224), .Z(out[829]) );
  XOR U3599 ( .A(n1674), .B(n1675), .Z(n1224) );
  ANDN U3600 ( .B(n1676), .A(n1504), .Z(n1673) );
  IV U3601 ( .A(n1677), .Z(n1504) );
  XNOR U3602 ( .A(n1678), .B(n1229), .Z(out[828]) );
  XOR U3603 ( .A(n1679), .B(n1680), .Z(n1229) );
  ANDN U3604 ( .B(n1681), .A(n1682), .Z(n1678) );
  XNOR U3605 ( .A(n1683), .B(n1233), .Z(out[827]) );
  IV U3606 ( .A(n1509), .Z(n1233) );
  XNOR U3607 ( .A(n1684), .B(n1685), .Z(n1509) );
  ANDN U3608 ( .B(n1686), .A(n1508), .Z(n1683) );
  XNOR U3609 ( .A(n1687), .B(n1237), .Z(out[826]) );
  IV U3610 ( .A(n1512), .Z(n1237) );
  XOR U3611 ( .A(n1688), .B(n1689), .Z(n1512) );
  ANDN U3612 ( .B(n1690), .A(n1511), .Z(n1687) );
  XOR U3613 ( .A(n1691), .B(n1240), .Z(out[825]) );
  XNOR U3614 ( .A(n1692), .B(n1693), .Z(n1240) );
  ANDN U3615 ( .B(n1694), .A(n1695), .Z(n1691) );
  XNOR U3616 ( .A(n1696), .B(n1244), .Z(out[824]) );
  XOR U3617 ( .A(n1697), .B(n1698), .Z(n1244) );
  ANDN U3618 ( .B(n1699), .A(n1700), .Z(n1696) );
  XOR U3619 ( .A(n1701), .B(n1248), .Z(out[823]) );
  XOR U3620 ( .A(n1702), .B(n1703), .Z(n1248) );
  ANDN U3621 ( .B(n1704), .A(n1705), .Z(n1701) );
  XNOR U3622 ( .A(n1706), .B(n1253), .Z(out[822]) );
  XNOR U3623 ( .A(n1707), .B(n1708), .Z(n1253) );
  ANDN U3624 ( .B(n1709), .A(n1710), .Z(n1706) );
  XOR U3625 ( .A(n1711), .B(n1260), .Z(out[821]) );
  XNOR U3626 ( .A(n1712), .B(n1713), .Z(n1260) );
  ANDN U3627 ( .B(n1714), .A(n1715), .Z(n1711) );
  XNOR U3628 ( .A(n1716), .B(n1265), .Z(out[820]) );
  XNOR U3629 ( .A(n1717), .B(n1718), .Z(n1265) );
  ANDN U3630 ( .B(n1719), .A(n1720), .Z(n1716) );
  XOR U3631 ( .A(n1721), .B(n1722), .Z(out[81]) );
  NOR U3632 ( .A(n1723), .B(n1724), .Z(n1721) );
  XNOR U3633 ( .A(n1725), .B(n1269), .Z(out[819]) );
  XOR U3634 ( .A(n1726), .B(n1727), .Z(n1269) );
  ANDN U3635 ( .B(n1728), .A(n1530), .Z(n1725) );
  IV U3636 ( .A(n1729), .Z(n1530) );
  XNOR U3637 ( .A(n1730), .B(n1273), .Z(out[818]) );
  XOR U3638 ( .A(n1731), .B(n1732), .Z(n1273) );
  NOR U3639 ( .A(n1532), .B(n1733), .Z(n1730) );
  XOR U3640 ( .A(n1734), .B(n1276), .Z(out[817]) );
  XOR U3641 ( .A(n1735), .B(n1736), .Z(n1276) );
  ANDN U3642 ( .B(n1737), .A(n1738), .Z(n1734) );
  XNOR U3643 ( .A(n1739), .B(n1280), .Z(out[816]) );
  XOR U3644 ( .A(n1740), .B(n1741), .Z(n1280) );
  NOR U3645 ( .A(n1742), .B(n1536), .Z(n1739) );
  XNOR U3646 ( .A(n1743), .B(n1284), .Z(out[815]) );
  XOR U3647 ( .A(n1744), .B(n1745), .Z(n1284) );
  NOR U3648 ( .A(n1746), .B(n1542), .Z(n1743) );
  XOR U3649 ( .A(n1747), .B(n1545), .Z(out[814]) );
  XOR U3650 ( .A(n1748), .B(n1749), .Z(n1545) );
  ANDN U3651 ( .B(n1750), .A(n1751), .Z(n1747) );
  XNOR U3652 ( .A(n1752), .B(n1292), .Z(out[813]) );
  XOR U3653 ( .A(n1753), .B(n1754), .Z(n1292) );
  ANDN U3654 ( .B(n1547), .A(n1755), .Z(n1752) );
  XOR U3655 ( .A(n1756), .B(n1550), .Z(out[812]) );
  XOR U3656 ( .A(n1757), .B(n1758), .Z(n1550) );
  ANDN U3657 ( .B(n1759), .A(n1760), .Z(n1756) );
  XOR U3658 ( .A(n1761), .B(n1304), .Z(out[811]) );
  XOR U3659 ( .A(n1762), .B(n1763), .Z(n1304) );
  AND U3660 ( .A(n1552), .B(n1764), .Z(n1761) );
  XOR U3661 ( .A(n1765), .B(n1555), .Z(out[810]) );
  XOR U3662 ( .A(n1766), .B(n1767), .Z(n1555) );
  XOR U3663 ( .A(n1769), .B(n1770), .Z(out[80]) );
  NOR U3664 ( .A(n1771), .B(n1772), .Z(n1769) );
  XOR U3665 ( .A(n1773), .B(n1312), .Z(out[809]) );
  XNOR U3666 ( .A(n1774), .B(n1775), .Z(n1312) );
  ANDN U3667 ( .B(n1557), .A(n1776), .Z(n1773) );
  IV U3668 ( .A(n1777), .Z(n1557) );
  XOR U3669 ( .A(n1778), .B(n1560), .Z(out[808]) );
  XOR U3670 ( .A(n1779), .B(n1780), .Z(n1560) );
  ANDN U3671 ( .B(n1559), .A(n1781), .Z(n1778) );
  IV U3672 ( .A(n1782), .Z(n1559) );
  XOR U3673 ( .A(n1783), .B(n1563), .Z(out[807]) );
  XOR U3674 ( .A(n1784), .B(n1785), .Z(n1563) );
  ANDN U3675 ( .B(n1562), .A(n1786), .Z(n1783) );
  IV U3676 ( .A(n1787), .Z(n1562) );
  XNOR U3677 ( .A(n1788), .B(n1325), .Z(out[806]) );
  XOR U3678 ( .A(n1789), .B(n1790), .Z(n1325) );
  ANDN U3679 ( .B(n1791), .A(n1565), .Z(n1788) );
  XNOR U3680 ( .A(n1792), .B(n1329), .Z(out[805]) );
  XOR U3681 ( .A(n1793), .B(n1794), .Z(n1329) );
  ANDN U3682 ( .B(n1795), .A(n1796), .Z(n1792) );
  XOR U3683 ( .A(n1797), .B(n1332), .Z(out[804]) );
  XOR U3684 ( .A(n1798), .B(n1799), .Z(n1332) );
  ANDN U3685 ( .B(n1800), .A(n1801), .Z(n1797) );
  XOR U3686 ( .A(n1802), .B(n1336), .Z(out[803]) );
  XOR U3687 ( .A(n1803), .B(n1804), .Z(n1336) );
  AND U3688 ( .A(n1575), .B(n1805), .Z(n1802) );
  XOR U3689 ( .A(n1806), .B(n1340), .Z(out[802]) );
  XOR U3690 ( .A(n1807), .B(n1808), .Z(n1340) );
  ANDN U3691 ( .B(n1577), .A(n1809), .Z(n1806) );
  XOR U3692 ( .A(n1810), .B(n1348), .Z(out[801]) );
  XNOR U3693 ( .A(n1811), .B(n1812), .Z(n1348) );
  AND U3694 ( .A(n1579), .B(n1813), .Z(n1810) );
  XOR U3695 ( .A(n1814), .B(n1352), .Z(out[800]) );
  XOR U3696 ( .A(n1815), .B(n1816), .Z(n1352) );
  ANDN U3697 ( .B(n1817), .A(n1818), .Z(n1814) );
  XNOR U3698 ( .A(n1819), .B(n1820), .Z(out[7]) );
  NOR U3699 ( .A(n1821), .B(n1822), .Z(n1819) );
  XOR U3700 ( .A(n1823), .B(n1824), .Z(out[79]) );
  NOR U3701 ( .A(n1825), .B(n1826), .Z(n1823) );
  XNOR U3702 ( .A(n1827), .B(n1357), .Z(out[799]) );
  XOR U3703 ( .A(n1828), .B(n1829), .Z(n1357) );
  AND U3704 ( .A(n1583), .B(n1830), .Z(n1827) );
  XNOR U3705 ( .A(n1831), .B(n1361), .Z(out[798]) );
  XOR U3706 ( .A(n1832), .B(n1833), .Z(n1361) );
  ANDN U3707 ( .B(n1834), .A(n1835), .Z(n1831) );
  XOR U3708 ( .A(n1836), .B(n1364), .Z(out[797]) );
  XNOR U3709 ( .A(n1837), .B(n1838), .Z(n1364) );
  ANDN U3710 ( .B(n1839), .A(n1587), .Z(n1836) );
  XOR U3711 ( .A(n1840), .B(n1368), .Z(out[796]) );
  XOR U3712 ( .A(n1841), .B(n1842), .Z(n1368) );
  ANDN U3713 ( .B(n1843), .A(n1844), .Z(n1840) );
  XOR U3714 ( .A(n1845), .B(n1372), .Z(out[795]) );
  XNOR U3715 ( .A(n1846), .B(n1847), .Z(n1372) );
  XOR U3716 ( .A(n1849), .B(n1376), .Z(out[794]) );
  XNOR U3717 ( .A(n1850), .B(n1851), .Z(n1376) );
  XOR U3718 ( .A(n1853), .B(n1380), .Z(out[793]) );
  XOR U3719 ( .A(n1854), .B(n1855), .Z(n1380) );
  ANDN U3720 ( .B(n1856), .A(n1599), .Z(n1853) );
  XNOR U3721 ( .A(n1857), .B(n1384), .Z(out[792]) );
  XOR U3722 ( .A(n1858), .B(n1859), .Z(n1384) );
  ANDN U3723 ( .B(n1860), .A(n1601), .Z(n1857) );
  XOR U3724 ( .A(n1861), .B(n1392), .Z(out[791]) );
  XOR U3725 ( .A(n1862), .B(n1863), .Z(n1392) );
  NOR U3726 ( .A(n1864), .B(n1603), .Z(n1861) );
  XOR U3727 ( .A(n1865), .B(n1396), .Z(out[790]) );
  XNOR U3728 ( .A(n1866), .B(n1867), .Z(n1396) );
  NOR U3729 ( .A(n1868), .B(n1605), .Z(n1865) );
  XNOR U3730 ( .A(n1869), .B(n1870), .Z(out[78]) );
  ANDN U3731 ( .B(n1871), .A(n1872), .Z(n1869) );
  XOR U3732 ( .A(n1873), .B(n1400), .Z(out[789]) );
  XNOR U3733 ( .A(n1874), .B(n1875), .Z(n1400) );
  ANDN U3734 ( .B(n1876), .A(n1607), .Z(n1873) );
  XNOR U3735 ( .A(n1877), .B(n1405), .Z(out[788]) );
  XOR U3736 ( .A(n1878), .B(n1879), .Z(n1405) );
  ANDN U3737 ( .B(n1880), .A(n1609), .Z(n1877) );
  XNOR U3738 ( .A(n1881), .B(n1408), .Z(out[787]) );
  XOR U3739 ( .A(n1882), .B(n1883), .Z(n1408) );
  NOR U3740 ( .A(n1884), .B(n1611), .Z(n1881) );
  XNOR U3741 ( .A(n1885), .B(n1413), .Z(out[786]) );
  XOR U3742 ( .A(n1886), .B(n1887), .Z(n1413) );
  ANDN U3743 ( .B(n1888), .A(n1889), .Z(n1885) );
  XOR U3744 ( .A(n1890), .B(n1416), .Z(out[785]) );
  XOR U3745 ( .A(n1891), .B(n1892), .Z(n1416) );
  ANDN U3746 ( .B(n1619), .A(n1893), .Z(n1890) );
  XOR U3747 ( .A(n1894), .B(n1420), .Z(out[784]) );
  XNOR U3748 ( .A(n1895), .B(n1896), .Z(n1420) );
  ANDN U3749 ( .B(n1621), .A(n1897), .Z(n1894) );
  XOR U3750 ( .A(n1898), .B(n1424), .Z(out[783]) );
  XNOR U3751 ( .A(n1899), .B(n1900), .Z(n1424) );
  XOR U3752 ( .A(n1902), .B(n1428), .Z(out[782]) );
  XOR U3753 ( .A(n1903), .B(n1904), .Z(n1428) );
  ANDN U3754 ( .B(n1905), .A(n1625), .Z(n1902) );
  XNOR U3755 ( .A(n1906), .B(n1437), .Z(out[781]) );
  XOR U3756 ( .A(n1907), .B(n1908), .Z(n1437) );
  AND U3757 ( .A(n1627), .B(n1909), .Z(n1906) );
  XOR U3758 ( .A(n1910), .B(n1440), .Z(out[780]) );
  XNOR U3759 ( .A(n1911), .B(n1912), .Z(n1440) );
  XNOR U3760 ( .A(n1914), .B(n1915), .Z(out[77]) );
  XNOR U3761 ( .A(n1918), .B(n1444), .Z(out[779]) );
  XOR U3762 ( .A(n1919), .B(n1920), .Z(n1444) );
  ANDN U3763 ( .B(n1631), .A(n1921), .Z(n1918) );
  XNOR U3764 ( .A(n1922), .B(n1449), .Z(out[778]) );
  XOR U3765 ( .A(n1923), .B(n1924), .Z(n1449) );
  ANDN U3766 ( .B(n1925), .A(n1926), .Z(n1922) );
  XOR U3767 ( .A(n1927), .B(n1452), .Z(out[777]) );
  XOR U3768 ( .A(n1928), .B(n1929), .Z(n1452) );
  ANDN U3769 ( .B(n1930), .A(n1635), .Z(n1927) );
  XOR U3770 ( .A(n1931), .B(n1456), .Z(out[776]) );
  XOR U3771 ( .A(n1932), .B(n1933), .Z(n1456) );
  ANDN U3772 ( .B(n1934), .A(n1935), .Z(n1931) );
  XOR U3773 ( .A(n1936), .B(n1460), .Z(out[775]) );
  XOR U3774 ( .A(n1937), .B(n1938), .Z(n1460) );
  ANDN U3775 ( .B(n1939), .A(n1643), .Z(n1936) );
  XNOR U3776 ( .A(n1940), .B(n1465), .Z(out[774]) );
  XNOR U3777 ( .A(n1941), .B(n1942), .Z(n1465) );
  ANDN U3778 ( .B(n1943), .A(n1944), .Z(n1940) );
  XOR U3779 ( .A(n1945), .B(n1468), .Z(out[773]) );
  XNOR U3780 ( .A(n1946), .B(n1947), .Z(n1468) );
  ANDN U3781 ( .B(n1948), .A(n1949), .Z(n1945) );
  XNOR U3782 ( .A(n1950), .B(n1473), .Z(out[772]) );
  IV U3783 ( .A(n1650), .Z(n1473) );
  XNOR U3784 ( .A(n1951), .B(n1952), .Z(n1650) );
  NOR U3785 ( .A(n1953), .B(n1649), .Z(n1950) );
  XOR U3786 ( .A(n1954), .B(n1484), .Z(out[771]) );
  XOR U3787 ( .A(n1955), .B(n1956), .Z(n1484) );
  ANDN U3788 ( .B(n1957), .A(n1958), .Z(n1954) );
  XNOR U3789 ( .A(n1959), .B(n1489), .Z(out[770]) );
  IV U3790 ( .A(n1655), .Z(n1489) );
  XOR U3791 ( .A(n1960), .B(n1961), .Z(n1655) );
  ANDN U3792 ( .B(n1962), .A(n1654), .Z(n1959) );
  XNOR U3793 ( .A(n1963), .B(n1964), .Z(out[76]) );
  ANDN U3794 ( .B(n1965), .A(n1966), .Z(n1963) );
  XNOR U3795 ( .A(n1967), .B(n1493), .Z(out[769]) );
  XOR U3796 ( .A(n1968), .B(n1969), .Z(n1493) );
  ANDN U3797 ( .B(n1970), .A(n1657), .Z(n1967) );
  XNOR U3798 ( .A(n1971), .B(n1497), .Z(out[768]) );
  XOR U3799 ( .A(n1972), .B(n1973), .Z(n1497) );
  NOR U3800 ( .A(n1974), .B(n1659), .Z(n1971) );
  XNOR U3801 ( .A(n1975), .B(n1664), .Z(out[767]) );
  XOR U3802 ( .A(n1976), .B(n1977), .Z(n1664) );
  NOR U3803 ( .A(n1215), .B(n1663), .Z(n1975) );
  XOR U3804 ( .A(n1978), .B(n1502), .Z(out[766]) );
  XOR U3805 ( .A(n1979), .B(n1980), .Z(n1502) );
  ANDN U3806 ( .B(n1668), .A(n1219), .Z(n1978) );
  XNOR U3807 ( .A(n1981), .B(n1677), .Z(out[765]) );
  XOR U3808 ( .A(n1982), .B(n1983), .Z(n1677) );
  NOR U3809 ( .A(n1223), .B(n1676), .Z(n1981) );
  XNOR U3810 ( .A(n1984), .B(n1506), .Z(out[764]) );
  IV U3811 ( .A(n1682), .Z(n1506) );
  XNOR U3812 ( .A(n1985), .B(n1986), .Z(n1682) );
  NOR U3813 ( .A(n1681), .B(n1227), .Z(n1984) );
  XOR U3814 ( .A(n1987), .B(n1508), .Z(out[763]) );
  XOR U3815 ( .A(n1988), .B(n1989), .Z(n1508) );
  NOR U3816 ( .A(n1686), .B(n1231), .Z(n1987) );
  XOR U3817 ( .A(n1990), .B(n1511), .Z(out[762]) );
  XNOR U3818 ( .A(n1991), .B(n1992), .Z(n1511) );
  NOR U3819 ( .A(n1690), .B(n1235), .Z(n1990) );
  XNOR U3820 ( .A(n1993), .B(n1518), .Z(out[761]) );
  IV U3821 ( .A(n1695), .Z(n1518) );
  XOR U3822 ( .A(n1994), .B(n1995), .Z(n1695) );
  NOR U3823 ( .A(n1694), .B(n1239), .Z(n1993) );
  XNOR U3824 ( .A(n1996), .B(n1520), .Z(out[760]) );
  IV U3825 ( .A(n1700), .Z(n1520) );
  XNOR U3826 ( .A(n1997), .B(n1998), .Z(n1700) );
  XOR U3827 ( .A(n1999), .B(n2000), .Z(out[75]) );
  NOR U3828 ( .A(n2001), .B(n2002), .Z(n1999) );
  XNOR U3829 ( .A(n2003), .B(n1522), .Z(out[759]) );
  IV U3830 ( .A(n1705), .Z(n1522) );
  XOR U3831 ( .A(n2004), .B(n2005), .Z(n1705) );
  NOR U3832 ( .A(n1704), .B(n1247), .Z(n2003) );
  IV U3833 ( .A(n2006), .Z(n1704) );
  XNOR U3834 ( .A(n2007), .B(n1524), .Z(out[758]) );
  IV U3835 ( .A(n1710), .Z(n1524) );
  XOR U3836 ( .A(n2008), .B(n2009), .Z(n1710) );
  NOR U3837 ( .A(n1709), .B(n1251), .Z(n2007) );
  XNOR U3838 ( .A(n2010), .B(n1526), .Z(out[757]) );
  IV U3839 ( .A(n1715), .Z(n1526) );
  XNOR U3840 ( .A(n2011), .B(n2012), .Z(n1715) );
  NOR U3841 ( .A(n1714), .B(n1259), .Z(n2010) );
  XNOR U3842 ( .A(n2013), .B(n1528), .Z(out[756]) );
  IV U3843 ( .A(n1720), .Z(n1528) );
  XNOR U3844 ( .A(n2014), .B(n2015), .Z(n1720) );
  NOR U3845 ( .A(n1719), .B(n1263), .Z(n2013) );
  IV U3846 ( .A(n2016), .Z(n1719) );
  XNOR U3847 ( .A(n2017), .B(n1729), .Z(out[755]) );
  XOR U3848 ( .A(n2018), .B(n2019), .Z(n1729) );
  NOR U3849 ( .A(n1728), .B(n1267), .Z(n2017) );
  XOR U3850 ( .A(n2020), .B(n1532), .Z(out[754]) );
  XNOR U3851 ( .A(n2021), .B(n2022), .Z(n1532) );
  ANDN U3852 ( .B(n1733), .A(n1271), .Z(n2020) );
  XNOR U3853 ( .A(n2023), .B(n1534), .Z(out[753]) );
  IV U3854 ( .A(n1738), .Z(n1534) );
  XOR U3855 ( .A(n2024), .B(n2025), .Z(n1738) );
  NOR U3856 ( .A(n1737), .B(n1275), .Z(n2023) );
  XOR U3857 ( .A(n2026), .B(n1536), .Z(out[752]) );
  XOR U3858 ( .A(n2027), .B(n2028), .Z(n1536) );
  XOR U3859 ( .A(n2029), .B(n1542), .Z(out[751]) );
  XNOR U3860 ( .A(n2030), .B(n2031), .Z(n1542) );
  XNOR U3861 ( .A(n2032), .B(n1544), .Z(out[750]) );
  IV U3862 ( .A(n1751), .Z(n1544) );
  XOR U3863 ( .A(n2033), .B(n2034), .Z(n1751) );
  ANDN U3864 ( .B(n1287), .A(n1750), .Z(n2032) );
  XOR U3865 ( .A(n2035), .B(n2036), .Z(out[74]) );
  ANDN U3866 ( .B(n2037), .A(n2038), .Z(n2035) );
  XNOR U3867 ( .A(n2039), .B(n1547), .Z(out[749]) );
  XOR U3868 ( .A(n2040), .B(n2041), .Z(n1547) );
  ANDN U3869 ( .B(n1291), .A(n2042), .Z(n2039) );
  XNOR U3870 ( .A(n2043), .B(n1549), .Z(out[748]) );
  IV U3871 ( .A(n1760), .Z(n1549) );
  XNOR U3872 ( .A(n2044), .B(n2045), .Z(n1760) );
  NOR U3873 ( .A(n2046), .B(n1759), .Z(n2043) );
  XNOR U3874 ( .A(n2047), .B(n1552), .Z(out[747]) );
  XNOR U3875 ( .A(n2048), .B(n2049), .Z(n1552) );
  NOR U3876 ( .A(n2050), .B(n1764), .Z(n2047) );
  XNOR U3877 ( .A(n2051), .B(n1554), .Z(out[746]) );
  XOR U3878 ( .A(n2052), .B(n2053), .Z(n1554) );
  ANDN U3879 ( .B(n1307), .A(n1768), .Z(n2051) );
  XOR U3880 ( .A(n2054), .B(n1777), .Z(out[745]) );
  XOR U3881 ( .A(n2055), .B(n2056), .Z(n1777) );
  ANDN U3882 ( .B(n1776), .A(n1311), .Z(n2054) );
  XOR U3883 ( .A(n2057), .B(n1782), .Z(out[744]) );
  XOR U3884 ( .A(n2058), .B(n2059), .Z(n1782) );
  ANDN U3885 ( .B(n1781), .A(n2060), .Z(n2057) );
  XOR U3886 ( .A(n2061), .B(n1787), .Z(out[743]) );
  XOR U3887 ( .A(n2062), .B(n2063), .Z(n1787) );
  XOR U3888 ( .A(n2064), .B(n1565), .Z(out[742]) );
  XNOR U3889 ( .A(n2065), .B(n2066), .Z(n1565) );
  NOR U3890 ( .A(n1791), .B(n1323), .Z(n2064) );
  XNOR U3891 ( .A(n2067), .B(n1571), .Z(out[741]) );
  IV U3892 ( .A(n1796), .Z(n1571) );
  XOR U3893 ( .A(n2068), .B(n2069), .Z(n1796) );
  NOR U3894 ( .A(n1795), .B(n1327), .Z(n2067) );
  XNOR U3895 ( .A(n2070), .B(n1573), .Z(out[740]) );
  IV U3896 ( .A(n1801), .Z(n1573) );
  XNOR U3897 ( .A(n2071), .B(n2072), .Z(n1801) );
  NOR U3898 ( .A(n2073), .B(n1800), .Z(n2070) );
  XNOR U3899 ( .A(n2074), .B(n2075), .Z(out[73]) );
  ANDN U3900 ( .B(n1031), .A(n1032), .Z(n2074) );
  IV U3901 ( .A(n2076), .Z(n1032) );
  XNOR U3902 ( .A(n2077), .B(n1575), .Z(out[739]) );
  XNOR U3903 ( .A(n2078), .B(n2079), .Z(n1575) );
  NOR U3904 ( .A(n1805), .B(n1335), .Z(n2077) );
  XNOR U3905 ( .A(n2080), .B(n1577), .Z(out[738]) );
  XOR U3906 ( .A(n2081), .B(n2082), .Z(n1577) );
  ANDN U3907 ( .B(n1339), .A(n2083), .Z(n2080) );
  XNOR U3908 ( .A(n2084), .B(n1579), .Z(out[737]) );
  XNOR U3909 ( .A(n2085), .B(n2086), .Z(n1579) );
  ANDN U3910 ( .B(n1347), .A(n1813), .Z(n2084) );
  XNOR U3911 ( .A(n2087), .B(n1581), .Z(out[736]) );
  IV U3912 ( .A(n1818), .Z(n1581) );
  XOR U3913 ( .A(n2088), .B(n2089), .Z(n1818) );
  XNOR U3914 ( .A(n2090), .B(n1583), .Z(out[735]) );
  XNOR U3915 ( .A(n2091), .B(n2092), .Z(n1583) );
  NOR U3916 ( .A(n1830), .B(n1355), .Z(n2090) );
  XNOR U3917 ( .A(n2093), .B(n1585), .Z(out[734]) );
  IV U3918 ( .A(n1835), .Z(n1585) );
  XNOR U3919 ( .A(n2094), .B(n2095), .Z(n1835) );
  NOR U3920 ( .A(n1834), .B(n1359), .Z(n2093) );
  XOR U3921 ( .A(n2096), .B(n1587), .Z(out[733]) );
  XNOR U3922 ( .A(n2097), .B(n2098), .Z(n1587) );
  NOR U3923 ( .A(n1363), .B(n1839), .Z(n2096) );
  XNOR U3924 ( .A(n2099), .B(n1589), .Z(out[732]) );
  IV U3925 ( .A(n1844), .Z(n1589) );
  XNOR U3926 ( .A(n2100), .B(n2101), .Z(n1844) );
  NOR U3927 ( .A(n2102), .B(n1843), .Z(n2099) );
  XNOR U3928 ( .A(n2103), .B(n1595), .Z(out[731]) );
  XOR U3929 ( .A(n2104), .B(n2105), .Z(n1595) );
  NOR U3930 ( .A(n2106), .B(n1848), .Z(n2103) );
  XNOR U3931 ( .A(n2107), .B(n1597), .Z(out[730]) );
  XOR U3932 ( .A(n2108), .B(n2109), .Z(n1597) );
  NOR U3933 ( .A(n1375), .B(n1852), .Z(n2107) );
  XOR U3934 ( .A(n2110), .B(n2111), .Z(out[72]) );
  ANDN U3935 ( .B(n1477), .A(n1475), .Z(n2110) );
  XOR U3936 ( .A(n2112), .B(n1599), .Z(out[729]) );
  XOR U3937 ( .A(n2113), .B(n2114), .Z(n1599) );
  NOR U3938 ( .A(n1856), .B(n1379), .Z(n2112) );
  XOR U3939 ( .A(n2115), .B(n1601), .Z(out[728]) );
  XNOR U3940 ( .A(n2116), .B(n2117), .Z(n1601) );
  NOR U3941 ( .A(n2118), .B(n1860), .Z(n2115) );
  XOR U3942 ( .A(n2119), .B(n1603), .Z(out[727]) );
  XNOR U3943 ( .A(n2120), .B(n2121), .Z(n1603) );
  NOR U3944 ( .A(n2122), .B(n1391), .Z(n2119) );
  XOR U3945 ( .A(n2123), .B(n1605), .Z(out[726]) );
  XNOR U3946 ( .A(n2124), .B(n2125), .Z(n1605) );
  ANDN U3947 ( .B(n1868), .A(n1395), .Z(n2123) );
  IV U3948 ( .A(n2126), .Z(n1395) );
  XOR U3949 ( .A(n2127), .B(n1607), .Z(out[725]) );
  XNOR U3950 ( .A(n2128), .B(n2129), .Z(n1607) );
  NOR U3951 ( .A(n1399), .B(n1876), .Z(n2127) );
  XOR U3952 ( .A(n2130), .B(n1609), .Z(out[724]) );
  XNOR U3953 ( .A(n2131), .B(n2132), .Z(n1609) );
  NOR U3954 ( .A(n1880), .B(n1403), .Z(n2130) );
  XOR U3955 ( .A(n2133), .B(n1611), .Z(out[723]) );
  XOR U3956 ( .A(n2134), .B(n2135), .Z(n1611) );
  ANDN U3957 ( .B(n1407), .A(n2136), .Z(n2133) );
  XNOR U3958 ( .A(n2137), .B(n1613), .Z(out[722]) );
  IV U3959 ( .A(n1889), .Z(n1613) );
  XNOR U3960 ( .A(n2138), .B(n2139), .Z(n1889) );
  NOR U3961 ( .A(n1888), .B(n1411), .Z(n2137) );
  XNOR U3962 ( .A(n2140), .B(n1619), .Z(out[721]) );
  XOR U3963 ( .A(n2141), .B(n2142), .Z(n1619) );
  ANDN U3964 ( .B(n1415), .A(n2143), .Z(n2140) );
  XNOR U3965 ( .A(n2144), .B(n1621), .Z(out[720]) );
  XNOR U3966 ( .A(n2145), .B(n2146), .Z(n1621) );
  NOR U3967 ( .A(n2147), .B(n1419), .Z(n2144) );
  XNOR U3968 ( .A(n2148), .B(n2149), .Z(out[71]) );
  XNOR U3969 ( .A(n2150), .B(n1623), .Z(out[719]) );
  XNOR U3970 ( .A(n2151), .B(n2152), .Z(n1623) );
  NOR U3971 ( .A(n1901), .B(n1423), .Z(n2150) );
  XOR U3972 ( .A(n2153), .B(n1625), .Z(out[718]) );
  XOR U3973 ( .A(n2154), .B(n2155), .Z(n1625) );
  NOR U3974 ( .A(n1427), .B(n1905), .Z(n2153) );
  XNOR U3975 ( .A(n2156), .B(n1627), .Z(out[717]) );
  XNOR U3976 ( .A(n2157), .B(n2158), .Z(n1627) );
  NOR U3977 ( .A(n1435), .B(n1909), .Z(n2156) );
  XNOR U3978 ( .A(n2159), .B(n1629), .Z(out[716]) );
  XNOR U3979 ( .A(n2160), .B(n2161), .Z(n1629) );
  NOR U3980 ( .A(n1913), .B(n1439), .Z(n2159) );
  XNOR U3981 ( .A(n2162), .B(n1631), .Z(out[715]) );
  XNOR U3982 ( .A(n2163), .B(n2164), .Z(n1631) );
  ANDN U3983 ( .B(n1921), .A(n2165), .Z(n2162) );
  IV U3984 ( .A(n2166), .Z(n1921) );
  XNOR U3985 ( .A(n2167), .B(n1633), .Z(out[714]) );
  IV U3986 ( .A(n1926), .Z(n1633) );
  XOR U3987 ( .A(n2168), .B(n2169), .Z(n1926) );
  ANDN U3988 ( .B(n1447), .A(n1925), .Z(n2167) );
  XOR U3989 ( .A(n2170), .B(n1635), .Z(out[713]) );
  XNOR U3990 ( .A(n2171), .B(n2172), .Z(n1635) );
  NOR U3991 ( .A(n1930), .B(n1451), .Z(n2170) );
  XNOR U3992 ( .A(n2173), .B(n1637), .Z(out[712]) );
  IV U3993 ( .A(n1935), .Z(n1637) );
  XOR U3994 ( .A(n2174), .B(n2175), .Z(n1935) );
  ANDN U3995 ( .B(n1455), .A(n1934), .Z(n2173) );
  XOR U3996 ( .A(n2176), .B(n1643), .Z(out[711]) );
  XNOR U3997 ( .A(n2177), .B(n2178), .Z(n1643) );
  NOR U3998 ( .A(n1939), .B(n1459), .Z(n2176) );
  XNOR U3999 ( .A(n2179), .B(n1645), .Z(out[710]) );
  IV U4000 ( .A(n1944), .Z(n1645) );
  XOR U4001 ( .A(n2180), .B(n2181), .Z(n1944) );
  NOR U4002 ( .A(n1943), .B(n1463), .Z(n2179) );
  XNOR U4003 ( .A(n2182), .B(n2183), .Z(out[70]) );
  AND U4004 ( .A(n2184), .B(n2185), .Z(n2182) );
  XNOR U4005 ( .A(n2186), .B(n1647), .Z(out[709]) );
  IV U4006 ( .A(n1949), .Z(n1647) );
  XNOR U4007 ( .A(n2187), .B(n2188), .Z(n1949) );
  NOR U4008 ( .A(n1948), .B(n1467), .Z(n2186) );
  XOR U4009 ( .A(n2189), .B(n1649), .Z(out[708]) );
  XNOR U4010 ( .A(n2190), .B(n2191), .Z(n1649) );
  XNOR U4011 ( .A(n2192), .B(n1652), .Z(out[707]) );
  IV U4012 ( .A(n1958), .Z(n1652) );
  XOR U4013 ( .A(n2193), .B(n2194), .Z(n1958) );
  NOR U4014 ( .A(n1483), .B(n1957), .Z(n2192) );
  XOR U4015 ( .A(n2195), .B(n1654), .Z(out[706]) );
  XOR U4016 ( .A(n2196), .B(n2197), .Z(n1654) );
  NOR U4017 ( .A(n1487), .B(n1962), .Z(n2195) );
  XOR U4018 ( .A(n2198), .B(n1657), .Z(out[705]) );
  XNOR U4019 ( .A(n2199), .B(n2200), .Z(n1657) );
  NOR U4020 ( .A(n1970), .B(n1491), .Z(n2198) );
  XOR U4021 ( .A(n2201), .B(n1659), .Z(out[704]) );
  XNOR U4022 ( .A(n2202), .B(n2203), .Z(n1659) );
  NOR U4023 ( .A(n2204), .B(n1495), .Z(n2201) );
  XOR U4024 ( .A(n2205), .B(n1663), .Z(out[703]) );
  XNOR U4025 ( .A(n2206), .B(n2207), .Z(n1663) );
  ANDN U4026 ( .B(n1215), .A(n1216), .Z(n2205) );
  XOR U4027 ( .A(n2208), .B(n2209), .Z(n1216) );
  XOR U4028 ( .A(n2210), .B(n2211), .Z(n1215) );
  XNOR U4029 ( .A(n2212), .B(n1668), .Z(out[702]) );
  XOR U4030 ( .A(n2213), .B(n2214), .Z(n1668) );
  ANDN U4031 ( .B(n1219), .A(n1220), .Z(n2212) );
  XOR U4032 ( .A(n2215), .B(n2216), .Z(n1220) );
  XNOR U4033 ( .A(n2217), .B(n2218), .Z(n1219) );
  XOR U4034 ( .A(n2219), .B(n1676), .Z(out[701]) );
  AND U4035 ( .A(n1225), .B(n1223), .Z(n2219) );
  XOR U4036 ( .A(n2222), .B(n2223), .Z(n1223) );
  XOR U4037 ( .A(n2224), .B(n2225), .Z(n1225) );
  XOR U4038 ( .A(n2226), .B(n1681), .Z(out[700]) );
  XNOR U4039 ( .A(n2227), .B(n2228), .Z(n1681) );
  ANDN U4040 ( .B(n1227), .A(n1228), .Z(n2226) );
  XOR U4041 ( .A(n2229), .B(n2230), .Z(n1228) );
  XOR U4042 ( .A(n2231), .B(n2232), .Z(n1227) );
  XNOR U4043 ( .A(n2233), .B(n2185), .Z(out[6]) );
  NOR U4044 ( .A(n2234), .B(n2184), .Z(n2233) );
  XOR U4045 ( .A(n2235), .B(n2236), .Z(out[69]) );
  NOR U4046 ( .A(n2237), .B(n2238), .Z(n2235) );
  XOR U4047 ( .A(n2239), .B(n1686), .Z(out[699]) );
  XNOR U4048 ( .A(n2240), .B(n2241), .Z(n1686) );
  ANDN U4049 ( .B(n1231), .A(n1232), .Z(n2239) );
  XNOR U4050 ( .A(n2242), .B(n2243), .Z(n1232) );
  XNOR U4051 ( .A(n2244), .B(n2245), .Z(n1231) );
  XOR U4052 ( .A(n2246), .B(n1690), .Z(out[698]) );
  XOR U4053 ( .A(n2247), .B(n2248), .Z(n1690) );
  ANDN U4054 ( .B(n1235), .A(n1236), .Z(n2246) );
  XOR U4055 ( .A(n2249), .B(n2250), .Z(n1236) );
  XNOR U4056 ( .A(n2251), .B(n2252), .Z(n1235) );
  XOR U4057 ( .A(n2253), .B(n1694), .Z(out[697]) );
  XOR U4058 ( .A(n2254), .B(n2255), .Z(n1694) );
  ANDN U4059 ( .B(n1239), .A(n1241), .Z(n2253) );
  XOR U4060 ( .A(n2256), .B(n2257), .Z(n1241) );
  XOR U4061 ( .A(n2258), .B(n2259), .Z(n1239) );
  XOR U4062 ( .A(n2260), .B(n1699), .Z(out[696]) );
  XOR U4063 ( .A(n2261), .B(n2262), .Z(n1699) );
  ANDN U4064 ( .B(n1245), .A(n1243), .Z(n2260) );
  XOR U4065 ( .A(n2263), .B(n2264), .Z(n1243) );
  XOR U4066 ( .A(n2265), .B(n2266), .Z(n1245) );
  XNOR U4067 ( .A(n2267), .B(n2006), .Z(out[695]) );
  XOR U4068 ( .A(n2268), .B(n2269), .Z(n2006) );
  ANDN U4069 ( .B(n1247), .A(n1249), .Z(n2267) );
  XOR U4070 ( .A(n2270), .B(n2271), .Z(n1249) );
  XOR U4071 ( .A(n2272), .B(n2273), .Z(n1247) );
  XOR U4072 ( .A(n2274), .B(n1709), .Z(out[694]) );
  XOR U4073 ( .A(n2275), .B(n2276), .Z(n1709) );
  ANDN U4074 ( .B(n1251), .A(n1252), .Z(n2274) );
  XOR U4075 ( .A(n2277), .B(n2278), .Z(n1252) );
  XOR U4076 ( .A(n2279), .B(n2280), .Z(n1251) );
  XOR U4077 ( .A(n2281), .B(n1714), .Z(out[693]) );
  XNOR U4078 ( .A(n2282), .B(n2283), .Z(n1714) );
  ANDN U4079 ( .B(n1259), .A(n1261), .Z(n2281) );
  XNOR U4080 ( .A(n2284), .B(n2285), .Z(n1261) );
  XOR U4081 ( .A(n2286), .B(n2287), .Z(n1259) );
  XNOR U4082 ( .A(n2288), .B(n2016), .Z(out[692]) );
  XOR U4083 ( .A(n2289), .B(n2290), .Z(n2016) );
  ANDN U4084 ( .B(n1263), .A(n1264), .Z(n2288) );
  XNOR U4085 ( .A(n2291), .B(n2292), .Z(n1264) );
  XOR U4086 ( .A(n2293), .B(n2294), .Z(n1263) );
  XOR U4087 ( .A(n2295), .B(n1728), .Z(out[691]) );
  XOR U4088 ( .A(n2296), .B(n2297), .Z(n1728) );
  ANDN U4089 ( .B(n1267), .A(n1268), .Z(n2295) );
  XNOR U4090 ( .A(n2298), .B(n2299), .Z(n1268) );
  XOR U4091 ( .A(n2300), .B(n2301), .Z(n1267) );
  XNOR U4092 ( .A(n2302), .B(n1733), .Z(out[690]) );
  XOR U4093 ( .A(n2303), .B(n2304), .Z(n1733) );
  ANDN U4094 ( .B(n1271), .A(n1272), .Z(n2302) );
  XOR U4095 ( .A(n2305), .B(n2306), .Z(n1272) );
  XNOR U4096 ( .A(n2307), .B(n2308), .Z(n1271) );
  XNOR U4097 ( .A(n2309), .B(n2310), .Z(out[68]) );
  AND U4098 ( .A(n2311), .B(n2312), .Z(n2309) );
  XOR U4099 ( .A(n2313), .B(n1737), .Z(out[689]) );
  XOR U4100 ( .A(n2314), .B(n2315), .Z(n1737) );
  ANDN U4101 ( .B(n1275), .A(n1277), .Z(n2313) );
  XOR U4102 ( .A(n2316), .B(n2317), .Z(n1277) );
  XOR U4103 ( .A(n2318), .B(n2319), .Z(n1275) );
  XNOR U4104 ( .A(n2320), .B(n1742), .Z(out[688]) );
  XNOR U4105 ( .A(n2321), .B(n2322), .Z(n1742) );
  ANDN U4106 ( .B(n1281), .A(n1279), .Z(n2320) );
  XOR U4107 ( .A(n2323), .B(n2324), .Z(n1279) );
  XNOR U4108 ( .A(n2325), .B(n2326), .Z(n1281) );
  XNOR U4109 ( .A(n2327), .B(n1746), .Z(out[687]) );
  XOR U4110 ( .A(n2328), .B(n2329), .Z(n1746) );
  ANDN U4111 ( .B(n1285), .A(n1283), .Z(n2327) );
  XOR U4112 ( .A(n2330), .B(n2331), .Z(n1283) );
  XOR U4113 ( .A(n2332), .B(n2333), .Z(n1285) );
  XOR U4114 ( .A(n2334), .B(n1750), .Z(out[686]) );
  XOR U4115 ( .A(n2335), .B(n2336), .Z(n1750) );
  ANDN U4116 ( .B(n1289), .A(n1287), .Z(n2334) );
  XOR U4117 ( .A(n2337), .B(n2338), .Z(n1287) );
  XOR U4118 ( .A(n2339), .B(n2340), .Z(n1289) );
  XNOR U4119 ( .A(n2341), .B(n1755), .Z(out[685]) );
  IV U4120 ( .A(n2042), .Z(n1755) );
  XOR U4121 ( .A(n2342), .B(n2343), .Z(n2042) );
  ANDN U4122 ( .B(n1293), .A(n1291), .Z(n2341) );
  XNOR U4123 ( .A(n2344), .B(n2345), .Z(n1291) );
  XOR U4124 ( .A(n2346), .B(n2347), .Z(n1293) );
  XOR U4125 ( .A(n2348), .B(n1759), .Z(out[684]) );
  XOR U4126 ( .A(n2349), .B(n2350), .Z(n1759) );
  ANDN U4127 ( .B(n1297), .A(n1295), .Z(n2348) );
  IV U4128 ( .A(n2046), .Z(n1295) );
  XOR U4129 ( .A(n2351), .B(n2352), .Z(n2046) );
  XOR U4130 ( .A(n2353), .B(n2354), .Z(n1297) );
  XOR U4131 ( .A(n2355), .B(n1764), .Z(out[683]) );
  XOR U4132 ( .A(n2356), .B(n2357), .Z(n1764) );
  ANDN U4133 ( .B(n1305), .A(n1303), .Z(n2355) );
  IV U4134 ( .A(n2050), .Z(n1303) );
  XOR U4135 ( .A(n2358), .B(n2359), .Z(n2050) );
  XNOR U4136 ( .A(n2360), .B(n2361), .Z(n1305) );
  XOR U4137 ( .A(n2362), .B(n1768), .Z(out[682]) );
  XOR U4138 ( .A(n2363), .B(n2364), .Z(n1768) );
  ANDN U4139 ( .B(n1309), .A(n1307), .Z(n2362) );
  XOR U4140 ( .A(n2365), .B(n2366), .Z(n1307) );
  XOR U4141 ( .A(n2367), .B(n2368), .Z(n1309) );
  XNOR U4142 ( .A(n2369), .B(n1776), .Z(out[681]) );
  XOR U4143 ( .A(n2370), .B(n2371), .Z(n1776) );
  AND U4144 ( .A(n1313), .B(n1311), .Z(n2369) );
  XNOR U4145 ( .A(n2372), .B(n2373), .Z(n1311) );
  XOR U4146 ( .A(n2374), .B(n2375), .Z(n1313) );
  XNOR U4147 ( .A(n2376), .B(n1781), .Z(out[680]) );
  XOR U4148 ( .A(n2377), .B(n2378), .Z(n1781) );
  ANDN U4149 ( .B(n1317), .A(n1315), .Z(n2376) );
  IV U4150 ( .A(n2060), .Z(n1315) );
  XOR U4151 ( .A(n2379), .B(n2380), .Z(n2060) );
  XNOR U4152 ( .A(n2381), .B(n2382), .Z(n1317) );
  XNOR U4153 ( .A(n2383), .B(n2384), .Z(out[67]) );
  ANDN U4154 ( .B(n2385), .A(n2386), .Z(n2383) );
  XNOR U4155 ( .A(n2387), .B(n1786), .Z(out[679]) );
  XOR U4156 ( .A(n2388), .B(n2389), .Z(n1786) );
  ANDN U4157 ( .B(n1321), .A(n1319), .Z(n2387) );
  XOR U4158 ( .A(n2390), .B(n2391), .Z(n1319) );
  XOR U4159 ( .A(n2392), .B(n2393), .Z(n1321) );
  XOR U4160 ( .A(n2394), .B(n1791), .Z(out[678]) );
  XOR U4161 ( .A(n2395), .B(n2396), .Z(n1791) );
  ANDN U4162 ( .B(n1323), .A(n1324), .Z(n2394) );
  XOR U4163 ( .A(n2397), .B(n2398), .Z(n1324) );
  XOR U4164 ( .A(n2399), .B(n2400), .Z(n1323) );
  XOR U4165 ( .A(n2401), .B(n1795), .Z(out[677]) );
  XNOR U4166 ( .A(n2402), .B(n2403), .Z(n1795) );
  ANDN U4167 ( .B(n1327), .A(n1328), .Z(n2401) );
  XOR U4168 ( .A(n2404), .B(n2405), .Z(n1328) );
  XOR U4169 ( .A(n2406), .B(n2407), .Z(n1327) );
  XOR U4170 ( .A(n2408), .B(n1800), .Z(out[676]) );
  XNOR U4171 ( .A(n2409), .B(n2410), .Z(n1800) );
  ANDN U4172 ( .B(n1333), .A(n1331), .Z(n2408) );
  IV U4173 ( .A(n2073), .Z(n1331) );
  XOR U4174 ( .A(n2411), .B(n2412), .Z(n2073) );
  XOR U4175 ( .A(n2413), .B(n2414), .Z(n1333) );
  XOR U4176 ( .A(n2415), .B(n1805), .Z(out[675]) );
  XNOR U4177 ( .A(n2416), .B(n2417), .Z(n1805) );
  ANDN U4178 ( .B(n1335), .A(n1337), .Z(n2415) );
  XOR U4179 ( .A(n2418), .B(n2419), .Z(n1337) );
  XNOR U4180 ( .A(n2420), .B(n2421), .Z(n1335) );
  XNOR U4181 ( .A(n2422), .B(n1809), .Z(out[674]) );
  IV U4182 ( .A(n2083), .Z(n1809) );
  XOR U4183 ( .A(n2423), .B(n2424), .Z(n2083) );
  ANDN U4184 ( .B(n1341), .A(n1339), .Z(n2422) );
  XNOR U4185 ( .A(n2425), .B(n2426), .Z(n1339) );
  XNOR U4186 ( .A(n2427), .B(n2428), .Z(n1341) );
  XOR U4187 ( .A(n2429), .B(n1813), .Z(out[673]) );
  XNOR U4188 ( .A(n2430), .B(n2431), .Z(n1813) );
  ANDN U4189 ( .B(n1349), .A(n1347), .Z(n2429) );
  XNOR U4190 ( .A(n2432), .B(n2433), .Z(n1347) );
  XNOR U4191 ( .A(n2434), .B(n2435), .Z(n1349) );
  XOR U4192 ( .A(n2436), .B(n1817), .Z(out[672]) );
  XOR U4193 ( .A(n2437), .B(n2438), .Z(n1817) );
  ANDN U4194 ( .B(n1353), .A(n1351), .Z(n2436) );
  XOR U4195 ( .A(n2439), .B(n2440), .Z(n1351) );
  XOR U4196 ( .A(n2441), .B(n2442), .Z(n1353) );
  XOR U4197 ( .A(n2443), .B(n1830), .Z(out[671]) );
  XOR U4198 ( .A(n2444), .B(n2445), .Z(n1830) );
  AND U4199 ( .A(n1356), .B(n1355), .Z(n2443) );
  XOR U4200 ( .A(n2446), .B(n2447), .Z(n1355) );
  XOR U4201 ( .A(n2448), .B(n2449), .Z(n1356) );
  XOR U4202 ( .A(n2450), .B(n1834), .Z(out[670]) );
  XOR U4203 ( .A(n2451), .B(n2452), .Z(n1834) );
  AND U4204 ( .A(n1360), .B(n1359), .Z(n2450) );
  XOR U4205 ( .A(n2453), .B(n2454), .Z(n1359) );
  XOR U4206 ( .A(n2455), .B(n2456), .Z(n1360) );
  XOR U4207 ( .A(n2457), .B(n2458), .Z(out[66]) );
  NOR U4208 ( .A(n2459), .B(n2460), .Z(n2457) );
  XOR U4209 ( .A(n2461), .B(n1839), .Z(out[669]) );
  XNOR U4210 ( .A(n2462), .B(n2463), .Z(n1839) );
  AND U4211 ( .A(n1365), .B(n1363), .Z(n2461) );
  XNOR U4212 ( .A(n2464), .B(n2465), .Z(n1363) );
  XOR U4213 ( .A(n2466), .B(n2467), .Z(n1365) );
  XOR U4214 ( .A(n2468), .B(n1843), .Z(out[668]) );
  XNOR U4215 ( .A(n2469), .B(n2470), .Z(n1843) );
  ANDN U4216 ( .B(n1369), .A(n1367), .Z(n2468) );
  IV U4217 ( .A(n2102), .Z(n1367) );
  XOR U4218 ( .A(n2471), .B(n2472), .Z(n2102) );
  XNOR U4219 ( .A(n2473), .B(n2474), .Z(n1369) );
  XOR U4220 ( .A(n2475), .B(n1848), .Z(out[667]) );
  XNOR U4221 ( .A(n2476), .B(n2477), .Z(n1848) );
  ANDN U4222 ( .B(n1373), .A(n1371), .Z(n2475) );
  IV U4223 ( .A(n2106), .Z(n1371) );
  XOR U4224 ( .A(n2478), .B(n2479), .Z(n2106) );
  XNOR U4225 ( .A(n2480), .B(n2481), .Z(n1373) );
  XOR U4226 ( .A(n2482), .B(n1852), .Z(out[666]) );
  XNOR U4227 ( .A(n2483), .B(n2484), .Z(n1852) );
  AND U4228 ( .A(n1377), .B(n1375), .Z(n2482) );
  XNOR U4229 ( .A(n2485), .B(n2486), .Z(n1375) );
  XOR U4230 ( .A(n2487), .B(n2488), .Z(n1377) );
  XOR U4231 ( .A(n2489), .B(n1856), .Z(out[665]) );
  XOR U4232 ( .A(n2490), .B(n2491), .Z(n1856) );
  ANDN U4233 ( .B(n1379), .A(n1381), .Z(n2489) );
  XNOR U4234 ( .A(n2492), .B(n2493), .Z(n1381) );
  XOR U4235 ( .A(n2494), .B(n2495), .Z(n1379) );
  XOR U4236 ( .A(n2496), .B(n1860), .Z(out[664]) );
  XNOR U4237 ( .A(n2497), .B(n2498), .Z(n1860) );
  ANDN U4238 ( .B(n1385), .A(n1383), .Z(n2496) );
  IV U4239 ( .A(n2118), .Z(n1383) );
  XOR U4240 ( .A(n2499), .B(n2500), .Z(n2118) );
  XNOR U4241 ( .A(n2501), .B(n2502), .Z(n1385) );
  XNOR U4242 ( .A(n2503), .B(n1864), .Z(out[663]) );
  IV U4243 ( .A(n2122), .Z(n1864) );
  XNOR U4244 ( .A(n2504), .B(n2505), .Z(n2122) );
  ANDN U4245 ( .B(n1391), .A(n1393), .Z(n2503) );
  XNOR U4246 ( .A(n2506), .B(n2507), .Z(n1393) );
  XNOR U4247 ( .A(n2508), .B(n2509), .Z(n1391) );
  XNOR U4248 ( .A(n2510), .B(n1868), .Z(out[662]) );
  XNOR U4249 ( .A(n2511), .B(n2512), .Z(n1868) );
  NOR U4250 ( .A(n2126), .B(n1397), .Z(n2510) );
  XOR U4251 ( .A(n2513), .B(n2514), .Z(n1397) );
  XNOR U4252 ( .A(n2515), .B(n2516), .Z(n2126) );
  XOR U4253 ( .A(n2517), .B(n1876), .Z(out[661]) );
  XOR U4254 ( .A(n2518), .B(n2519), .Z(n1876) );
  ANDN U4255 ( .B(n1399), .A(n1401), .Z(n2517) );
  XNOR U4256 ( .A(n2520), .B(n2521), .Z(n1401) );
  XOR U4257 ( .A(n2522), .B(n2523), .Z(n1399) );
  XOR U4258 ( .A(n2524), .B(n1880), .Z(out[660]) );
  XOR U4259 ( .A(n2525), .B(n2526), .Z(n1880) );
  ANDN U4260 ( .B(n1403), .A(n1404), .Z(n2524) );
  XNOR U4261 ( .A(n2527), .B(n2528), .Z(n1404) );
  XNOR U4262 ( .A(n2529), .B(n2530), .Z(n1403) );
  XNOR U4263 ( .A(n2531), .B(n2532), .Z(out[65]) );
  NOR U4264 ( .A(n2533), .B(n2534), .Z(n2531) );
  XNOR U4265 ( .A(n2535), .B(n1884), .Z(out[659]) );
  IV U4266 ( .A(n2136), .Z(n1884) );
  XNOR U4267 ( .A(n2536), .B(n2537), .Z(n2136) );
  ANDN U4268 ( .B(n1409), .A(n1407), .Z(n2535) );
  XOR U4269 ( .A(n2538), .B(n2539), .Z(n1407) );
  XNOR U4270 ( .A(n2540), .B(n2541), .Z(n1409) );
  XOR U4271 ( .A(n2542), .B(n1888), .Z(out[658]) );
  XOR U4272 ( .A(n2543), .B(n2544), .Z(n1888) );
  ANDN U4273 ( .B(n1411), .A(n1412), .Z(n2542) );
  XNOR U4274 ( .A(n2545), .B(n2546), .Z(n1412) );
  XOR U4275 ( .A(n2547), .B(n2548), .Z(n1411) );
  XNOR U4276 ( .A(n2549), .B(n1893), .Z(out[657]) );
  IV U4277 ( .A(n2143), .Z(n1893) );
  XNOR U4278 ( .A(n2550), .B(n2551), .Z(n2143) );
  ANDN U4279 ( .B(n1417), .A(n1415), .Z(n2549) );
  XOR U4280 ( .A(n2552), .B(n2553), .Z(n1415) );
  XOR U4281 ( .A(n2554), .B(n2555), .Z(n1417) );
  XNOR U4282 ( .A(n2556), .B(n1897), .Z(out[656]) );
  IV U4283 ( .A(n2147), .Z(n1897) );
  XOR U4284 ( .A(n2557), .B(n2558), .Z(n2147) );
  ANDN U4285 ( .B(n1419), .A(n1421), .Z(n2556) );
  XNOR U4286 ( .A(n2559), .B(n2560), .Z(n1421) );
  XOR U4287 ( .A(n2561), .B(n2562), .Z(n1419) );
  XOR U4288 ( .A(n2563), .B(n1901), .Z(out[655]) );
  XOR U4289 ( .A(n2564), .B(n2565), .Z(n1901) );
  ANDN U4290 ( .B(n1423), .A(n1425), .Z(n2563) );
  XNOR U4291 ( .A(n2566), .B(n2567), .Z(n1425) );
  XNOR U4292 ( .A(n2568), .B(n2569), .Z(n1423) );
  XOR U4293 ( .A(n2570), .B(n1905), .Z(out[654]) );
  XOR U4294 ( .A(n2571), .B(n2572), .Z(n1905) );
  ANDN U4295 ( .B(n1427), .A(n1429), .Z(n2570) );
  XNOR U4296 ( .A(n2573), .B(n2574), .Z(n1429) );
  XNOR U4297 ( .A(n2575), .B(n2576), .Z(n1427) );
  XOR U4298 ( .A(n2577), .B(n1909), .Z(out[653]) );
  XOR U4299 ( .A(n2578), .B(n2579), .Z(n1909) );
  ANDN U4300 ( .B(n1435), .A(n1436), .Z(n2577) );
  XNOR U4301 ( .A(n2580), .B(n2581), .Z(n1436) );
  XNOR U4302 ( .A(n2582), .B(n2583), .Z(n1435) );
  XOR U4303 ( .A(n2584), .B(n1913), .Z(out[652]) );
  XOR U4304 ( .A(n2585), .B(n2586), .Z(n1913) );
  ANDN U4305 ( .B(n1439), .A(n1441), .Z(n2584) );
  XNOR U4306 ( .A(n2587), .B(n2588), .Z(n1441) );
  XOR U4307 ( .A(n2589), .B(n2590), .Z(n1439) );
  XOR U4308 ( .A(n2591), .B(n2166), .Z(out[651]) );
  XOR U4309 ( .A(n2592), .B(n2593), .Z(n2166) );
  ANDN U4310 ( .B(n1445), .A(n1443), .Z(n2591) );
  IV U4311 ( .A(n2165), .Z(n1443) );
  XNOR U4312 ( .A(n2594), .B(n2595), .Z(n2165) );
  XOR U4313 ( .A(n2596), .B(n2597), .Z(n1445) );
  XOR U4314 ( .A(n2598), .B(n1925), .Z(out[650]) );
  XOR U4315 ( .A(n2599), .B(n2600), .Z(n1925) );
  NOR U4316 ( .A(n1447), .B(n1448), .Z(n2598) );
  XNOR U4317 ( .A(n2601), .B(n2602), .Z(n1448) );
  XOR U4318 ( .A(n2603), .B(n2604), .Z(n1447) );
  XOR U4319 ( .A(n2605), .B(n2606), .Z(out[64]) );
  NOR U4320 ( .A(n2607), .B(n2608), .Z(n2605) );
  XOR U4321 ( .A(n2609), .B(n1930), .Z(out[649]) );
  XNOR U4322 ( .A(n2610), .B(n2611), .Z(n1930) );
  ANDN U4323 ( .B(n1451), .A(n1453), .Z(n2609) );
  XNOR U4324 ( .A(n2612), .B(n2613), .Z(n1453) );
  XOR U4325 ( .A(n2614), .B(n2615), .Z(n1451) );
  XOR U4326 ( .A(n2616), .B(n1934), .Z(out[648]) );
  XOR U4327 ( .A(n2617), .B(n2618), .Z(n1934) );
  NOR U4328 ( .A(n1457), .B(n1455), .Z(n2616) );
  XOR U4329 ( .A(n2619), .B(n2620), .Z(n1455) );
  XNOR U4330 ( .A(n2621), .B(n2622), .Z(n1457) );
  XOR U4331 ( .A(n2623), .B(n1939), .Z(out[647]) );
  XOR U4332 ( .A(n2624), .B(n2625), .Z(n1939) );
  ANDN U4333 ( .B(n1459), .A(n1461), .Z(n2623) );
  XOR U4334 ( .A(n2626), .B(n2627), .Z(n1461) );
  XNOR U4335 ( .A(n2628), .B(n2629), .Z(n1459) );
  XOR U4336 ( .A(n2630), .B(n1943), .Z(out[646]) );
  XNOR U4337 ( .A(n2631), .B(n2632), .Z(n1943) );
  ANDN U4338 ( .B(n1463), .A(n1464), .Z(n2630) );
  XNOR U4339 ( .A(n2633), .B(n2634), .Z(n1464) );
  XOR U4340 ( .A(n2635), .B(n2636), .Z(n1463) );
  XOR U4341 ( .A(n2637), .B(n1948), .Z(out[645]) );
  XOR U4342 ( .A(n2638), .B(n2639), .Z(n1948) );
  ANDN U4343 ( .B(n1467), .A(n1469), .Z(n2637) );
  XOR U4344 ( .A(n2640), .B(n2641), .Z(n1469) );
  XOR U4345 ( .A(n2642), .B(n2643), .Z(n1467) );
  XNOR U4346 ( .A(n2644), .B(n1953), .Z(out[644]) );
  XOR U4347 ( .A(n2645), .B(n2646), .Z(n1953) );
  ANDN U4348 ( .B(n1471), .A(n1472), .Z(n2644) );
  XOR U4349 ( .A(n2647), .B(n2648), .Z(n1472) );
  XOR U4350 ( .A(n2649), .B(n2650), .Z(n1471) );
  XOR U4351 ( .A(n2651), .B(n1957), .Z(out[643]) );
  XNOR U4352 ( .A(n2652), .B(n2653), .Z(n1957) );
  ANDN U4353 ( .B(n1483), .A(n1485), .Z(n2651) );
  XOR U4354 ( .A(n2654), .B(n2655), .Z(n1485) );
  XOR U4355 ( .A(n2656), .B(n2657), .Z(n1483) );
  XOR U4356 ( .A(n2658), .B(n1962), .Z(out[642]) );
  XOR U4357 ( .A(n2659), .B(n2660), .Z(n1962) );
  ANDN U4358 ( .B(n1487), .A(n1488), .Z(n2658) );
  XOR U4359 ( .A(n2661), .B(n2662), .Z(n1488) );
  XOR U4360 ( .A(n2663), .B(n2664), .Z(n1487) );
  XOR U4361 ( .A(n2665), .B(n1970), .Z(out[641]) );
  XOR U4362 ( .A(n2666), .B(n2667), .Z(n1970) );
  ANDN U4363 ( .B(n1491), .A(n1492), .Z(n2665) );
  XNOR U4364 ( .A(n2668), .B(n2669), .Z(n1492) );
  XNOR U4365 ( .A(n2670), .B(n2671), .Z(n1491) );
  XNOR U4366 ( .A(n2672), .B(n1974), .Z(out[640]) );
  IV U4367 ( .A(n2204), .Z(n1974) );
  XOR U4368 ( .A(n2673), .B(n2674), .Z(n2204) );
  ANDN U4369 ( .B(n1495), .A(n1496), .Z(n2672) );
  XOR U4370 ( .A(n2675), .B(n2676), .Z(n1496) );
  XOR U4371 ( .A(n2677), .B(n2678), .Z(n1495) );
  XNOR U4372 ( .A(n2679), .B(n2680), .Z(out[63]) );
  ANDN U4373 ( .B(n2681), .A(n2682), .Z(n2679) );
  XOR U4374 ( .A(n2683), .B(n2684), .Z(out[639]) );
  NOR U4375 ( .A(n2685), .B(n2686), .Z(n2683) );
  XOR U4376 ( .A(n2687), .B(n2688), .Z(out[638]) );
  ANDN U4377 ( .B(n2689), .A(n2690), .Z(n2687) );
  XNOR U4378 ( .A(n2691), .B(n2692), .Z(out[637]) );
  AND U4379 ( .A(n2693), .B(n2694), .Z(n2691) );
  XNOR U4380 ( .A(n2695), .B(n2696), .Z(out[636]) );
  NOR U4381 ( .A(n2697), .B(n2698), .Z(n2695) );
  XOR U4382 ( .A(n2699), .B(n2700), .Z(out[635]) );
  ANDN U4383 ( .B(n2701), .A(n2702), .Z(n2699) );
  XNOR U4384 ( .A(n2703), .B(n2704), .Z(out[634]) );
  NOR U4385 ( .A(n2705), .B(n2706), .Z(n2703) );
  XNOR U4386 ( .A(n2707), .B(n2708), .Z(out[633]) );
  NOR U4387 ( .A(n2709), .B(n2710), .Z(n2707) );
  XOR U4388 ( .A(n2711), .B(n2712), .Z(out[632]) );
  XOR U4389 ( .A(n2715), .B(n2716), .Z(out[631]) );
  ANDN U4390 ( .B(n2717), .A(n2718), .Z(n2715) );
  XNOR U4391 ( .A(n2719), .B(n2720), .Z(out[630]) );
  NOR U4392 ( .A(n2721), .B(n2722), .Z(n2719) );
  XNOR U4393 ( .A(n2723), .B(n2724), .Z(out[62]) );
  AND U4394 ( .A(n2725), .B(n2726), .Z(n2723) );
  XNOR U4395 ( .A(n2727), .B(n2728), .Z(out[629]) );
  NOR U4396 ( .A(n2729), .B(n2730), .Z(n2727) );
  XNOR U4397 ( .A(n2731), .B(n2732), .Z(out[628]) );
  ANDN U4398 ( .B(n2733), .A(n2734), .Z(n2731) );
  XNOR U4399 ( .A(n2735), .B(n2736), .Z(out[627]) );
  ANDN U4400 ( .B(n2737), .A(n2738), .Z(n2735) );
  XNOR U4401 ( .A(n2739), .B(n2740), .Z(out[626]) );
  AND U4402 ( .A(n2741), .B(n2742), .Z(n2739) );
  XOR U4403 ( .A(n2743), .B(n2744), .Z(out[625]) );
  AND U4404 ( .A(n2745), .B(n2746), .Z(n2743) );
  XOR U4405 ( .A(n2747), .B(n2748), .Z(out[624]) );
  NOR U4406 ( .A(n2749), .B(n2750), .Z(n2747) );
  XNOR U4407 ( .A(n2751), .B(n2752), .Z(out[623]) );
  ANDN U4408 ( .B(n2753), .A(n2754), .Z(n2751) );
  XOR U4409 ( .A(n2755), .B(n2756), .Z(out[622]) );
  XOR U4410 ( .A(n2759), .B(n2760), .Z(out[621]) );
  NOR U4411 ( .A(n2761), .B(n2762), .Z(n2759) );
  XNOR U4412 ( .A(n2763), .B(n2764), .Z(out[620]) );
  ANDN U4413 ( .B(n2765), .A(n2766), .Z(n2763) );
  XOR U4414 ( .A(n2767), .B(n2768), .Z(out[61]) );
  AND U4415 ( .A(n2769), .B(n2770), .Z(n2767) );
  XNOR U4416 ( .A(n2771), .B(n2772), .Z(out[619]) );
  ANDN U4417 ( .B(n2773), .A(n2774), .Z(n2771) );
  XNOR U4418 ( .A(n2775), .B(n2776), .Z(out[618]) );
  NOR U4419 ( .A(n2777), .B(n2778), .Z(n2775) );
  XNOR U4420 ( .A(n2779), .B(n2780), .Z(out[617]) );
  AND U4421 ( .A(n2781), .B(n2782), .Z(n2779) );
  XNOR U4422 ( .A(n2783), .B(n2784), .Z(out[616]) );
  AND U4423 ( .A(n2785), .B(n2786), .Z(n2783) );
  XOR U4424 ( .A(n2787), .B(n2788), .Z(out[615]) );
  XNOR U4425 ( .A(n2791), .B(n2792), .Z(out[614]) );
  NOR U4426 ( .A(n2793), .B(n2794), .Z(n2791) );
  XNOR U4427 ( .A(n2795), .B(n2796), .Z(out[613]) );
  ANDN U4428 ( .B(n2797), .A(n2798), .Z(n2795) );
  XNOR U4429 ( .A(n2799), .B(n2800), .Z(out[612]) );
  NOR U4430 ( .A(n2801), .B(n2802), .Z(n2799) );
  XNOR U4431 ( .A(n2803), .B(n2804), .Z(out[611]) );
  ANDN U4432 ( .B(n2805), .A(n2806), .Z(n2803) );
  XNOR U4433 ( .A(n2807), .B(n2808), .Z(out[610]) );
  AND U4434 ( .A(n2809), .B(n2810), .Z(n2807) );
  XOR U4435 ( .A(n2811), .B(n2812), .Z(out[60]) );
  XOR U4436 ( .A(n2815), .B(n2816), .Z(out[609]) );
  NOR U4437 ( .A(n2817), .B(n2818), .Z(n2815) );
  XNOR U4438 ( .A(n2819), .B(n2820), .Z(out[608]) );
  NOR U4439 ( .A(n2821), .B(n2822), .Z(n2819) );
  XNOR U4440 ( .A(n2823), .B(n2824), .Z(out[607]) );
  AND U4441 ( .A(n2825), .B(n2826), .Z(n2823) );
  XNOR U4442 ( .A(n2827), .B(n2828), .Z(out[606]) );
  ANDN U4443 ( .B(n2829), .A(n2830), .Z(n2827) );
  XNOR U4444 ( .A(n2831), .B(n2832), .Z(out[605]) );
  AND U4445 ( .A(n2833), .B(n2834), .Z(n2831) );
  XOR U4446 ( .A(n2835), .B(n2836), .Z(out[604]) );
  NOR U4447 ( .A(n2837), .B(n2838), .Z(n2835) );
  XOR U4448 ( .A(n2839), .B(n2840), .Z(out[603]) );
  NOR U4449 ( .A(n2841), .B(n2842), .Z(n2839) );
  XNOR U4450 ( .A(n2843), .B(n2844), .Z(out[602]) );
  NOR U4451 ( .A(n2845), .B(n2846), .Z(n2843) );
  XNOR U4452 ( .A(n2847), .B(n2848), .Z(out[601]) );
  ANDN U4453 ( .B(n2849), .A(n2850), .Z(n2847) );
  NOR U4454 ( .A(n2853), .B(n2854), .Z(n2851) );
  XOR U4455 ( .A(n2855), .B(n2238), .Z(out[5]) );
  ANDN U4456 ( .B(n2856), .A(n2857), .Z(n2855) );
  XOR U4457 ( .A(n2858), .B(n2859), .Z(out[59]) );
  AND U4458 ( .A(n2860), .B(n2861), .Z(n2858) );
  XOR U4459 ( .A(n2862), .B(n2863), .Z(out[599]) );
  NOR U4460 ( .A(n2864), .B(n2865), .Z(n2862) );
  XOR U4461 ( .A(n2866), .B(n2867), .Z(out[598]) );
  NOR U4462 ( .A(n2868), .B(n2869), .Z(n2866) );
  XNOR U4463 ( .A(n2870), .B(n2871), .Z(out[597]) );
  NOR U4464 ( .A(n2872), .B(n2873), .Z(n2870) );
  XOR U4465 ( .A(n2874), .B(n2875), .Z(out[596]) );
  NOR U4466 ( .A(n2876), .B(n2877), .Z(n2874) );
  XNOR U4467 ( .A(n2878), .B(n2879), .Z(out[595]) );
  AND U4468 ( .A(n2880), .B(n2881), .Z(n2878) );
  XNOR U4469 ( .A(n2882), .B(n2883), .Z(out[594]) );
  AND U4470 ( .A(n2884), .B(n2885), .Z(n2882) );
  XNOR U4471 ( .A(n2886), .B(n2887), .Z(out[593]) );
  ANDN U4472 ( .B(n2888), .A(n2889), .Z(n2886) );
  XNOR U4473 ( .A(n2890), .B(n2891), .Z(out[592]) );
  AND U4474 ( .A(n2892), .B(n2893), .Z(n2890) );
  XOR U4475 ( .A(n2894), .B(n2895), .Z(out[591]) );
  NOR U4476 ( .A(n2896), .B(n2897), .Z(n2894) );
  XNOR U4477 ( .A(n2898), .B(n2899), .Z(out[590]) );
  ANDN U4478 ( .B(n2900), .A(n2901), .Z(n2898) );
  XOR U4479 ( .A(n2902), .B(n2903), .Z(out[58]) );
  XOR U4480 ( .A(n2906), .B(n2907), .Z(out[589]) );
  NOR U4481 ( .A(n2908), .B(n2909), .Z(n2906) );
  NOR U4482 ( .A(n2912), .B(n2913), .Z(n2910) );
  XNOR U4483 ( .A(n2914), .B(n2915), .Z(out[587]) );
  AND U4484 ( .A(n2916), .B(n2917), .Z(n2914) );
  XOR U4485 ( .A(n2918), .B(n2919), .Z(out[586]) );
  NOR U4486 ( .A(n2920), .B(n2921), .Z(n2918) );
  XNOR U4487 ( .A(n2922), .B(n2923), .Z(out[585]) );
  AND U4488 ( .A(n2924), .B(n2925), .Z(n2922) );
  XNOR U4489 ( .A(n2926), .B(n2927), .Z(out[584]) );
  ANDN U4490 ( .B(n2928), .A(n2929), .Z(n2926) );
  XNOR U4491 ( .A(n2930), .B(n2931), .Z(out[583]) );
  ANDN U4492 ( .B(n2932), .A(n2933), .Z(n2930) );
  XNOR U4493 ( .A(n2934), .B(n2935), .Z(out[582]) );
  ANDN U4494 ( .B(n2936), .A(n2937), .Z(n2934) );
  XNOR U4495 ( .A(n2938), .B(n2939), .Z(out[581]) );
  AND U4496 ( .A(n2940), .B(n2941), .Z(n2938) );
  XOR U4497 ( .A(n2942), .B(n2943), .Z(out[580]) );
  ANDN U4498 ( .B(n2944), .A(n2945), .Z(n2942) );
  XNOR U4499 ( .A(n2946), .B(n2947), .Z(out[57]) );
  ANDN U4500 ( .B(n2948), .A(n2949), .Z(n2946) );
  XOR U4501 ( .A(n2950), .B(n2951), .Z(out[579]) );
  ANDN U4502 ( .B(n2952), .A(n2953), .Z(n2950) );
  XOR U4503 ( .A(n2954), .B(n2955), .Z(out[578]) );
  ANDN U4504 ( .B(n2956), .A(n2957), .Z(n2954) );
  XNOR U4505 ( .A(n2958), .B(n2959), .Z(out[577]) );
  ANDN U4506 ( .B(n2960), .A(n2961), .Z(n2958) );
  XOR U4507 ( .A(n2962), .B(n2963), .Z(out[576]) );
  AND U4508 ( .A(n2964), .B(n2965), .Z(n2962) );
  XOR U4509 ( .A(n2966), .B(n2686), .Z(out[575]) );
  ANDN U4510 ( .B(n2685), .A(n2967), .Z(n2966) );
  XNOR U4511 ( .A(n2968), .B(n2689), .Z(out[574]) );
  ANDN U4512 ( .B(n2690), .A(n2969), .Z(n2968) );
  XNOR U4513 ( .A(n2970), .B(n2694), .Z(out[573]) );
  NOR U4514 ( .A(n2971), .B(n2693), .Z(n2970) );
  XOR U4515 ( .A(n2972), .B(n2698), .Z(out[572]) );
  ANDN U4516 ( .B(n2697), .A(n2973), .Z(n2972) );
  IV U4517 ( .A(n2974), .Z(n2697) );
  XNOR U4518 ( .A(n2975), .B(n2701), .Z(out[571]) );
  ANDN U4519 ( .B(n2702), .A(n2976), .Z(n2975) );
  XOR U4520 ( .A(n2977), .B(n2706), .Z(out[570]) );
  ANDN U4521 ( .B(n2705), .A(n2978), .Z(n2977) );
  IV U4522 ( .A(n2979), .Z(n2705) );
  XNOR U4523 ( .A(n2980), .B(n2981), .Z(out[56]) );
  ANDN U4524 ( .B(n2982), .A(n2983), .Z(n2980) );
  XOR U4525 ( .A(n2984), .B(n2710), .Z(out[569]) );
  AND U4526 ( .A(n2709), .B(n2985), .Z(n2984) );
  XOR U4527 ( .A(n2986), .B(n2713), .Z(out[568]) );
  ANDN U4528 ( .B(n2987), .A(n2714), .Z(n2986) );
  XNOR U4529 ( .A(n2988), .B(n2717), .Z(out[567]) );
  ANDN U4530 ( .B(n2989), .A(n2990), .Z(n2988) );
  XOR U4531 ( .A(n2991), .B(n2722), .Z(out[566]) );
  ANDN U4532 ( .B(n2992), .A(n2993), .Z(n2991) );
  XOR U4533 ( .A(n2994), .B(n2729), .Z(out[565]) );
  AND U4534 ( .A(n2730), .B(n2995), .Z(n2994) );
  XNOR U4535 ( .A(n2996), .B(n2733), .Z(out[564]) );
  ANDN U4536 ( .B(n2997), .A(n2998), .Z(n2996) );
  XNOR U4537 ( .A(n2999), .B(n2737), .Z(out[563]) );
  AND U4538 ( .A(n2738), .B(n3000), .Z(n2999) );
  XNOR U4539 ( .A(n3001), .B(n2742), .Z(out[562]) );
  ANDN U4540 ( .B(n3002), .A(n2741), .Z(n3001) );
  XNOR U4541 ( .A(n3003), .B(n2746), .Z(out[561]) );
  ANDN U4542 ( .B(n3004), .A(n2745), .Z(n3003) );
  XOR U4543 ( .A(n3005), .B(n2750), .Z(out[560]) );
  ANDN U4544 ( .B(n3006), .A(n3007), .Z(n3005) );
  XNOR U4545 ( .A(n3008), .B(n3009), .Z(out[55]) );
  XNOR U4546 ( .A(n3012), .B(n2753), .Z(out[559]) );
  XOR U4547 ( .A(n3014), .B(n2757), .Z(out[558]) );
  ANDN U4548 ( .B(n3015), .A(n2758), .Z(n3014) );
  XOR U4549 ( .A(n3016), .B(n2762), .Z(out[557]) );
  ANDN U4550 ( .B(n3017), .A(n3018), .Z(n3016) );
  XNOR U4551 ( .A(n3019), .B(n2765), .Z(out[556]) );
  XNOR U4552 ( .A(n3021), .B(n2773), .Z(out[555]) );
  AND U4553 ( .A(n2774), .B(n3022), .Z(n3021) );
  XOR U4554 ( .A(n3023), .B(n2778), .Z(out[554]) );
  AND U4555 ( .A(n2777), .B(n3024), .Z(n3023) );
  XNOR U4556 ( .A(n3025), .B(n2782), .Z(out[553]) );
  ANDN U4557 ( .B(n3026), .A(n2781), .Z(n3025) );
  XNOR U4558 ( .A(n3027), .B(n2786), .Z(out[552]) );
  ANDN U4559 ( .B(n3028), .A(n2785), .Z(n3027) );
  XOR U4560 ( .A(n3029), .B(n2789), .Z(out[551]) );
  ANDN U4561 ( .B(n3030), .A(n2790), .Z(n3029) );
  XOR U4562 ( .A(n3031), .B(n2794), .Z(out[550]) );
  XNOR U4563 ( .A(n3033), .B(n3034), .Z(out[54]) );
  ANDN U4564 ( .B(n3035), .A(n3036), .Z(n3033) );
  XNOR U4565 ( .A(n3037), .B(n2797), .Z(out[549]) );
  ANDN U4566 ( .B(n3038), .A(n3039), .Z(n3037) );
  XOR U4567 ( .A(n3040), .B(n2802), .Z(out[548]) );
  AND U4568 ( .A(n2801), .B(n3041), .Z(n3040) );
  XNOR U4569 ( .A(n3042), .B(n2805), .Z(out[547]) );
  ANDN U4570 ( .B(n3043), .A(n3044), .Z(n3042) );
  XNOR U4571 ( .A(n3045), .B(n2810), .Z(out[546]) );
  ANDN U4572 ( .B(n3046), .A(n2809), .Z(n3045) );
  XOR U4573 ( .A(n3047), .B(n2818), .Z(out[545]) );
  AND U4574 ( .A(n2817), .B(n3048), .Z(n3047) );
  XOR U4575 ( .A(n3049), .B(n2822), .Z(out[544]) );
  XNOR U4576 ( .A(n3051), .B(n2826), .Z(out[543]) );
  NOR U4577 ( .A(n3052), .B(n2825), .Z(n3051) );
  XNOR U4578 ( .A(n3053), .B(n2829), .Z(out[542]) );
  ANDN U4579 ( .B(n3054), .A(n3055), .Z(n3053) );
  XNOR U4580 ( .A(n3056), .B(n2834), .Z(out[541]) );
  ANDN U4581 ( .B(n3057), .A(n2833), .Z(n3056) );
  XOR U4582 ( .A(n3058), .B(n2838), .Z(out[540]) );
  ANDN U4583 ( .B(n2837), .A(n3059), .Z(n3058) );
  XOR U4584 ( .A(n3060), .B(n3061), .Z(out[53]) );
  ANDN U4585 ( .B(n3062), .A(n3063), .Z(n3060) );
  XOR U4586 ( .A(n3064), .B(n2842), .Z(out[539]) );
  ANDN U4587 ( .B(n3065), .A(n3066), .Z(n3064) );
  XOR U4588 ( .A(n3067), .B(n2846), .Z(out[538]) );
  ANDN U4589 ( .B(n3068), .A(n3069), .Z(n3067) );
  XNOR U4590 ( .A(n3070), .B(n2849), .Z(out[537]) );
  ANDN U4591 ( .B(n2850), .A(n3071), .Z(n3070) );
  XOR U4592 ( .A(n3072), .B(n2854), .Z(out[536]) );
  ANDN U4593 ( .B(n2853), .A(n3073), .Z(n3072) );
  XOR U4594 ( .A(n3074), .B(n2865), .Z(out[535]) );
  ANDN U4595 ( .B(n3075), .A(n3076), .Z(n3074) );
  XOR U4596 ( .A(n3077), .B(n2869), .Z(out[534]) );
  ANDN U4597 ( .B(n2868), .A(n3078), .Z(n3077) );
  IV U4598 ( .A(n3079), .Z(n2868) );
  XOR U4599 ( .A(n3080), .B(n2873), .Z(out[533]) );
  XOR U4600 ( .A(n3082), .B(n2877), .Z(out[532]) );
  ANDN U4601 ( .B(n3083), .A(n3084), .Z(n3082) );
  XNOR U4602 ( .A(n3085), .B(n2881), .Z(out[531]) );
  ANDN U4603 ( .B(n3086), .A(n2880), .Z(n3085) );
  XNOR U4604 ( .A(n3087), .B(n2885), .Z(out[530]) );
  ANDN U4605 ( .B(n3088), .A(n2884), .Z(n3087) );
  XNOR U4606 ( .A(n3089), .B(n3090), .Z(out[52]) );
  ANDN U4607 ( .B(n3091), .A(n3092), .Z(n3089) );
  XNOR U4608 ( .A(n3093), .B(n2888), .Z(out[529]) );
  ANDN U4609 ( .B(n2889), .A(n3094), .Z(n3093) );
  XNOR U4610 ( .A(n3095), .B(n2893), .Z(out[528]) );
  NOR U4611 ( .A(n3096), .B(n2892), .Z(n3095) );
  XOR U4612 ( .A(n3097), .B(n2897), .Z(out[527]) );
  XNOR U4613 ( .A(n3099), .B(n2900), .Z(out[526]) );
  ANDN U4614 ( .B(n2901), .A(n3100), .Z(n3099) );
  XOR U4615 ( .A(n3101), .B(n2909), .Z(out[525]) );
  ANDN U4616 ( .B(n2908), .A(n3102), .Z(n3101) );
  IV U4617 ( .A(n3103), .Z(n2908) );
  XOR U4618 ( .A(n3104), .B(n2913), .Z(out[524]) );
  ANDN U4619 ( .B(n3105), .A(n3106), .Z(n3104) );
  XNOR U4620 ( .A(n3107), .B(n2917), .Z(out[523]) );
  NOR U4621 ( .A(n3108), .B(n2916), .Z(n3107) );
  XOR U4622 ( .A(n3109), .B(n2921), .Z(out[522]) );
  ANDN U4623 ( .B(n2920), .A(n3110), .Z(n3109) );
  IV U4624 ( .A(n3111), .Z(n2920) );
  XNOR U4625 ( .A(n3112), .B(n2925), .Z(out[521]) );
  NOR U4626 ( .A(n3113), .B(n2924), .Z(n3112) );
  XNOR U4627 ( .A(n3114), .B(n2928), .Z(out[520]) );
  ANDN U4628 ( .B(n2929), .A(n3115), .Z(n3114) );
  XOR U4629 ( .A(n3116), .B(n3117), .Z(out[51]) );
  ANDN U4630 ( .B(n3118), .A(n3119), .Z(n3116) );
  XNOR U4631 ( .A(n3120), .B(n2932), .Z(out[519]) );
  ANDN U4632 ( .B(n2933), .A(n3121), .Z(n3120) );
  XNOR U4633 ( .A(n3122), .B(n2936), .Z(out[518]) );
  ANDN U4634 ( .B(n2937), .A(n3123), .Z(n3122) );
  XNOR U4635 ( .A(n3124), .B(n2941), .Z(out[517]) );
  ANDN U4636 ( .B(n3125), .A(n2940), .Z(n3124) );
  XOR U4637 ( .A(n3126), .B(n2945), .Z(out[516]) );
  NOR U4638 ( .A(n3127), .B(n2944), .Z(n3126) );
  XNOR U4639 ( .A(n3128), .B(n2952), .Z(out[515]) );
  ANDN U4640 ( .B(n2953), .A(n3129), .Z(n3128) );
  XNOR U4641 ( .A(n3130), .B(n2956), .Z(out[514]) );
  ANDN U4642 ( .B(n2957), .A(n3131), .Z(n3130) );
  XNOR U4643 ( .A(n3132), .B(n2960), .Z(out[513]) );
  ANDN U4644 ( .B(n2961), .A(n3133), .Z(n3132) );
  XNOR U4645 ( .A(n3134), .B(n2965), .Z(out[512]) );
  NOR U4646 ( .A(n3135), .B(n2964), .Z(n3134) );
  XNOR U4647 ( .A(n3136), .B(n2685), .Z(out[511]) );
  ANDN U4648 ( .B(n3138), .A(n3139), .Z(n3136) );
  XNOR U4649 ( .A(n3140), .B(n2690), .Z(out[510]) );
  XOR U4650 ( .A(n3141), .B(n3142), .Z(n2690) );
  ANDN U4651 ( .B(n3143), .A(n3144), .Z(n3140) );
  XNOR U4652 ( .A(n3145), .B(n3146), .Z(out[50]) );
  ANDN U4653 ( .B(n3147), .A(n3148), .Z(n3145) );
  XOR U4654 ( .A(n3149), .B(n2693), .Z(out[509]) );
  ANDN U4655 ( .B(n2971), .A(n3151), .Z(n3149) );
  XOR U4656 ( .A(n3152), .B(n2974), .Z(out[508]) );
  XOR U4657 ( .A(n3153), .B(n3154), .Z(n2974) );
  AND U4658 ( .A(n2973), .B(n3155), .Z(n3152) );
  XNOR U4659 ( .A(n3156), .B(n2702), .Z(out[507]) );
  XOR U4660 ( .A(n3157), .B(n3158), .Z(n2702) );
  ANDN U4661 ( .B(n3159), .A(n3160), .Z(n3156) );
  XOR U4662 ( .A(n3161), .B(n2979), .Z(out[506]) );
  XOR U4663 ( .A(n3162), .B(n3163), .Z(n2979) );
  AND U4664 ( .A(n2978), .B(n3164), .Z(n3161) );
  XNOR U4665 ( .A(n3165), .B(n2709), .Z(out[505]) );
  XOR U4666 ( .A(n3166), .B(n2324), .Z(n2709) );
  ANDN U4667 ( .B(n3167), .A(n2985), .Z(n3165) );
  XOR U4668 ( .A(n3168), .B(n2714), .Z(out[504]) );
  XOR U4669 ( .A(n3169), .B(n2331), .Z(n2714) );
  ANDN U4670 ( .B(n3170), .A(n2987), .Z(n3168) );
  XNOR U4671 ( .A(n3171), .B(n2718), .Z(out[503]) );
  IV U4672 ( .A(n2990), .Z(n2718) );
  XOR U4673 ( .A(n3172), .B(n3173), .Z(n2990) );
  NOR U4674 ( .A(n3174), .B(n2989), .Z(n3171) );
  XNOR U4675 ( .A(n3175), .B(n2721), .Z(out[502]) );
  IV U4676 ( .A(n2993), .Z(n2721) );
  XNOR U4677 ( .A(n3176), .B(n2345), .Z(n2993) );
  ANDN U4678 ( .B(n3177), .A(n2992), .Z(n3175) );
  XNOR U4679 ( .A(n3178), .B(n2730), .Z(out[501]) );
  XOR U4680 ( .A(n3179), .B(n2352), .Z(n2730) );
  ANDN U4681 ( .B(n3180), .A(n2995), .Z(n3178) );
  XNOR U4682 ( .A(n3181), .B(n2734), .Z(out[500]) );
  IV U4683 ( .A(n2998), .Z(n2734) );
  XNOR U4684 ( .A(n3182), .B(n2359), .Z(n2998) );
  NOR U4685 ( .A(n3183), .B(n2997), .Z(n3181) );
  XNOR U4686 ( .A(n3184), .B(n2312), .Z(out[4]) );
  NOR U4687 ( .A(n3185), .B(n2311), .Z(n3184) );
  XNOR U4688 ( .A(n3186), .B(n3187), .Z(out[49]) );
  ANDN U4689 ( .B(n3188), .A(n3189), .Z(n3186) );
  XNOR U4690 ( .A(n3190), .B(n2738), .Z(out[499]) );
  XOR U4691 ( .A(n3191), .B(n3192), .Z(n2738) );
  ANDN U4692 ( .B(n3193), .A(n3000), .Z(n3190) );
  XOR U4693 ( .A(n3194), .B(n2741), .Z(out[498]) );
  XNOR U4694 ( .A(n3195), .B(n3196), .Z(n2741) );
  ANDN U4695 ( .B(n3197), .A(n3002), .Z(n3194) );
  XOR U4696 ( .A(n3198), .B(n2745), .Z(out[497]) );
  XNOR U4697 ( .A(n3199), .B(n2380), .Z(n2745) );
  NOR U4698 ( .A(n3200), .B(n3004), .Z(n3198) );
  XNOR U4699 ( .A(n3201), .B(n2749), .Z(out[496]) );
  IV U4700 ( .A(n3007), .Z(n2749) );
  XOR U4701 ( .A(n3202), .B(n2391), .Z(n3007) );
  ANDN U4702 ( .B(n3203), .A(n3006), .Z(n3201) );
  XNOR U4703 ( .A(n3204), .B(n2754), .Z(out[495]) );
  XOR U4704 ( .A(n3205), .B(n3206), .Z(n2754) );
  ANDN U4705 ( .B(n3207), .A(n3013), .Z(n3204) );
  XOR U4706 ( .A(n3208), .B(n2758), .Z(out[494]) );
  XOR U4707 ( .A(n3209), .B(n3210), .Z(n2758) );
  NOR U4708 ( .A(n3211), .B(n3015), .Z(n3208) );
  XNOR U4709 ( .A(n3212), .B(n2761), .Z(out[493]) );
  IV U4710 ( .A(n3018), .Z(n2761) );
  XNOR U4711 ( .A(n3213), .B(n2412), .Z(n3018) );
  NOR U4712 ( .A(n3214), .B(n3017), .Z(n3212) );
  XNOR U4713 ( .A(n3215), .B(n2766), .Z(out[492]) );
  XOR U4714 ( .A(n3216), .B(n3217), .Z(n2766) );
  NOR U4715 ( .A(n3218), .B(n3020), .Z(n3215) );
  XNOR U4716 ( .A(n3219), .B(n2774), .Z(out[491]) );
  XOR U4717 ( .A(n2425), .B(n3220), .Z(n2774) );
  NOR U4718 ( .A(n3221), .B(n3022), .Z(n3219) );
  XNOR U4719 ( .A(n3222), .B(n2777), .Z(out[490]) );
  XOR U4720 ( .A(n2432), .B(n3223), .Z(n2777) );
  ANDN U4721 ( .B(n3224), .A(n3024), .Z(n3222) );
  XNOR U4722 ( .A(n3225), .B(n3226), .Z(out[48]) );
  AND U4723 ( .A(n3227), .B(n3228), .Z(n3225) );
  XOR U4724 ( .A(n3229), .B(n2781), .Z(out[489]) );
  XNOR U4725 ( .A(n3230), .B(n2440), .Z(n2781) );
  NOR U4726 ( .A(n3231), .B(n3026), .Z(n3229) );
  XOR U4727 ( .A(n3232), .B(n2785), .Z(out[488]) );
  XNOR U4728 ( .A(n3233), .B(n3234), .Z(n2785) );
  ANDN U4729 ( .B(n3235), .A(n3028), .Z(n3232) );
  XOR U4730 ( .A(n3236), .B(n2790), .Z(out[487]) );
  XOR U4731 ( .A(n3237), .B(n3238), .Z(n2790) );
  NOR U4732 ( .A(n3239), .B(n3030), .Z(n3236) );
  XNOR U4733 ( .A(n3240), .B(n2793), .Z(out[486]) );
  XOR U4734 ( .A(n3241), .B(n2465), .Z(n2793) );
  NOR U4735 ( .A(n3242), .B(n3032), .Z(n3240) );
  XNOR U4736 ( .A(n3243), .B(n2798), .Z(out[485]) );
  IV U4737 ( .A(n3039), .Z(n2798) );
  XNOR U4738 ( .A(n3244), .B(n2472), .Z(n3039) );
  NOR U4739 ( .A(n3245), .B(n3038), .Z(n3243) );
  XNOR U4740 ( .A(n3246), .B(n2801), .Z(out[484]) );
  XOR U4741 ( .A(n3247), .B(n2479), .Z(n2801) );
  ANDN U4742 ( .B(n3248), .A(n3041), .Z(n3246) );
  XNOR U4743 ( .A(n3249), .B(n2806), .Z(out[483]) );
  IV U4744 ( .A(n3044), .Z(n2806) );
  XOR U4745 ( .A(n3250), .B(n2486), .Z(n3044) );
  ANDN U4746 ( .B(n3251), .A(n3043), .Z(n3249) );
  XOR U4747 ( .A(n3252), .B(n2809), .Z(out[482]) );
  XOR U4748 ( .A(n3253), .B(n3254), .Z(n2809) );
  ANDN U4749 ( .B(n3255), .A(n3046), .Z(n3252) );
  XNOR U4750 ( .A(n3256), .B(n2817), .Z(out[481]) );
  XOR U4751 ( .A(n3257), .B(n2500), .Z(n2817) );
  NOR U4752 ( .A(n3258), .B(n3048), .Z(n3256) );
  XNOR U4753 ( .A(n3259), .B(n2821), .Z(out[480]) );
  XOR U4754 ( .A(n3260), .B(n3261), .Z(n2821) );
  ANDN U4755 ( .B(n3262), .A(n3050), .Z(n3259) );
  IV U4756 ( .A(n3263), .Z(n3050) );
  XNOR U4757 ( .A(n3264), .B(n3265), .Z(out[47]) );
  NOR U4758 ( .A(n3266), .B(n3267), .Z(n3264) );
  XOR U4759 ( .A(n3268), .B(n2825), .Z(out[479]) );
  XNOR U4760 ( .A(n3269), .B(n2516), .Z(n2825) );
  ANDN U4761 ( .B(n3270), .A(n3271), .Z(n3268) );
  XNOR U4762 ( .A(n3272), .B(n2830), .Z(out[478]) );
  IV U4763 ( .A(n3055), .Z(n2830) );
  XNOR U4764 ( .A(n3273), .B(n2523), .Z(n3055) );
  NOR U4765 ( .A(n3274), .B(n3054), .Z(n3272) );
  XOR U4766 ( .A(n3275), .B(n2833), .Z(out[477]) );
  XOR U4767 ( .A(n3276), .B(n3277), .Z(n2833) );
  NOR U4768 ( .A(n3278), .B(n3057), .Z(n3275) );
  XNOR U4769 ( .A(n3279), .B(n2837), .Z(out[476]) );
  XOR U4770 ( .A(n3280), .B(n3281), .Z(n2837) );
  ANDN U4771 ( .B(n3282), .A(n3283), .Z(n3279) );
  XNOR U4772 ( .A(n3284), .B(n2841), .Z(out[475]) );
  IV U4773 ( .A(n3066), .Z(n2841) );
  XNOR U4774 ( .A(n3285), .B(n2548), .Z(n3066) );
  ANDN U4775 ( .B(n3286), .A(n3065), .Z(n3284) );
  XNOR U4776 ( .A(n3287), .B(n2845), .Z(out[474]) );
  IV U4777 ( .A(n3069), .Z(n2845) );
  XOR U4778 ( .A(n3288), .B(n2553), .Z(n3069) );
  ANDN U4779 ( .B(n3289), .A(n3068), .Z(n3287) );
  IV U4780 ( .A(n3290), .Z(n3068) );
  XNOR U4781 ( .A(n3291), .B(n2850), .Z(out[473]) );
  XOR U4782 ( .A(n3292), .B(n2562), .Z(n2850) );
  ANDN U4783 ( .B(n3071), .A(n3293), .Z(n3291) );
  XNOR U4784 ( .A(n3294), .B(n2853), .Z(out[472]) );
  XOR U4785 ( .A(n3295), .B(n3296), .Z(n2853) );
  ANDN U4786 ( .B(n3073), .A(n3297), .Z(n3294) );
  IV U4787 ( .A(n3298), .Z(n3073) );
  XNOR U4788 ( .A(n3299), .B(n2864), .Z(out[471]) );
  IV U4789 ( .A(n3076), .Z(n2864) );
  XOR U4790 ( .A(n3300), .B(n2576), .Z(n3076) );
  ANDN U4791 ( .B(n3301), .A(n3075), .Z(n3299) );
  XOR U4792 ( .A(n3302), .B(n3079), .Z(out[470]) );
  XOR U4793 ( .A(n3303), .B(n2583), .Z(n3079) );
  ANDN U4794 ( .B(n3078), .A(n3304), .Z(n3302) );
  IV U4795 ( .A(n3305), .Z(n3078) );
  XNOR U4796 ( .A(n3306), .B(n3307), .Z(out[46]) );
  ANDN U4797 ( .B(n3308), .A(n3309), .Z(n3306) );
  XNOR U4798 ( .A(n3310), .B(n2872), .Z(out[469]) );
  XOR U4799 ( .A(n3311), .B(n3312), .Z(n2872) );
  ANDN U4800 ( .B(n3313), .A(n3081), .Z(n3310) );
  XNOR U4801 ( .A(n3314), .B(n2876), .Z(out[468]) );
  IV U4802 ( .A(n3084), .Z(n2876) );
  XOR U4803 ( .A(n3315), .B(n2595), .Z(n3084) );
  ANDN U4804 ( .B(n3316), .A(n3083), .Z(n3314) );
  XOR U4805 ( .A(n3317), .B(n2880), .Z(out[467]) );
  XOR U4806 ( .A(n3318), .B(n2604), .Z(n2880) );
  ANDN U4807 ( .B(n3319), .A(n3086), .Z(n3317) );
  XOR U4808 ( .A(n3320), .B(n2884), .Z(out[466]) );
  XOR U4809 ( .A(n3321), .B(n3322), .Z(n2884) );
  NOR U4810 ( .A(n3323), .B(n3088), .Z(n3320) );
  XNOR U4811 ( .A(n3324), .B(n2889), .Z(out[465]) );
  XOR U4812 ( .A(n2619), .B(n3325), .Z(n2889) );
  XOR U4813 ( .A(n3328), .B(n2892), .Z(out[464]) );
  XNOR U4814 ( .A(n3329), .B(n3330), .Z(n2892) );
  XNOR U4815 ( .A(n3332), .B(n2896), .Z(out[463]) );
  XOR U4816 ( .A(n3333), .B(n3334), .Z(n2896) );
  NOR U4817 ( .A(n3335), .B(n3098), .Z(n3332) );
  XNOR U4818 ( .A(n3336), .B(n2901), .Z(out[462]) );
  XOR U4819 ( .A(n3337), .B(n3338), .Z(n2901) );
  XOR U4820 ( .A(n3340), .B(n3103), .Z(out[461]) );
  XOR U4821 ( .A(n3341), .B(n2650), .Z(n3103) );
  ANDN U4822 ( .B(n3342), .A(n3343), .Z(n3340) );
  XNOR U4823 ( .A(n3344), .B(n2912), .Z(out[460]) );
  IV U4824 ( .A(n3106), .Z(n2912) );
  XOR U4825 ( .A(n3345), .B(n2657), .Z(n3106) );
  NOR U4826 ( .A(n3346), .B(n3105), .Z(n3344) );
  XNOR U4827 ( .A(n3347), .B(n3348), .Z(out[45]) );
  AND U4828 ( .A(n3349), .B(n3350), .Z(n3347) );
  XOR U4829 ( .A(n3351), .B(n2916), .Z(out[459]) );
  XNOR U4830 ( .A(n3352), .B(n2664), .Z(n2916) );
  AND U4831 ( .A(n3108), .B(n3353), .Z(n3351) );
  XOR U4832 ( .A(n3354), .B(n3111), .Z(out[458]) );
  XOR U4833 ( .A(n3355), .B(n3356), .Z(n3111) );
  ANDN U4834 ( .B(n3110), .A(n3357), .Z(n3354) );
  XOR U4835 ( .A(n3358), .B(n2924), .Z(out[457]) );
  XNOR U4836 ( .A(n3359), .B(n2678), .Z(n2924) );
  XNOR U4837 ( .A(n3362), .B(n2929), .Z(out[456]) );
  XOR U4838 ( .A(n3363), .B(n3364), .Z(n2929) );
  ANDN U4839 ( .B(n3115), .A(n3365), .Z(n3362) );
  IV U4840 ( .A(n3366), .Z(n3115) );
  XNOR U4841 ( .A(n3367), .B(n2933), .Z(out[455]) );
  XNOR U4842 ( .A(n2217), .B(n3368), .Z(n2933) );
  ANDN U4843 ( .B(n3121), .A(n3369), .Z(n3367) );
  XNOR U4844 ( .A(n3370), .B(n2937), .Z(out[454]) );
  XOR U4845 ( .A(n3371), .B(n3372), .Z(n2937) );
  ANDN U4846 ( .B(n3373), .A(n3374), .Z(n3370) );
  XOR U4847 ( .A(n3375), .B(n2940), .Z(out[453]) );
  XNOR U4848 ( .A(n2231), .B(n3376), .Z(n2940) );
  ANDN U4849 ( .B(n3377), .A(n3125), .Z(n3375) );
  XOR U4850 ( .A(n3378), .B(n2944), .Z(out[452]) );
  XOR U4851 ( .A(n2244), .B(n3379), .Z(n2944) );
  ANDN U4852 ( .B(n3380), .A(n3381), .Z(n3378) );
  XNOR U4853 ( .A(n3382), .B(n2953), .Z(out[451]) );
  XOR U4854 ( .A(n3383), .B(n3384), .Z(n2953) );
  ANDN U4855 ( .B(n3385), .A(n3386), .Z(n3382) );
  XNOR U4856 ( .A(n3387), .B(n2957), .Z(out[450]) );
  XOR U4857 ( .A(n3388), .B(n2259), .Z(n2957) );
  ANDN U4858 ( .B(n3389), .A(n3390), .Z(n3387) );
  XNOR U4859 ( .A(n3391), .B(n3392), .Z(out[44]) );
  ANDN U4860 ( .B(n3393), .A(n3394), .Z(n3391) );
  XNOR U4861 ( .A(n3395), .B(n2961), .Z(out[449]) );
  XOR U4862 ( .A(n3396), .B(n3397), .Z(n2961) );
  ANDN U4863 ( .B(n3133), .A(n3398), .Z(n3395) );
  XOR U4864 ( .A(n3399), .B(n2964), .Z(out[448]) );
  XNOR U4865 ( .A(n3400), .B(n3401), .Z(n2964) );
  AND U4866 ( .A(n3135), .B(n3402), .Z(n3399) );
  XNOR U4867 ( .A(n3403), .B(n2967), .Z(out[447]) );
  IV U4868 ( .A(n3139), .Z(n2967) );
  XOR U4869 ( .A(n3404), .B(n2278), .Z(n3139) );
  ANDN U4870 ( .B(n2684), .A(n3138), .Z(n3403) );
  IV U4871 ( .A(n3405), .Z(n3138) );
  XNOR U4872 ( .A(n3406), .B(n2969), .Z(out[446]) );
  IV U4873 ( .A(n3144), .Z(n2969) );
  XOR U4874 ( .A(n3407), .B(n2285), .Z(n3144) );
  ANDN U4875 ( .B(n2688), .A(n3143), .Z(n3406) );
  XNOR U4876 ( .A(n3408), .B(n2971), .Z(out[445]) );
  XOR U4877 ( .A(n3409), .B(n2292), .Z(n2971) );
  XNOR U4878 ( .A(n3410), .B(n2973), .Z(out[444]) );
  XOR U4879 ( .A(n3411), .B(n2299), .Z(n2973) );
  NOR U4880 ( .A(n2696), .B(n3155), .Z(n3410) );
  IV U4881 ( .A(n3412), .Z(n2696) );
  XNOR U4882 ( .A(n3413), .B(n2976), .Z(out[443]) );
  IV U4883 ( .A(n3160), .Z(n2976) );
  XOR U4884 ( .A(n3414), .B(n2306), .Z(n3160) );
  ANDN U4885 ( .B(n2700), .A(n3159), .Z(n3413) );
  IV U4886 ( .A(n3415), .Z(n3159) );
  XNOR U4887 ( .A(n3416), .B(n2978), .Z(out[442]) );
  XOR U4888 ( .A(n3417), .B(n2317), .Z(n2978) );
  NOR U4889 ( .A(n2704), .B(n3164), .Z(n3416) );
  IV U4890 ( .A(n3418), .Z(n2704) );
  XOR U4891 ( .A(n3419), .B(n2985), .Z(out[441]) );
  XOR U4892 ( .A(n3420), .B(n3421), .Z(n2985) );
  NOR U4893 ( .A(n2708), .B(n3167), .Z(n3419) );
  IV U4894 ( .A(n3422), .Z(n2708) );
  XOR U4895 ( .A(n3423), .B(n2987), .Z(out[440]) );
  XOR U4896 ( .A(n2332), .B(n3424), .Z(n2987) );
  ANDN U4897 ( .B(n2712), .A(n3170), .Z(n3423) );
  XNOR U4898 ( .A(n3425), .B(n3426), .Z(out[43]) );
  XOR U4899 ( .A(n3429), .B(n2989), .Z(out[439]) );
  XOR U4900 ( .A(n2339), .B(n3430), .Z(n2989) );
  AND U4901 ( .A(n3174), .B(n2716), .Z(n3429) );
  XOR U4902 ( .A(n3431), .B(n2992), .Z(out[438]) );
  XOR U4903 ( .A(n2346), .B(n3432), .Z(n2992) );
  NOR U4904 ( .A(n2720), .B(n3177), .Z(n3431) );
  IV U4905 ( .A(n3433), .Z(n2720) );
  XOR U4906 ( .A(n3434), .B(n2995), .Z(out[437]) );
  XNOR U4907 ( .A(n3435), .B(n3436), .Z(n2995) );
  NOR U4908 ( .A(n2728), .B(n3180), .Z(n3434) );
  XOR U4909 ( .A(n3437), .B(n2997), .Z(out[436]) );
  XOR U4910 ( .A(n3438), .B(n3439), .Z(n2997) );
  XOR U4911 ( .A(n3440), .B(n3000), .Z(out[435]) );
  XNOR U4912 ( .A(n3441), .B(n3442), .Z(n3000) );
  NOR U4913 ( .A(n2736), .B(n3193), .Z(n3440) );
  XOR U4914 ( .A(n3443), .B(n3002), .Z(out[434]) );
  XNOR U4915 ( .A(n3444), .B(n3445), .Z(n3002) );
  NOR U4916 ( .A(n2740), .B(n3197), .Z(n3443) );
  XOR U4917 ( .A(n3446), .B(n3004), .Z(out[433]) );
  XOR U4918 ( .A(n3447), .B(n3448), .Z(n3004) );
  ANDN U4919 ( .B(n2744), .A(n3449), .Z(n3446) );
  XOR U4920 ( .A(n3450), .B(n3006), .Z(out[432]) );
  XOR U4921 ( .A(n3451), .B(n3452), .Z(n3006) );
  ANDN U4922 ( .B(n2748), .A(n3203), .Z(n3450) );
  XOR U4923 ( .A(n3453), .B(n3013), .Z(out[431]) );
  XOR U4924 ( .A(n3454), .B(n2398), .Z(n3013) );
  NOR U4925 ( .A(n2752), .B(n3207), .Z(n3453) );
  XOR U4926 ( .A(n3455), .B(n3015), .Z(out[430]) );
  XNOR U4927 ( .A(n3456), .B(n2405), .Z(n3015) );
  XNOR U4928 ( .A(n3457), .B(n3458), .Z(out[42]) );
  XOR U4929 ( .A(n3461), .B(n3017), .Z(out[429]) );
  XNOR U4930 ( .A(n3462), .B(n3463), .Z(n3017) );
  ANDN U4931 ( .B(n3214), .A(n3464), .Z(n3461) );
  XOR U4932 ( .A(n3465), .B(n3020), .Z(out[428]) );
  XNOR U4933 ( .A(n2418), .B(n3466), .Z(n3020) );
  ANDN U4934 ( .B(n3218), .A(n2764), .Z(n3465) );
  IV U4935 ( .A(n3467), .Z(n2764) );
  XOR U4936 ( .A(n3468), .B(n3022), .Z(out[427]) );
  XOR U4937 ( .A(n3469), .B(n3470), .Z(n3022) );
  ANDN U4938 ( .B(n3221), .A(n2772), .Z(n3468) );
  XOR U4939 ( .A(n3471), .B(n3024), .Z(out[426]) );
  XNOR U4940 ( .A(n2434), .B(n3472), .Z(n3024) );
  NOR U4941 ( .A(n2776), .B(n3224), .Z(n3471) );
  XOR U4942 ( .A(n3473), .B(n3026), .Z(out[425]) );
  XOR U4943 ( .A(n2441), .B(n3474), .Z(n3026) );
  NOR U4944 ( .A(n3475), .B(n2780), .Z(n3473) );
  XOR U4945 ( .A(n3476), .B(n3028), .Z(out[424]) );
  XNOR U4946 ( .A(n3477), .B(n3478), .Z(n3028) );
  NOR U4947 ( .A(n3235), .B(n2784), .Z(n3476) );
  XOR U4948 ( .A(n3479), .B(n3030), .Z(out[423]) );
  XOR U4949 ( .A(n2455), .B(n3480), .Z(n3030) );
  XOR U4950 ( .A(n3481), .B(n3032), .Z(out[422]) );
  XOR U4951 ( .A(n2466), .B(n3482), .Z(n3032) );
  ANDN U4952 ( .B(n3242), .A(n2792), .Z(n3481) );
  IV U4953 ( .A(n3483), .Z(n2792) );
  XOR U4954 ( .A(n3484), .B(n3038), .Z(out[421]) );
  XOR U4955 ( .A(n3485), .B(n3486), .Z(n3038) );
  ANDN U4956 ( .B(n3245), .A(n2796), .Z(n3484) );
  IV U4957 ( .A(n3487), .Z(n2796) );
  XOR U4958 ( .A(n3488), .B(n3041), .Z(out[420]) );
  XOR U4959 ( .A(n3489), .B(n3490), .Z(n3041) );
  NOR U4960 ( .A(n2800), .B(n3248), .Z(n3488) );
  IV U4961 ( .A(n3491), .Z(n2800) );
  XOR U4962 ( .A(n3492), .B(n3493), .Z(out[41]) );
  ANDN U4963 ( .B(n3494), .A(n3495), .Z(n3492) );
  XOR U4964 ( .A(n3496), .B(n3043), .Z(out[419]) );
  XOR U4965 ( .A(n2487), .B(n3497), .Z(n3043) );
  NOR U4966 ( .A(n2804), .B(n3251), .Z(n3496) );
  XOR U4967 ( .A(n3498), .B(n3046), .Z(out[418]) );
  XOR U4968 ( .A(n2492), .B(n3499), .Z(n3046) );
  NOR U4969 ( .A(n3255), .B(n2808), .Z(n3498) );
  XOR U4970 ( .A(n3500), .B(n3048), .Z(out[417]) );
  XNOR U4971 ( .A(n3501), .B(n2502), .Z(n3048) );
  ANDN U4972 ( .B(n2816), .A(n3502), .Z(n3500) );
  XNOR U4973 ( .A(n3503), .B(n3263), .Z(out[416]) );
  XOR U4974 ( .A(n2506), .B(n3504), .Z(n3263) );
  NOR U4975 ( .A(n2820), .B(n3262), .Z(n3503) );
  IV U4976 ( .A(n3505), .Z(n2820) );
  XNOR U4977 ( .A(n3506), .B(n3052), .Z(out[415]) );
  IV U4978 ( .A(n3271), .Z(n3052) );
  XOR U4979 ( .A(n2513), .B(n3507), .Z(n3271) );
  NOR U4980 ( .A(n2824), .B(n3270), .Z(n3506) );
  XOR U4981 ( .A(n3508), .B(n3054), .Z(out[414]) );
  XNOR U4982 ( .A(n2520), .B(n3509), .Z(n3054) );
  NOR U4983 ( .A(n3510), .B(n2828), .Z(n3508) );
  XOR U4984 ( .A(n3511), .B(n3057), .Z(out[413]) );
  XNOR U4985 ( .A(n2527), .B(n3512), .Z(n3057) );
  XNOR U4986 ( .A(n3513), .B(n3059), .Z(out[412]) );
  IV U4987 ( .A(n3283), .Z(n3059) );
  XOR U4988 ( .A(n3514), .B(n3515), .Z(n3283) );
  XOR U4989 ( .A(n3516), .B(n3065), .Z(out[411]) );
  XOR U4990 ( .A(n3517), .B(n3518), .Z(n3065) );
  NOR U4991 ( .A(n3519), .B(n3286), .Z(n3516) );
  XNOR U4992 ( .A(n3520), .B(n3290), .Z(out[410]) );
  XOR U4993 ( .A(n3521), .B(n3522), .Z(n3290) );
  NOR U4994 ( .A(n2844), .B(n3289), .Z(n3520) );
  XNOR U4995 ( .A(n3523), .B(n3524), .Z(out[40]) );
  ANDN U4996 ( .B(n3525), .A(n3526), .Z(n3523) );
  XNOR U4997 ( .A(n3527), .B(n3071), .Z(out[409]) );
  XNOR U4998 ( .A(n3528), .B(n2560), .Z(n3071) );
  NOR U4999 ( .A(n3529), .B(n2848), .Z(n3527) );
  XOR U5000 ( .A(n3530), .B(n3298), .Z(out[408]) );
  XOR U5001 ( .A(n3531), .B(n2567), .Z(n3298) );
  ANDN U5002 ( .B(n2852), .A(n3532), .Z(n3530) );
  XOR U5003 ( .A(n3533), .B(n3075), .Z(out[407]) );
  XOR U5004 ( .A(n3534), .B(n2574), .Z(n3075) );
  XOR U5005 ( .A(n3535), .B(n3305), .Z(out[406]) );
  XOR U5006 ( .A(n3536), .B(n2581), .Z(n3305) );
  ANDN U5007 ( .B(n3304), .A(n3537), .Z(n3535) );
  XOR U5008 ( .A(n3538), .B(n3081), .Z(out[405]) );
  XOR U5009 ( .A(n3539), .B(n2588), .Z(n3081) );
  NOR U5010 ( .A(n2871), .B(n3313), .Z(n3538) );
  IV U5011 ( .A(n3540), .Z(n2871) );
  XOR U5012 ( .A(n3541), .B(n3083), .Z(out[404]) );
  XNOR U5013 ( .A(n3542), .B(n3543), .Z(n3083) );
  XOR U5014 ( .A(n3544), .B(n3086), .Z(out[403]) );
  XNOR U5015 ( .A(n3545), .B(n3546), .Z(n3086) );
  NOR U5016 ( .A(n3319), .B(n2879), .Z(n3544) );
  XOR U5017 ( .A(n3547), .B(n3088), .Z(out[402]) );
  XOR U5018 ( .A(n3548), .B(n2613), .Z(n3088) );
  NOR U5019 ( .A(n3549), .B(n2883), .Z(n3547) );
  XNOR U5020 ( .A(n3550), .B(n3094), .Z(out[401]) );
  IV U5021 ( .A(n3326), .Z(n3094) );
  XNOR U5022 ( .A(n3551), .B(n2622), .Z(n3326) );
  ANDN U5023 ( .B(n3327), .A(n2887), .Z(n3550) );
  IV U5024 ( .A(n3552), .Z(n2887) );
  XNOR U5025 ( .A(n3553), .B(n3096), .Z(out[400]) );
  XOR U5026 ( .A(n3554), .B(n2627), .Z(n3096) );
  NOR U5027 ( .A(n3331), .B(n2891), .Z(n3553) );
  XOR U5028 ( .A(n3555), .B(n2386), .Z(out[3]) );
  NOR U5029 ( .A(n3556), .B(n2385), .Z(n3555) );
  XNOR U5030 ( .A(n3557), .B(n3558), .Z(out[39]) );
  ANDN U5031 ( .B(n3559), .A(n3560), .Z(n3557) );
  XOR U5032 ( .A(n3561), .B(n3098), .Z(out[399]) );
  XOR U5033 ( .A(n3562), .B(n2634), .Z(n3098) );
  ANDN U5034 ( .B(n3335), .A(n3563), .Z(n3561) );
  XNOR U5035 ( .A(n3564), .B(n3100), .Z(out[398]) );
  XOR U5036 ( .A(n3565), .B(n2641), .Z(n3100) );
  NOR U5037 ( .A(n3339), .B(n2899), .Z(n3564) );
  XNOR U5038 ( .A(n3566), .B(n3102), .Z(out[397]) );
  IV U5039 ( .A(n3343), .Z(n3102) );
  XNOR U5040 ( .A(n3567), .B(n2648), .Z(n3343) );
  ANDN U5041 ( .B(n2907), .A(n3342), .Z(n3566) );
  XOR U5042 ( .A(n3568), .B(n3105), .Z(out[396]) );
  XNOR U5043 ( .A(n3569), .B(n2655), .Z(n3105) );
  XNOR U5044 ( .A(n3570), .B(n3108), .Z(out[395]) );
  XNOR U5045 ( .A(n3571), .B(n2662), .Z(n3108) );
  NOR U5046 ( .A(n3353), .B(n2915), .Z(n3570) );
  XNOR U5047 ( .A(n3572), .B(n3110), .Z(out[394]) );
  XOR U5048 ( .A(n3573), .B(n2669), .Z(n3110) );
  ANDN U5049 ( .B(n3357), .A(n3574), .Z(n3572) );
  XNOR U5050 ( .A(n3575), .B(n3113), .Z(out[393]) );
  IV U5051 ( .A(n3360), .Z(n3113) );
  XNOR U5052 ( .A(n3576), .B(n2676), .Z(n3360) );
  ANDN U5053 ( .B(n3361), .A(n2923), .Z(n3575) );
  IV U5054 ( .A(n3577), .Z(n2923) );
  XOR U5055 ( .A(n3578), .B(n3366), .Z(out[392]) );
  XOR U5056 ( .A(n3579), .B(n2209), .Z(n3366) );
  XNOR U5057 ( .A(n3580), .B(n3121), .Z(out[391]) );
  XOR U5058 ( .A(n3581), .B(n2216), .Z(n3121) );
  XNOR U5059 ( .A(n3582), .B(n3123), .Z(out[390]) );
  IV U5060 ( .A(n3374), .Z(n3123) );
  XOR U5061 ( .A(n3583), .B(n2225), .Z(n3374) );
  NOR U5062 ( .A(n2935), .B(n3373), .Z(n3582) );
  XNOR U5063 ( .A(n3584), .B(n3585), .Z(out[38]) );
  XOR U5064 ( .A(n3588), .B(n3125), .Z(out[389]) );
  XNOR U5065 ( .A(n3589), .B(n2230), .Z(n3125) );
  NOR U5066 ( .A(n2939), .B(n3377), .Z(n3588) );
  XNOR U5067 ( .A(n3590), .B(n3127), .Z(out[388]) );
  IV U5068 ( .A(n3381), .Z(n3127) );
  XOR U5069 ( .A(n3591), .B(n2243), .Z(n3381) );
  ANDN U5070 ( .B(n2943), .A(n3380), .Z(n3590) );
  IV U5071 ( .A(n3592), .Z(n3380) );
  XNOR U5072 ( .A(n3593), .B(n3129), .Z(out[387]) );
  IV U5073 ( .A(n3386), .Z(n3129) );
  XNOR U5074 ( .A(n3594), .B(n2250), .Z(n3386) );
  ANDN U5075 ( .B(n2951), .A(n3385), .Z(n3593) );
  XNOR U5076 ( .A(n3595), .B(n3131), .Z(out[386]) );
  IV U5077 ( .A(n3390), .Z(n3131) );
  XNOR U5078 ( .A(n3596), .B(n2257), .Z(n3390) );
  ANDN U5079 ( .B(n2955), .A(n3389), .Z(n3595) );
  XNOR U5080 ( .A(n3597), .B(n3133), .Z(out[385]) );
  XOR U5081 ( .A(n3598), .B(n2266), .Z(n3133) );
  NOR U5082 ( .A(n3599), .B(n2959), .Z(n3597) );
  XNOR U5083 ( .A(n3600), .B(n3135), .Z(out[384]) );
  XOR U5084 ( .A(n3601), .B(n2271), .Z(n3135) );
  ANDN U5085 ( .B(n2963), .A(n3402), .Z(n3600) );
  XNOR U5086 ( .A(n3602), .B(n3405), .Z(out[383]) );
  XOR U5087 ( .A(n1815), .B(n3603), .Z(n3405) );
  ANDN U5088 ( .B(n2686), .A(n2684), .Z(n3602) );
  XOR U5089 ( .A(n3604), .B(n2045), .Z(n2684) );
  XNOR U5090 ( .A(n3605), .B(n3606), .Z(n2686) );
  XOR U5091 ( .A(n3607), .B(n3143), .Z(out[382]) );
  XNOR U5092 ( .A(n1828), .B(n3608), .Z(n3143) );
  NOR U5093 ( .A(n2689), .B(n2688), .Z(n3607) );
  XOR U5094 ( .A(n3609), .B(n2049), .Z(n2688) );
  XNOR U5095 ( .A(n3610), .B(n2350), .Z(n2689) );
  XNOR U5096 ( .A(n3611), .B(n3151), .Z(out[381]) );
  XOR U5097 ( .A(n1832), .B(n3612), .Z(n3151) );
  ANDN U5098 ( .B(n2692), .A(n2694), .Z(n3611) );
  XOR U5099 ( .A(n3613), .B(n3614), .Z(n2694) );
  XNOR U5100 ( .A(n3615), .B(n2053), .Z(n2692) );
  XOR U5101 ( .A(n3616), .B(n3155), .Z(out[380]) );
  XNOR U5102 ( .A(n1837), .B(n3617), .Z(n3155) );
  ANDN U5103 ( .B(n2698), .A(n3412), .Z(n3616) );
  XOR U5104 ( .A(n3618), .B(n2056), .Z(n3412) );
  XOR U5105 ( .A(n3619), .B(n3620), .Z(n2698) );
  XNOR U5106 ( .A(n3621), .B(n3622), .Z(out[37]) );
  ANDN U5107 ( .B(n3623), .A(n3624), .Z(n3621) );
  XNOR U5108 ( .A(n3625), .B(n3415), .Z(out[379]) );
  XOR U5109 ( .A(n3626), .B(n3627), .Z(n3415) );
  NOR U5110 ( .A(n2701), .B(n2700), .Z(n3625) );
  XNOR U5111 ( .A(n3628), .B(n2059), .Z(n2700) );
  XOR U5112 ( .A(n3629), .B(n2371), .Z(n2701) );
  XOR U5113 ( .A(n3630), .B(n3164), .Z(out[378]) );
  XNOR U5114 ( .A(n1846), .B(n3631), .Z(n3164) );
  ANDN U5115 ( .B(n2706), .A(n3418), .Z(n3630) );
  XOR U5116 ( .A(n3632), .B(n2063), .Z(n3418) );
  XNOR U5117 ( .A(n3633), .B(n3634), .Z(n2706) );
  XOR U5118 ( .A(n3635), .B(n3167), .Z(out[377]) );
  XNOR U5119 ( .A(n1850), .B(n3636), .Z(n3167) );
  ANDN U5120 ( .B(n2710), .A(n3422), .Z(n3635) );
  XOR U5121 ( .A(n3637), .B(n2066), .Z(n3422) );
  XOR U5122 ( .A(n3638), .B(n3639), .Z(n2710) );
  XOR U5123 ( .A(n3640), .B(n3170), .Z(out[376]) );
  XNOR U5124 ( .A(n3641), .B(n3642), .Z(n3170) );
  ANDN U5125 ( .B(n2713), .A(n2712), .Z(n3640) );
  XOR U5126 ( .A(n3643), .B(n2069), .Z(n2712) );
  XOR U5127 ( .A(n3644), .B(n2396), .Z(n2713) );
  XNOR U5128 ( .A(n3645), .B(n3174), .Z(out[375]) );
  XOR U5129 ( .A(n1858), .B(n3646), .Z(n3174) );
  NOR U5130 ( .A(n2717), .B(n2716), .Z(n3645) );
  XOR U5131 ( .A(n3647), .B(n2072), .Z(n2716) );
  XOR U5132 ( .A(n3648), .B(n2403), .Z(n2717) );
  XOR U5133 ( .A(n3649), .B(n3177), .Z(out[374]) );
  XOR U5134 ( .A(n1862), .B(n3650), .Z(n3177) );
  ANDN U5135 ( .B(n2722), .A(n3433), .Z(n3649) );
  XNOR U5136 ( .A(n3651), .B(n2079), .Z(n3433) );
  XOR U5137 ( .A(n3653), .B(n3180), .Z(out[373]) );
  XNOR U5138 ( .A(n1866), .B(n3654), .Z(n3180) );
  AND U5139 ( .A(n2729), .B(n2728), .Z(n3653) );
  XOR U5140 ( .A(n3655), .B(n2082), .Z(n2728) );
  XOR U5141 ( .A(n3656), .B(n3657), .Z(n2729) );
  XNOR U5142 ( .A(n3658), .B(n3183), .Z(out[372]) );
  XOR U5143 ( .A(n1874), .B(n3659), .Z(n3183) );
  ANDN U5144 ( .B(n2732), .A(n2733), .Z(n3658) );
  XOR U5145 ( .A(n3660), .B(n2424), .Z(n2733) );
  XNOR U5146 ( .A(n3661), .B(n2086), .Z(n2732) );
  XOR U5147 ( .A(n3662), .B(n3193), .Z(out[371]) );
  XNOR U5148 ( .A(n1878), .B(n3663), .Z(n3193) );
  ANDN U5149 ( .B(n2736), .A(n2737), .Z(n3662) );
  XOR U5150 ( .A(n3664), .B(n2431), .Z(n2737) );
  XNOR U5151 ( .A(n3665), .B(n2089), .Z(n2736) );
  XOR U5152 ( .A(n3666), .B(n3197), .Z(out[370]) );
  XNOR U5153 ( .A(n1882), .B(n3667), .Z(n3197) );
  ANDN U5154 ( .B(n2740), .A(n2742), .Z(n3666) );
  XOR U5155 ( .A(n3669), .B(n2092), .Z(n2740) );
  XNOR U5156 ( .A(n3670), .B(n3671), .Z(out[36]) );
  XNOR U5157 ( .A(n3674), .B(n3200), .Z(out[369]) );
  IV U5158 ( .A(n3449), .Z(n3200) );
  XOR U5159 ( .A(n3675), .B(n3676), .Z(n3449) );
  NOR U5160 ( .A(n2746), .B(n2744), .Z(n3674) );
  XNOR U5161 ( .A(n3677), .B(n2095), .Z(n2744) );
  XOR U5162 ( .A(n3679), .B(n3203), .Z(out[368]) );
  XOR U5163 ( .A(n1891), .B(n3680), .Z(n3203) );
  ANDN U5164 ( .B(n2750), .A(n2748), .Z(n3679) );
  XNOR U5165 ( .A(n3681), .B(n2098), .Z(n2748) );
  XNOR U5166 ( .A(n3682), .B(n3683), .Z(n2750) );
  XOR U5167 ( .A(n3684), .B(n3207), .Z(out[367]) );
  XOR U5168 ( .A(n1895), .B(n3685), .Z(n3207) );
  ANDN U5169 ( .B(n2752), .A(n2753), .Z(n3684) );
  XOR U5170 ( .A(n3686), .B(n2463), .Z(n2753) );
  XOR U5171 ( .A(n3687), .B(n2101), .Z(n2752) );
  XNOR U5172 ( .A(n3688), .B(n3211), .Z(out[366]) );
  XOR U5173 ( .A(n1899), .B(n3689), .Z(n3211) );
  ANDN U5174 ( .B(n2757), .A(n2756), .Z(n3688) );
  XOR U5175 ( .A(n3690), .B(n3691), .Z(n2756) );
  XOR U5176 ( .A(n3692), .B(n3693), .Z(n2757) );
  XNOR U5177 ( .A(n3694), .B(n3214), .Z(out[365]) );
  XOR U5178 ( .A(n3695), .B(n3696), .Z(n3214) );
  ANDN U5179 ( .B(n2762), .A(n2760), .Z(n3694) );
  IV U5180 ( .A(n3464), .Z(n2760) );
  XOR U5181 ( .A(n2108), .B(n3697), .Z(n3464) );
  XOR U5182 ( .A(n3698), .B(n2477), .Z(n2762) );
  XNOR U5183 ( .A(n3699), .B(n3218), .Z(out[364]) );
  XOR U5184 ( .A(n1907), .B(n3700), .Z(n3218) );
  NOR U5185 ( .A(n3467), .B(n2765), .Z(n3699) );
  XOR U5186 ( .A(n3701), .B(n2484), .Z(n2765) );
  XOR U5187 ( .A(n3702), .B(n2114), .Z(n3467) );
  XNOR U5188 ( .A(n3703), .B(n3221), .Z(out[363]) );
  XOR U5189 ( .A(n1911), .B(n3704), .Z(n3221) );
  ANDN U5190 ( .B(n2772), .A(n2773), .Z(n3703) );
  XOR U5191 ( .A(n3705), .B(n2491), .Z(n2773) );
  XOR U5192 ( .A(n2116), .B(n3706), .Z(n2772) );
  XOR U5193 ( .A(n3707), .B(n3224), .Z(out[362]) );
  XOR U5194 ( .A(n3708), .B(n3709), .Z(n3224) );
  AND U5195 ( .A(n2776), .B(n2778), .Z(n3707) );
  XOR U5196 ( .A(n3710), .B(n3711), .Z(n2778) );
  XOR U5197 ( .A(n2120), .B(n3712), .Z(n2776) );
  XNOR U5198 ( .A(n3713), .B(n3231), .Z(out[361]) );
  IV U5199 ( .A(n3475), .Z(n3231) );
  XOR U5200 ( .A(n3714), .B(n3715), .Z(n3475) );
  ANDN U5201 ( .B(n2780), .A(n2782), .Z(n3713) );
  XOR U5202 ( .A(n3716), .B(n2505), .Z(n2782) );
  XOR U5203 ( .A(n2124), .B(n3717), .Z(n2780) );
  XOR U5204 ( .A(n3718), .B(n3235), .Z(out[360]) );
  XNOR U5205 ( .A(n3719), .B(n3720), .Z(n3235) );
  ANDN U5206 ( .B(n2784), .A(n2786), .Z(n3718) );
  XNOR U5207 ( .A(n3721), .B(n2512), .Z(n2786) );
  XOR U5208 ( .A(n2128), .B(n3722), .Z(n2784) );
  XNOR U5209 ( .A(n3723), .B(n1036), .Z(out[35]) );
  XNOR U5210 ( .A(n3725), .B(n3239), .Z(out[359]) );
  XOR U5211 ( .A(n3726), .B(n3727), .Z(n3239) );
  ANDN U5212 ( .B(n2789), .A(n2788), .Z(n3725) );
  XOR U5213 ( .A(n3728), .B(n3729), .Z(n2788) );
  XOR U5214 ( .A(n3730), .B(n3731), .Z(n2789) );
  XNOR U5215 ( .A(n3732), .B(n3242), .Z(out[358]) );
  XOR U5216 ( .A(n3733), .B(n3734), .Z(n3242) );
  ANDN U5217 ( .B(n2794), .A(n3483), .Z(n3732) );
  XOR U5218 ( .A(n2134), .B(n3735), .Z(n3483) );
  XOR U5219 ( .A(n3736), .B(n2526), .Z(n2794) );
  XNOR U5220 ( .A(n3737), .B(n3245), .Z(out[357]) );
  XNOR U5221 ( .A(n1941), .B(n3738), .Z(n3245) );
  NOR U5222 ( .A(n3487), .B(n2797), .Z(n3737) );
  XOR U5223 ( .A(n3739), .B(n2537), .Z(n2797) );
  XOR U5224 ( .A(n3740), .B(n2139), .Z(n3487) );
  XOR U5225 ( .A(n3741), .B(n3248), .Z(out[356]) );
  XNOR U5226 ( .A(n1946), .B(n3742), .Z(n3248) );
  ANDN U5227 ( .B(n2802), .A(n3491), .Z(n3741) );
  XNOR U5228 ( .A(n3743), .B(n2142), .Z(n3491) );
  XNOR U5229 ( .A(n3744), .B(n2544), .Z(n2802) );
  XOR U5230 ( .A(n3745), .B(n3251), .Z(out[355]) );
  XNOR U5231 ( .A(n1951), .B(n3746), .Z(n3251) );
  ANDN U5232 ( .B(n2804), .A(n2805), .Z(n3745) );
  XOR U5233 ( .A(n3747), .B(n2551), .Z(n2805) );
  XNOR U5234 ( .A(n3748), .B(n2146), .Z(n2804) );
  XOR U5235 ( .A(n3749), .B(n3255), .Z(out[354]) );
  XNOR U5236 ( .A(n1955), .B(n3750), .Z(n3255) );
  ANDN U5237 ( .B(n2808), .A(n2810), .Z(n3749) );
  XNOR U5238 ( .A(n3751), .B(n2558), .Z(n2810) );
  XOR U5239 ( .A(n3752), .B(n2152), .Z(n2808) );
  XNOR U5240 ( .A(n3753), .B(n3258), .Z(out[353]) );
  IV U5241 ( .A(n3502), .Z(n3258) );
  XOR U5242 ( .A(n3754), .B(n1961), .Z(n3502) );
  ANDN U5243 ( .B(n2818), .A(n2816), .Z(n3753) );
  XOR U5244 ( .A(n3755), .B(n2155), .Z(n2816) );
  XNOR U5245 ( .A(n3756), .B(n3757), .Z(n2818) );
  XOR U5246 ( .A(n3758), .B(n3262), .Z(out[352]) );
  XNOR U5247 ( .A(n3759), .B(n1969), .Z(n3262) );
  ANDN U5248 ( .B(n2822), .A(n3505), .Z(n3758) );
  XOR U5249 ( .A(n3760), .B(n2158), .Z(n3505) );
  XOR U5250 ( .A(n3761), .B(n3762), .Z(n2822) );
  XOR U5251 ( .A(n3763), .B(n3270), .Z(out[351]) );
  XNOR U5252 ( .A(n3764), .B(n1973), .Z(n3270) );
  ANDN U5253 ( .B(n2824), .A(n2826), .Z(n3763) );
  XNOR U5254 ( .A(n3765), .B(n2579), .Z(n2826) );
  XNOR U5255 ( .A(n3766), .B(n2161), .Z(n2824) );
  XNOR U5256 ( .A(n3767), .B(n3274), .Z(out[350]) );
  IV U5257 ( .A(n3510), .Z(n3274) );
  XOR U5258 ( .A(n3768), .B(n1662), .Z(n3510) );
  ANDN U5259 ( .B(n2828), .A(n2829), .Z(n3767) );
  XNOR U5260 ( .A(n2585), .B(n3769), .Z(n2829) );
  XNOR U5261 ( .A(n3770), .B(n2164), .Z(n2828) );
  XNOR U5262 ( .A(n3771), .B(n1081), .Z(out[34]) );
  ANDN U5263 ( .B(n3772), .A(n1080), .Z(n3771) );
  XNOR U5264 ( .A(n3773), .B(n3278), .Z(out[349]) );
  XOR U5265 ( .A(n3774), .B(n1667), .Z(n3278) );
  ANDN U5266 ( .B(n2832), .A(n2834), .Z(n3773) );
  XNOR U5267 ( .A(n2592), .B(n3775), .Z(n2834) );
  XNOR U5268 ( .A(n3776), .B(n2169), .Z(n2832) );
  XOR U5269 ( .A(n3777), .B(n3282), .Z(out[348]) );
  XOR U5270 ( .A(n3778), .B(n1675), .Z(n3282) );
  ANDN U5271 ( .B(n2838), .A(n2836), .Z(n3777) );
  XOR U5272 ( .A(n3779), .B(n3780), .Z(n2836) );
  XOR U5273 ( .A(n2599), .B(n3781), .Z(n2838) );
  XOR U5274 ( .A(n3782), .B(n3286), .Z(out[347]) );
  XOR U5275 ( .A(n3783), .B(n1680), .Z(n3286) );
  ANDN U5276 ( .B(n2842), .A(n2840), .Z(n3782) );
  IV U5277 ( .A(n3519), .Z(n2840) );
  XNOR U5278 ( .A(n3784), .B(n2175), .Z(n3519) );
  XNOR U5279 ( .A(n3785), .B(n2611), .Z(n2842) );
  XOR U5280 ( .A(n3786), .B(n3289), .Z(out[346]) );
  XNOR U5281 ( .A(n3787), .B(n1685), .Z(n3289) );
  AND U5282 ( .A(n2844), .B(n2846), .Z(n3786) );
  XNOR U5283 ( .A(n3788), .B(n3789), .Z(n2846) );
  XOR U5284 ( .A(n3790), .B(n3791), .Z(n2844) );
  XNOR U5285 ( .A(n3792), .B(n3293), .Z(out[345]) );
  IV U5286 ( .A(n3529), .Z(n3293) );
  XOR U5287 ( .A(n3793), .B(n1689), .Z(n3529) );
  ANDN U5288 ( .B(n2848), .A(n2849), .Z(n3792) );
  XNOR U5289 ( .A(n3794), .B(n3795), .Z(n2849) );
  XNOR U5290 ( .A(n3796), .B(n2181), .Z(n2848) );
  XNOR U5291 ( .A(n3797), .B(n3297), .Z(out[344]) );
  IV U5292 ( .A(n3532), .Z(n3297) );
  XNOR U5293 ( .A(n3798), .B(n1693), .Z(n3532) );
  ANDN U5294 ( .B(n2854), .A(n2852), .Z(n3797) );
  XOR U5295 ( .A(n3799), .B(n2188), .Z(n2852) );
  XOR U5296 ( .A(n3800), .B(n3801), .Z(n2854) );
  XOR U5297 ( .A(n3802), .B(n3301), .Z(out[343]) );
  XNOR U5298 ( .A(n3803), .B(n1698), .Z(n3301) );
  ANDN U5299 ( .B(n2865), .A(n2863), .Z(n3802) );
  XOR U5300 ( .A(n3804), .B(n3805), .Z(n2863) );
  XOR U5301 ( .A(n3806), .B(n2639), .Z(n2865) );
  XNOR U5302 ( .A(n3807), .B(n3304), .Z(out[342]) );
  XNOR U5303 ( .A(n3808), .B(n1703), .Z(n3304) );
  ANDN U5304 ( .B(n2869), .A(n2867), .Z(n3807) );
  IV U5305 ( .A(n3537), .Z(n2867) );
  XNOR U5306 ( .A(n3809), .B(n2194), .Z(n3537) );
  XOR U5307 ( .A(n3810), .B(n3811), .Z(n2869) );
  XOR U5308 ( .A(n3812), .B(n3313), .Z(out[341]) );
  XNOR U5309 ( .A(n3813), .B(n1708), .Z(n3313) );
  ANDN U5310 ( .B(n2873), .A(n3540), .Z(n3812) );
  XOR U5311 ( .A(n3814), .B(n2197), .Z(n3540) );
  XNOR U5312 ( .A(n3815), .B(n2653), .Z(n2873) );
  XOR U5313 ( .A(n3816), .B(n3316), .Z(out[340]) );
  XOR U5314 ( .A(n3817), .B(n3818), .Z(n3316) );
  ANDN U5315 ( .B(n2877), .A(n2875), .Z(n3816) );
  XOR U5316 ( .A(n3819), .B(n3820), .Z(n2875) );
  XOR U5317 ( .A(n3821), .B(n3822), .Z(n2877) );
  XNOR U5318 ( .A(n3823), .B(n1125), .Z(out[33]) );
  ANDN U5319 ( .B(n3824), .A(n1124), .Z(n3823) );
  XOR U5320 ( .A(n3825), .B(n3319), .Z(out[339]) );
  XOR U5321 ( .A(n3826), .B(n1718), .Z(n3319) );
  ANDN U5322 ( .B(n2879), .A(n2881), .Z(n3825) );
  XOR U5323 ( .A(n3827), .B(n3828), .Z(n2881) );
  XOR U5324 ( .A(n3829), .B(n2203), .Z(n2879) );
  XNOR U5325 ( .A(n3830), .B(n3323), .Z(out[338]) );
  IV U5326 ( .A(n3549), .Z(n3323) );
  XOR U5327 ( .A(n3831), .B(n1727), .Z(n3549) );
  ANDN U5328 ( .B(n2883), .A(n2885), .Z(n3830) );
  XOR U5329 ( .A(n3832), .B(n2674), .Z(n2885) );
  XNOR U5330 ( .A(n3833), .B(n3834), .Z(n2883) );
  XNOR U5331 ( .A(n3835), .B(n3327), .Z(out[337]) );
  XOR U5332 ( .A(n3836), .B(n1732), .Z(n3327) );
  NOR U5333 ( .A(n3552), .B(n2888), .Z(n3835) );
  XNOR U5334 ( .A(n3837), .B(n2207), .Z(n2888) );
  XOR U5335 ( .A(n3838), .B(n1980), .Z(n3552) );
  XOR U5336 ( .A(n3839), .B(n3331), .Z(out[336]) );
  XOR U5337 ( .A(n3840), .B(n1736), .Z(n3331) );
  ANDN U5338 ( .B(n2891), .A(n2893), .Z(n3839) );
  XOR U5339 ( .A(n3841), .B(n2214), .Z(n2893) );
  XNOR U5340 ( .A(n3842), .B(n3843), .Z(n2891) );
  XNOR U5341 ( .A(n3844), .B(n3335), .Z(out[335]) );
  XOR U5342 ( .A(n3845), .B(n1741), .Z(n3335) );
  ANDN U5343 ( .B(n2897), .A(n2895), .Z(n3844) );
  IV U5344 ( .A(n3563), .Z(n2895) );
  XOR U5345 ( .A(n3846), .B(n1986), .Z(n3563) );
  XOR U5346 ( .A(n3847), .B(n2221), .Z(n2897) );
  XOR U5347 ( .A(n3848), .B(n3339), .Z(out[334]) );
  XOR U5348 ( .A(n3849), .B(n1745), .Z(n3339) );
  ANDN U5349 ( .B(n2899), .A(n2900), .Z(n3848) );
  XOR U5350 ( .A(n3850), .B(n2228), .Z(n2900) );
  XNOR U5351 ( .A(n3851), .B(n1989), .Z(n2899) );
  XOR U5352 ( .A(n3852), .B(n3342), .Z(out[333]) );
  XOR U5353 ( .A(n3853), .B(n1749), .Z(n3342) );
  ANDN U5354 ( .B(n2909), .A(n2907), .Z(n3852) );
  XNOR U5355 ( .A(n3854), .B(n1992), .Z(n2907) );
  XOR U5356 ( .A(n3855), .B(n2241), .Z(n2909) );
  XNOR U5357 ( .A(n3856), .B(n3346), .Z(out[332]) );
  XOR U5358 ( .A(n3857), .B(n1754), .Z(n3346) );
  ANDN U5359 ( .B(n2913), .A(n2911), .Z(n3856) );
  XOR U5360 ( .A(n3858), .B(n1995), .Z(n2911) );
  XOR U5361 ( .A(n3859), .B(n2248), .Z(n2913) );
  XOR U5362 ( .A(n3860), .B(n3353), .Z(out[331]) );
  XNOR U5363 ( .A(n3861), .B(n3862), .Z(n3353) );
  ANDN U5364 ( .B(n2915), .A(n2917), .Z(n3860) );
  XNOR U5365 ( .A(n3863), .B(n2255), .Z(n2917) );
  XOR U5366 ( .A(n3864), .B(n1998), .Z(n2915) );
  XNOR U5367 ( .A(n3865), .B(n3357), .Z(out[330]) );
  XOR U5368 ( .A(n3866), .B(n3867), .Z(n3357) );
  ANDN U5369 ( .B(n2921), .A(n2919), .Z(n3865) );
  IV U5370 ( .A(n3574), .Z(n2919) );
  XOR U5371 ( .A(n3868), .B(n2005), .Z(n3574) );
  XOR U5372 ( .A(n3869), .B(n3870), .Z(n2921) );
  XOR U5373 ( .A(n3871), .B(n1169), .Z(out[32]) );
  ANDN U5374 ( .B(n1168), .A(n3872), .Z(n3871) );
  IV U5375 ( .A(n3873), .Z(n1168) );
  XNOR U5376 ( .A(n3874), .B(n3361), .Z(out[329]) );
  XOR U5377 ( .A(n3875), .B(n1767), .Z(n3361) );
  NOR U5378 ( .A(n3577), .B(n2925), .Z(n3874) );
  XNOR U5379 ( .A(n3876), .B(n2269), .Z(n2925) );
  XOR U5380 ( .A(n3877), .B(n2009), .Z(n3577) );
  XNOR U5381 ( .A(n3878), .B(n3365), .Z(out[328]) );
  XOR U5382 ( .A(n3879), .B(n1775), .Z(n3365) );
  ANDN U5383 ( .B(n2927), .A(n2928), .Z(n3878) );
  XOR U5384 ( .A(n3880), .B(n2276), .Z(n2928) );
  IV U5385 ( .A(n3881), .Z(n2276) );
  XNOR U5386 ( .A(n3882), .B(n2012), .Z(n2927) );
  XNOR U5387 ( .A(n3883), .B(n3369), .Z(out[327]) );
  XOR U5388 ( .A(n3884), .B(n1780), .Z(n3369) );
  ANDN U5389 ( .B(n2931), .A(n2932), .Z(n3883) );
  XOR U5390 ( .A(n3885), .B(n2283), .Z(n2932) );
  XNOR U5391 ( .A(n3886), .B(n2015), .Z(n2931) );
  XOR U5392 ( .A(n3887), .B(n3373), .Z(out[326]) );
  XNOR U5393 ( .A(n3888), .B(n1785), .Z(n3373) );
  ANDN U5394 ( .B(n2935), .A(n2936), .Z(n3887) );
  XNOR U5395 ( .A(n3889), .B(n2290), .Z(n2936) );
  XOR U5396 ( .A(n3890), .B(n2019), .Z(n2935) );
  XOR U5397 ( .A(n3891), .B(n3377), .Z(out[325]) );
  XNOR U5398 ( .A(n3892), .B(n1790), .Z(n3377) );
  ANDN U5399 ( .B(n2939), .A(n2941), .Z(n3891) );
  XNOR U5400 ( .A(n3894), .B(n2022), .Z(n2939) );
  XNOR U5401 ( .A(n3895), .B(n3592), .Z(out[324]) );
  XOR U5402 ( .A(n3896), .B(n1794), .Z(n3592) );
  ANDN U5403 ( .B(n2945), .A(n2943), .Z(n3895) );
  XOR U5404 ( .A(n3897), .B(n2025), .Z(n2943) );
  XOR U5405 ( .A(n3898), .B(n3899), .Z(n2945) );
  XOR U5406 ( .A(n3900), .B(n3385), .Z(out[323]) );
  XOR U5407 ( .A(n1798), .B(n3901), .Z(n3385) );
  NOR U5408 ( .A(n2952), .B(n2951), .Z(n3900) );
  XOR U5409 ( .A(n3902), .B(n2028), .Z(n2951) );
  XNOR U5410 ( .A(n3903), .B(n2315), .Z(n2952) );
  XOR U5411 ( .A(n3904), .B(n3389), .Z(out[322]) );
  XOR U5412 ( .A(n3905), .B(n1804), .Z(n3389) );
  NOR U5413 ( .A(n2956), .B(n2955), .Z(n3904) );
  XNOR U5414 ( .A(n3906), .B(n2031), .Z(n2955) );
  XNOR U5415 ( .A(n3907), .B(n2322), .Z(n2956) );
  IV U5416 ( .A(n3908), .Z(n2322) );
  XNOR U5417 ( .A(n3909), .B(n3398), .Z(out[321]) );
  IV U5418 ( .A(n3599), .Z(n3398) );
  XOR U5419 ( .A(n1807), .B(n3910), .Z(n3599) );
  ANDN U5420 ( .B(n2959), .A(n2960), .Z(n3909) );
  XOR U5421 ( .A(n3911), .B(n2329), .Z(n2960) );
  XNOR U5422 ( .A(n3912), .B(n2034), .Z(n2959) );
  XOR U5423 ( .A(n3913), .B(n3402), .Z(out[320]) );
  XNOR U5424 ( .A(n1811), .B(n3914), .Z(n3402) );
  NOR U5425 ( .A(n2965), .B(n2963), .Z(n3913) );
  XOR U5426 ( .A(n3915), .B(n2041), .Z(n2963) );
  XNOR U5427 ( .A(n3916), .B(n2336), .Z(n2965) );
  XNOR U5428 ( .A(n3917), .B(n1213), .Z(out[31]) );
  XOR U5429 ( .A(n3919), .B(n2682), .Z(out[319]) );
  NOR U5430 ( .A(n3920), .B(n2681), .Z(n3919) );
  XNOR U5431 ( .A(n3921), .B(n2726), .Z(out[318]) );
  ANDN U5432 ( .B(n3922), .A(n2725), .Z(n3921) );
  XNOR U5433 ( .A(n3923), .B(n2770), .Z(out[317]) );
  ANDN U5434 ( .B(n3924), .A(n2769), .Z(n3923) );
  XNOR U5435 ( .A(n3925), .B(n2814), .Z(out[316]) );
  NOR U5436 ( .A(n3926), .B(n2813), .Z(n3925) );
  XNOR U5437 ( .A(n3927), .B(n2861), .Z(out[315]) );
  ANDN U5438 ( .B(n3928), .A(n2860), .Z(n3927) );
  XNOR U5439 ( .A(n3929), .B(n2905), .Z(out[314]) );
  ANDN U5440 ( .B(n3930), .A(n2904), .Z(n3929) );
  XNOR U5441 ( .A(n3931), .B(n2948), .Z(out[313]) );
  XNOR U5442 ( .A(n3933), .B(n2982), .Z(out[312]) );
  XNOR U5443 ( .A(n3935), .B(n3011), .Z(out[311]) );
  ANDN U5444 ( .B(n3936), .A(n3010), .Z(n3935) );
  XNOR U5445 ( .A(n3937), .B(n3035), .Z(out[310]) );
  XOR U5446 ( .A(n3939), .B(n1257), .Z(out[30]) );
  ANDN U5447 ( .B(n1256), .A(n3940), .Z(n3939) );
  XOR U5448 ( .A(n3941), .B(n3063), .Z(out[309]) );
  ANDN U5449 ( .B(n3942), .A(n3062), .Z(n3941) );
  XOR U5450 ( .A(n3943), .B(n3092), .Z(out[308]) );
  ANDN U5451 ( .B(n3944), .A(n3091), .Z(n3943) );
  XOR U5452 ( .A(n3945), .B(n3119), .Z(out[307]) );
  NOR U5453 ( .A(n3946), .B(n3118), .Z(n3945) );
  XNOR U5454 ( .A(n3947), .B(n3147), .Z(out[306]) );
  XOR U5455 ( .A(n3949), .B(n3189), .Z(out[305]) );
  NOR U5456 ( .A(n3950), .B(n3188), .Z(n3949) );
  XNOR U5457 ( .A(n3951), .B(n3228), .Z(out[304]) );
  ANDN U5458 ( .B(n3952), .A(n3227), .Z(n3951) );
  XOR U5459 ( .A(n3953), .B(n3267), .Z(out[303]) );
  ANDN U5460 ( .B(n3954), .A(n3955), .Z(n3953) );
  XNOR U5461 ( .A(n3956), .B(n3308), .Z(out[302]) );
  AND U5462 ( .A(n3309), .B(n3957), .Z(n3956) );
  XNOR U5463 ( .A(n3958), .B(n3350), .Z(out[301]) );
  ANDN U5464 ( .B(n3959), .A(n3349), .Z(n3958) );
  XNOR U5465 ( .A(n3960), .B(n3393), .Z(out[300]) );
  ANDN U5466 ( .B(n3961), .A(n3962), .Z(n3960) );
  XOR U5467 ( .A(n3963), .B(n2460), .Z(out[2]) );
  ANDN U5468 ( .B(n3964), .A(n3965), .Z(n3963) );
  XNOR U5469 ( .A(n3966), .B(n1301), .Z(out[29]) );
  NOR U5470 ( .A(n3967), .B(n1300), .Z(n3966) );
  XNOR U5471 ( .A(n3968), .B(n3428), .Z(out[299]) );
  NOR U5472 ( .A(n3969), .B(n3427), .Z(n3968) );
  XNOR U5473 ( .A(n3970), .B(n3460), .Z(out[298]) );
  ANDN U5474 ( .B(n3971), .A(n3459), .Z(n3970) );
  XOR U5475 ( .A(n3972), .B(n3495), .Z(out[297]) );
  ANDN U5476 ( .B(n3973), .A(n3494), .Z(n3972) );
  XOR U5477 ( .A(n3974), .B(n3526), .Z(out[296]) );
  NOR U5478 ( .A(n3975), .B(n3525), .Z(n3974) );
  XOR U5479 ( .A(n3976), .B(n3560), .Z(out[295]) );
  NOR U5480 ( .A(n3977), .B(n3559), .Z(n3976) );
  XNOR U5481 ( .A(n3978), .B(n3587), .Z(out[294]) );
  ANDN U5482 ( .B(n3979), .A(n3586), .Z(n3978) );
  XOR U5483 ( .A(n3980), .B(n3624), .Z(out[293]) );
  ANDN U5484 ( .B(n3981), .A(n3623), .Z(n3980) );
  XNOR U5485 ( .A(n3982), .B(n3673), .Z(out[292]) );
  NOR U5486 ( .A(n3983), .B(n3672), .Z(n3982) );
  XNOR U5487 ( .A(n3984), .B(n1037), .Z(out[291]) );
  XOR U5488 ( .A(n3438), .B(n3985), .Z(n1037) );
  IV U5489 ( .A(n2360), .Z(n3438) );
  ANDN U5490 ( .B(n3986), .A(n3724), .Z(n3984) );
  XOR U5491 ( .A(n3987), .B(n1080), .Z(out[290]) );
  XOR U5492 ( .A(n3441), .B(n3988), .Z(n1080) );
  ANDN U5493 ( .B(n3989), .A(n3772), .Z(n3987) );
  XNOR U5494 ( .A(n3990), .B(n1344), .Z(out[28]) );
  XOR U5495 ( .A(n3992), .B(n1124), .Z(out[289]) );
  XOR U5496 ( .A(n2374), .B(n3993), .Z(n1124) );
  IV U5497 ( .A(n3444), .Z(n2374) );
  NOR U5498 ( .A(n3994), .B(n3824), .Z(n3992) );
  XOR U5499 ( .A(n3995), .B(n3873), .Z(out[288]) );
  XOR U5500 ( .A(n3447), .B(n3996), .Z(n3873) );
  ANDN U5501 ( .B(n3872), .A(n3997), .Z(n3995) );
  XOR U5502 ( .A(n3998), .B(n1212), .Z(out[287]) );
  XOR U5503 ( .A(n3451), .B(n3999), .Z(n1212) );
  IV U5504 ( .A(n2392), .Z(n3451) );
  ANDN U5505 ( .B(n4000), .A(n3918), .Z(n3998) );
  XNOR U5506 ( .A(n4001), .B(n1256), .Z(out[286]) );
  XNOR U5507 ( .A(n4002), .B(n2398), .Z(n1256) );
  ANDN U5508 ( .B(n3940), .A(n4003), .Z(n4001) );
  IV U5509 ( .A(n4004), .Z(n3940) );
  XOR U5510 ( .A(n4005), .B(n1300), .Z(out[285]) );
  XNOR U5511 ( .A(n4006), .B(n2405), .Z(n1300) );
  XNOR U5512 ( .A(n4008), .B(n1345), .Z(out[284]) );
  XOR U5513 ( .A(n3462), .B(n4009), .Z(n1345) );
  IV U5514 ( .A(n2413), .Z(n3462) );
  NOR U5515 ( .A(n4010), .B(n3991), .Z(n4008) );
  XNOR U5516 ( .A(n4011), .B(n1389), .Z(out[283]) );
  XOR U5517 ( .A(n4014), .B(n1433), .Z(out[282]) );
  ANDN U5518 ( .B(n4015), .A(n4016), .Z(n4014) );
  XOR U5519 ( .A(n4017), .B(n1480), .Z(out[281]) );
  ANDN U5520 ( .B(n4018), .A(n4019), .Z(n4017) );
  XOR U5521 ( .A(n4020), .B(n1515), .Z(out[280]) );
  ANDN U5522 ( .B(n4021), .A(n4022), .Z(n4020) );
  XNOR U5523 ( .A(n4023), .B(n1388), .Z(out[27]) );
  ANDN U5524 ( .B(n1389), .A(n4012), .Z(n4023) );
  XOR U5525 ( .A(n2418), .B(n4024), .Z(n1389) );
  XOR U5526 ( .A(n4025), .B(n1540), .Z(out[279]) );
  AND U5527 ( .A(n4026), .B(n4027), .Z(n4025) );
  XOR U5528 ( .A(n4028), .B(n1569), .Z(out[278]) );
  AND U5529 ( .A(n4029), .B(n4030), .Z(n4028) );
  XOR U5530 ( .A(n4031), .B(n1593), .Z(out[277]) );
  ANDN U5531 ( .B(n4032), .A(n4033), .Z(n4031) );
  XOR U5532 ( .A(n4034), .B(n1616), .Z(out[276]) );
  ANDN U5533 ( .B(n4035), .A(n4036), .Z(n4034) );
  XOR U5534 ( .A(n4037), .B(n1640), .Z(out[275]) );
  ANDN U5535 ( .B(n4038), .A(n4039), .Z(n4037) );
  XOR U5536 ( .A(n4040), .B(n1671), .Z(out[274]) );
  ANDN U5537 ( .B(n4041), .A(n4042), .Z(n4040) );
  XNOR U5538 ( .A(n4043), .B(n1723), .Z(out[273]) );
  ANDN U5539 ( .B(n4044), .A(n4045), .Z(n4043) );
  XNOR U5540 ( .A(n4046), .B(n1771), .Z(out[272]) );
  IV U5541 ( .A(n4047), .Z(n1771) );
  ANDN U5542 ( .B(n4048), .A(n4049), .Z(n4046) );
  XNOR U5543 ( .A(n4050), .B(n1826), .Z(out[271]) );
  NOR U5544 ( .A(n4051), .B(n4052), .Z(n4050) );
  XOR U5545 ( .A(n4053), .B(n4054), .Z(out[270]) );
  ANDN U5546 ( .B(n4055), .A(n4056), .Z(n4053) );
  XOR U5547 ( .A(n4057), .B(n1432), .Z(out[26]) );
  NOR U5548 ( .A(n1433), .B(n4015), .Z(n4057) );
  XOR U5549 ( .A(n3469), .B(n4058), .Z(n1433) );
  IV U5550 ( .A(n2427), .Z(n3469) );
  XOR U5551 ( .A(n4059), .B(n1916), .Z(out[269]) );
  AND U5552 ( .A(n4060), .B(n4061), .Z(n4059) );
  XOR U5553 ( .A(n4062), .B(n1965), .Z(out[268]) );
  ANDN U5554 ( .B(n4063), .A(n4064), .Z(n4062) );
  XNOR U5555 ( .A(n4065), .B(n2002), .Z(out[267]) );
  ANDN U5556 ( .B(n4066), .A(n4067), .Z(n4065) );
  XOR U5557 ( .A(n4068), .B(n2037), .Z(out[266]) );
  ANDN U5558 ( .B(n4069), .A(n4070), .Z(n4068) );
  XOR U5559 ( .A(n4071), .B(n2076), .Z(out[265]) );
  XOR U5560 ( .A(n3521), .B(n4072), .Z(n2076) );
  XOR U5561 ( .A(n4074), .B(n1477), .Z(out[264]) );
  XOR U5562 ( .A(n4075), .B(n2560), .Z(n1477) );
  ANDN U5563 ( .B(n4076), .A(n1476), .Z(n4074) );
  XOR U5564 ( .A(n4077), .B(n1822), .Z(out[263]) );
  XOR U5565 ( .A(n4078), .B(n2567), .Z(n1822) );
  IV U5566 ( .A(n4080), .Z(n1821) );
  XOR U5567 ( .A(n4081), .B(n2184), .Z(out[262]) );
  XOR U5568 ( .A(n4082), .B(n2574), .Z(n2184) );
  ANDN U5569 ( .B(n4083), .A(n4084), .Z(n4081) );
  XNOR U5570 ( .A(n4085), .B(n2237), .Z(out[261]) );
  IV U5571 ( .A(n2857), .Z(n2237) );
  XNOR U5572 ( .A(n4086), .B(n2581), .Z(n2857) );
  NOR U5573 ( .A(n4087), .B(n2856), .Z(n4085) );
  XOR U5574 ( .A(n4088), .B(n2311), .Z(out[260]) );
  XOR U5575 ( .A(n4089), .B(n2588), .Z(n2311) );
  XNOR U5576 ( .A(n4091), .B(n1481), .Z(out[25]) );
  ANDN U5577 ( .B(n4019), .A(n1480), .Z(n4091) );
  XOR U5578 ( .A(n4093), .B(n2385), .Z(out[259]) );
  XNOR U5579 ( .A(n4094), .B(n3543), .Z(n2385) );
  XNOR U5580 ( .A(n4096), .B(n2459), .Z(out[258]) );
  IV U5581 ( .A(n3965), .Z(n2459) );
  XOR U5582 ( .A(n4097), .B(n2602), .Z(n3965) );
  NOR U5583 ( .A(n4098), .B(n3964), .Z(n4096) );
  XNOR U5584 ( .A(n4099), .B(n2533), .Z(out[257]) );
  IV U5585 ( .A(n4100), .Z(n2533) );
  ANDN U5586 ( .B(n4101), .A(n4102), .Z(n4099) );
  XNOR U5587 ( .A(n4103), .B(n2607), .Z(out[256]) );
  ANDN U5588 ( .B(n4104), .A(n4105), .Z(n4103) );
  XOR U5589 ( .A(n4106), .B(n2681), .Z(out[255]) );
  XOR U5590 ( .A(n4107), .B(n4108), .Z(n2681) );
  ANDN U5591 ( .B(n3920), .A(n4109), .Z(n4106) );
  XOR U5592 ( .A(n4110), .B(n2725), .Z(out[254]) );
  XOR U5593 ( .A(n1815), .B(n4111), .Z(n2725) );
  XOR U5594 ( .A(n4113), .B(n2769), .Z(out[253]) );
  XNOR U5595 ( .A(n1828), .B(n4114), .Z(n2769) );
  NOR U5596 ( .A(n4115), .B(n3924), .Z(n4113) );
  XOR U5597 ( .A(n4116), .B(n2813), .Z(out[252]) );
  XOR U5598 ( .A(n4117), .B(n4118), .Z(n2813) );
  ANDN U5599 ( .B(n4119), .A(n4120), .Z(n4116) );
  XOR U5600 ( .A(n4121), .B(n2860), .Z(out[251]) );
  XNOR U5601 ( .A(n1837), .B(n4122), .Z(n2860) );
  ANDN U5602 ( .B(n4123), .A(n3928), .Z(n4121) );
  XOR U5603 ( .A(n4124), .B(n2904), .Z(out[250]) );
  XOR U5604 ( .A(n1841), .B(n4125), .Z(n2904) );
  ANDN U5605 ( .B(n4126), .A(n3930), .Z(n4124) );
  XNOR U5606 ( .A(n4127), .B(n1516), .Z(out[24]) );
  NOR U5607 ( .A(n4021), .B(n1515), .Z(n4127) );
  XNOR U5608 ( .A(n4128), .B(n4129), .Z(n1515) );
  XNOR U5609 ( .A(n4130), .B(n2949), .Z(out[249]) );
  XOR U5610 ( .A(n1846), .B(n4131), .Z(n2949) );
  ANDN U5611 ( .B(n4132), .A(n3932), .Z(n4130) );
  XNOR U5612 ( .A(n4133), .B(n2983), .Z(out[248]) );
  XOR U5613 ( .A(n1850), .B(n4134), .Z(n2983) );
  ANDN U5614 ( .B(n4135), .A(n3934), .Z(n4133) );
  XOR U5615 ( .A(n4136), .B(n3010), .Z(out[247]) );
  XNOR U5616 ( .A(n3641), .B(n4137), .Z(n3010) );
  ANDN U5617 ( .B(n4138), .A(n3936), .Z(n4136) );
  XNOR U5618 ( .A(n4139), .B(n3036), .Z(out[246]) );
  XOR U5619 ( .A(n1858), .B(n4140), .Z(n3036) );
  ANDN U5620 ( .B(n4141), .A(n3938), .Z(n4139) );
  XOR U5621 ( .A(n4142), .B(n3062), .Z(out[245]) );
  XOR U5622 ( .A(n1862), .B(n4143), .Z(n3062) );
  NOR U5623 ( .A(n4144), .B(n3942), .Z(n4142) );
  XOR U5624 ( .A(n4145), .B(n3091), .Z(out[244]) );
  XNOR U5625 ( .A(n1866), .B(n4146), .Z(n3091) );
  ANDN U5626 ( .B(n4147), .A(n3944), .Z(n4145) );
  XOR U5627 ( .A(n4148), .B(n3118), .Z(out[243]) );
  XNOR U5628 ( .A(n1874), .B(n4149), .Z(n3118) );
  XNOR U5629 ( .A(n4151), .B(n3148), .Z(out[242]) );
  XOR U5630 ( .A(n1878), .B(n4152), .Z(n3148) );
  ANDN U5631 ( .B(n4153), .A(n3948), .Z(n4151) );
  XOR U5632 ( .A(n4154), .B(n3188), .Z(out[241]) );
  XNOR U5633 ( .A(n1882), .B(n4155), .Z(n3188) );
  ANDN U5634 ( .B(n4156), .A(n4157), .Z(n4154) );
  XOR U5635 ( .A(n4158), .B(n3227), .Z(out[240]) );
  XOR U5636 ( .A(n3675), .B(n4159), .Z(n3227) );
  NOR U5637 ( .A(n4160), .B(n3952), .Z(n4158) );
  XNOR U5638 ( .A(n4161), .B(n1539), .Z(out[23]) );
  NOR U5639 ( .A(n1540), .B(n4027), .Z(n4161) );
  XOR U5640 ( .A(n2448), .B(n4162), .Z(n1540) );
  XNOR U5641 ( .A(n4163), .B(n3266), .Z(out[239]) );
  IV U5642 ( .A(n3955), .Z(n3266) );
  XOR U5643 ( .A(n1891), .B(n4164), .Z(n3955) );
  ANDN U5644 ( .B(n4165), .A(n3954), .Z(n4163) );
  XNOR U5645 ( .A(n4166), .B(n3309), .Z(out[238]) );
  XOR U5646 ( .A(n1895), .B(n4167), .Z(n3309) );
  ANDN U5647 ( .B(n4168), .A(n3957), .Z(n4166) );
  XOR U5648 ( .A(n4169), .B(n3349), .Z(out[237]) );
  XNOR U5649 ( .A(n1899), .B(n4170), .Z(n3349) );
  ANDN U5650 ( .B(n4171), .A(n3959), .Z(n4169) );
  XNOR U5651 ( .A(n4172), .B(n3394), .Z(out[236]) );
  IV U5652 ( .A(n3962), .Z(n3394) );
  XOR U5653 ( .A(n1903), .B(n4173), .Z(n3962) );
  ANDN U5654 ( .B(n4174), .A(n3961), .Z(n4172) );
  XOR U5655 ( .A(n4175), .B(n3427), .Z(out[235]) );
  XOR U5656 ( .A(n4176), .B(n4177), .Z(n3427) );
  ANDN U5657 ( .B(n3969), .A(n4178), .Z(n4175) );
  IV U5658 ( .A(n4179), .Z(n3969) );
  XOR U5659 ( .A(n4180), .B(n3459), .Z(out[234]) );
  XOR U5660 ( .A(n4181), .B(n4182), .Z(n3459) );
  ANDN U5661 ( .B(n4183), .A(n3971), .Z(n4180) );
  XOR U5662 ( .A(n4184), .B(n3494), .Z(out[233]) );
  XOR U5663 ( .A(n3708), .B(n4185), .Z(n3494) );
  ANDN U5664 ( .B(n4186), .A(n3973), .Z(n4184) );
  XOR U5665 ( .A(n4187), .B(n3525), .Z(out[232]) );
  XOR U5666 ( .A(n3714), .B(n4188), .Z(n3525) );
  ANDN U5667 ( .B(n3975), .A(n4189), .Z(n4187) );
  XOR U5668 ( .A(n4190), .B(n3559), .Z(out[231]) );
  XOR U5669 ( .A(n1928), .B(n4191), .Z(n3559) );
  ANDN U5670 ( .B(n4192), .A(n4193), .Z(n4190) );
  XOR U5671 ( .A(n4194), .B(n3586), .Z(out[230]) );
  XOR U5672 ( .A(n1932), .B(n4195), .Z(n3586) );
  NOR U5673 ( .A(n4196), .B(n3979), .Z(n4194) );
  XNOR U5674 ( .A(n4197), .B(n1568), .Z(out[22]) );
  NOR U5675 ( .A(n1569), .B(n4030), .Z(n4197) );
  XOR U5676 ( .A(n2455), .B(n4198), .Z(n1569) );
  IV U5677 ( .A(n4199), .Z(n2455) );
  XOR U5678 ( .A(n4200), .B(n3623), .Z(out[229]) );
  XOR U5679 ( .A(n1937), .B(n4201), .Z(n3623) );
  ANDN U5680 ( .B(n4202), .A(n3981), .Z(n4200) );
  XOR U5681 ( .A(n4203), .B(n3672), .Z(out[228]) );
  XOR U5682 ( .A(n1941), .B(n4204), .Z(n3672) );
  ANDN U5683 ( .B(n3983), .A(n4205), .Z(n4203) );
  XOR U5684 ( .A(n4206), .B(n3724), .Z(out[227]) );
  XNOR U5685 ( .A(n1946), .B(n4207), .Z(n3724) );
  NOR U5686 ( .A(n1035), .B(n3986), .Z(n4206) );
  XOR U5687 ( .A(n4208), .B(n3772), .Z(out[226]) );
  XNOR U5688 ( .A(n1951), .B(n4209), .Z(n3772) );
  NOR U5689 ( .A(n3989), .B(n1079), .Z(n4208) );
  XOR U5690 ( .A(n4210), .B(n3824), .Z(out[225]) );
  XNOR U5691 ( .A(n1955), .B(n4211), .Z(n3824) );
  NOR U5692 ( .A(n4212), .B(n1123), .Z(n4210) );
  XNOR U5693 ( .A(n4213), .B(n3872), .Z(out[224]) );
  XOR U5694 ( .A(n4214), .B(n4215), .Z(n3872) );
  ANDN U5695 ( .B(n3997), .A(n4216), .Z(n4213) );
  XOR U5696 ( .A(n4217), .B(n3918), .Z(out[223]) );
  XOR U5697 ( .A(n4218), .B(n4219), .Z(n3918) );
  NOR U5698 ( .A(n4000), .B(n1211), .Z(n4217) );
  XOR U5699 ( .A(n4220), .B(n4004), .Z(out[222]) );
  XOR U5700 ( .A(n4221), .B(n4222), .Z(n4004) );
  ANDN U5701 ( .B(n4003), .A(n4223), .Z(n4220) );
  IV U5702 ( .A(n4224), .Z(n4003) );
  XNOR U5703 ( .A(n4225), .B(n3967), .Z(out[221]) );
  NOR U5704 ( .A(n4007), .B(n1299), .Z(n4225) );
  XOR U5705 ( .A(n4227), .B(n3991), .Z(out[220]) );
  XNOR U5706 ( .A(n4228), .B(n1667), .Z(n3991) );
  ANDN U5707 ( .B(n4010), .A(n1343), .Z(n4227) );
  IV U5708 ( .A(n4229), .Z(n1343) );
  XOR U5709 ( .A(n4230), .B(n1592), .Z(out[21]) );
  ANDN U5710 ( .B(n4033), .A(n1593), .Z(n4230) );
  XOR U5711 ( .A(n2466), .B(n4231), .Z(n1593) );
  XNOR U5712 ( .A(n4232), .B(n4012), .Z(out[219]) );
  XOR U5713 ( .A(n4233), .B(n4234), .Z(n4012) );
  NOR U5714 ( .A(n4013), .B(n1387), .Z(n4232) );
  XNOR U5715 ( .A(n4235), .B(n4015), .Z(out[218]) );
  XNOR U5716 ( .A(n4236), .B(n4237), .Z(n4015) );
  ANDN U5717 ( .B(n4016), .A(n4238), .Z(n4235) );
  XOR U5718 ( .A(n4239), .B(n4019), .Z(out[217]) );
  XNOR U5719 ( .A(n4240), .B(n1685), .Z(n4019) );
  NOR U5720 ( .A(n4018), .B(n1479), .Z(n4239) );
  XNOR U5721 ( .A(n4241), .B(n4021), .Z(out[216]) );
  XNOR U5722 ( .A(n4242), .B(n1689), .Z(n4021) );
  NOR U5723 ( .A(n4243), .B(n1514), .Z(n4241) );
  XNOR U5724 ( .A(n4244), .B(n4027), .Z(out[215]) );
  XOR U5725 ( .A(n4245), .B(n1693), .Z(n4027) );
  NOR U5726 ( .A(n1538), .B(n4026), .Z(n4244) );
  IV U5727 ( .A(n4246), .Z(n1538) );
  XNOR U5728 ( .A(n4247), .B(n4030), .Z(out[214]) );
  XNOR U5729 ( .A(n4248), .B(n4249), .Z(n4030) );
  NOR U5730 ( .A(n4029), .B(n1567), .Z(n4247) );
  XOR U5731 ( .A(n4250), .B(n4033), .Z(out[213]) );
  XOR U5732 ( .A(n4251), .B(n1703), .Z(n4033) );
  ANDN U5733 ( .B(n1591), .A(n4032), .Z(n4250) );
  XNOR U5734 ( .A(n4252), .B(n4035), .Z(out[212]) );
  NOR U5735 ( .A(n4253), .B(n1615), .Z(n4252) );
  XNOR U5736 ( .A(n4254), .B(n4038), .Z(out[211]) );
  NOR U5737 ( .A(n4255), .B(n1639), .Z(n4254) );
  XNOR U5738 ( .A(n4256), .B(n4041), .Z(out[210]) );
  XNOR U5739 ( .A(n4257), .B(n1617), .Z(out[20]) );
  NOR U5740 ( .A(n4035), .B(n1616), .Z(n4257) );
  XOR U5741 ( .A(n3485), .B(n4258), .Z(n1616) );
  XNOR U5742 ( .A(n4259), .B(n1708), .Z(n4035) );
  XNOR U5743 ( .A(n4260), .B(n4044), .Z(out[209]) );
  XNOR U5744 ( .A(n4261), .B(n4262), .Z(out[208]) );
  XOR U5745 ( .A(n4263), .B(n4051), .Z(out[207]) );
  ANDN U5746 ( .B(n4052), .A(n4264), .Z(n4263) );
  XNOR U5747 ( .A(n4265), .B(n4055), .Z(out[206]) );
  NOR U5748 ( .A(n4266), .B(n1870), .Z(n4265) );
  XNOR U5749 ( .A(n4267), .B(n4061), .Z(out[205]) );
  NOR U5750 ( .A(n4060), .B(n1915), .Z(n4267) );
  XNOR U5751 ( .A(n4268), .B(n4063), .Z(out[204]) );
  NOR U5752 ( .A(n4269), .B(n1964), .Z(n4268) );
  XNOR U5753 ( .A(n4270), .B(n4066), .Z(out[203]) );
  ANDN U5754 ( .B(n2000), .A(n4271), .Z(n4270) );
  XNOR U5755 ( .A(n4272), .B(n4069), .Z(out[202]) );
  ANDN U5756 ( .B(n2036), .A(n4273), .Z(n4272) );
  XNOR U5757 ( .A(n4274), .B(n1033), .Z(out[201]) );
  XOR U5758 ( .A(n3866), .B(n4275), .Z(n1033) );
  NOR U5759 ( .A(n4073), .B(n2075), .Z(n4274) );
  XOR U5760 ( .A(n4276), .B(n1476), .Z(out[200]) );
  XOR U5761 ( .A(n4277), .B(n1767), .Z(n1476) );
  XOR U5762 ( .A(n4278), .B(n2534), .Z(out[1]) );
  ANDN U5763 ( .B(n4102), .A(n4100), .Z(n4278) );
  XOR U5764 ( .A(n4279), .B(n2613), .Z(n4100) );
  IV U5765 ( .A(n4280), .Z(n4102) );
  XNOR U5766 ( .A(n4281), .B(n1641), .Z(out[19]) );
  NOR U5767 ( .A(n4038), .B(n1640), .Z(n4281) );
  XOR U5768 ( .A(n3489), .B(n4282), .Z(n1640) );
  XOR U5769 ( .A(n4283), .B(n1713), .Z(n4038) );
  XOR U5770 ( .A(n4284), .B(n4080), .Z(out[199]) );
  XOR U5771 ( .A(n4285), .B(n1775), .Z(n4080) );
  NOR U5772 ( .A(n4079), .B(n2149), .Z(n4284) );
  XNOR U5773 ( .A(n4286), .B(n2234), .Z(out[198]) );
  IV U5774 ( .A(n4084), .Z(n2234) );
  XOR U5775 ( .A(n4287), .B(n1780), .Z(n4084) );
  NOR U5776 ( .A(n2183), .B(n4083), .Z(n4286) );
  XOR U5777 ( .A(n4288), .B(n2856), .Z(out[197]) );
  XNOR U5778 ( .A(n4289), .B(n1785), .Z(n2856) );
  IV U5779 ( .A(n4290), .Z(n4087) );
  XNOR U5780 ( .A(n4291), .B(n3185), .Z(out[196]) );
  XOR U5781 ( .A(n4292), .B(n1790), .Z(n3185) );
  IV U5782 ( .A(n4293), .Z(n1790) );
  NOR U5783 ( .A(n2310), .B(n4090), .Z(n4291) );
  XNOR U5784 ( .A(n4294), .B(n3556), .Z(out[195]) );
  XOR U5785 ( .A(n4295), .B(n1794), .Z(n3556) );
  NOR U5786 ( .A(n4095), .B(n2384), .Z(n4294) );
  XOR U5787 ( .A(n4296), .B(n3964), .Z(out[194]) );
  XOR U5788 ( .A(n1798), .B(n4297), .Z(n3964) );
  ANDN U5789 ( .B(n2458), .A(n4298), .Z(n4296) );
  XNOR U5790 ( .A(n4299), .B(n4280), .Z(out[193]) );
  XNOR U5791 ( .A(n4300), .B(n1804), .Z(n4280) );
  NOR U5792 ( .A(n2532), .B(n4101), .Z(n4299) );
  IV U5793 ( .A(n4301), .Z(n2532) );
  XOR U5794 ( .A(n4302), .B(n4105), .Z(out[192]) );
  NOR U5795 ( .A(n4303), .B(n4104), .Z(n4302) );
  XNOR U5796 ( .A(n4304), .B(n3920), .Z(out[191]) );
  XNOR U5797 ( .A(n4305), .B(n2089), .Z(n3920) );
  ANDN U5798 ( .B(n4109), .A(n2680), .Z(n4304) );
  IV U5799 ( .A(n4306), .Z(n2680) );
  IV U5800 ( .A(n4307), .Z(n4109) );
  XOR U5801 ( .A(n4308), .B(n3922), .Z(out[190]) );
  XOR U5802 ( .A(n4309), .B(n2092), .Z(n3922) );
  NOR U5803 ( .A(n4112), .B(n2724), .Z(n4308) );
  XOR U5804 ( .A(n4310), .B(n1672), .Z(out[18]) );
  NOR U5805 ( .A(n4041), .B(n1671), .Z(n4310) );
  XOR U5806 ( .A(n2487), .B(n4311), .Z(n1671) );
  XNOR U5807 ( .A(n4312), .B(n1718), .Z(n4041) );
  XOR U5808 ( .A(n4313), .B(n3924), .Z(out[189]) );
  XNOR U5809 ( .A(n4314), .B(n2095), .Z(n3924) );
  ANDN U5810 ( .B(n2768), .A(n4315), .Z(n4313) );
  XNOR U5811 ( .A(n4316), .B(n3926), .Z(out[188]) );
  IV U5812 ( .A(n4120), .Z(n3926) );
  XNOR U5813 ( .A(n4317), .B(n2098), .Z(n4120) );
  ANDN U5814 ( .B(n2812), .A(n4119), .Z(n4316) );
  XOR U5815 ( .A(n4318), .B(n3928), .Z(out[187]) );
  XNOR U5816 ( .A(n4319), .B(n2101), .Z(n3928) );
  ANDN U5817 ( .B(n2859), .A(n4123), .Z(n4318) );
  XOR U5818 ( .A(n4320), .B(n3930), .Z(out[186]) );
  XNOR U5819 ( .A(n2104), .B(n4321), .Z(n3930) );
  ANDN U5820 ( .B(n2903), .A(n4126), .Z(n4320) );
  XOR U5821 ( .A(n4322), .B(n3932), .Z(out[185]) );
  XOR U5822 ( .A(n4323), .B(n4324), .Z(n3932) );
  NOR U5823 ( .A(n2947), .B(n4132), .Z(n4322) );
  XOR U5824 ( .A(n4325), .B(n3934), .Z(out[184]) );
  XOR U5825 ( .A(n4326), .B(n2114), .Z(n3934) );
  NOR U5826 ( .A(n2981), .B(n4135), .Z(n4325) );
  XOR U5827 ( .A(n4327), .B(n3936), .Z(out[183]) );
  XOR U5828 ( .A(n4328), .B(n4329), .Z(n3936) );
  NOR U5829 ( .A(n4138), .B(n3009), .Z(n4327) );
  XOR U5830 ( .A(n4330), .B(n3938), .Z(out[182]) );
  XOR U5831 ( .A(n4331), .B(n4332), .Z(n3938) );
  NOR U5832 ( .A(n4141), .B(n3034), .Z(n4330) );
  XOR U5833 ( .A(n4333), .B(n3942), .Z(out[181]) );
  XNOR U5834 ( .A(n2124), .B(n4334), .Z(n3942) );
  ANDN U5835 ( .B(n3061), .A(n4335), .Z(n4333) );
  XOR U5836 ( .A(n4336), .B(n3944), .Z(out[180]) );
  XNOR U5837 ( .A(n2128), .B(n4337), .Z(n3944) );
  NOR U5838 ( .A(n3090), .B(n4147), .Z(n4336) );
  XOR U5839 ( .A(n4338), .B(n1724), .Z(out[17]) );
  ANDN U5840 ( .B(n1723), .A(n4044), .Z(n4338) );
  XNOR U5841 ( .A(n4339), .B(n1727), .Z(n4044) );
  XNOR U5842 ( .A(n2492), .B(n4340), .Z(n1723) );
  XNOR U5843 ( .A(n4341), .B(n3946), .Z(out[179]) );
  XOR U5844 ( .A(n2131), .B(n4342), .Z(n3946) );
  XOR U5845 ( .A(n4343), .B(n3948), .Z(out[178]) );
  XOR U5846 ( .A(n2134), .B(n4344), .Z(n3948) );
  NOR U5847 ( .A(n3146), .B(n4153), .Z(n4343) );
  XNOR U5848 ( .A(n4345), .B(n3950), .Z(out[177]) );
  IV U5849 ( .A(n4157), .Z(n3950) );
  XOR U5850 ( .A(n4346), .B(n2139), .Z(n4157) );
  NOR U5851 ( .A(n3187), .B(n4156), .Z(n4345) );
  XOR U5852 ( .A(n4347), .B(n3952), .Z(out[176]) );
  XNOR U5853 ( .A(n4348), .B(n2142), .Z(n3952) );
  ANDN U5854 ( .B(n4160), .A(n3226), .Z(n4347) );
  XOR U5855 ( .A(n4349), .B(n3954), .Z(out[175]) );
  XOR U5856 ( .A(n4350), .B(n2146), .Z(n3954) );
  NOR U5857 ( .A(n3265), .B(n4165), .Z(n4349) );
  XOR U5858 ( .A(n4351), .B(n3957), .Z(out[174]) );
  XOR U5859 ( .A(n4352), .B(n2152), .Z(n3957) );
  NOR U5860 ( .A(n4168), .B(n3307), .Z(n4351) );
  XOR U5861 ( .A(n4353), .B(n3959), .Z(out[173]) );
  XOR U5862 ( .A(n4354), .B(n2155), .Z(n3959) );
  NOR U5863 ( .A(n4171), .B(n3348), .Z(n4353) );
  XOR U5864 ( .A(n4355), .B(n3961), .Z(out[172]) );
  XOR U5865 ( .A(n4356), .B(n2158), .Z(n3961) );
  NOR U5866 ( .A(n3392), .B(n4174), .Z(n4355) );
  XOR U5867 ( .A(n4357), .B(n4179), .Z(out[171]) );
  XOR U5868 ( .A(n4358), .B(n2161), .Z(n4179) );
  XOR U5869 ( .A(n4359), .B(n3971), .Z(out[170]) );
  XOR U5870 ( .A(n4360), .B(n2164), .Z(n3971) );
  NOR U5871 ( .A(n3458), .B(n4183), .Z(n4359) );
  XOR U5872 ( .A(n4361), .B(n1772), .Z(out[16]) );
  ANDN U5873 ( .B(n4049), .A(n4047), .Z(n4361) );
  XNOR U5874 ( .A(n4362), .B(n2502), .Z(n4047) );
  IV U5875 ( .A(n4262), .Z(n4049) );
  XOR U5876 ( .A(n4363), .B(n1732), .Z(n4262) );
  XOR U5877 ( .A(n4364), .B(n3973), .Z(out[169]) );
  XOR U5878 ( .A(n4365), .B(n2169), .Z(n3973) );
  ANDN U5879 ( .B(n3493), .A(n4186), .Z(n4364) );
  XNOR U5880 ( .A(n4366), .B(n3975), .Z(out[168]) );
  XOR U5881 ( .A(n4367), .B(n2172), .Z(n3975) );
  IV U5882 ( .A(n3780), .Z(n2172) );
  NOR U5883 ( .A(n4368), .B(n3524), .Z(n4366) );
  XNOR U5884 ( .A(n4369), .B(n3977), .Z(out[167]) );
  IV U5885 ( .A(n4193), .Z(n3977) );
  XOR U5886 ( .A(n4370), .B(n2175), .Z(n4193) );
  NOR U5887 ( .A(n3558), .B(n4192), .Z(n4369) );
  XOR U5888 ( .A(n4371), .B(n3979), .Z(out[166]) );
  XOR U5889 ( .A(n4372), .B(n2178), .Z(n3979) );
  NOR U5890 ( .A(n4373), .B(n3585), .Z(n4371) );
  XOR U5891 ( .A(n4374), .B(n3981), .Z(out[165]) );
  XOR U5892 ( .A(n4375), .B(n2181), .Z(n3981) );
  NOR U5893 ( .A(n3622), .B(n4202), .Z(n4374) );
  IV U5894 ( .A(n4376), .Z(n3622) );
  XNOR U5895 ( .A(n4377), .B(n3983), .Z(out[164]) );
  XNOR U5896 ( .A(n4378), .B(n2188), .Z(n3983) );
  NOR U5897 ( .A(n4379), .B(n3671), .Z(n4377) );
  XOR U5898 ( .A(n4380), .B(n3986), .Z(out[163]) );
  XNOR U5899 ( .A(n4381), .B(n2191), .Z(n3986) );
  IV U5900 ( .A(n3805), .Z(n2191) );
  ANDN U5901 ( .B(n1035), .A(n1036), .Z(n4380) );
  XOR U5902 ( .A(n2425), .B(n4382), .Z(n1036) );
  XOR U5903 ( .A(n2585), .B(n4383), .Z(n1035) );
  XOR U5904 ( .A(n4384), .B(n3989), .Z(out[162]) );
  XOR U5905 ( .A(n4385), .B(n2194), .Z(n3989) );
  ANDN U5906 ( .B(n1079), .A(n1081), .Z(n4384) );
  XNOR U5907 ( .A(n2432), .B(n4386), .Z(n1081) );
  XOR U5908 ( .A(n4387), .B(n4388), .Z(n1079) );
  XNOR U5909 ( .A(n4389), .B(n3994), .Z(out[161]) );
  IV U5910 ( .A(n4212), .Z(n3994) );
  XOR U5911 ( .A(n4390), .B(n2197), .Z(n4212) );
  ANDN U5912 ( .B(n1123), .A(n1125), .Z(n4389) );
  XOR U5913 ( .A(n4391), .B(n2440), .Z(n1125) );
  XOR U5914 ( .A(n2599), .B(n4392), .Z(n1123) );
  XNOR U5915 ( .A(n4393), .B(n3997), .Z(out[160]) );
  XOR U5916 ( .A(n4394), .B(n2200), .Z(n3997) );
  IV U5917 ( .A(n3820), .Z(n2200) );
  ANDN U5918 ( .B(n1169), .A(n1167), .Z(n4393) );
  IV U5919 ( .A(n4216), .Z(n1167) );
  XOR U5920 ( .A(n4395), .B(n2611), .Z(n4216) );
  XOR U5921 ( .A(n4396), .B(n2447), .Z(n1169) );
  XOR U5922 ( .A(n4397), .B(n1825), .Z(out[15]) );
  AND U5923 ( .A(n4051), .B(n1826), .Z(n4397) );
  XOR U5924 ( .A(n2506), .B(n4398), .Z(n1826) );
  XOR U5925 ( .A(n4399), .B(n1736), .Z(n4051) );
  XOR U5926 ( .A(n4400), .B(n4000), .Z(out[159]) );
  XOR U5927 ( .A(n4401), .B(n2203), .Z(n4000) );
  ANDN U5928 ( .B(n1211), .A(n1213), .Z(n4400) );
  XNOR U5929 ( .A(n4402), .B(n3238), .Z(n1213) );
  XOR U5930 ( .A(n4403), .B(n3789), .Z(n1211) );
  XOR U5931 ( .A(n4404), .B(n4405), .Z(out[1599]) );
  XOR U5932 ( .A(n4406), .B(n4407), .Z(n4405) );
  AND U5933 ( .A(n4408), .B(n4409), .Z(n4406) );
  XNOR U5934 ( .A(n4410), .B(n4411), .Z(out[1598]) );
  XNOR U5935 ( .A(n4414), .B(n4415), .Z(out[1597]) );
  ANDN U5936 ( .B(n4416), .A(n4417), .Z(n4414) );
  XOR U5937 ( .A(n4418), .B(n4419), .Z(out[1596]) );
  AND U5938 ( .A(n4420), .B(n4421), .Z(n4418) );
  XNOR U5939 ( .A(n4422), .B(n4423), .Z(out[1595]) );
  AND U5940 ( .A(n4424), .B(n4425), .Z(n4422) );
  XNOR U5941 ( .A(n4426), .B(n4427), .Z(out[1594]) );
  AND U5942 ( .A(n4428), .B(n4429), .Z(n4426) );
  XNOR U5943 ( .A(n4430), .B(n4431), .Z(out[1593]) );
  AND U5944 ( .A(n4432), .B(n4433), .Z(n4430) );
  XOR U5945 ( .A(n4434), .B(n4435), .Z(out[1592]) );
  ANDN U5946 ( .B(n4436), .A(n4437), .Z(n4434) );
  XOR U5947 ( .A(n4438), .B(n4439), .Z(out[1591]) );
  NOR U5948 ( .A(n4440), .B(n4441), .Z(n4438) );
  XOR U5949 ( .A(n4442), .B(n4443), .Z(out[1590]) );
  XOR U5950 ( .A(n4446), .B(n4224), .Z(out[158]) );
  XOR U5951 ( .A(n4447), .B(n1977), .Z(n4224) );
  ANDN U5952 ( .B(n1257), .A(n1255), .Z(n4446) );
  IV U5953 ( .A(n4223), .Z(n1255) );
  XOR U5954 ( .A(n4448), .B(n3795), .Z(n4223) );
  XNOR U5955 ( .A(n4449), .B(n4450), .Z(n1257) );
  XOR U5956 ( .A(n4451), .B(n4452), .Z(out[1589]) );
  ANDN U5957 ( .B(n4453), .A(n4454), .Z(n4451) );
  XOR U5958 ( .A(n4455), .B(n4456), .Z(out[1588]) );
  ANDN U5959 ( .B(n4457), .A(n4458), .Z(n4455) );
  XOR U5960 ( .A(n4459), .B(n4460), .Z(out[1587]) );
  XOR U5961 ( .A(n4463), .B(n4464), .Z(out[1586]) );
  ANDN U5962 ( .B(n4465), .A(n4466), .Z(n4463) );
  XNOR U5963 ( .A(n4467), .B(n4468), .Z(out[1585]) );
  AND U5964 ( .A(n4469), .B(n4470), .Z(n4467) );
  XOR U5965 ( .A(n4471), .B(n4472), .Z(out[1584]) );
  ANDN U5966 ( .B(n4473), .A(n4474), .Z(n4471) );
  XOR U5967 ( .A(n4475), .B(n4476), .Z(out[1583]) );
  ANDN U5968 ( .B(n4477), .A(n4478), .Z(n4475) );
  XNOR U5969 ( .A(n4479), .B(n4480), .Z(out[1582]) );
  AND U5970 ( .A(n4481), .B(n4482), .Z(n4479) );
  XNOR U5971 ( .A(n4483), .B(n4484), .Z(out[1581]) );
  ANDN U5972 ( .B(n4485), .A(n4486), .Z(n4483) );
  XOR U5973 ( .A(n4487), .B(n4488), .Z(out[1580]) );
  AND U5974 ( .A(n4489), .B(n4490), .Z(n4487) );
  XOR U5975 ( .A(n4491), .B(n4007), .Z(out[157]) );
  XOR U5976 ( .A(n4492), .B(n1980), .Z(n4007) );
  ANDN U5977 ( .B(n1299), .A(n1301), .Z(n4491) );
  XNOR U5978 ( .A(n4493), .B(n2472), .Z(n1301) );
  XNOR U5979 ( .A(n4494), .B(n3801), .Z(n1299) );
  XOR U5980 ( .A(n4495), .B(n4496), .Z(out[1579]) );
  AND U5981 ( .A(n4497), .B(n4498), .Z(n4495) );
  XOR U5982 ( .A(n4499), .B(n4500), .Z(out[1578]) );
  AND U5983 ( .A(n4501), .B(n4502), .Z(n4499) );
  XOR U5984 ( .A(n4503), .B(n4504), .Z(out[1577]) );
  XNOR U5985 ( .A(n4507), .B(n4508), .Z(out[1576]) );
  XNOR U5986 ( .A(n4511), .B(n4512), .Z(out[1575]) );
  XOR U5987 ( .A(n4515), .B(n4516), .Z(out[1574]) );
  XOR U5988 ( .A(n4519), .B(n4520), .Z(out[1573]) );
  ANDN U5989 ( .B(n4521), .A(n4522), .Z(n4519) );
  XNOR U5990 ( .A(n4523), .B(n4524), .Z(out[1572]) );
  ANDN U5991 ( .B(n4525), .A(n4526), .Z(n4523) );
  XNOR U5992 ( .A(n4527), .B(n4528), .Z(out[1571]) );
  ANDN U5993 ( .B(n4529), .A(n4530), .Z(n4527) );
  XNOR U5994 ( .A(n4531), .B(n4532), .Z(out[1570]) );
  AND U5995 ( .A(n4533), .B(n4534), .Z(n4531) );
  XNOR U5996 ( .A(n4535), .B(n4010), .Z(out[156]) );
  XOR U5997 ( .A(n4536), .B(n1983), .Z(n4010) );
  NOR U5998 ( .A(n4229), .B(n1344), .Z(n4535) );
  XOR U5999 ( .A(n4537), .B(n2479), .Z(n1344) );
  XOR U6000 ( .A(n4538), .B(n2639), .Z(n4229) );
  XOR U6001 ( .A(n4539), .B(n4540), .Z(out[1569]) );
  NOR U6002 ( .A(n4541), .B(n4542), .Z(n4539) );
  XNOR U6003 ( .A(n4543), .B(n4544), .Z(out[1568]) );
  AND U6004 ( .A(n4545), .B(n4546), .Z(n4543) );
  XNOR U6005 ( .A(n4547), .B(n4548), .Z(out[1567]) );
  XNOR U6006 ( .A(n4549), .B(n4550), .Z(n4548) );
  XOR U6007 ( .A(n4553), .B(n4554), .Z(out[1566]) );
  ANDN U6008 ( .B(n4555), .A(n4556), .Z(n4553) );
  XNOR U6009 ( .A(n4557), .B(n4558), .Z(out[1565]) );
  ANDN U6010 ( .B(n4559), .A(n4560), .Z(n4557) );
  XOR U6011 ( .A(n4561), .B(n4562), .Z(out[1564]) );
  ANDN U6012 ( .B(n4563), .A(n4564), .Z(n4561) );
  XNOR U6013 ( .A(n4565), .B(n4566), .Z(out[1563]) );
  XNOR U6014 ( .A(n4569), .B(n4570), .Z(out[1562]) );
  ANDN U6015 ( .B(n4571), .A(n4572), .Z(n4569) );
  XNOR U6016 ( .A(n4573), .B(n4574), .Z(out[1561]) );
  ANDN U6017 ( .B(n4575), .A(n4576), .Z(n4573) );
  XNOR U6018 ( .A(n4577), .B(n4578), .Z(out[1560]) );
  AND U6019 ( .A(n4579), .B(n4580), .Z(n4577) );
  XOR U6020 ( .A(n4581), .B(n4013), .Z(out[155]) );
  XNOR U6021 ( .A(n4582), .B(n1986), .Z(n4013) );
  ANDN U6022 ( .B(n1387), .A(n1388), .Z(n4581) );
  XOR U6023 ( .A(n4583), .B(n2486), .Z(n1388) );
  XNOR U6024 ( .A(n4584), .B(n3811), .Z(n1387) );
  XNOR U6025 ( .A(n4585), .B(n4586), .Z(out[1559]) );
  XOR U6026 ( .A(n4589), .B(n4590), .Z(out[1558]) );
  AND U6027 ( .A(n4591), .B(n4592), .Z(n4589) );
  XNOR U6028 ( .A(n4593), .B(n4594), .Z(out[1557]) );
  ANDN U6029 ( .B(n4595), .A(n4596), .Z(n4593) );
  XNOR U6030 ( .A(n4597), .B(n4598), .Z(out[1556]) );
  ANDN U6031 ( .B(n4599), .A(n4600), .Z(n4597) );
  XNOR U6032 ( .A(n4601), .B(n4602), .Z(out[1555]) );
  AND U6033 ( .A(n4603), .B(n4604), .Z(n4601) );
  XNOR U6034 ( .A(n4605), .B(n4606), .Z(out[1554]) );
  XOR U6035 ( .A(n4609), .B(n4610), .Z(out[1553]) );
  ANDN U6036 ( .B(n4611), .A(n4612), .Z(n4609) );
  XNOR U6037 ( .A(n4613), .B(n4614), .Z(out[1552]) );
  XNOR U6038 ( .A(n4617), .B(n4618), .Z(out[1551]) );
  XOR U6039 ( .A(n4619), .B(n4620), .Z(n4618) );
  AND U6040 ( .A(n4621), .B(n4622), .Z(n4619) );
  XNOR U6041 ( .A(n4623), .B(n4624), .Z(out[1550]) );
  XNOR U6042 ( .A(n4627), .B(n4016), .Z(out[154]) );
  XNOR U6043 ( .A(n4628), .B(n1989), .Z(n4016) );
  ANDN U6044 ( .B(n1432), .A(n1431), .Z(n4627) );
  IV U6045 ( .A(n4238), .Z(n1431) );
  XOR U6046 ( .A(n4629), .B(n2653), .Z(n4238) );
  XNOR U6047 ( .A(n4630), .B(n2495), .Z(n1432) );
  XNOR U6048 ( .A(n4631), .B(n4632), .Z(out[1549]) );
  XNOR U6049 ( .A(n4635), .B(n4636), .Z(out[1548]) );
  XNOR U6050 ( .A(n4639), .B(n4640), .Z(out[1547]) );
  AND U6051 ( .A(n4641), .B(n4642), .Z(n4639) );
  XNOR U6052 ( .A(n4643), .B(n4644), .Z(out[1546]) );
  ANDN U6053 ( .B(n4645), .A(n4646), .Z(n4643) );
  XNOR U6054 ( .A(n4647), .B(n4648), .Z(out[1545]) );
  ANDN U6055 ( .B(n4649), .A(n4650), .Z(n4647) );
  XOR U6056 ( .A(n4651), .B(n4652), .Z(out[1544]) );
  AND U6057 ( .A(n4653), .B(n4654), .Z(n4651) );
  XNOR U6058 ( .A(n4655), .B(n4656), .Z(out[1543]) );
  AND U6059 ( .A(n4657), .B(n4658), .Z(n4655) );
  XOR U6060 ( .A(n4659), .B(n4660), .Z(out[1542]) );
  AND U6061 ( .A(n4661), .B(n4662), .Z(n4659) );
  XNOR U6062 ( .A(n4663), .B(n4664), .Z(out[1541]) );
  ANDN U6063 ( .B(n4665), .A(n4666), .Z(n4663) );
  XOR U6064 ( .A(n4667), .B(n4668), .Z(out[1540]) );
  XOR U6065 ( .A(n4671), .B(n4018), .Z(out[153]) );
  XOR U6066 ( .A(n4672), .B(n1992), .Z(n4018) );
  ANDN U6067 ( .B(n1479), .A(n1481), .Z(n4671) );
  XOR U6068 ( .A(n4673), .B(n2500), .Z(n1481) );
  XOR U6069 ( .A(n4674), .B(n3822), .Z(n1479) );
  XOR U6070 ( .A(n4675), .B(n4676), .Z(out[1539]) );
  XOR U6071 ( .A(n4677), .B(n4678), .Z(n4676) );
  XOR U6072 ( .A(n4681), .B(n4682), .Z(out[1538]) );
  AND U6073 ( .A(n4683), .B(n4684), .Z(n4681) );
  XOR U6074 ( .A(n4685), .B(n4686), .Z(out[1537]) );
  XNOR U6075 ( .A(n4687), .B(n4688), .Z(n4686) );
  AND U6076 ( .A(n4689), .B(n4690), .Z(n4688) );
  XOR U6077 ( .A(n4691), .B(n4692), .Z(out[1536]) );
  XOR U6078 ( .A(n4693), .B(n4694), .Z(n4692) );
  XNOR U6079 ( .A(n4697), .B(n4408), .Z(out[1535]) );
  NOR U6080 ( .A(n4698), .B(n4409), .Z(n4697) );
  XNOR U6081 ( .A(n4699), .B(n4413), .Z(out[1534]) );
  ANDN U6082 ( .B(n4700), .A(n4412), .Z(n4699) );
  XNOR U6083 ( .A(n4701), .B(n4416), .Z(out[1533]) );
  ANDN U6084 ( .B(n4702), .A(n4703), .Z(n4701) );
  XNOR U6085 ( .A(n4704), .B(n4421), .Z(out[1532]) );
  ANDN U6086 ( .B(n4705), .A(n4420), .Z(n4704) );
  XNOR U6087 ( .A(n4706), .B(n4425), .Z(out[1531]) );
  ANDN U6088 ( .B(n4707), .A(n4424), .Z(n4706) );
  XNOR U6089 ( .A(n4708), .B(n4429), .Z(out[1530]) );
  ANDN U6090 ( .B(n4709), .A(n4428), .Z(n4708) );
  XNOR U6091 ( .A(n4710), .B(n4022), .Z(out[152]) );
  IV U6092 ( .A(n4243), .Z(n4022) );
  XNOR U6093 ( .A(n4711), .B(n1995), .Z(n4243) );
  ANDN U6094 ( .B(n1514), .A(n1516), .Z(n4710) );
  XOR U6095 ( .A(n4712), .B(n3261), .Z(n1516) );
  XOR U6096 ( .A(n4713), .B(n3828), .Z(n1514) );
  XNOR U6097 ( .A(n4714), .B(n4433), .Z(out[1529]) );
  ANDN U6098 ( .B(n4715), .A(n4432), .Z(n4714) );
  XOR U6099 ( .A(n4716), .B(n4437), .Z(out[1528]) );
  ANDN U6100 ( .B(n4717), .A(n4436), .Z(n4716) );
  XOR U6101 ( .A(n4718), .B(n4441), .Z(out[1527]) );
  ANDN U6102 ( .B(n4440), .A(n4719), .Z(n4718) );
  XNOR U6103 ( .A(n4720), .B(n4445), .Z(out[1526]) );
  NOR U6104 ( .A(n4721), .B(n4444), .Z(n4720) );
  XOR U6105 ( .A(n4722), .B(n4454), .Z(out[1525]) );
  NOR U6106 ( .A(n4723), .B(n4453), .Z(n4722) );
  XOR U6107 ( .A(n4724), .B(n4458), .Z(out[1524]) );
  NOR U6108 ( .A(n4725), .B(n4457), .Z(n4724) );
  XNOR U6109 ( .A(n4726), .B(n4462), .Z(out[1523]) );
  XOR U6110 ( .A(n4728), .B(n4466), .Z(out[1522]) );
  ANDN U6111 ( .B(n4729), .A(n4465), .Z(n4728) );
  XNOR U6112 ( .A(n4730), .B(n4470), .Z(out[1521]) );
  NOR U6113 ( .A(n4731), .B(n4469), .Z(n4730) );
  XOR U6114 ( .A(n4732), .B(n4474), .Z(out[1520]) );
  NOR U6115 ( .A(n4733), .B(n4473), .Z(n4732) );
  XOR U6116 ( .A(n4734), .B(n4026), .Z(out[151]) );
  XNOR U6117 ( .A(n4735), .B(n1998), .Z(n4026) );
  NOR U6118 ( .A(n4246), .B(n1539), .Z(n4734) );
  XNOR U6119 ( .A(n4736), .B(n2516), .Z(n1539) );
  XOR U6120 ( .A(n4737), .B(n2674), .Z(n4246) );
  XOR U6121 ( .A(n4738), .B(n4478), .Z(out[1519]) );
  NOR U6122 ( .A(n4739), .B(n4477), .Z(n4738) );
  XNOR U6123 ( .A(n4740), .B(n4482), .Z(out[1518]) );
  ANDN U6124 ( .B(n4741), .A(n4481), .Z(n4740) );
  XNOR U6125 ( .A(n4742), .B(n4485), .Z(out[1517]) );
  XNOR U6126 ( .A(n4744), .B(n4490), .Z(out[1516]) );
  ANDN U6127 ( .B(n4745), .A(n4489), .Z(n4744) );
  XNOR U6128 ( .A(n4746), .B(n4498), .Z(out[1515]) );
  ANDN U6129 ( .B(n4747), .A(n4497), .Z(n4746) );
  XNOR U6130 ( .A(n4748), .B(n4502), .Z(out[1514]) );
  ANDN U6131 ( .B(n4749), .A(n4501), .Z(n4748) );
  XNOR U6132 ( .A(n4750), .B(n4505), .Z(out[1513]) );
  ANDN U6133 ( .B(n4751), .A(n4506), .Z(n4750) );
  XNOR U6134 ( .A(n4752), .B(n4509), .Z(out[1512]) );
  ANDN U6135 ( .B(n4753), .A(n4510), .Z(n4752) );
  XNOR U6136 ( .A(n4754), .B(n4514), .Z(out[1511]) );
  ANDN U6137 ( .B(n4755), .A(n4513), .Z(n4754) );
  XNOR U6138 ( .A(n4756), .B(n4518), .Z(out[1510]) );
  ANDN U6139 ( .B(n4757), .A(n4517), .Z(n4756) );
  XOR U6140 ( .A(n4758), .B(n4029), .Z(out[150]) );
  XOR U6141 ( .A(n4759), .B(n2005), .Z(n4029) );
  ANDN U6142 ( .B(n1567), .A(n1568), .Z(n4758) );
  XOR U6143 ( .A(n4760), .B(n2523), .Z(n1568) );
  XNOR U6144 ( .A(n4761), .B(n4762), .Z(n1567) );
  XNOR U6145 ( .A(n4763), .B(n4521), .Z(out[1509]) );
  ANDN U6146 ( .B(n4522), .A(n4764), .Z(n4763) );
  IV U6147 ( .A(n4765), .Z(n4522) );
  XOR U6148 ( .A(n4766), .B(n4526), .Z(out[1508]) );
  ANDN U6149 ( .B(n4767), .A(n4525), .Z(n4766) );
  XNOR U6150 ( .A(n4768), .B(n4529), .Z(out[1507]) );
  ANDN U6151 ( .B(n4530), .A(n4769), .Z(n4768) );
  XNOR U6152 ( .A(n4770), .B(n4534), .Z(out[1506]) );
  ANDN U6153 ( .B(n4771), .A(n4533), .Z(n4770) );
  XOR U6154 ( .A(n4772), .B(n4542), .Z(out[1505]) );
  XNOR U6155 ( .A(n4774), .B(n4546), .Z(out[1504]) );
  ANDN U6156 ( .B(n4775), .A(n4545), .Z(n4774) );
  XOR U6157 ( .A(n4776), .B(n4551), .Z(out[1503]) );
  ANDN U6158 ( .B(n4777), .A(n4552), .Z(n4776) );
  XOR U6159 ( .A(n4778), .B(n4556), .Z(out[1502]) );
  ANDN U6160 ( .B(n4779), .A(n4555), .Z(n4778) );
  XNOR U6161 ( .A(n4780), .B(n4559), .Z(out[1501]) );
  ANDN U6162 ( .B(n4781), .A(n4782), .Z(n4780) );
  XOR U6163 ( .A(n4783), .B(n4564), .Z(out[1500]) );
  ANDN U6164 ( .B(n4784), .A(n4563), .Z(n4783) );
  XNOR U6165 ( .A(n4785), .B(n1871), .Z(out[14]) );
  ANDN U6166 ( .B(n1872), .A(n4055), .Z(n4785) );
  XOR U6167 ( .A(n4786), .B(n1741), .Z(n4055) );
  IV U6168 ( .A(n4054), .Z(n1872) );
  XOR U6169 ( .A(n2513), .B(n4787), .Z(n4054) );
  XOR U6170 ( .A(n4788), .B(n4032), .Z(out[149]) );
  XOR U6171 ( .A(n4789), .B(n2009), .Z(n4032) );
  ANDN U6172 ( .B(n1592), .A(n1591), .Z(n4788) );
  XOR U6173 ( .A(n4790), .B(n4791), .Z(n1591) );
  XOR U6174 ( .A(n4792), .B(n2530), .Z(n1592) );
  XOR U6175 ( .A(n4793), .B(n4567), .Z(out[1499]) );
  ANDN U6176 ( .B(n4794), .A(n4568), .Z(n4793) );
  XNOR U6177 ( .A(n4795), .B(n4571), .Z(out[1498]) );
  ANDN U6178 ( .B(n4796), .A(n4797), .Z(n4795) );
  XOR U6179 ( .A(n4798), .B(n4576), .Z(out[1497]) );
  ANDN U6180 ( .B(n4799), .A(n4575), .Z(n4798) );
  XNOR U6181 ( .A(n4800), .B(n4580), .Z(out[1496]) );
  ANDN U6182 ( .B(n4801), .A(n4579), .Z(n4800) );
  XNOR U6183 ( .A(n4802), .B(n4587), .Z(out[1495]) );
  ANDN U6184 ( .B(n4803), .A(n4588), .Z(n4802) );
  XNOR U6185 ( .A(n4804), .B(n4592), .Z(out[1494]) );
  ANDN U6186 ( .B(n4805), .A(n4591), .Z(n4804) );
  XOR U6187 ( .A(n4806), .B(n4596), .Z(out[1493]) );
  NOR U6188 ( .A(n4807), .B(n4595), .Z(n4806) );
  XOR U6189 ( .A(n4808), .B(n4600), .Z(out[1492]) );
  ANDN U6190 ( .B(n4809), .A(n4599), .Z(n4808) );
  XNOR U6191 ( .A(n4810), .B(n4603), .Z(out[1491]) );
  NOR U6192 ( .A(n4811), .B(n4604), .Z(n4810) );
  XNOR U6193 ( .A(n4812), .B(n4608), .Z(out[1490]) );
  NOR U6194 ( .A(n4813), .B(n4607), .Z(n4812) );
  XNOR U6195 ( .A(n4814), .B(n4036), .Z(out[148]) );
  IV U6196 ( .A(n4253), .Z(n4036) );
  XNOR U6197 ( .A(n4815), .B(n2012), .Z(n4253) );
  ANDN U6198 ( .B(n1615), .A(n1617), .Z(n4814) );
  XOR U6199 ( .A(n4816), .B(n3281), .Z(n1617) );
  XOR U6200 ( .A(n4817), .B(n2221), .Z(n1615) );
  XOR U6201 ( .A(n4818), .B(n4612), .Z(out[1489]) );
  ANDN U6202 ( .B(n4819), .A(n4611), .Z(n4818) );
  XNOR U6203 ( .A(n4820), .B(n4616), .Z(out[1488]) );
  NOR U6204 ( .A(n4821), .B(n4615), .Z(n4820) );
  XNOR U6205 ( .A(n4822), .B(n4622), .Z(out[1487]) );
  NOR U6206 ( .A(n4823), .B(n4621), .Z(n4822) );
  XOR U6207 ( .A(n4824), .B(n4625), .Z(out[1486]) );
  XNOR U6208 ( .A(n4826), .B(n4633), .Z(out[1485]) );
  ANDN U6209 ( .B(n4634), .A(n4827), .Z(n4826) );
  XNOR U6210 ( .A(n4828), .B(n4638), .Z(out[1484]) );
  ANDN U6211 ( .B(n4829), .A(n4637), .Z(n4828) );
  XNOR U6212 ( .A(n4830), .B(n4641), .Z(out[1483]) );
  NOR U6213 ( .A(n4831), .B(n4642), .Z(n4830) );
  XNOR U6214 ( .A(n4832), .B(n4645), .Z(out[1482]) );
  ANDN U6215 ( .B(n4833), .A(n4834), .Z(n4832) );
  XOR U6216 ( .A(n4835), .B(n4650), .Z(out[1481]) );
  ANDN U6217 ( .B(n4836), .A(n4649), .Z(n4835) );
  XNOR U6218 ( .A(n4837), .B(n4653), .Z(out[1480]) );
  NOR U6219 ( .A(n4838), .B(n4654), .Z(n4837) );
  XNOR U6220 ( .A(n4839), .B(n4039), .Z(out[147]) );
  IV U6221 ( .A(n4255), .Z(n4039) );
  XNOR U6222 ( .A(n4840), .B(n2015), .Z(n4255) );
  ANDN U6223 ( .B(n1639), .A(n1641), .Z(n4839) );
  XOR U6224 ( .A(n4841), .B(n2548), .Z(n1641) );
  XOR U6225 ( .A(n4842), .B(n2228), .Z(n1639) );
  IV U6226 ( .A(n4843), .Z(n2228) );
  XNOR U6227 ( .A(n4844), .B(n4658), .Z(out[1479]) );
  NOR U6228 ( .A(n4845), .B(n4657), .Z(n4844) );
  XNOR U6229 ( .A(n4846), .B(n4661), .Z(out[1478]) );
  NOR U6230 ( .A(n4847), .B(n4662), .Z(n4846) );
  XNOR U6231 ( .A(n4848), .B(n4665), .Z(out[1477]) );
  ANDN U6232 ( .B(n4666), .A(n4849), .Z(n4848) );
  XNOR U6233 ( .A(n4850), .B(n4670), .Z(out[1476]) );
  NOR U6234 ( .A(n4851), .B(n4669), .Z(n4850) );
  XNOR U6235 ( .A(n4852), .B(n4679), .Z(out[1475]) );
  ANDN U6236 ( .B(n4680), .A(n4853), .Z(n4852) );
  XNOR U6237 ( .A(n4854), .B(n4683), .Z(out[1474]) );
  NOR U6238 ( .A(n4855), .B(n4684), .Z(n4854) );
  XNOR U6239 ( .A(n4856), .B(n4689), .Z(out[1473]) );
  ANDN U6240 ( .B(n4857), .A(n4690), .Z(n4856) );
  XNOR U6241 ( .A(n4858), .B(n4696), .Z(out[1472]) );
  ANDN U6242 ( .B(n4859), .A(n4695), .Z(n4858) );
  IV U6243 ( .A(n4860), .Z(n4695) );
  XOR U6244 ( .A(n4861), .B(n4409), .Z(out[1471]) );
  XNOR U6245 ( .A(n4862), .B(n4863), .Z(n4409) );
  ANDN U6246 ( .B(n4864), .A(n4865), .Z(n4861) );
  XOR U6247 ( .A(n4866), .B(n4412), .Z(out[1470]) );
  XOR U6248 ( .A(n2492), .B(n4867), .Z(n4412) );
  NOR U6249 ( .A(n4868), .B(n4700), .Z(n4866) );
  XNOR U6250 ( .A(n4869), .B(n4042), .Z(out[146]) );
  XOR U6251 ( .A(n4870), .B(n2019), .Z(n4042) );
  IV U6252 ( .A(n4871), .Z(n2019) );
  ANDN U6253 ( .B(n1672), .A(n1670), .Z(n4869) );
  XOR U6254 ( .A(n4873), .B(n2553), .Z(n1672) );
  XNOR U6255 ( .A(n4874), .B(n4417), .Z(out[1469]) );
  IV U6256 ( .A(n4703), .Z(n4417) );
  XNOR U6257 ( .A(n4875), .B(n2502), .Z(n4703) );
  NOR U6258 ( .A(n4876), .B(n4702), .Z(n4874) );
  XOR U6259 ( .A(n4877), .B(n4420), .Z(out[1468]) );
  XNOR U6260 ( .A(n4878), .B(n4879), .Z(n4420) );
  ANDN U6261 ( .B(n4880), .A(n4705), .Z(n4877) );
  XOR U6262 ( .A(n4881), .B(n4424), .Z(out[1467]) );
  XOR U6263 ( .A(n2513), .B(n4882), .Z(n4424) );
  ANDN U6264 ( .B(n4883), .A(n4707), .Z(n4881) );
  XOR U6265 ( .A(n4884), .B(n4428), .Z(out[1466]) );
  XNOR U6266 ( .A(n4885), .B(n4886), .Z(n4428) );
  ANDN U6267 ( .B(n4887), .A(n4709), .Z(n4884) );
  XOR U6268 ( .A(n4888), .B(n4432), .Z(out[1465]) );
  XOR U6269 ( .A(n4889), .B(n4890), .Z(n4432) );
  ANDN U6270 ( .B(n4891), .A(n4715), .Z(n4888) );
  XOR U6271 ( .A(n4892), .B(n4436), .Z(out[1464]) );
  XOR U6272 ( .A(n3514), .B(n4893), .Z(n4436) );
  NOR U6273 ( .A(n4894), .B(n4717), .Z(n4892) );
  XNOR U6274 ( .A(n4895), .B(n4440), .Z(out[1463]) );
  XNOR U6275 ( .A(n3517), .B(n4896), .Z(n4440) );
  ANDN U6276 ( .B(n4719), .A(n4897), .Z(n4895) );
  IV U6277 ( .A(n4898), .Z(n4719) );
  XOR U6278 ( .A(n4899), .B(n4444), .Z(out[1462]) );
  XOR U6279 ( .A(n2554), .B(n4900), .Z(n4444) );
  ANDN U6280 ( .B(n4721), .A(n4901), .Z(n4899) );
  XOR U6281 ( .A(n4902), .B(n4453), .Z(out[1461]) );
  XNOR U6282 ( .A(n4903), .B(n2560), .Z(n4453) );
  ANDN U6283 ( .B(n4723), .A(n4904), .Z(n4902) );
  IV U6284 ( .A(n4905), .Z(n4723) );
  XOR U6285 ( .A(n4906), .B(n4457), .Z(out[1460]) );
  XOR U6286 ( .A(n4907), .B(n2567), .Z(n4457) );
  ANDN U6287 ( .B(n4725), .A(n4908), .Z(n4906) );
  XNOR U6288 ( .A(n4909), .B(n4045), .Z(out[145]) );
  XOR U6289 ( .A(n4910), .B(n2022), .Z(n4045) );
  ANDN U6290 ( .B(n1724), .A(n1722), .Z(n4909) );
  XOR U6291 ( .A(n4911), .B(n2248), .Z(n1722) );
  XOR U6292 ( .A(n4912), .B(n4913), .Z(n1724) );
  XOR U6293 ( .A(n4914), .B(n4461), .Z(out[1459]) );
  XOR U6294 ( .A(n4915), .B(n2574), .Z(n4461) );
  ANDN U6295 ( .B(n4916), .A(n4727), .Z(n4914) );
  XOR U6296 ( .A(n4917), .B(n4465), .Z(out[1458]) );
  XOR U6297 ( .A(n4918), .B(n2581), .Z(n4465) );
  ANDN U6298 ( .B(n4919), .A(n4729), .Z(n4917) );
  XOR U6299 ( .A(n4920), .B(n4469), .Z(out[1457]) );
  XOR U6300 ( .A(n4921), .B(n2588), .Z(n4469) );
  XOR U6301 ( .A(n4923), .B(n4473), .Z(out[1456]) );
  XOR U6302 ( .A(n4924), .B(n2597), .Z(n4473) );
  ANDN U6303 ( .B(n4733), .A(n4925), .Z(n4923) );
  IV U6304 ( .A(n4926), .Z(n4733) );
  XOR U6305 ( .A(n4927), .B(n4477), .Z(out[1455]) );
  XOR U6306 ( .A(n4928), .B(n2602), .Z(n4477) );
  ANDN U6307 ( .B(n4739), .A(n4929), .Z(n4927) );
  IV U6308 ( .A(n4930), .Z(n4739) );
  XOR U6309 ( .A(n4931), .B(n4481), .Z(out[1454]) );
  XOR U6310 ( .A(n4932), .B(n2613), .Z(n4481) );
  XNOR U6311 ( .A(n4934), .B(n4486), .Z(out[1453]) );
  XOR U6312 ( .A(n4935), .B(n2622), .Z(n4486) );
  ANDN U6313 ( .B(n4936), .A(n4743), .Z(n4934) );
  XOR U6314 ( .A(n4937), .B(n4489), .Z(out[1452]) );
  XOR U6315 ( .A(n4938), .B(n4939), .Z(n4489) );
  ANDN U6316 ( .B(n4940), .A(n4745), .Z(n4937) );
  XOR U6317 ( .A(n4941), .B(n4497), .Z(out[1451]) );
  XOR U6318 ( .A(n4942), .B(n2634), .Z(n4497) );
  NOR U6319 ( .A(n4943), .B(n4747), .Z(n4941) );
  XOR U6320 ( .A(n4944), .B(n4501), .Z(out[1450]) );
  XNOR U6321 ( .A(n4945), .B(n2641), .Z(n4501) );
  ANDN U6322 ( .B(n4946), .A(n4749), .Z(n4944) );
  XOR U6323 ( .A(n4947), .B(n4048), .Z(out[144]) );
  XOR U6324 ( .A(n4948), .B(n2025), .Z(n4048) );
  ANDN U6325 ( .B(n1772), .A(n1770), .Z(n4947) );
  XOR U6326 ( .A(n4949), .B(n2255), .Z(n1770) );
  XOR U6327 ( .A(n4950), .B(n2569), .Z(n1772) );
  XOR U6328 ( .A(n4951), .B(n4506), .Z(out[1449]) );
  XNOR U6329 ( .A(n4952), .B(n2648), .Z(n4506) );
  ANDN U6330 ( .B(n4953), .A(n4751), .Z(n4951) );
  XOR U6331 ( .A(n4954), .B(n4510), .Z(out[1448]) );
  XNOR U6332 ( .A(n4955), .B(n2655), .Z(n4510) );
  NOR U6333 ( .A(n4956), .B(n4753), .Z(n4954) );
  XOR U6334 ( .A(n4957), .B(n4513), .Z(out[1447]) );
  XOR U6335 ( .A(n4958), .B(n2662), .Z(n4513) );
  XOR U6336 ( .A(n4960), .B(n4517), .Z(out[1446]) );
  XNOR U6337 ( .A(n4961), .B(n2669), .Z(n4517) );
  ANDN U6338 ( .B(n4962), .A(n4757), .Z(n4960) );
  XOR U6339 ( .A(n4963), .B(n4765), .Z(out[1445]) );
  XNOR U6340 ( .A(n4964), .B(n2676), .Z(n4765) );
  XOR U6341 ( .A(n4966), .B(n4525), .Z(out[1444]) );
  XOR U6342 ( .A(n4967), .B(n4968), .Z(n4525) );
  XNOR U6343 ( .A(n4970), .B(n4530), .Z(out[1443]) );
  XOR U6344 ( .A(n4971), .B(n2216), .Z(n4530) );
  ANDN U6345 ( .B(n4972), .A(n4973), .Z(n4970) );
  XOR U6346 ( .A(n4974), .B(n4533), .Z(out[1442]) );
  XOR U6347 ( .A(n4975), .B(n2225), .Z(n4533) );
  XNOR U6348 ( .A(n4977), .B(n4541), .Z(out[1441]) );
  XOR U6349 ( .A(n4978), .B(n2230), .Z(n4541) );
  ANDN U6350 ( .B(n4979), .A(n4773), .Z(n4977) );
  IV U6351 ( .A(n4980), .Z(n4773) );
  XOR U6352 ( .A(n4981), .B(n4545), .Z(out[1440]) );
  XOR U6353 ( .A(n4982), .B(n2243), .Z(n4545) );
  NOR U6354 ( .A(n4983), .B(n4775), .Z(n4981) );
  XNOR U6355 ( .A(n4984), .B(n4052), .Z(out[143]) );
  XNOR U6356 ( .A(n4985), .B(n2028), .Z(n4052) );
  ANDN U6357 ( .B(n1825), .A(n1824), .Z(n4984) );
  IV U6358 ( .A(n4264), .Z(n1824) );
  XOR U6359 ( .A(n4986), .B(n2262), .Z(n4264) );
  IV U6360 ( .A(n3870), .Z(n2262) );
  XOR U6361 ( .A(n4987), .B(n4988), .Z(n1825) );
  XOR U6362 ( .A(n4989), .B(n4552), .Z(out[1439]) );
  XNOR U6363 ( .A(n4990), .B(n2250), .Z(n4552) );
  ANDN U6364 ( .B(n4991), .A(n4777), .Z(n4989) );
  XOR U6365 ( .A(n4992), .B(n4555), .Z(out[1438]) );
  XNOR U6366 ( .A(n4993), .B(n2257), .Z(n4555) );
  NOR U6367 ( .A(n4994), .B(n4779), .Z(n4992) );
  XNOR U6368 ( .A(n4995), .B(n4560), .Z(out[1437]) );
  IV U6369 ( .A(n4782), .Z(n4560) );
  XNOR U6370 ( .A(n4996), .B(n2266), .Z(n4782) );
  NOR U6371 ( .A(n4997), .B(n4781), .Z(n4995) );
  XOR U6372 ( .A(n4998), .B(n4563), .Z(out[1436]) );
  XNOR U6373 ( .A(n4999), .B(n2271), .Z(n4563) );
  NOR U6374 ( .A(n5000), .B(n4784), .Z(n4998) );
  XOR U6375 ( .A(n5001), .B(n4568), .Z(out[1435]) );
  XOR U6376 ( .A(n5002), .B(n2278), .Z(n4568) );
  ANDN U6377 ( .B(n5003), .A(n4794), .Z(n5001) );
  XNOR U6378 ( .A(n5004), .B(n4572), .Z(out[1434]) );
  IV U6379 ( .A(n4797), .Z(n4572) );
  XOR U6380 ( .A(n5005), .B(n2285), .Z(n4797) );
  ANDN U6381 ( .B(n5006), .A(n4796), .Z(n5004) );
  XOR U6382 ( .A(n5007), .B(n4575), .Z(out[1433]) );
  XNOR U6383 ( .A(n5008), .B(n2292), .Z(n4575) );
  XOR U6384 ( .A(n5010), .B(n4579), .Z(out[1432]) );
  XOR U6385 ( .A(n5011), .B(n2299), .Z(n4579) );
  NOR U6386 ( .A(n5012), .B(n4801), .Z(n5010) );
  XOR U6387 ( .A(n5013), .B(n4588), .Z(out[1431]) );
  XNOR U6388 ( .A(n5014), .B(n2306), .Z(n4588) );
  NOR U6389 ( .A(n5015), .B(n4803), .Z(n5013) );
  XOR U6390 ( .A(n5016), .B(n4591), .Z(out[1430]) );
  XNOR U6391 ( .A(n5017), .B(n2317), .Z(n4591) );
  ANDN U6392 ( .B(n5018), .A(n4805), .Z(n5016) );
  XNOR U6393 ( .A(n5019), .B(n4056), .Z(out[142]) );
  IV U6394 ( .A(n4266), .Z(n4056) );
  XNOR U6395 ( .A(n5020), .B(n2031), .Z(n4266) );
  ANDN U6396 ( .B(n1870), .A(n1871), .Z(n5019) );
  XNOR U6397 ( .A(n5021), .B(n2583), .Z(n1871) );
  XOR U6398 ( .A(n5022), .B(n2269), .Z(n1870) );
  IV U6399 ( .A(n5023), .Z(n2269) );
  XOR U6400 ( .A(n5024), .B(n4595), .Z(out[1429]) );
  XNOR U6401 ( .A(n2325), .B(n5025), .Z(n4595) );
  XOR U6402 ( .A(n5027), .B(n4599), .Z(out[1428]) );
  XOR U6403 ( .A(n2332), .B(n5028), .Z(n4599) );
  ANDN U6404 ( .B(n5029), .A(n4809), .Z(n5027) );
  XOR U6405 ( .A(n5030), .B(n4604), .Z(out[1427]) );
  XOR U6406 ( .A(n2339), .B(n5031), .Z(n4604) );
  ANDN U6407 ( .B(n4811), .A(n5032), .Z(n5030) );
  XOR U6408 ( .A(n5033), .B(n4607), .Z(out[1426]) );
  XOR U6409 ( .A(n2346), .B(n5034), .Z(n4607) );
  XOR U6410 ( .A(n5036), .B(n4611), .Z(out[1425]) );
  XOR U6411 ( .A(n2353), .B(n5037), .Z(n4611) );
  ANDN U6412 ( .B(n5038), .A(n4819), .Z(n5036) );
  XOR U6413 ( .A(n5039), .B(n4615), .Z(out[1424]) );
  XNOR U6414 ( .A(n2360), .B(n5040), .Z(n4615) );
  ANDN U6415 ( .B(n5041), .A(n5042), .Z(n5039) );
  XOR U6416 ( .A(n5043), .B(n4621), .Z(out[1423]) );
  XOR U6417 ( .A(n2367), .B(n5044), .Z(n4621) );
  ANDN U6418 ( .B(n5045), .A(n5046), .Z(n5043) );
  XNOR U6419 ( .A(n5047), .B(n4626), .Z(out[1422]) );
  XOR U6420 ( .A(n3444), .B(n5048), .Z(n4626) );
  ANDN U6421 ( .B(n5049), .A(n4825), .Z(n5047) );
  XNOR U6422 ( .A(n5050), .B(n4634), .Z(out[1421]) );
  XOR U6423 ( .A(n2381), .B(n5051), .Z(n4634) );
  XOR U6424 ( .A(n5053), .B(n4637), .Z(out[1420]) );
  XNOR U6425 ( .A(n2392), .B(n5054), .Z(n4637) );
  ANDN U6426 ( .B(n5055), .A(n4829), .Z(n5053) );
  XOR U6427 ( .A(n5056), .B(n4060), .Z(out[141]) );
  XOR U6428 ( .A(n5057), .B(n2034), .Z(n4060) );
  ANDN U6429 ( .B(n1915), .A(n1917), .Z(n5056) );
  XNOR U6430 ( .A(n5058), .B(n3881), .Z(n1915) );
  XOR U6431 ( .A(n5059), .B(n4642), .Z(out[1419]) );
  XOR U6432 ( .A(n5060), .B(n2398), .Z(n4642) );
  ANDN U6433 ( .B(n5061), .A(n5062), .Z(n5059) );
  XNOR U6434 ( .A(n5063), .B(n4646), .Z(out[1418]) );
  IV U6435 ( .A(n4834), .Z(n4646) );
  XNOR U6436 ( .A(n5064), .B(n2405), .Z(n4834) );
  ANDN U6437 ( .B(n5065), .A(n4833), .Z(n5063) );
  XOR U6438 ( .A(n5066), .B(n4649), .Z(out[1417]) );
  XOR U6439 ( .A(n2413), .B(n5067), .Z(n4649) );
  ANDN U6440 ( .B(n5068), .A(n4836), .Z(n5066) );
  XOR U6441 ( .A(n5069), .B(n4654), .Z(out[1416]) );
  XOR U6442 ( .A(n5070), .B(n5071), .Z(n4654) );
  ANDN U6443 ( .B(n5072), .A(n5073), .Z(n5069) );
  XOR U6444 ( .A(n5074), .B(n4657), .Z(out[1415]) );
  XNOR U6445 ( .A(n2427), .B(n5075), .Z(n4657) );
  XOR U6446 ( .A(n5077), .B(n4662), .Z(out[1414]) );
  XNOR U6447 ( .A(n2434), .B(n5078), .Z(n4662) );
  ANDN U6448 ( .B(n4847), .A(n5079), .Z(n5077) );
  XNOR U6449 ( .A(n5080), .B(n4666), .Z(out[1413]) );
  XOR U6450 ( .A(n4128), .B(n5081), .Z(n4666) );
  IV U6451 ( .A(n2441), .Z(n4128) );
  XOR U6452 ( .A(n5083), .B(n4669), .Z(out[1412]) );
  XNOR U6453 ( .A(n3477), .B(n5084), .Z(n4669) );
  ANDN U6454 ( .B(n4851), .A(n5085), .Z(n5083) );
  XNOR U6455 ( .A(n5086), .B(n4680), .Z(out[1411]) );
  XOR U6456 ( .A(n4199), .B(n5087), .Z(n4680) );
  XOR U6457 ( .A(n5089), .B(n4684), .Z(out[1410]) );
  XNOR U6458 ( .A(n5090), .B(n5091), .Z(n4684) );
  ANDN U6459 ( .B(n4855), .A(n5092), .Z(n5089) );
  XNOR U6460 ( .A(n5093), .B(n4064), .Z(out[140]) );
  IV U6461 ( .A(n4269), .Z(n4064) );
  XNOR U6462 ( .A(n5094), .B(n2041), .Z(n4269) );
  AND U6463 ( .A(n1966), .B(n1964), .Z(n5093) );
  XOR U6464 ( .A(n5095), .B(n5096), .Z(n1964) );
  XOR U6465 ( .A(n5097), .B(n4690), .Z(out[1409]) );
  XNOR U6466 ( .A(n2473), .B(n5098), .Z(n4690) );
  ANDN U6467 ( .B(n5099), .A(n4857), .Z(n5097) );
  XNOR U6468 ( .A(n5100), .B(n4860), .Z(out[1408]) );
  XOR U6469 ( .A(n2480), .B(n5101), .Z(n4860) );
  ANDN U6470 ( .B(n5102), .A(n4859), .Z(n5100) );
  XNOR U6471 ( .A(n5103), .B(n4698), .Z(out[1407]) );
  IV U6472 ( .A(n4865), .Z(n4698) );
  XNOR U6473 ( .A(n1955), .B(n5104), .Z(n4865) );
  ANDN U6474 ( .B(n4404), .A(n4864), .Z(n5103) );
  XOR U6475 ( .A(n5105), .B(n4700), .Z(out[1406]) );
  XNOR U6476 ( .A(n5106), .B(n4215), .Z(n4700) );
  NOR U6477 ( .A(n5107), .B(n4411), .Z(n5105) );
  XOR U6478 ( .A(n5108), .B(n4702), .Z(out[1405]) );
  XNOR U6479 ( .A(n5109), .B(n1969), .Z(n4702) );
  ANDN U6480 ( .B(n4876), .A(n4415), .Z(n5108) );
  XOR U6481 ( .A(n5110), .B(n4705), .Z(out[1404]) );
  XOR U6482 ( .A(n5111), .B(n4222), .Z(n4705) );
  ANDN U6483 ( .B(n4419), .A(n4880), .Z(n5110) );
  XOR U6484 ( .A(n5112), .B(n4707), .Z(out[1403]) );
  XOR U6485 ( .A(n5113), .B(n1662), .Z(n4707) );
  NOR U6486 ( .A(n4883), .B(n4423), .Z(n5112) );
  XOR U6487 ( .A(n5114), .B(n4709), .Z(out[1402]) );
  XNOR U6488 ( .A(n5115), .B(n1667), .Z(n4709) );
  NOR U6489 ( .A(n4887), .B(n4427), .Z(n5114) );
  XOR U6490 ( .A(n5116), .B(n4715), .Z(out[1401]) );
  XOR U6491 ( .A(n5117), .B(n1675), .Z(n4715) );
  NOR U6492 ( .A(n4891), .B(n4431), .Z(n5116) );
  XOR U6493 ( .A(n5118), .B(n4717), .Z(out[1400]) );
  XNOR U6494 ( .A(n5119), .B(n1680), .Z(n4717) );
  XNOR U6495 ( .A(n5120), .B(n1917), .Z(out[13]) );
  XOR U6496 ( .A(n5121), .B(n3312), .Z(n1917) );
  NOR U6497 ( .A(n4061), .B(n1916), .Z(n5120) );
  XNOR U6498 ( .A(n2520), .B(n5122), .Z(n1916) );
  XOR U6499 ( .A(n5123), .B(n1745), .Z(n4061) );
  XNOR U6500 ( .A(n5124), .B(n4067), .Z(out[139]) );
  IV U6501 ( .A(n4271), .Z(n4067) );
  XNOR U6502 ( .A(n5125), .B(n2045), .Z(n4271) );
  XNOR U6503 ( .A(n5126), .B(n5127), .Z(n2000) );
  XOR U6504 ( .A(n5128), .B(n4898), .Z(out[1399]) );
  XNOR U6505 ( .A(n5129), .B(n1685), .Z(n4898) );
  ANDN U6506 ( .B(n4439), .A(n5130), .Z(n5128) );
  XNOR U6507 ( .A(n5131), .B(n4721), .Z(out[1398]) );
  XNOR U6508 ( .A(n5132), .B(n1689), .Z(n4721) );
  ANDN U6509 ( .B(n4443), .A(n5133), .Z(n5131) );
  XOR U6510 ( .A(n5134), .B(n4905), .Z(out[1397]) );
  XNOR U6511 ( .A(n5135), .B(n1693), .Z(n4905) );
  IV U6512 ( .A(n5136), .Z(n4904) );
  XNOR U6513 ( .A(n5137), .B(n4725), .Z(out[1396]) );
  XOR U6514 ( .A(n5138), .B(n1698), .Z(n4725) );
  ANDN U6515 ( .B(n4456), .A(n5139), .Z(n5137) );
  XOR U6516 ( .A(n5140), .B(n4727), .Z(out[1395]) );
  XOR U6517 ( .A(n5141), .B(n1703), .Z(n4727) );
  ANDN U6518 ( .B(n4460), .A(n4916), .Z(n5140) );
  XOR U6519 ( .A(n5142), .B(n4729), .Z(out[1394]) );
  XOR U6520 ( .A(n5143), .B(n1708), .Z(n4729) );
  ANDN U6521 ( .B(n4464), .A(n4919), .Z(n5142) );
  XNOR U6522 ( .A(n5144), .B(n4731), .Z(out[1393]) );
  XOR U6523 ( .A(n5145), .B(n3818), .Z(n4731) );
  NOR U6524 ( .A(n4922), .B(n4468), .Z(n5144) );
  XOR U6525 ( .A(n5146), .B(n4926), .Z(out[1392]) );
  XNOR U6526 ( .A(n5147), .B(n1718), .Z(n4926) );
  XOR U6527 ( .A(n5148), .B(n4930), .Z(out[1391]) );
  XNOR U6528 ( .A(n5149), .B(n1727), .Z(n4930) );
  XOR U6529 ( .A(n5150), .B(n4741), .Z(out[1390]) );
  XNOR U6530 ( .A(n5151), .B(n1732), .Z(n4741) );
  NOR U6531 ( .A(n4933), .B(n4480), .Z(n5150) );
  XNOR U6532 ( .A(n5152), .B(n4070), .Z(out[138]) );
  IV U6533 ( .A(n4273), .Z(n4070) );
  XOR U6534 ( .A(n5153), .B(n2049), .Z(n4273) );
  ANDN U6535 ( .B(n2038), .A(n2036), .Z(n5152) );
  XOR U6536 ( .A(n5154), .B(n2297), .Z(n2036) );
  XOR U6537 ( .A(n5155), .B(n4743), .Z(out[1389]) );
  XOR U6538 ( .A(n5156), .B(n1736), .Z(n4743) );
  NOR U6539 ( .A(n4936), .B(n4484), .Z(n5155) );
  XOR U6540 ( .A(n5157), .B(n4745), .Z(out[1388]) );
  XNOR U6541 ( .A(n5158), .B(n1741), .Z(n4745) );
  ANDN U6542 ( .B(n4488), .A(n4940), .Z(n5157) );
  XOR U6543 ( .A(n5159), .B(n4747), .Z(out[1387]) );
  XNOR U6544 ( .A(n5160), .B(n1745), .Z(n4747) );
  ANDN U6545 ( .B(n4496), .A(n5161), .Z(n5159) );
  XOR U6546 ( .A(n5162), .B(n4749), .Z(out[1386]) );
  XOR U6547 ( .A(n5163), .B(n1749), .Z(n4749) );
  ANDN U6548 ( .B(n4500), .A(n4946), .Z(n5162) );
  XOR U6549 ( .A(n5164), .B(n4751), .Z(out[1385]) );
  XNOR U6550 ( .A(n5165), .B(n1754), .Z(n4751) );
  ANDN U6551 ( .B(n4504), .A(n4953), .Z(n5164) );
  XOR U6552 ( .A(n5166), .B(n4753), .Z(out[1384]) );
  XNOR U6553 ( .A(n5167), .B(n3862), .Z(n4753) );
  NOR U6554 ( .A(n5168), .B(n4508), .Z(n5166) );
  XOR U6555 ( .A(n5169), .B(n4755), .Z(out[1383]) );
  XNOR U6556 ( .A(n3866), .B(n5170), .Z(n4755) );
  IV U6557 ( .A(n1762), .Z(n3866) );
  NOR U6558 ( .A(n4959), .B(n4512), .Z(n5169) );
  XOR U6559 ( .A(n5171), .B(n4757), .Z(out[1382]) );
  XOR U6560 ( .A(n5172), .B(n1767), .Z(n4757) );
  IV U6561 ( .A(n5173), .Z(n1767) );
  ANDN U6562 ( .B(n4516), .A(n4962), .Z(n5171) );
  XNOR U6563 ( .A(n5174), .B(n4764), .Z(out[1381]) );
  XOR U6564 ( .A(n5175), .B(n1775), .Z(n4764) );
  IV U6565 ( .A(n5176), .Z(n1775) );
  ANDN U6566 ( .B(n4520), .A(n4965), .Z(n5174) );
  XOR U6567 ( .A(n5177), .B(n4767), .Z(out[1380]) );
  XOR U6568 ( .A(n5178), .B(n1780), .Z(n4767) );
  IV U6569 ( .A(n5179), .Z(n1780) );
  NOR U6570 ( .A(n4969), .B(n4524), .Z(n5177) );
  XOR U6571 ( .A(n5180), .B(n4073), .Z(out[137]) );
  XNOR U6572 ( .A(n5181), .B(n2053), .Z(n4073) );
  IV U6573 ( .A(n5182), .Z(n2053) );
  ANDN U6574 ( .B(n2075), .A(n1031), .Z(n5180) );
  XOR U6575 ( .A(n5183), .B(n2619), .Z(n1031) );
  XOR U6576 ( .A(n5184), .B(n2304), .Z(n2075) );
  XNOR U6577 ( .A(n5185), .B(n4769), .Z(out[1379]) );
  IV U6578 ( .A(n4973), .Z(n4769) );
  XOR U6579 ( .A(n5186), .B(n1785), .Z(n4973) );
  IV U6580 ( .A(n5187), .Z(n1785) );
  NOR U6581 ( .A(n4972), .B(n4528), .Z(n5185) );
  XOR U6582 ( .A(n5188), .B(n4771), .Z(out[1378]) );
  XOR U6583 ( .A(n5189), .B(n4293), .Z(n4771) );
  NOR U6584 ( .A(n4976), .B(n4532), .Z(n5188) );
  XNOR U6585 ( .A(n5190), .B(n4980), .Z(out[1377]) );
  XOR U6586 ( .A(n5191), .B(n1794), .Z(n4980) );
  IV U6587 ( .A(n5192), .Z(n1794) );
  ANDN U6588 ( .B(n4540), .A(n4979), .Z(n5190) );
  IV U6589 ( .A(n5193), .Z(n4979) );
  XOR U6590 ( .A(n5194), .B(n4775), .Z(out[1376]) );
  XNOR U6591 ( .A(n5195), .B(n5196), .Z(n4775) );
  NOR U6592 ( .A(n5197), .B(n4544), .Z(n5194) );
  XOR U6593 ( .A(n5198), .B(n4777), .Z(out[1375]) );
  XNOR U6594 ( .A(n5199), .B(n1804), .Z(n4777) );
  ANDN U6595 ( .B(n4547), .A(n4991), .Z(n5198) );
  XOR U6596 ( .A(n5200), .B(n4779), .Z(out[1374]) );
  XNOR U6597 ( .A(n5201), .B(n5202), .Z(n4779) );
  XOR U6598 ( .A(n5203), .B(n4781), .Z(out[1373]) );
  XOR U6599 ( .A(n4107), .B(n5204), .Z(n4781) );
  XOR U6600 ( .A(n5205), .B(n4784), .Z(out[1372]) );
  XNOR U6601 ( .A(n5206), .B(n5207), .Z(n4784) );
  XOR U6602 ( .A(n5208), .B(n4794), .Z(out[1371]) );
  XOR U6603 ( .A(n5209), .B(n5210), .Z(n4794) );
  NOR U6604 ( .A(n4566), .B(n5003), .Z(n5208) );
  XOR U6605 ( .A(n5211), .B(n4796), .Z(out[1370]) );
  XOR U6606 ( .A(n4117), .B(n5212), .Z(n4796) );
  NOR U6607 ( .A(n4570), .B(n5006), .Z(n5211) );
  XOR U6608 ( .A(n5213), .B(n4076), .Z(out[136]) );
  XNOR U6609 ( .A(n5214), .B(n5215), .Z(n4076) );
  ANDN U6610 ( .B(n1475), .A(n2111), .Z(n5213) );
  XOR U6611 ( .A(n5216), .B(n2315), .Z(n2111) );
  XOR U6612 ( .A(n5217), .B(n3330), .Z(n1475) );
  IV U6613 ( .A(n2629), .Z(n3330) );
  XOR U6614 ( .A(n5218), .B(n4799), .Z(out[1369]) );
  XNOR U6615 ( .A(n1837), .B(n5219), .Z(n4799) );
  NOR U6616 ( .A(n5009), .B(n4574), .Z(n5218) );
  XOR U6617 ( .A(n5220), .B(n4801), .Z(out[1368]) );
  XNOR U6618 ( .A(n3626), .B(n5221), .Z(n4801) );
  ANDN U6619 ( .B(n5012), .A(n4578), .Z(n5220) );
  XOR U6620 ( .A(n5222), .B(n4803), .Z(out[1367]) );
  XOR U6621 ( .A(n5223), .B(n5224), .Z(n4803) );
  NOR U6622 ( .A(n5225), .B(n4586), .Z(n5222) );
  XOR U6623 ( .A(n5226), .B(n4805), .Z(out[1366]) );
  XOR U6624 ( .A(n5227), .B(n5228), .Z(n4805) );
  ANDN U6625 ( .B(n4590), .A(n5018), .Z(n5226) );
  XNOR U6626 ( .A(n5229), .B(n4807), .Z(out[1365]) );
  XOR U6627 ( .A(n3641), .B(n5230), .Z(n4807) );
  NOR U6628 ( .A(n4594), .B(n5026), .Z(n5229) );
  XOR U6629 ( .A(n5231), .B(n4809), .Z(out[1364]) );
  XOR U6630 ( .A(n5232), .B(n5233), .Z(n4809) );
  NOR U6631 ( .A(n4598), .B(n5029), .Z(n5231) );
  IV U6632 ( .A(n5234), .Z(n4598) );
  XNOR U6633 ( .A(n5235), .B(n4811), .Z(out[1363]) );
  XNOR U6634 ( .A(n1862), .B(n5236), .Z(n4811) );
  NOR U6635 ( .A(n5237), .B(n4602), .Z(n5235) );
  XNOR U6636 ( .A(n5238), .B(n4813), .Z(out[1362]) );
  XNOR U6637 ( .A(n5239), .B(n5240), .Z(n4813) );
  NOR U6638 ( .A(n5035), .B(n4606), .Z(n5238) );
  XOR U6639 ( .A(n5241), .B(n4819), .Z(out[1361]) );
  XOR U6640 ( .A(n5242), .B(n5243), .Z(n4819) );
  ANDN U6641 ( .B(n4610), .A(n5038), .Z(n5241) );
  XNOR U6642 ( .A(n5244), .B(n4821), .Z(out[1360]) );
  IV U6643 ( .A(n5042), .Z(n4821) );
  XOR U6644 ( .A(n5245), .B(n5246), .Z(n5042) );
  NOR U6645 ( .A(n4614), .B(n5041), .Z(n5244) );
  XOR U6646 ( .A(n5247), .B(n4079), .Z(out[135]) );
  XOR U6647 ( .A(n5248), .B(n2059), .Z(n4079) );
  ANDN U6648 ( .B(n2149), .A(n1820), .Z(n5247) );
  XOR U6649 ( .A(n5249), .B(n3334), .Z(n1820) );
  XOR U6650 ( .A(n5250), .B(n3908), .Z(n2149) );
  XNOR U6651 ( .A(n5251), .B(n4823), .Z(out[1359]) );
  IV U6652 ( .A(n5046), .Z(n4823) );
  XOR U6653 ( .A(n5252), .B(n5253), .Z(n5046) );
  NOR U6654 ( .A(n5254), .B(n5045), .Z(n5251) );
  XOR U6655 ( .A(n5255), .B(n4825), .Z(out[1358]) );
  XOR U6656 ( .A(n1886), .B(n5256), .Z(n4825) );
  NOR U6657 ( .A(n5049), .B(n4624), .Z(n5255) );
  XNOR U6658 ( .A(n5257), .B(n4827), .Z(out[1357]) );
  XOR U6659 ( .A(n5258), .B(n5259), .Z(n4827) );
  NOR U6660 ( .A(n5052), .B(n4632), .Z(n5257) );
  IV U6661 ( .A(n5260), .Z(n5052) );
  XOR U6662 ( .A(n5261), .B(n4829), .Z(out[1356]) );
  XOR U6663 ( .A(n5262), .B(n5263), .Z(n4829) );
  NOR U6664 ( .A(n5055), .B(n4636), .Z(n5261) );
  XNOR U6665 ( .A(n5264), .B(n4831), .Z(out[1355]) );
  IV U6666 ( .A(n5062), .Z(n4831) );
  XOR U6667 ( .A(n5265), .B(n5266), .Z(n5062) );
  NOR U6668 ( .A(n4640), .B(n5061), .Z(n5264) );
  XOR U6669 ( .A(n5267), .B(n4833), .Z(out[1354]) );
  XNOR U6670 ( .A(n3695), .B(n5268), .Z(n4833) );
  NOR U6671 ( .A(n5065), .B(n4644), .Z(n5267) );
  XOR U6672 ( .A(n5269), .B(n4836), .Z(out[1353]) );
  XOR U6673 ( .A(n4176), .B(n5270), .Z(n4836) );
  NOR U6674 ( .A(n5068), .B(n4648), .Z(n5269) );
  XNOR U6675 ( .A(n5271), .B(n4838), .Z(out[1352]) );
  IV U6676 ( .A(n5073), .Z(n4838) );
  XOR U6677 ( .A(n4181), .B(n5272), .Z(n5073) );
  ANDN U6678 ( .B(n4652), .A(n5072), .Z(n5271) );
  XNOR U6679 ( .A(n5273), .B(n4845), .Z(out[1351]) );
  XOR U6680 ( .A(n1919), .B(n5274), .Z(n4845) );
  NOR U6681 ( .A(n5076), .B(n4656), .Z(n5273) );
  XNOR U6682 ( .A(n5275), .B(n4847), .Z(out[1350]) );
  XOR U6683 ( .A(n1923), .B(n5276), .Z(n4847) );
  XOR U6684 ( .A(n5277), .B(n4083), .Z(out[134]) );
  XOR U6685 ( .A(n5278), .B(n2063), .Z(n4083) );
  IV U6686 ( .A(n5279), .Z(n2063) );
  ANDN U6687 ( .B(n2183), .A(n2185), .Z(n5277) );
  XOR U6688 ( .A(n5280), .B(n2643), .Z(n2185) );
  IV U6689 ( .A(n3338), .Z(n2643) );
  XOR U6690 ( .A(n5281), .B(n2329), .Z(n2183) );
  XNOR U6691 ( .A(n5282), .B(n4849), .Z(out[1349]) );
  XOR U6692 ( .A(n3719), .B(n5283), .Z(n4849) );
  NOR U6693 ( .A(n5082), .B(n4664), .Z(n5282) );
  XNOR U6694 ( .A(n5284), .B(n4851), .Z(out[1348]) );
  XOR U6695 ( .A(n3726), .B(n5285), .Z(n4851) );
  XNOR U6696 ( .A(n5286), .B(n4853), .Z(out[1347]) );
  XOR U6697 ( .A(n3733), .B(n5287), .Z(n4853) );
  NOR U6698 ( .A(n5088), .B(n4675), .Z(n5286) );
  XNOR U6699 ( .A(n5288), .B(n4855), .Z(out[1346]) );
  XNOR U6700 ( .A(n1941), .B(n5289), .Z(n4855) );
  ANDN U6701 ( .B(n4682), .A(n5290), .Z(n5288) );
  XOR U6702 ( .A(n5291), .B(n4857), .Z(out[1345]) );
  XNOR U6703 ( .A(n1946), .B(n5292), .Z(n4857) );
  ANDN U6704 ( .B(n4685), .A(n5099), .Z(n5291) );
  XOR U6705 ( .A(n5293), .B(n4859), .Z(out[1344]) );
  XNOR U6706 ( .A(n1951), .B(n5294), .Z(n4859) );
  ANDN U6707 ( .B(n4691), .A(n5102), .Z(n5293) );
  XOR U6708 ( .A(n5295), .B(n4864), .Z(out[1343]) );
  XOR U6709 ( .A(n5296), .B(n1995), .Z(n4864) );
  NOR U6710 ( .A(n4408), .B(n4404), .Z(n5295) );
  XOR U6711 ( .A(n5297), .B(n2551), .Z(n4404) );
  XNOR U6712 ( .A(n5298), .B(n2530), .Z(n4408) );
  XNOR U6713 ( .A(n5299), .B(n4868), .Z(out[1342]) );
  IV U6714 ( .A(n5107), .Z(n4868) );
  XNOR U6715 ( .A(n5300), .B(n1998), .Z(n5107) );
  ANDN U6716 ( .B(n4411), .A(n4413), .Z(n5299) );
  XOR U6717 ( .A(n5301), .B(n3281), .Z(n4413) );
  IV U6718 ( .A(n2539), .Z(n3281) );
  XOR U6719 ( .A(n5302), .B(n2558), .Z(n4411) );
  XNOR U6720 ( .A(n5303), .B(n4876), .Z(out[1341]) );
  XNOR U6721 ( .A(n5304), .B(n2005), .Z(n4876) );
  ANDN U6722 ( .B(n4415), .A(n4416), .Z(n5303) );
  XOR U6723 ( .A(n5305), .B(n2548), .Z(n4416) );
  XNOR U6724 ( .A(n5306), .B(n2565), .Z(n4415) );
  XOR U6725 ( .A(n5307), .B(n4880), .Z(out[1340]) );
  XOR U6726 ( .A(n5308), .B(n2009), .Z(n4880) );
  NOR U6727 ( .A(n4421), .B(n4419), .Z(n5307) );
  XOR U6728 ( .A(n5309), .B(n3762), .Z(n4419) );
  XOR U6729 ( .A(n5310), .B(n2553), .Z(n4421) );
  XOR U6730 ( .A(n5311), .B(n4290), .Z(out[133]) );
  XOR U6731 ( .A(n5312), .B(n2066), .Z(n4290) );
  ANDN U6732 ( .B(n2238), .A(n2236), .Z(n5311) );
  XOR U6733 ( .A(n5313), .B(n2336), .Z(n2236) );
  XOR U6734 ( .A(n5314), .B(n2650), .Z(n2238) );
  IV U6735 ( .A(n5315), .Z(n2650) );
  XOR U6736 ( .A(n5316), .B(n4883), .Z(out[1339]) );
  XOR U6737 ( .A(n5317), .B(n2012), .Z(n4883) );
  ANDN U6738 ( .B(n4423), .A(n4425), .Z(n5316) );
  XNOR U6739 ( .A(n5318), .B(n2562), .Z(n4425) );
  XOR U6740 ( .A(n5319), .B(n2579), .Z(n4423) );
  XOR U6741 ( .A(n5320), .B(n4887), .Z(out[1338]) );
  XOR U6742 ( .A(n5321), .B(n2015), .Z(n4887) );
  ANDN U6743 ( .B(n4427), .A(n4429), .Z(n5320) );
  XNOR U6744 ( .A(n5322), .B(n3296), .Z(n4429) );
  IV U6745 ( .A(n2569), .Z(n3296) );
  XNOR U6746 ( .A(n2585), .B(n5323), .Z(n4427) );
  IV U6747 ( .A(n5324), .Z(n2585) );
  XOR U6748 ( .A(n5325), .B(n4891), .Z(out[1337]) );
  XOR U6749 ( .A(n5326), .B(n4871), .Z(n4891) );
  ANDN U6750 ( .B(n4431), .A(n4433), .Z(n5325) );
  XOR U6751 ( .A(n5327), .B(n2576), .Z(n4433) );
  IV U6752 ( .A(n4988), .Z(n2576) );
  XOR U6753 ( .A(n2592), .B(n5328), .Z(n4431) );
  IV U6754 ( .A(n4387), .Z(n2592) );
  XNOR U6755 ( .A(n5329), .B(n4894), .Z(out[1336]) );
  XOR U6756 ( .A(n5330), .B(n2022), .Z(n4894) );
  IV U6757 ( .A(n5331), .Z(n2022) );
  ANDN U6758 ( .B(n4437), .A(n4435), .Z(n5329) );
  XOR U6759 ( .A(n2599), .B(n5332), .Z(n4435) );
  IV U6760 ( .A(n5333), .Z(n2599) );
  XOR U6761 ( .A(n5334), .B(n2583), .Z(n4437) );
  IV U6762 ( .A(n5335), .Z(n2583) );
  XNOR U6763 ( .A(n5336), .B(n4897), .Z(out[1335]) );
  IV U6764 ( .A(n5130), .Z(n4897) );
  XNOR U6765 ( .A(n5337), .B(n2025), .Z(n5130) );
  ANDN U6766 ( .B(n4441), .A(n4439), .Z(n5336) );
  XNOR U6767 ( .A(n5338), .B(n2611), .Z(n4439) );
  XOR U6768 ( .A(n5339), .B(n3312), .Z(n4441) );
  IV U6769 ( .A(n2590), .Z(n3312) );
  XNOR U6770 ( .A(n5340), .B(n4901), .Z(out[1334]) );
  IV U6771 ( .A(n5133), .Z(n4901) );
  XNOR U6772 ( .A(n5341), .B(n2028), .Z(n5133) );
  NOR U6773 ( .A(n4445), .B(n4443), .Z(n5340) );
  XOR U6774 ( .A(n5342), .B(n3789), .Z(n4443) );
  XOR U6775 ( .A(n5343), .B(n2595), .Z(n4445) );
  XOR U6776 ( .A(n5344), .B(n5136), .Z(out[1333]) );
  XOR U6777 ( .A(n5345), .B(n2031), .Z(n5136) );
  ANDN U6778 ( .B(n4454), .A(n4452), .Z(n5344) );
  XOR U6779 ( .A(n5346), .B(n2625), .Z(n4452) );
  XOR U6780 ( .A(n5347), .B(n5348), .Z(n4454) );
  XNOR U6781 ( .A(n5349), .B(n4908), .Z(out[1332]) );
  IV U6782 ( .A(n5139), .Z(n4908) );
  XNOR U6783 ( .A(n5350), .B(n2034), .Z(n5139) );
  ANDN U6784 ( .B(n4458), .A(n4456), .Z(n5349) );
  XOR U6785 ( .A(n5351), .B(n3801), .Z(n4456) );
  IV U6786 ( .A(n2632), .Z(n3801) );
  XOR U6787 ( .A(n5352), .B(n2615), .Z(n4458) );
  XOR U6788 ( .A(n5353), .B(n4916), .Z(out[1331]) );
  XNOR U6789 ( .A(n5354), .B(n2041), .Z(n4916) );
  NOR U6790 ( .A(n4462), .B(n4460), .Z(n5353) );
  XOR U6791 ( .A(n5355), .B(n2639), .Z(n4460) );
  XOR U6792 ( .A(n2619), .B(n5356), .Z(n4462) );
  IV U6793 ( .A(n5357), .Z(n2619) );
  XOR U6794 ( .A(n5358), .B(n4919), .Z(out[1330]) );
  XOR U6795 ( .A(n5359), .B(n2045), .Z(n4919) );
  ANDN U6796 ( .B(n4466), .A(n4464), .Z(n5358) );
  XOR U6797 ( .A(n5360), .B(n3811), .Z(n4464) );
  XOR U6798 ( .A(n5361), .B(n2629), .Z(n4466) );
  XOR U6799 ( .A(n5362), .B(n4090), .Z(out[132]) );
  XNOR U6800 ( .A(n5363), .B(n2069), .Z(n4090) );
  ANDN U6801 ( .B(n2310), .A(n2312), .Z(n5362) );
  XOR U6802 ( .A(n5364), .B(n2657), .Z(n2312) );
  XNOR U6803 ( .A(n5365), .B(n2343), .Z(n2310) );
  XOR U6804 ( .A(n5366), .B(n4922), .Z(out[1329]) );
  XNOR U6805 ( .A(n5367), .B(n2049), .Z(n4922) );
  ANDN U6806 ( .B(n4468), .A(n4470), .Z(n5366) );
  XNOR U6807 ( .A(n5368), .B(n3334), .Z(n4470) );
  IV U6808 ( .A(n2636), .Z(n3334) );
  XNOR U6809 ( .A(n5369), .B(n2653), .Z(n4468) );
  XNOR U6810 ( .A(n5370), .B(n4925), .Z(out[1328]) );
  XOR U6811 ( .A(n5371), .B(n5182), .Z(n4925) );
  ANDN U6812 ( .B(n4474), .A(n4472), .Z(n5370) );
  XNOR U6813 ( .A(n5372), .B(n3822), .Z(n4472) );
  XOR U6814 ( .A(n5373), .B(n3338), .Z(n4474) );
  XNOR U6815 ( .A(n5374), .B(n4929), .Z(out[1327]) );
  XOR U6816 ( .A(n5375), .B(n2056), .Z(n4929) );
  ANDN U6817 ( .B(n4478), .A(n4476), .Z(n5374) );
  XOR U6818 ( .A(n5376), .B(n2667), .Z(n4476) );
  XOR U6819 ( .A(n5377), .B(n5315), .Z(n4478) );
  XOR U6820 ( .A(n5378), .B(n4933), .Z(out[1326]) );
  XOR U6821 ( .A(n5379), .B(n2059), .Z(n4933) );
  IV U6822 ( .A(n5380), .Z(n2059) );
  ANDN U6823 ( .B(n4480), .A(n4482), .Z(n5378) );
  XOR U6824 ( .A(n5381), .B(n2657), .Z(n4482) );
  IV U6825 ( .A(n5382), .Z(n2657) );
  XOR U6826 ( .A(n5383), .B(n2674), .Z(n4480) );
  XOR U6827 ( .A(n5384), .B(n4936), .Z(out[1325]) );
  XNOR U6828 ( .A(n5385), .B(n5279), .Z(n4936) );
  ANDN U6829 ( .B(n4484), .A(n4485), .Z(n5384) );
  XNOR U6830 ( .A(n5386), .B(n2664), .Z(n4485) );
  XOR U6831 ( .A(n5387), .B(n2207), .Z(n4484) );
  XOR U6832 ( .A(n5388), .B(n4940), .Z(out[1324]) );
  XOR U6833 ( .A(n5389), .B(n2066), .Z(n4940) );
  IV U6834 ( .A(n5390), .Z(n2066) );
  NOR U6835 ( .A(n4490), .B(n4488), .Z(n5388) );
  XOR U6836 ( .A(n5391), .B(n4791), .Z(n4488) );
  IV U6837 ( .A(n2214), .Z(n4791) );
  XOR U6838 ( .A(n5392), .B(n3356), .Z(n4490) );
  XNOR U6839 ( .A(n5393), .B(n4943), .Z(out[1323]) );
  IV U6840 ( .A(n5161), .Z(n4943) );
  XOR U6841 ( .A(n5394), .B(n2069), .Z(n5161) );
  NOR U6842 ( .A(n4498), .B(n4496), .Z(n5393) );
  XOR U6843 ( .A(n5395), .B(n2221), .Z(n4496) );
  XOR U6844 ( .A(n5396), .B(n2678), .Z(n4498) );
  XOR U6845 ( .A(n5397), .B(n4946), .Z(out[1322]) );
  XNOR U6846 ( .A(n5398), .B(n2072), .Z(n4946) );
  NOR U6847 ( .A(n4502), .B(n4500), .Z(n5397) );
  XOR U6848 ( .A(n5399), .B(n4843), .Z(n4500) );
  XNOR U6849 ( .A(n2210), .B(n5400), .Z(n4502) );
  XOR U6850 ( .A(n5401), .B(n4953), .Z(out[1321]) );
  XOR U6851 ( .A(n5402), .B(n2079), .Z(n4953) );
  NOR U6852 ( .A(n4505), .B(n4504), .Z(n5401) );
  XOR U6853 ( .A(n5403), .B(n2241), .Z(n4504) );
  XNOR U6854 ( .A(n2217), .B(n5404), .Z(n4505) );
  XNOR U6855 ( .A(n5405), .B(n4956), .Z(out[1320]) );
  IV U6856 ( .A(n5168), .Z(n4956) );
  XNOR U6857 ( .A(n5406), .B(n2082), .Z(n5168) );
  ANDN U6858 ( .B(n4508), .A(n4509), .Z(n5405) );
  XOR U6859 ( .A(n2222), .B(n5407), .Z(n4509) );
  XOR U6860 ( .A(n5409), .B(n4095), .Z(out[131]) );
  XNOR U6861 ( .A(n5410), .B(n2072), .Z(n4095) );
  AND U6862 ( .A(n2386), .B(n2384), .Z(n5409) );
  XOR U6863 ( .A(n5411), .B(n5412), .Z(n2384) );
  XOR U6864 ( .A(n5413), .B(n2664), .Z(n2386) );
  IV U6865 ( .A(n5414), .Z(n2664) );
  XOR U6866 ( .A(n5415), .B(n4959), .Z(out[1319]) );
  XOR U6867 ( .A(n5416), .B(n2086), .Z(n4959) );
  ANDN U6868 ( .B(n4512), .A(n4514), .Z(n5415) );
  XOR U6869 ( .A(n2231), .B(n5417), .Z(n4514) );
  XNOR U6870 ( .A(n5418), .B(n2255), .Z(n4512) );
  IV U6871 ( .A(n5419), .Z(n2255) );
  XOR U6872 ( .A(n5420), .B(n4962), .Z(out[1318]) );
  XOR U6873 ( .A(n5421), .B(n2089), .Z(n4962) );
  NOR U6874 ( .A(n4518), .B(n4516), .Z(n5420) );
  XOR U6875 ( .A(n5422), .B(n3870), .Z(n4516) );
  XOR U6876 ( .A(n2244), .B(n5423), .Z(n4518) );
  XOR U6877 ( .A(n5424), .B(n4965), .Z(out[1317]) );
  XNOR U6878 ( .A(n5425), .B(n2092), .Z(n4965) );
  NOR U6879 ( .A(n4521), .B(n4520), .Z(n5424) );
  XOR U6880 ( .A(n5426), .B(n5023), .Z(n4520) );
  XOR U6881 ( .A(n5427), .B(n3384), .Z(n4521) );
  XOR U6882 ( .A(n5428), .B(n4969), .Z(out[1316]) );
  XNOR U6883 ( .A(n5429), .B(n2095), .Z(n4969) );
  AND U6884 ( .A(n4526), .B(n4524), .Z(n5428) );
  XOR U6885 ( .A(n5430), .B(n3881), .Z(n4524) );
  XOR U6886 ( .A(n5431), .B(n5432), .Z(n4526) );
  XOR U6887 ( .A(n5433), .B(n4972), .Z(out[1315]) );
  XOR U6888 ( .A(n5434), .B(n2098), .Z(n4972) );
  ANDN U6889 ( .B(n4528), .A(n4529), .Z(n5433) );
  XNOR U6890 ( .A(n5435), .B(n2264), .Z(n4529) );
  XNOR U6891 ( .A(n5436), .B(n2283), .Z(n4528) );
  XOR U6892 ( .A(n5437), .B(n4976), .Z(out[1314]) );
  XNOR U6893 ( .A(n5438), .B(n2101), .Z(n4976) );
  ANDN U6894 ( .B(n4532), .A(n4534), .Z(n5437) );
  XOR U6895 ( .A(n5439), .B(n3401), .Z(n4534) );
  XNOR U6896 ( .A(n5440), .B(n2290), .Z(n4532) );
  IV U6897 ( .A(n5127), .Z(n2290) );
  XNOR U6898 ( .A(n5441), .B(n5193), .Z(out[1313]) );
  XOR U6899 ( .A(n3690), .B(n5442), .Z(n5193) );
  ANDN U6900 ( .B(n4542), .A(n4540), .Z(n5441) );
  XOR U6901 ( .A(n5443), .B(n2297), .Z(n4540) );
  XOR U6902 ( .A(n5444), .B(n2280), .Z(n4542) );
  XNOR U6903 ( .A(n5445), .B(n4983), .Z(out[1312]) );
  IV U6904 ( .A(n5197), .Z(n4983) );
  XOR U6905 ( .A(n4323), .B(n5446), .Z(n5197) );
  ANDN U6906 ( .B(n4544), .A(n4546), .Z(n5445) );
  XNOR U6907 ( .A(n5447), .B(n2287), .Z(n4546) );
  IV U6908 ( .A(n3142), .Z(n2287) );
  XNOR U6909 ( .A(n5448), .B(n3899), .Z(n4544) );
  XOR U6910 ( .A(n5449), .B(n4991), .Z(out[1311]) );
  XOR U6911 ( .A(n5450), .B(n2114), .Z(n4991) );
  ANDN U6912 ( .B(n4551), .A(n4547), .Z(n5449) );
  XOR U6913 ( .A(n5451), .B(n2315), .Z(n4547) );
  IV U6914 ( .A(n5452), .Z(n2315) );
  XNOR U6915 ( .A(n5453), .B(n2294), .Z(n4551) );
  XNOR U6916 ( .A(n5454), .B(n4994), .Z(out[1310]) );
  XOR U6917 ( .A(n4328), .B(n5455), .Z(n4994) );
  ANDN U6918 ( .B(n4556), .A(n4554), .Z(n5454) );
  XNOR U6919 ( .A(n5456), .B(n3908), .Z(n4554) );
  XNOR U6920 ( .A(n5457), .B(n2301), .Z(n4556) );
  XNOR U6921 ( .A(n5458), .B(n4098), .Z(out[130]) );
  IV U6922 ( .A(n4298), .Z(n4098) );
  XOR U6923 ( .A(n5459), .B(n2079), .Z(n4298) );
  ANDN U6924 ( .B(n2460), .A(n2458), .Z(n5458) );
  XOR U6925 ( .A(n5460), .B(n2357), .Z(n2458) );
  XNOR U6926 ( .A(n5461), .B(n3356), .Z(n2460) );
  IV U6927 ( .A(n2671), .Z(n3356) );
  XNOR U6928 ( .A(n5462), .B(n4997), .Z(out[1309]) );
  XOR U6929 ( .A(n4331), .B(n5463), .Z(n4997) );
  ANDN U6930 ( .B(n4558), .A(n4559), .Z(n5462) );
  XOR U6931 ( .A(n5464), .B(n3158), .Z(n4559) );
  XOR U6932 ( .A(n5465), .B(n2329), .Z(n4558) );
  IV U6933 ( .A(n5466), .Z(n2329) );
  XNOR U6934 ( .A(n5467), .B(n5000), .Z(out[1308]) );
  XOR U6935 ( .A(n5468), .B(n5469), .Z(n5000) );
  ANDN U6936 ( .B(n4564), .A(n4562), .Z(n5467) );
  XOR U6937 ( .A(n5470), .B(n2336), .Z(n4562) );
  IV U6938 ( .A(n5471), .Z(n2336) );
  XNOR U6939 ( .A(n5472), .B(n2319), .Z(n4564) );
  XOR U6940 ( .A(n5473), .B(n5003), .Z(out[1307]) );
  XNOR U6941 ( .A(n2128), .B(n5474), .Z(n5003) );
  AND U6942 ( .A(n4566), .B(n4567), .Z(n5473) );
  XOR U6943 ( .A(n5475), .B(n5476), .Z(n4567) );
  XOR U6944 ( .A(n5477), .B(n2343), .Z(n4566) );
  XOR U6945 ( .A(n5478), .B(n5006), .Z(out[1306]) );
  XOR U6946 ( .A(n2131), .B(n5479), .Z(n5006) );
  IV U6947 ( .A(n3728), .Z(n2131) );
  ANDN U6948 ( .B(n4570), .A(n4571), .Z(n5478) );
  XNOR U6949 ( .A(n5480), .B(n2331), .Z(n4571) );
  IV U6950 ( .A(n5481), .Z(n2331) );
  XNOR U6951 ( .A(n5482), .B(n2350), .Z(n4570) );
  IV U6952 ( .A(n5412), .Z(n2350) );
  XOR U6953 ( .A(n5483), .B(n5009), .Z(out[1305]) );
  XNOR U6954 ( .A(n2134), .B(n5484), .Z(n5009) );
  AND U6955 ( .A(n4576), .B(n4574), .Z(n5483) );
  XOR U6956 ( .A(n5485), .B(n3614), .Z(n4574) );
  IV U6957 ( .A(n2357), .Z(n3614) );
  XOR U6958 ( .A(n5486), .B(n2338), .Z(n4576) );
  XNOR U6959 ( .A(n5487), .B(n5012), .Z(out[1304]) );
  XNOR U6960 ( .A(n5488), .B(n2139), .Z(n5012) );
  ANDN U6961 ( .B(n4578), .A(n4580), .Z(n5487) );
  XOR U6962 ( .A(n5489), .B(n2345), .Z(n4580) );
  XOR U6963 ( .A(n5490), .B(n2364), .Z(n4578) );
  XNOR U6964 ( .A(n5491), .B(n5015), .Z(out[1303]) );
  IV U6965 ( .A(n5225), .Z(n5015) );
  XNOR U6966 ( .A(n5492), .B(n2142), .Z(n5225) );
  ANDN U6967 ( .B(n4586), .A(n4587), .Z(n5491) );
  XNOR U6968 ( .A(n5493), .B(n2352), .Z(n4587) );
  XNOR U6969 ( .A(n5494), .B(n2371), .Z(n4586) );
  XOR U6970 ( .A(n5495), .B(n5018), .Z(out[1302]) );
  XOR U6971 ( .A(n5496), .B(n2146), .Z(n5018) );
  NOR U6972 ( .A(n4592), .B(n4590), .Z(n5495) );
  XNOR U6973 ( .A(n5497), .B(n3634), .Z(n4590) );
  XOR U6974 ( .A(n5498), .B(n2359), .Z(n4592) );
  XOR U6975 ( .A(n5499), .B(n5026), .Z(out[1301]) );
  XOR U6976 ( .A(n5500), .B(n2152), .Z(n5026) );
  AND U6977 ( .A(n4596), .B(n4594), .Z(n5499) );
  XNOR U6978 ( .A(n5501), .B(n2389), .Z(n4594) );
  XOR U6979 ( .A(n5502), .B(n2366), .Z(n4596) );
  XOR U6980 ( .A(n5503), .B(n5029), .Z(out[1300]) );
  XOR U6981 ( .A(n5504), .B(n2155), .Z(n5029) );
  ANDN U6982 ( .B(n4600), .A(n5234), .Z(n5503) );
  XOR U6983 ( .A(n5505), .B(n2396), .Z(n5234) );
  XOR U6984 ( .A(n5506), .B(n2373), .Z(n4600) );
  XOR U6985 ( .A(n5507), .B(n1966), .Z(out[12]) );
  XNOR U6986 ( .A(n5508), .B(n2595), .Z(n1966) );
  NOR U6987 ( .A(n4063), .B(n1965), .Z(n5507) );
  XNOR U6988 ( .A(n2527), .B(n5509), .Z(n1965) );
  XNOR U6989 ( .A(n5510), .B(n1749), .Z(n4063) );
  XOR U6990 ( .A(n5511), .B(n4101), .Z(out[129]) );
  XNOR U6991 ( .A(n5512), .B(n2082), .Z(n4101) );
  ANDN U6992 ( .B(n2534), .A(n4301), .Z(n5511) );
  XOR U6993 ( .A(n5513), .B(n2364), .Z(n4301) );
  IV U6994 ( .A(n3620), .Z(n2364) );
  XNOR U6995 ( .A(n5514), .B(n2678), .Z(n2534) );
  IV U6996 ( .A(n5515), .Z(n2678) );
  XNOR U6997 ( .A(n5516), .B(n5032), .Z(out[1299]) );
  IV U6998 ( .A(n5237), .Z(n5032) );
  XOR U6999 ( .A(n5517), .B(n2158), .Z(n5237) );
  ANDN U7000 ( .B(n4602), .A(n4603), .Z(n5516) );
  XOR U7001 ( .A(n5518), .B(n2380), .Z(n4603) );
  XOR U7002 ( .A(n5519), .B(n2403), .Z(n4602) );
  XOR U7003 ( .A(n5520), .B(n5035), .Z(out[1298]) );
  XOR U7004 ( .A(n5521), .B(n2161), .Z(n5035) );
  ANDN U7005 ( .B(n4606), .A(n4608), .Z(n5520) );
  XNOR U7006 ( .A(n5522), .B(n2391), .Z(n4608) );
  XOR U7007 ( .A(n5523), .B(n2410), .Z(n4606) );
  XOR U7008 ( .A(n5524), .B(n5038), .Z(out[1297]) );
  XOR U7009 ( .A(n5525), .B(n2164), .Z(n5038) );
  ANDN U7010 ( .B(n4612), .A(n4610), .Z(n5524) );
  XNOR U7011 ( .A(n5526), .B(n2417), .Z(n4610) );
  XOR U7012 ( .A(n5527), .B(n2400), .Z(n4612) );
  XOR U7013 ( .A(n5528), .B(n5041), .Z(out[1296]) );
  XOR U7014 ( .A(n5529), .B(n2169), .Z(n5041) );
  ANDN U7015 ( .B(n4614), .A(n4616), .Z(n5528) );
  XOR U7016 ( .A(n5530), .B(n2407), .Z(n4616) );
  XNOR U7017 ( .A(n5531), .B(n2424), .Z(n4614) );
  XOR U7018 ( .A(n5532), .B(n5045), .Z(out[1295]) );
  XOR U7019 ( .A(n5533), .B(n3780), .Z(n5045) );
  NOR U7020 ( .A(n4617), .B(n4622), .Z(n5532) );
  XOR U7021 ( .A(n5534), .B(n2412), .Z(n4622) );
  IV U7022 ( .A(n5254), .Z(n4617) );
  XOR U7023 ( .A(n5535), .B(n2431), .Z(n5254) );
  XOR U7024 ( .A(n5536), .B(n5049), .Z(out[1294]) );
  XOR U7025 ( .A(n5537), .B(n2175), .Z(n5049) );
  AND U7026 ( .A(n4625), .B(n4624), .Z(n5536) );
  XNOR U7027 ( .A(n5538), .B(n2438), .Z(n4624) );
  XOR U7028 ( .A(n5539), .B(n2421), .Z(n4625) );
  XNOR U7029 ( .A(n5540), .B(n5260), .Z(out[1293]) );
  XOR U7030 ( .A(n5541), .B(n2178), .Z(n5260) );
  IV U7031 ( .A(n3791), .Z(n2178) );
  ANDN U7032 ( .B(n4632), .A(n4633), .Z(n5540) );
  XOR U7033 ( .A(n2425), .B(n5542), .Z(n4633) );
  IV U7034 ( .A(n5543), .Z(n2425) );
  XNOR U7035 ( .A(n5544), .B(n2445), .Z(n4632) );
  XOR U7036 ( .A(n5545), .B(n5055), .Z(out[1292]) );
  XNOR U7037 ( .A(n5546), .B(n2181), .Z(n5055) );
  ANDN U7038 ( .B(n4636), .A(n4638), .Z(n5545) );
  XOR U7039 ( .A(n2432), .B(n5547), .Z(n4638) );
  XNOR U7040 ( .A(n5548), .B(n2452), .Z(n4636) );
  XOR U7041 ( .A(n5549), .B(n5061), .Z(out[1291]) );
  XOR U7042 ( .A(n5550), .B(n2188), .Z(n5061) );
  ANDN U7043 ( .B(n4640), .A(n4641), .Z(n5549) );
  XOR U7044 ( .A(n5551), .B(n2440), .Z(n4641) );
  XOR U7045 ( .A(n5552), .B(n2463), .Z(n4640) );
  XOR U7046 ( .A(n5553), .B(n5065), .Z(out[1290]) );
  XOR U7047 ( .A(n5554), .B(n3805), .Z(n5065) );
  ANDN U7048 ( .B(n4644), .A(n4645), .Z(n5553) );
  XNOR U7049 ( .A(n5555), .B(n2447), .Z(n4645) );
  XOR U7050 ( .A(n5556), .B(n2470), .Z(n4644) );
  XOR U7051 ( .A(n5557), .B(n4104), .Z(out[128]) );
  XOR U7052 ( .A(n5558), .B(n2086), .Z(n4104) );
  ANDN U7053 ( .B(n2608), .A(n2606), .Z(n5557) );
  IV U7054 ( .A(n4303), .Z(n2606) );
  XOR U7055 ( .A(n5559), .B(n2371), .Z(n4303) );
  IV U7056 ( .A(n5560), .Z(n2371) );
  XOR U7057 ( .A(n5561), .B(n5068), .Z(out[1289]) );
  XOR U7058 ( .A(n5562), .B(n2194), .Z(n5068) );
  AND U7059 ( .A(n4650), .B(n4648), .Z(n5561) );
  XOR U7060 ( .A(n5563), .B(n5564), .Z(n4648) );
  XOR U7061 ( .A(n5565), .B(n2454), .Z(n4650) );
  XOR U7062 ( .A(n5566), .B(n5072), .Z(out[1288]) );
  XOR U7063 ( .A(n5567), .B(n2197), .Z(n5072) );
  NOR U7064 ( .A(n4653), .B(n4652), .Z(n5566) );
  XOR U7065 ( .A(n5568), .B(n2484), .Z(n4652) );
  XOR U7066 ( .A(n5569), .B(n4450), .Z(n4653) );
  IV U7067 ( .A(n2465), .Z(n4450) );
  XOR U7068 ( .A(n5570), .B(n5076), .Z(out[1287]) );
  XOR U7069 ( .A(n5571), .B(n3820), .Z(n5076) );
  ANDN U7070 ( .B(n4656), .A(n4658), .Z(n5570) );
  XOR U7071 ( .A(n5572), .B(n2472), .Z(n4658) );
  XOR U7072 ( .A(n5573), .B(n2491), .Z(n4656) );
  XNOR U7073 ( .A(n5574), .B(n5079), .Z(out[1286]) );
  XOR U7074 ( .A(n5575), .B(n2203), .Z(n5079) );
  NOR U7075 ( .A(n4661), .B(n4660), .Z(n5574) );
  XNOR U7076 ( .A(n5576), .B(n3711), .Z(n4660) );
  IV U7077 ( .A(n2498), .Z(n3711) );
  XOR U7078 ( .A(n5577), .B(n2479), .Z(n4661) );
  XOR U7079 ( .A(n5578), .B(n5082), .Z(out[1285]) );
  XOR U7080 ( .A(n5579), .B(n3834), .Z(n5082) );
  ANDN U7081 ( .B(n4664), .A(n4665), .Z(n5578) );
  XOR U7082 ( .A(n5580), .B(n2486), .Z(n4665) );
  XOR U7083 ( .A(n5581), .B(n2505), .Z(n4664) );
  XNOR U7084 ( .A(n5582), .B(n5085), .Z(out[1284]) );
  XOR U7085 ( .A(n5583), .B(n5584), .Z(n5085) );
  NOR U7086 ( .A(n4670), .B(n4668), .Z(n5582) );
  XOR U7087 ( .A(n5585), .B(n2512), .Z(n4668) );
  XOR U7088 ( .A(n5586), .B(n2495), .Z(n4670) );
  XOR U7089 ( .A(n5587), .B(n5088), .Z(out[1283]) );
  XOR U7090 ( .A(n5588), .B(n3843), .Z(n5088) );
  ANDN U7091 ( .B(n4675), .A(n4679), .Z(n5587) );
  XNOR U7092 ( .A(n5589), .B(n2500), .Z(n4679) );
  XOR U7093 ( .A(n5590), .B(n3731), .Z(n4675) );
  XNOR U7094 ( .A(n5591), .B(n5092), .Z(out[1282]) );
  IV U7095 ( .A(n5290), .Z(n5092) );
  XNOR U7096 ( .A(n5592), .B(n1986), .Z(n5290) );
  NOR U7097 ( .A(n4683), .B(n4682), .Z(n5591) );
  XNOR U7098 ( .A(n5593), .B(n2526), .Z(n4682) );
  XOR U7099 ( .A(n5594), .B(n2509), .Z(n4683) );
  IV U7100 ( .A(n3261), .Z(n2509) );
  XOR U7101 ( .A(n5595), .B(n5099), .Z(out[1281]) );
  XOR U7102 ( .A(n5596), .B(n1989), .Z(n5099) );
  NOR U7103 ( .A(n4689), .B(n4685), .Z(n5595) );
  XOR U7104 ( .A(n5597), .B(n2537), .Z(n4685) );
  XOR U7105 ( .A(n5598), .B(n2516), .Z(n4689) );
  XOR U7106 ( .A(n5599), .B(n5102), .Z(out[1280]) );
  XOR U7107 ( .A(n5600), .B(n1992), .Z(n5102) );
  NOR U7108 ( .A(n4696), .B(n4691), .Z(n5599) );
  XNOR U7109 ( .A(n5601), .B(n2544), .Z(n4691) );
  XNOR U7110 ( .A(n5602), .B(n2523), .Z(n4696) );
  XOR U7111 ( .A(n5603), .B(n4307), .Z(out[127]) );
  XOR U7112 ( .A(n5604), .B(n2378), .Z(n4307) );
  ANDN U7113 ( .B(n2682), .A(n4306), .Z(n5603) );
  XNOR U7114 ( .A(n2217), .B(n5605), .Z(n4306) );
  XNOR U7115 ( .A(n5606), .B(n4939), .Z(n2682) );
  XOR U7116 ( .A(n5607), .B(n5608), .Z(out[1279]) );
  ANDN U7117 ( .B(n5609), .A(n5610), .Z(n5607) );
  XNOR U7118 ( .A(n5611), .B(n5612), .Z(out[1278]) );
  ANDN U7119 ( .B(n5613), .A(n5614), .Z(n5611) );
  XOR U7120 ( .A(n5615), .B(n5616), .Z(out[1277]) );
  XNOR U7121 ( .A(n5619), .B(n5620), .Z(out[1276]) );
  XOR U7122 ( .A(n5623), .B(n5624), .Z(out[1275]) );
  AND U7123 ( .A(n5625), .B(n5626), .Z(n5623) );
  XOR U7124 ( .A(n5627), .B(n5628), .Z(out[1274]) );
  ANDN U7125 ( .B(n5629), .A(n5630), .Z(n5627) );
  XOR U7126 ( .A(n5631), .B(n5632), .Z(out[1273]) );
  ANDN U7127 ( .B(n5633), .A(n5634), .Z(n5631) );
  XOR U7128 ( .A(n5635), .B(n5636), .Z(out[1272]) );
  ANDN U7129 ( .B(n5637), .A(n5638), .Z(n5635) );
  XOR U7130 ( .A(n5639), .B(n5640), .Z(out[1271]) );
  ANDN U7131 ( .B(n5641), .A(n5642), .Z(n5639) );
  XNOR U7132 ( .A(n5643), .B(n5644), .Z(out[1270]) );
  ANDN U7133 ( .B(n5645), .A(n5646), .Z(n5643) );
  XOR U7134 ( .A(n5647), .B(n4112), .Z(out[126]) );
  XOR U7135 ( .A(n5648), .B(n2389), .Z(n4112) );
  IV U7136 ( .A(n3639), .Z(n2389) );
  ANDN U7137 ( .B(n2724), .A(n2726), .Z(n5647) );
  XNOR U7138 ( .A(n5649), .B(n2634), .Z(n2726) );
  XOR U7139 ( .A(n2222), .B(n5650), .Z(n2724) );
  IV U7140 ( .A(n3371), .Z(n2222) );
  XOR U7141 ( .A(n5651), .B(n5652), .Z(out[1269]) );
  ANDN U7142 ( .B(n5653), .A(n5654), .Z(n5651) );
  XNOR U7143 ( .A(n5655), .B(n5656), .Z(out[1268]) );
  ANDN U7144 ( .B(n5657), .A(n5658), .Z(n5655) );
  XOR U7145 ( .A(n5659), .B(n5660), .Z(out[1267]) );
  ANDN U7146 ( .B(n5661), .A(n5662), .Z(n5659) );
  XNOR U7147 ( .A(n5663), .B(n5664), .Z(out[1266]) );
  ANDN U7148 ( .B(n5665), .A(n5666), .Z(n5663) );
  XOR U7149 ( .A(n5667), .B(n5668), .Z(out[1265]) );
  ANDN U7150 ( .B(n5669), .A(n5670), .Z(n5667) );
  XOR U7151 ( .A(n5671), .B(n5672), .Z(out[1264]) );
  ANDN U7152 ( .B(n5673), .A(n5674), .Z(n5671) );
  XOR U7153 ( .A(n5675), .B(n5676), .Z(out[1263]) );
  ANDN U7154 ( .B(n5677), .A(n5678), .Z(n5675) );
  XNOR U7155 ( .A(n5679), .B(n5680), .Z(out[1262]) );
  AND U7156 ( .A(n5681), .B(n5682), .Z(n5679) );
  XOR U7157 ( .A(n5683), .B(n5684), .Z(out[1261]) );
  ANDN U7158 ( .B(n5685), .A(n5686), .Z(n5683) );
  XNOR U7159 ( .A(n5687), .B(n5688), .Z(out[1260]) );
  XNOR U7160 ( .A(n5691), .B(n4115), .Z(out[125]) );
  IV U7161 ( .A(n4315), .Z(n4115) );
  XOR U7162 ( .A(n5692), .B(n2396), .Z(n4315) );
  NOR U7163 ( .A(n2770), .B(n2768), .Z(n5691) );
  XNOR U7164 ( .A(n2231), .B(n5693), .Z(n2768) );
  IV U7165 ( .A(n5694), .Z(n2231) );
  XOR U7166 ( .A(n5695), .B(n2641), .Z(n2770) );
  XNOR U7167 ( .A(n5696), .B(n5697), .Z(out[1259]) );
  ANDN U7168 ( .B(n5698), .A(n5699), .Z(n5696) );
  XNOR U7169 ( .A(n5700), .B(n5701), .Z(out[1258]) );
  AND U7170 ( .A(n5702), .B(n5703), .Z(n5700) );
  XNOR U7171 ( .A(n5704), .B(n5705), .Z(out[1257]) );
  AND U7172 ( .A(n5706), .B(n5707), .Z(n5704) );
  XOR U7173 ( .A(n5708), .B(n5709), .Z(out[1256]) );
  AND U7174 ( .A(n5710), .B(n5711), .Z(n5708) );
  XOR U7175 ( .A(n5712), .B(n1041), .Z(out[1255]) );
  IV U7176 ( .A(n5713), .Z(n1040) );
  XOR U7177 ( .A(n5715), .B(n1045), .Z(out[1254]) );
  XOR U7178 ( .A(n5717), .B(n1048), .Z(out[1253]) );
  AND U7179 ( .A(n1049), .B(n5718), .Z(n5717) );
  XOR U7180 ( .A(n5719), .B(n1053), .Z(out[1252]) );
  ANDN U7181 ( .B(n5720), .A(n1052), .Z(n5719) );
  XOR U7182 ( .A(n5721), .B(n1057), .Z(out[1251]) );
  ANDN U7183 ( .B(n5722), .A(n1056), .Z(n5721) );
  XOR U7184 ( .A(n5723), .B(n1061), .Z(out[1250]) );
  IV U7185 ( .A(n5724), .Z(n1060) );
  XOR U7186 ( .A(n5726), .B(n4119), .Z(out[124]) );
  XOR U7187 ( .A(n5727), .B(n2403), .Z(n4119) );
  NOR U7188 ( .A(n2814), .B(n2812), .Z(n5726) );
  XNOR U7189 ( .A(n5728), .B(n5729), .Z(n2812) );
  XOR U7190 ( .A(n5730), .B(n2648), .Z(n2814) );
  XOR U7191 ( .A(n5731), .B(n1065), .Z(out[1249]) );
  ANDN U7192 ( .B(n5732), .A(n1064), .Z(n5731) );
  IV U7193 ( .A(n5733), .Z(n1064) );
  XNOR U7194 ( .A(n5734), .B(n1069), .Z(out[1248]) );
  ANDN U7195 ( .B(n5735), .A(n1068), .Z(n5734) );
  XNOR U7196 ( .A(n5736), .B(n1072), .Z(out[1247]) );
  ANDN U7197 ( .B(n5737), .A(n5738), .Z(n5736) );
  XOR U7198 ( .A(n5739), .B(n1076), .Z(out[1246]) );
  AND U7199 ( .A(n1077), .B(n5740), .Z(n5739) );
  XNOR U7200 ( .A(n5741), .B(n1085), .Z(out[1245]) );
  ANDN U7201 ( .B(n5742), .A(n1084), .Z(n5741) );
  XNOR U7202 ( .A(n5743), .B(n1089), .Z(out[1244]) );
  ANDN U7203 ( .B(n5744), .A(n1088), .Z(n5743) );
  XNOR U7204 ( .A(n5745), .B(n1093), .Z(out[1243]) );
  ANDN U7205 ( .B(n5746), .A(n1092), .Z(n5745) );
  XNOR U7206 ( .A(n5747), .B(n1096), .Z(out[1242]) );
  ANDN U7207 ( .B(n5748), .A(n5749), .Z(n5747) );
  XOR U7208 ( .A(n5750), .B(n1100), .Z(out[1241]) );
  AND U7209 ( .A(n1101), .B(n5751), .Z(n5750) );
  XOR U7210 ( .A(n5752), .B(n1105), .Z(out[1240]) );
  XOR U7211 ( .A(n5754), .B(n4123), .Z(out[123]) );
  XOR U7212 ( .A(n5755), .B(n2410), .Z(n4123) );
  NOR U7213 ( .A(n2861), .B(n2859), .Z(n5754) );
  XNOR U7214 ( .A(n5756), .B(n3384), .Z(n2859) );
  IV U7215 ( .A(n2252), .Z(n3384) );
  XOR U7216 ( .A(n5757), .B(n2655), .Z(n2861) );
  XNOR U7217 ( .A(n5758), .B(n1108), .Z(out[1239]) );
  ANDN U7218 ( .B(n5759), .A(n5760), .Z(n5758) );
  XOR U7219 ( .A(n5761), .B(n1112), .Z(out[1238]) );
  AND U7220 ( .A(n1113), .B(n5762), .Z(n5761) );
  XOR U7221 ( .A(n5763), .B(n1117), .Z(out[1237]) );
  ANDN U7222 ( .B(n5764), .A(n1116), .Z(n5763) );
  IV U7223 ( .A(n5765), .Z(n1116) );
  XOR U7224 ( .A(n5766), .B(n1120), .Z(out[1236]) );
  AND U7225 ( .A(n1121), .B(n5767), .Z(n5766) );
  XOR U7226 ( .A(n5768), .B(n1129), .Z(out[1235]) );
  ANDN U7227 ( .B(n5769), .A(n1128), .Z(n5768) );
  IV U7228 ( .A(n5770), .Z(n1128) );
  XOR U7229 ( .A(n5771), .B(n1132), .Z(out[1234]) );
  AND U7230 ( .A(n1133), .B(n5772), .Z(n5771) );
  XNOR U7231 ( .A(n5773), .B(n1136), .Z(out[1233]) );
  ANDN U7232 ( .B(n5774), .A(n5775), .Z(n5773) );
  XNOR U7233 ( .A(n5776), .B(n1140), .Z(out[1232]) );
  XOR U7234 ( .A(n5778), .B(n1144), .Z(out[1231]) );
  AND U7235 ( .A(n1145), .B(n5779), .Z(n5778) );
  XNOR U7236 ( .A(n5780), .B(n1148), .Z(out[1230]) );
  ANDN U7237 ( .B(n5781), .A(n5782), .Z(n5780) );
  XOR U7238 ( .A(n5783), .B(n4126), .Z(out[122]) );
  XOR U7239 ( .A(n5784), .B(n3657), .Z(n4126) );
  NOR U7240 ( .A(n2905), .B(n2903), .Z(n5783) );
  XOR U7241 ( .A(n5785), .B(n5432), .Z(n2903) );
  IV U7242 ( .A(n2259), .Z(n5432) );
  XOR U7243 ( .A(n5786), .B(n2662), .Z(n2905) );
  XOR U7244 ( .A(n5787), .B(n1153), .Z(out[1229]) );
  ANDN U7245 ( .B(n5788), .A(n1152), .Z(n5787) );
  XOR U7246 ( .A(n5789), .B(n1157), .Z(out[1228]) );
  ANDN U7247 ( .B(n5790), .A(n5791), .Z(n5789) );
  XOR U7248 ( .A(n5792), .B(n1161), .Z(out[1227]) );
  ANDN U7249 ( .B(n1160), .A(n5793), .Z(n5792) );
  XNOR U7250 ( .A(n5794), .B(n1165), .Z(out[1226]) );
  ANDN U7251 ( .B(n5795), .A(n1164), .Z(n5794) );
  XNOR U7252 ( .A(n5796), .B(n1172), .Z(out[1225]) );
  XNOR U7253 ( .A(n5798), .B(n1176), .Z(out[1224]) );
  ANDN U7254 ( .B(n1177), .A(n5799), .Z(n5798) );
  XNOR U7255 ( .A(n5800), .B(n1180), .Z(out[1223]) );
  ANDN U7256 ( .B(n5801), .A(n5802), .Z(n5800) );
  XNOR U7257 ( .A(n5803), .B(n1184), .Z(out[1222]) );
  ANDN U7258 ( .B(n5804), .A(n5805), .Z(n5803) );
  XOR U7259 ( .A(n5806), .B(n1189), .Z(out[1221]) );
  ANDN U7260 ( .B(n5807), .A(n5808), .Z(n5806) );
  XOR U7261 ( .A(n5809), .B(n1193), .Z(out[1220]) );
  ANDN U7262 ( .B(n5810), .A(n5811), .Z(n5809) );
  XOR U7263 ( .A(n5812), .B(n4132), .Z(out[121]) );
  XOR U7264 ( .A(n5813), .B(n2424), .Z(n4132) );
  IV U7265 ( .A(n5814), .Z(n2424) );
  ANDN U7266 ( .B(n2947), .A(n2948), .Z(n5812) );
  XOR U7267 ( .A(n5815), .B(n2669), .Z(n2948) );
  XNOR U7268 ( .A(n5816), .B(n2264), .Z(n2947) );
  IV U7269 ( .A(n3397), .Z(n2264) );
  XOR U7270 ( .A(n5817), .B(n1197), .Z(out[1219]) );
  ANDN U7271 ( .B(n5818), .A(n5819), .Z(n5817) );
  XNOR U7272 ( .A(n5820), .B(n1201), .Z(out[1218]) );
  ANDN U7273 ( .B(n5821), .A(n1200), .Z(n5820) );
  XNOR U7274 ( .A(n5822), .B(n1205), .Z(out[1217]) );
  ANDN U7275 ( .B(n5823), .A(n1204), .Z(n5822) );
  XOR U7276 ( .A(n5824), .B(n1209), .Z(out[1216]) );
  AND U7277 ( .A(n1208), .B(n5825), .Z(n5824) );
  XOR U7278 ( .A(n5826), .B(n5610), .Z(out[1215]) );
  ANDN U7279 ( .B(n5827), .A(n5609), .Z(n5826) );
  XOR U7280 ( .A(n5828), .B(n5614), .Z(out[1214]) );
  NOR U7281 ( .A(n5829), .B(n5613), .Z(n5828) );
  XNOR U7282 ( .A(n5830), .B(n5618), .Z(out[1213]) );
  ANDN U7283 ( .B(n5831), .A(n5617), .Z(n5830) );
  XNOR U7284 ( .A(n5832), .B(n5622), .Z(out[1212]) );
  ANDN U7285 ( .B(n5833), .A(n5621), .Z(n5832) );
  IV U7286 ( .A(n5834), .Z(n5621) );
  XNOR U7287 ( .A(n5835), .B(n5626), .Z(out[1211]) );
  ANDN U7288 ( .B(n5836), .A(n5625), .Z(n5835) );
  XOR U7289 ( .A(n5837), .B(n5630), .Z(out[1210]) );
  NOR U7290 ( .A(n5838), .B(n5629), .Z(n5837) );
  XOR U7291 ( .A(n5839), .B(n4135), .Z(out[120]) );
  XOR U7292 ( .A(n5840), .B(n2431), .Z(n4135) );
  ANDN U7293 ( .B(n2981), .A(n2982), .Z(n5839) );
  XOR U7294 ( .A(n5841), .B(n2676), .Z(n2982) );
  XOR U7295 ( .A(n5842), .B(n3401), .Z(n2981) );
  IV U7296 ( .A(n2273), .Z(n3401) );
  XOR U7297 ( .A(n5843), .B(n5634), .Z(out[1209]) );
  ANDN U7298 ( .B(n5844), .A(n5633), .Z(n5843) );
  XNOR U7299 ( .A(n5845), .B(n5637), .Z(out[1208]) );
  ANDN U7300 ( .B(n5846), .A(n5847), .Z(n5845) );
  XOR U7301 ( .A(n5848), .B(n5642), .Z(out[1207]) );
  ANDN U7302 ( .B(n5849), .A(n5641), .Z(n5848) );
  XOR U7303 ( .A(n5850), .B(n5646), .Z(out[1206]) );
  ANDN U7304 ( .B(n5851), .A(n5645), .Z(n5850) );
  XOR U7305 ( .A(n5852), .B(n5654), .Z(out[1205]) );
  ANDN U7306 ( .B(n5853), .A(n5653), .Z(n5852) );
  XOR U7307 ( .A(n5854), .B(n5658), .Z(out[1204]) );
  ANDN U7308 ( .B(n5855), .A(n5657), .Z(n5854) );
  XOR U7309 ( .A(n5856), .B(n5662), .Z(out[1203]) );
  ANDN U7310 ( .B(n5857), .A(n5661), .Z(n5856) );
  XOR U7311 ( .A(n5858), .B(n5666), .Z(out[1202]) );
  NOR U7312 ( .A(n5859), .B(n5665), .Z(n5858) );
  XOR U7313 ( .A(n5860), .B(n5670), .Z(out[1201]) );
  ANDN U7314 ( .B(n5861), .A(n5669), .Z(n5860) );
  XNOR U7315 ( .A(n5862), .B(n5673), .Z(out[1200]) );
  ANDN U7316 ( .B(n5863), .A(n5864), .Z(n5862) );
  XOR U7317 ( .A(n5865), .B(n2001), .Z(out[11]) );
  XOR U7318 ( .A(n5866), .B(n2604), .Z(n2001) );
  ANDN U7319 ( .B(n2002), .A(n4066), .Z(n5865) );
  XOR U7320 ( .A(n5867), .B(n1754), .Z(n4066) );
  XOR U7321 ( .A(n2540), .B(n5868), .Z(n2002) );
  IV U7322 ( .A(n3514), .Z(n2540) );
  XOR U7323 ( .A(n5869), .B(n4138), .Z(out[119]) );
  XOR U7324 ( .A(n5870), .B(n2438), .Z(n4138) );
  ANDN U7325 ( .B(n3009), .A(n3011), .Z(n5869) );
  XOR U7326 ( .A(n5871), .B(n2209), .Z(n3011) );
  XOR U7327 ( .A(n5872), .B(n2280), .Z(n3009) );
  XOR U7328 ( .A(n5873), .B(n5678), .Z(out[1199]) );
  ANDN U7329 ( .B(n5874), .A(n5677), .Z(n5873) );
  XNOR U7330 ( .A(n5875), .B(n5682), .Z(out[1198]) );
  ANDN U7331 ( .B(n5876), .A(n5681), .Z(n5875) );
  XOR U7332 ( .A(n5877), .B(n5686), .Z(out[1197]) );
  ANDN U7333 ( .B(n5878), .A(n5685), .Z(n5877) );
  XNOR U7334 ( .A(n5879), .B(n5690), .Z(out[1196]) );
  ANDN U7335 ( .B(n5880), .A(n5689), .Z(n5879) );
  XOR U7336 ( .A(n5881), .B(n5699), .Z(out[1195]) );
  ANDN U7337 ( .B(n5882), .A(n5698), .Z(n5881) );
  XNOR U7338 ( .A(n5883), .B(n5703), .Z(out[1194]) );
  NOR U7339 ( .A(n5884), .B(n5702), .Z(n5883) );
  XNOR U7340 ( .A(n5885), .B(n5707), .Z(out[1193]) );
  ANDN U7341 ( .B(n5886), .A(n5706), .Z(n5885) );
  XNOR U7342 ( .A(n5887), .B(n5711), .Z(out[1192]) );
  NOR U7343 ( .A(n5888), .B(n5710), .Z(n5887) );
  XNOR U7344 ( .A(n5889), .B(n5713), .Z(out[1191]) );
  XOR U7345 ( .A(n2104), .B(n5890), .Z(n5713) );
  IV U7346 ( .A(n3690), .Z(n2104) );
  XNOR U7347 ( .A(n5891), .B(n5892), .Z(n3690) );
  XNOR U7348 ( .A(n5894), .B(n1044), .Z(out[1190]) );
  XOR U7349 ( .A(n2108), .B(n5895), .Z(n1044) );
  IV U7350 ( .A(n4323), .Z(n2108) );
  XNOR U7351 ( .A(n5896), .B(n5897), .Z(n4323) );
  NOR U7352 ( .A(n5898), .B(n5716), .Z(n5894) );
  XOR U7353 ( .A(n5899), .B(n4141), .Z(out[118]) );
  XOR U7354 ( .A(n5900), .B(n2445), .Z(n4141) );
  ANDN U7355 ( .B(n3034), .A(n3035), .Z(n5899) );
  XOR U7356 ( .A(n5901), .B(n2216), .Z(n3035) );
  IV U7357 ( .A(n5902), .Z(n2216) );
  XOR U7358 ( .A(n5903), .B(n3142), .Z(n3034) );
  XNOR U7359 ( .A(n5904), .B(n1049), .Z(out[1189]) );
  XOR U7360 ( .A(n5905), .B(n2114), .Z(n1049) );
  XOR U7361 ( .A(n5906), .B(n5907), .Z(n2114) );
  NOR U7362 ( .A(n5908), .B(n5718), .Z(n5904) );
  XOR U7363 ( .A(n5909), .B(n1052), .Z(out[1188]) );
  XOR U7364 ( .A(n2116), .B(n5910), .Z(n1052) );
  IV U7365 ( .A(n4328), .Z(n2116) );
  XNOR U7366 ( .A(n5911), .B(n5912), .Z(n4328) );
  NOR U7367 ( .A(n5913), .B(n5720), .Z(n5909) );
  XOR U7368 ( .A(n5914), .B(n1056), .Z(out[1187]) );
  XOR U7369 ( .A(n2120), .B(n5915), .Z(n1056) );
  IV U7370 ( .A(n4331), .Z(n2120) );
  XNOR U7371 ( .A(n5916), .B(n5917), .Z(n4331) );
  NOR U7372 ( .A(n5918), .B(n5722), .Z(n5914) );
  XNOR U7373 ( .A(n5919), .B(n5724), .Z(out[1186]) );
  XOR U7374 ( .A(n2124), .B(n5920), .Z(n5724) );
  IV U7375 ( .A(n5468), .Z(n2124) );
  XNOR U7376 ( .A(n5921), .B(n5922), .Z(n5468) );
  XNOR U7377 ( .A(n5924), .B(n5733), .Z(out[1185]) );
  XOR U7378 ( .A(n2128), .B(n5925), .Z(n5733) );
  XNOR U7379 ( .A(n5926), .B(n5927), .Z(n2128) );
  ANDN U7380 ( .B(n5928), .A(n5732), .Z(n5924) );
  IV U7381 ( .A(n5929), .Z(n5732) );
  XOR U7382 ( .A(n5930), .B(n1068), .Z(out[1184]) );
  XOR U7383 ( .A(n3728), .B(n5931), .Z(n1068) );
  XNOR U7384 ( .A(n5932), .B(n5933), .Z(n3728) );
  ANDN U7385 ( .B(n5934), .A(n5735), .Z(n5930) );
  XNOR U7386 ( .A(n5935), .B(n1073), .Z(out[1183]) );
  IV U7387 ( .A(n5738), .Z(n1073) );
  XOR U7388 ( .A(n2134), .B(n5936), .Z(n5738) );
  XOR U7389 ( .A(n5937), .B(n5938), .Z(n2134) );
  NOR U7390 ( .A(n5939), .B(n5737), .Z(n5935) );
  XNOR U7391 ( .A(n5940), .B(n1077), .Z(out[1182]) );
  XNOR U7392 ( .A(n5941), .B(n2139), .Z(n1077) );
  XNOR U7393 ( .A(n5942), .B(n5943), .Z(n2139) );
  XOR U7394 ( .A(n5945), .B(n1084), .Z(out[1181]) );
  XNOR U7395 ( .A(n5946), .B(n2142), .Z(n1084) );
  XNOR U7396 ( .A(n5947), .B(n5948), .Z(n2142) );
  NOR U7397 ( .A(n5949), .B(n5742), .Z(n5945) );
  XOR U7398 ( .A(n5950), .B(n1088), .Z(out[1180]) );
  XNOR U7399 ( .A(n5951), .B(n2146), .Z(n1088) );
  XOR U7400 ( .A(n5952), .B(n5953), .Z(n2146) );
  ANDN U7401 ( .B(n5954), .A(n5744), .Z(n5950) );
  XNOR U7402 ( .A(n5955), .B(n4144), .Z(out[117]) );
  IV U7403 ( .A(n4335), .Z(n4144) );
  XOR U7404 ( .A(n5956), .B(n2452), .Z(n4335) );
  IV U7405 ( .A(n3683), .Z(n2452) );
  ANDN U7406 ( .B(n3063), .A(n3061), .Z(n5955) );
  XOR U7407 ( .A(n5957), .B(n2294), .Z(n3061) );
  XOR U7408 ( .A(n5958), .B(n2225), .Z(n3063) );
  IV U7409 ( .A(n5959), .Z(n2225) );
  XOR U7410 ( .A(n5960), .B(n1092), .Z(out[1179]) );
  XOR U7411 ( .A(n5961), .B(n2152), .Z(n1092) );
  XNOR U7412 ( .A(n5962), .B(n5963), .Z(n2152) );
  ANDN U7413 ( .B(n5964), .A(n5746), .Z(n5960) );
  XNOR U7414 ( .A(n5965), .B(n1097), .Z(out[1178]) );
  IV U7415 ( .A(n5749), .Z(n1097) );
  XOR U7416 ( .A(n5966), .B(n2155), .Z(n5749) );
  XNOR U7417 ( .A(n5967), .B(n5968), .Z(n2155) );
  ANDN U7418 ( .B(n5969), .A(n5748), .Z(n5965) );
  XNOR U7419 ( .A(n5970), .B(n1101), .Z(out[1177]) );
  XNOR U7420 ( .A(n5971), .B(n2158), .Z(n1101) );
  XNOR U7421 ( .A(n5972), .B(n5973), .Z(n2158) );
  NOR U7422 ( .A(n5974), .B(n5751), .Z(n5970) );
  XOR U7423 ( .A(n5975), .B(n1104), .Z(out[1176]) );
  XOR U7424 ( .A(n5976), .B(n2161), .Z(n1104) );
  XNOR U7425 ( .A(n5977), .B(n5978), .Z(n2161) );
  ANDN U7426 ( .B(n5753), .A(n5979), .Z(n5975) );
  XNOR U7427 ( .A(n5980), .B(n1109), .Z(out[1175]) );
  IV U7428 ( .A(n5760), .Z(n1109) );
  XOR U7429 ( .A(n5981), .B(n2164), .Z(n5760) );
  XNOR U7430 ( .A(n5982), .B(n5983), .Z(n2164) );
  NOR U7431 ( .A(n5984), .B(n5759), .Z(n5980) );
  XNOR U7432 ( .A(n5985), .B(n1113), .Z(out[1174]) );
  XNOR U7433 ( .A(n5986), .B(n2169), .Z(n1113) );
  XNOR U7434 ( .A(n5987), .B(n5988), .Z(n2169) );
  NOR U7435 ( .A(n5989), .B(n5762), .Z(n5985) );
  XNOR U7436 ( .A(n5990), .B(n5765), .Z(out[1173]) );
  XOR U7437 ( .A(n5991), .B(n3780), .Z(n5765) );
  XOR U7438 ( .A(n5992), .B(n5993), .Z(n3780) );
  NOR U7439 ( .A(n5994), .B(n5764), .Z(n5990) );
  XNOR U7440 ( .A(n5995), .B(n1121), .Z(out[1172]) );
  XNOR U7441 ( .A(n5996), .B(n2175), .Z(n1121) );
  XNOR U7442 ( .A(n5997), .B(n5998), .Z(n2175) );
  NOR U7443 ( .A(n5999), .B(n5767), .Z(n5995) );
  XNOR U7444 ( .A(n6000), .B(n5770), .Z(out[1171]) );
  XOR U7445 ( .A(n6001), .B(n3791), .Z(n5770) );
  ANDN U7446 ( .B(n6004), .A(n5769), .Z(n6000) );
  XNOR U7447 ( .A(n6005), .B(n1133), .Z(out[1170]) );
  XOR U7448 ( .A(n6006), .B(n2181), .Z(n1133) );
  XNOR U7449 ( .A(n6007), .B(n6008), .Z(n2181) );
  NOR U7450 ( .A(n6009), .B(n5772), .Z(n6005) );
  XOR U7451 ( .A(n6010), .B(n4147), .Z(out[116]) );
  XNOR U7452 ( .A(n6011), .B(n2463), .Z(n4147) );
  AND U7453 ( .A(n3090), .B(n3092), .Z(n6010) );
  XNOR U7454 ( .A(n6012), .B(n2230), .Z(n3092) );
  IV U7455 ( .A(n6013), .Z(n2230) );
  XOR U7456 ( .A(n6014), .B(n3154), .Z(n3090) );
  IV U7457 ( .A(n2301), .Z(n3154) );
  XNOR U7458 ( .A(n6015), .B(n1137), .Z(out[1169]) );
  IV U7459 ( .A(n5775), .Z(n1137) );
  XOR U7460 ( .A(n6016), .B(n2188), .Z(n5775) );
  XNOR U7461 ( .A(n6017), .B(n6018), .Z(n2188) );
  ANDN U7462 ( .B(n6019), .A(n5774), .Z(n6015) );
  XNOR U7463 ( .A(n6020), .B(n1141), .Z(out[1168]) );
  XOR U7464 ( .A(n6021), .B(n3805), .Z(n1141) );
  XOR U7465 ( .A(n6022), .B(n6023), .Z(n3805) );
  NOR U7466 ( .A(n6024), .B(n5777), .Z(n6020) );
  XNOR U7467 ( .A(n6025), .B(n1145), .Z(out[1167]) );
  XNOR U7468 ( .A(n6026), .B(n2194), .Z(n1145) );
  XNOR U7469 ( .A(n6027), .B(n6028), .Z(n2194) );
  ANDN U7470 ( .B(n6029), .A(n5779), .Z(n6025) );
  XNOR U7471 ( .A(n6030), .B(n1149), .Z(out[1166]) );
  IV U7472 ( .A(n5782), .Z(n1149) );
  XOR U7473 ( .A(n6031), .B(n2197), .Z(n5782) );
  XNOR U7474 ( .A(n6032), .B(n6033), .Z(n2197) );
  NOR U7475 ( .A(n6034), .B(n5781), .Z(n6030) );
  XOR U7476 ( .A(n6035), .B(n1152), .Z(out[1165]) );
  XOR U7477 ( .A(n6036), .B(n3820), .Z(n1152) );
  XOR U7478 ( .A(n6037), .B(n6038), .Z(n3820) );
  NOR U7479 ( .A(n6039), .B(n5788), .Z(n6035) );
  XNOR U7480 ( .A(n6040), .B(n1156), .Z(out[1164]) );
  IV U7481 ( .A(n5791), .Z(n1156) );
  ANDN U7482 ( .B(n6044), .A(n5790), .Z(n6040) );
  XNOR U7483 ( .A(n6045), .B(n1160), .Z(out[1163]) );
  XOR U7484 ( .A(n6046), .B(n1977), .Z(n1160) );
  IV U7485 ( .A(n3834), .Z(n1977) );
  ANDN U7486 ( .B(n6049), .A(n6050), .Z(n6045) );
  XOR U7487 ( .A(n6051), .B(n1164), .Z(out[1162]) );
  XOR U7488 ( .A(n6052), .B(n1980), .Z(n1164) );
  IV U7489 ( .A(n5584), .Z(n1980) );
  NOR U7490 ( .A(n6055), .B(n5795), .Z(n6051) );
  XNOR U7491 ( .A(n6056), .B(n1173), .Z(out[1161]) );
  XOR U7492 ( .A(n6057), .B(n1983), .Z(n1173) );
  IV U7493 ( .A(n3843), .Z(n1983) );
  ANDN U7494 ( .B(n6060), .A(n5797), .Z(n6056) );
  XNOR U7495 ( .A(n6061), .B(n1177), .Z(out[1160]) );
  XOR U7496 ( .A(n6062), .B(n1986), .Z(n1177) );
  XNOR U7497 ( .A(n6063), .B(n6064), .Z(n1986) );
  ANDN U7498 ( .B(n6065), .A(n6066), .Z(n6061) );
  XNOR U7499 ( .A(n6067), .B(n4150), .Z(out[115]) );
  XOR U7500 ( .A(n6068), .B(n2470), .Z(n4150) );
  ANDN U7501 ( .B(n3119), .A(n3117), .Z(n6067) );
  XOR U7502 ( .A(n6069), .B(n3158), .Z(n3117) );
  IV U7503 ( .A(n2308), .Z(n3158) );
  XNOR U7504 ( .A(n6070), .B(n2243), .Z(n3119) );
  XNOR U7505 ( .A(n6071), .B(n1181), .Z(out[1159]) );
  IV U7506 ( .A(n5802), .Z(n1181) );
  XOR U7507 ( .A(n6072), .B(n1989), .Z(n5802) );
  XOR U7508 ( .A(n6073), .B(n6074), .Z(n1989) );
  ANDN U7509 ( .B(n6075), .A(n5801), .Z(n6071) );
  XNOR U7510 ( .A(n6076), .B(n1185), .Z(out[1158]) );
  IV U7511 ( .A(n5805), .Z(n1185) );
  XNOR U7512 ( .A(n6077), .B(n1992), .Z(n5805) );
  XNOR U7513 ( .A(n6078), .B(n6079), .Z(n1992) );
  NOR U7514 ( .A(n6080), .B(n5804), .Z(n6076) );
  XNOR U7515 ( .A(n6081), .B(n1188), .Z(out[1157]) );
  IV U7516 ( .A(n5808), .Z(n1188) );
  XOR U7517 ( .A(n6082), .B(n1995), .Z(n5808) );
  XNOR U7518 ( .A(n6083), .B(n6084), .Z(n1995) );
  NOR U7519 ( .A(n6085), .B(n5807), .Z(n6081) );
  XNOR U7520 ( .A(n6086), .B(n1192), .Z(out[1156]) );
  IV U7521 ( .A(n5811), .Z(n1192) );
  XOR U7522 ( .A(n6087), .B(n1998), .Z(n5811) );
  XNOR U7523 ( .A(n6088), .B(n6089), .Z(n1998) );
  ANDN U7524 ( .B(n6090), .A(n5810), .Z(n6086) );
  XNOR U7525 ( .A(n6091), .B(n1196), .Z(out[1155]) );
  IV U7526 ( .A(n5819), .Z(n1196) );
  XOR U7527 ( .A(n6092), .B(n2005), .Z(n5819) );
  XNOR U7528 ( .A(n6093), .B(n6094), .Z(n2005) );
  ANDN U7529 ( .B(n6095), .A(n5818), .Z(n6091) );
  XOR U7530 ( .A(n6096), .B(n1200), .Z(out[1154]) );
  XOR U7531 ( .A(n6097), .B(n2009), .Z(n1200) );
  XNOR U7532 ( .A(n6098), .B(n6099), .Z(n2009) );
  ANDN U7533 ( .B(n6100), .A(n5821), .Z(n6096) );
  XOR U7534 ( .A(n6101), .B(n1204), .Z(out[1153]) );
  XOR U7535 ( .A(n6102), .B(n2012), .Z(n1204) );
  XNOR U7536 ( .A(n6103), .B(n6104), .Z(n2012) );
  NOR U7537 ( .A(n6105), .B(n5823), .Z(n6101) );
  XNOR U7538 ( .A(n6106), .B(n1208), .Z(out[1152]) );
  XOR U7539 ( .A(n6107), .B(n2015), .Z(n1208) );
  XNOR U7540 ( .A(n6108), .B(n6109), .Z(n2015) );
  ANDN U7541 ( .B(n6110), .A(n5825), .Z(n6106) );
  XOR U7542 ( .A(n6111), .B(n5609), .Z(out[1151]) );
  XNOR U7543 ( .A(n6112), .B(n3762), .Z(n5609) );
  IV U7544 ( .A(n2572), .Z(n3762) );
  ANDN U7545 ( .B(n6113), .A(n5827), .Z(n6111) );
  XOR U7546 ( .A(n6114), .B(n5613), .Z(out[1150]) );
  XOR U7547 ( .A(n6115), .B(n2579), .Z(n5613) );
  ANDN U7548 ( .B(n5829), .A(n6116), .Z(n6114) );
  XOR U7549 ( .A(n6117), .B(n4153), .Z(out[114]) );
  XOR U7550 ( .A(n6118), .B(n5564), .Z(n4153) );
  ANDN U7551 ( .B(n3146), .A(n3147), .Z(n6117) );
  XNOR U7552 ( .A(n6119), .B(n2250), .Z(n3147) );
  XOR U7553 ( .A(n6120), .B(n3163), .Z(n3146) );
  IV U7554 ( .A(n2319), .Z(n3163) );
  XOR U7555 ( .A(n6121), .B(n5617), .Z(out[1149]) );
  XNOR U7556 ( .A(n5324), .B(n6122), .Z(n5617) );
  XNOR U7557 ( .A(n6123), .B(n6124), .Z(n5324) );
  ANDN U7558 ( .B(n6125), .A(n5831), .Z(n6121) );
  XNOR U7559 ( .A(n6126), .B(n5834), .Z(out[1148]) );
  XOR U7560 ( .A(n4387), .B(n6127), .Z(n5834) );
  XNOR U7561 ( .A(n6128), .B(n6129), .Z(n4387) );
  ANDN U7562 ( .B(n6130), .A(n5833), .Z(n6126) );
  XOR U7563 ( .A(n6131), .B(n5625), .Z(out[1147]) );
  XNOR U7564 ( .A(n5333), .B(n6132), .Z(n5625) );
  XNOR U7565 ( .A(n6133), .B(n6134), .Z(n5333) );
  ANDN U7566 ( .B(n6135), .A(n5836), .Z(n6131) );
  XOR U7567 ( .A(n6136), .B(n5629), .Z(out[1146]) );
  XNOR U7568 ( .A(n6137), .B(n2611), .Z(n5629) );
  XNOR U7569 ( .A(n6138), .B(n6139), .Z(n2611) );
  XOR U7570 ( .A(n6141), .B(n5633), .Z(out[1145]) );
  XNOR U7571 ( .A(n6142), .B(n3789), .Z(n5633) );
  IV U7572 ( .A(n2618), .Z(n3789) );
  XOR U7573 ( .A(n6143), .B(n6144), .Z(n2618) );
  ANDN U7574 ( .B(n6145), .A(n5844), .Z(n6141) );
  XNOR U7575 ( .A(n6146), .B(n5638), .Z(out[1144]) );
  IV U7576 ( .A(n5847), .Z(n5638) );
  XOR U7577 ( .A(n6147), .B(n2625), .Z(n5847) );
  IV U7578 ( .A(n3795), .Z(n2625) );
  XOR U7579 ( .A(n6148), .B(n6149), .Z(n3795) );
  NOR U7580 ( .A(n6150), .B(n5846), .Z(n6146) );
  XOR U7581 ( .A(n6151), .B(n5641), .Z(out[1143]) );
  XNOR U7582 ( .A(n6152), .B(n2632), .Z(n5641) );
  XOR U7583 ( .A(n6153), .B(n6154), .Z(n2632) );
  ANDN U7584 ( .B(n6155), .A(n5849), .Z(n6151) );
  XOR U7585 ( .A(n6156), .B(n5645), .Z(out[1142]) );
  XOR U7586 ( .A(n6157), .B(n2639), .Z(n5645) );
  XNOR U7587 ( .A(n6158), .B(n6159), .Z(n2639) );
  ANDN U7588 ( .B(n6160), .A(n5851), .Z(n6156) );
  XOR U7589 ( .A(n6161), .B(n5653), .Z(out[1141]) );
  XOR U7590 ( .A(n6162), .B(n3811), .Z(n5653) );
  IV U7591 ( .A(n2646), .Z(n3811) );
  XOR U7592 ( .A(n6163), .B(n6164), .Z(n2646) );
  NOR U7593 ( .A(n6165), .B(n5853), .Z(n6161) );
  XOR U7594 ( .A(n6166), .B(n5657), .Z(out[1140]) );
  XNOR U7595 ( .A(n6167), .B(n2653), .Z(n5657) );
  XNOR U7596 ( .A(n6168), .B(n6169), .Z(n2653) );
  ANDN U7597 ( .B(n6170), .A(n5855), .Z(n6166) );
  IV U7598 ( .A(n6171), .Z(n5855) );
  XOR U7599 ( .A(n6172), .B(n4156), .Z(out[113]) );
  XNOR U7600 ( .A(n6173), .B(n2484), .Z(n4156) );
  AND U7601 ( .A(n3187), .B(n3189), .Z(n6172) );
  XNOR U7602 ( .A(n6174), .B(n2257), .Z(n3189) );
  XOR U7603 ( .A(n6175), .B(n2324), .Z(n3187) );
  IV U7604 ( .A(n5476), .Z(n2324) );
  XOR U7605 ( .A(n6176), .B(n5661), .Z(out[1139]) );
  XNOR U7606 ( .A(n6177), .B(n3822), .Z(n5661) );
  IV U7607 ( .A(n2660), .Z(n3822) );
  XOR U7608 ( .A(n6178), .B(n6179), .Z(n2660) );
  ANDN U7609 ( .B(n6180), .A(n5857), .Z(n6176) );
  XOR U7610 ( .A(n6181), .B(n5665), .Z(out[1138]) );
  XOR U7611 ( .A(n6182), .B(n2667), .Z(n5665) );
  IV U7612 ( .A(n3828), .Z(n2667) );
  XOR U7613 ( .A(n6183), .B(n6184), .Z(n3828) );
  XOR U7614 ( .A(n6186), .B(n5669), .Z(out[1137]) );
  XOR U7615 ( .A(n6187), .B(n2674), .Z(n5669) );
  XNOR U7616 ( .A(n6188), .B(n6189), .Z(n2674) );
  NOR U7617 ( .A(n6190), .B(n5861), .Z(n6186) );
  XNOR U7618 ( .A(n6191), .B(n5674), .Z(out[1136]) );
  IV U7619 ( .A(n5864), .Z(n5674) );
  XOR U7620 ( .A(n6192), .B(n4762), .Z(n5864) );
  IV U7621 ( .A(n2207), .Z(n4762) );
  XOR U7622 ( .A(n6193), .B(n6194), .Z(n2207) );
  NOR U7623 ( .A(n6195), .B(n5863), .Z(n6191) );
  XOR U7624 ( .A(n6196), .B(n5677), .Z(out[1135]) );
  XNOR U7625 ( .A(n6197), .B(n2214), .Z(n5677) );
  XOR U7626 ( .A(n6198), .B(n6199), .Z(n2214) );
  NOR U7627 ( .A(n6200), .B(n5874), .Z(n6196) );
  XOR U7628 ( .A(n6201), .B(n5681), .Z(out[1134]) );
  XNOR U7629 ( .A(n6202), .B(n2221), .Z(n5681) );
  XOR U7630 ( .A(n6203), .B(n6204), .Z(n2221) );
  NOR U7631 ( .A(n6205), .B(n5876), .Z(n6201) );
  XOR U7632 ( .A(n6206), .B(n5685), .Z(out[1133]) );
  XOR U7633 ( .A(n6207), .B(n4843), .Z(n5685) );
  XOR U7634 ( .A(n6208), .B(n6209), .Z(n4843) );
  NOR U7635 ( .A(n6210), .B(n5878), .Z(n6206) );
  XOR U7636 ( .A(n6211), .B(n5689), .Z(out[1132]) );
  XOR U7637 ( .A(n6212), .B(n2241), .Z(n5689) );
  XOR U7638 ( .A(n6213), .B(n6214), .Z(n2241) );
  NOR U7639 ( .A(n6215), .B(n5880), .Z(n6211) );
  XOR U7640 ( .A(n6216), .B(n5698), .Z(out[1131]) );
  XOR U7641 ( .A(n6217), .B(n2248), .Z(n5698) );
  XOR U7642 ( .A(n6218), .B(n6219), .Z(n2248) );
  ANDN U7643 ( .B(n6220), .A(n5882), .Z(n6216) );
  XOR U7644 ( .A(n6221), .B(n5702), .Z(out[1130]) );
  XOR U7645 ( .A(n6222), .B(n5419), .Z(n5702) );
  XOR U7646 ( .A(n6223), .B(n6224), .Z(n5419) );
  ANDN U7647 ( .B(n6225), .A(n6226), .Z(n6221) );
  XNOR U7648 ( .A(n6227), .B(n4160), .Z(out[112]) );
  XNOR U7649 ( .A(n6228), .B(n2491), .Z(n4160) );
  ANDN U7650 ( .B(n3226), .A(n3228), .Z(n6227) );
  XNOR U7651 ( .A(n6229), .B(n2266), .Z(n3228) );
  XNOR U7652 ( .A(n6230), .B(n5481), .Z(n3226) );
  XOR U7653 ( .A(n6231), .B(n5706), .Z(out[1129]) );
  XOR U7654 ( .A(n6232), .B(n3870), .Z(n5706) );
  XOR U7655 ( .A(n6233), .B(n6234), .Z(n3870) );
  ANDN U7656 ( .B(n6235), .A(n5886), .Z(n6231) );
  XOR U7657 ( .A(n6236), .B(n5710), .Z(out[1128]) );
  XNOR U7658 ( .A(n6237), .B(n5023), .Z(n5710) );
  XOR U7659 ( .A(n6238), .B(n6239), .Z(n5023) );
  XNOR U7660 ( .A(n6241), .B(n5714), .Z(out[1127]) );
  XOR U7661 ( .A(n6242), .B(n3881), .Z(n5714) );
  XOR U7662 ( .A(n6243), .B(n6244), .Z(n3881) );
  NOR U7663 ( .A(n5893), .B(n1039), .Z(n6241) );
  XOR U7664 ( .A(n6245), .B(n5716), .Z(out[1126]) );
  XNOR U7665 ( .A(n6246), .B(n2283), .Z(n5716) );
  IV U7666 ( .A(n5096), .Z(n2283) );
  XOR U7667 ( .A(n6247), .B(n6248), .Z(n5096) );
  IV U7668 ( .A(n6249), .Z(n5898) );
  XOR U7669 ( .A(n6250), .B(n5718), .Z(out[1125]) );
  XNOR U7670 ( .A(n6251), .B(n5127), .Z(n5718) );
  XOR U7671 ( .A(n6252), .B(n6253), .Z(n5127) );
  XOR U7672 ( .A(n6254), .B(n5720), .Z(out[1124]) );
  XOR U7673 ( .A(n6255), .B(n2297), .Z(n5720) );
  XNOR U7674 ( .A(n6256), .B(n6257), .Z(n2297) );
  XOR U7675 ( .A(n6258), .B(n5722), .Z(out[1123]) );
  XNOR U7676 ( .A(n6259), .B(n2304), .Z(n5722) );
  IV U7677 ( .A(n3899), .Z(n2304) );
  XNOR U7678 ( .A(n6260), .B(n6261), .Z(n3899) );
  XNOR U7679 ( .A(n6262), .B(n5725), .Z(out[1122]) );
  XOR U7680 ( .A(n6263), .B(n5452), .Z(n5725) );
  XNOR U7681 ( .A(n6264), .B(n6265), .Z(n5452) );
  NOR U7682 ( .A(n5923), .B(n1059), .Z(n6262) );
  XNOR U7683 ( .A(n6266), .B(n5929), .Z(out[1121]) );
  XOR U7684 ( .A(n6267), .B(n3908), .Z(n5929) );
  XNOR U7685 ( .A(n6268), .B(n6269), .Z(n3908) );
  NOR U7686 ( .A(n1063), .B(n5928), .Z(n6266) );
  XOR U7687 ( .A(n6270), .B(n5735), .Z(out[1120]) );
  XOR U7688 ( .A(n6271), .B(n5466), .Z(n5735) );
  XNOR U7689 ( .A(n6272), .B(n6273), .Z(n5466) );
  NOR U7690 ( .A(n5934), .B(n1067), .Z(n6270) );
  XOR U7691 ( .A(n6274), .B(n4165), .Z(out[111]) );
  XNOR U7692 ( .A(n6275), .B(n2498), .Z(n4165) );
  AND U7693 ( .A(n3265), .B(n3267), .Z(n6274) );
  XNOR U7694 ( .A(n6276), .B(n2271), .Z(n3267) );
  XOR U7695 ( .A(n6277), .B(n3173), .Z(n3265) );
  XOR U7696 ( .A(n6278), .B(n5737), .Z(out[1119]) );
  XOR U7697 ( .A(n6279), .B(n5471), .Z(n5737) );
  XNOR U7698 ( .A(n6280), .B(n6281), .Z(n5471) );
  ANDN U7699 ( .B(n5939), .A(n1071), .Z(n6278) );
  XOR U7700 ( .A(n6282), .B(n5740), .Z(out[1118]) );
  XOR U7701 ( .A(n6283), .B(n2343), .Z(n5740) );
  IV U7702 ( .A(n3606), .Z(n2343) );
  XNOR U7703 ( .A(n6284), .B(n6285), .Z(n3606) );
  NOR U7704 ( .A(n5944), .B(n1075), .Z(n6282) );
  XOR U7705 ( .A(n6286), .B(n5742), .Z(out[1117]) );
  XNOR U7706 ( .A(n6287), .B(n5412), .Z(n5742) );
  XNOR U7707 ( .A(n6288), .B(n6289), .Z(n5412) );
  NOR U7708 ( .A(n6290), .B(n1083), .Z(n6286) );
  XOR U7709 ( .A(n6291), .B(n5744), .Z(out[1116]) );
  XOR U7710 ( .A(n6292), .B(n2357), .Z(n5744) );
  XOR U7711 ( .A(n6293), .B(n6294), .Z(n2357) );
  ANDN U7712 ( .B(n1087), .A(n5954), .Z(n6291) );
  XOR U7713 ( .A(n6295), .B(n5746), .Z(out[1115]) );
  XOR U7714 ( .A(n6296), .B(n3620), .Z(n5746) );
  XOR U7715 ( .A(n6297), .B(n6298), .Z(n3620) );
  NOR U7716 ( .A(n5964), .B(n1091), .Z(n6295) );
  XOR U7717 ( .A(n6299), .B(n5748), .Z(out[1114]) );
  XOR U7718 ( .A(n6300), .B(n5560), .Z(n5748) );
  XOR U7719 ( .A(n6301), .B(n6302), .Z(n5560) );
  NOR U7720 ( .A(n1095), .B(n5969), .Z(n6299) );
  XOR U7721 ( .A(n6303), .B(n5751), .Z(out[1113]) );
  XOR U7722 ( .A(n6304), .B(n2378), .Z(n5751) );
  IV U7723 ( .A(n3634), .Z(n2378) );
  XOR U7724 ( .A(n6305), .B(n6306), .Z(n3634) );
  ANDN U7725 ( .B(n5974), .A(n1099), .Z(n6303) );
  XNOR U7726 ( .A(n6307), .B(n5753), .Z(out[1112]) );
  XOR U7727 ( .A(n6308), .B(n3639), .Z(n5753) );
  XOR U7728 ( .A(n6309), .B(n6310), .Z(n3639) );
  ANDN U7729 ( .B(n5979), .A(n1103), .Z(n6307) );
  XOR U7730 ( .A(n6311), .B(n5759), .Z(out[1111]) );
  XNOR U7731 ( .A(n6312), .B(n2396), .Z(n5759) );
  XOR U7732 ( .A(n6313), .B(n6314), .Z(n2396) );
  ANDN U7733 ( .B(n5984), .A(n1107), .Z(n6311) );
  XOR U7734 ( .A(n6315), .B(n5762), .Z(out[1110]) );
  XNOR U7735 ( .A(n6316), .B(n2403), .Z(n5762) );
  XNOR U7736 ( .A(n6317), .B(n6318), .Z(n2403) );
  XOR U7737 ( .A(n6319), .B(n4168), .Z(out[110]) );
  XNOR U7738 ( .A(n6320), .B(n2505), .Z(n4168) );
  ANDN U7739 ( .B(n3307), .A(n3308), .Z(n6319) );
  XOR U7740 ( .A(n6321), .B(n2278), .Z(n3308) );
  XOR U7741 ( .A(n6322), .B(n2345), .Z(n3307) );
  XOR U7742 ( .A(n6323), .B(n5764), .Z(out[1109]) );
  XNOR U7743 ( .A(n6324), .B(n2410), .Z(n5764) );
  XOR U7744 ( .A(n6325), .B(n6326), .Z(n2410) );
  NOR U7745 ( .A(n6327), .B(n1115), .Z(n6323) );
  XOR U7746 ( .A(n6328), .B(n5767), .Z(out[1108]) );
  XNOR U7747 ( .A(n6329), .B(n2417), .Z(n5767) );
  IV U7748 ( .A(n3657), .Z(n2417) );
  XOR U7749 ( .A(n6330), .B(n6331), .Z(n3657) );
  ANDN U7750 ( .B(n5999), .A(n1119), .Z(n6328) );
  XOR U7751 ( .A(n6332), .B(n5769), .Z(out[1107]) );
  XOR U7752 ( .A(n6333), .B(n5814), .Z(n5769) );
  XOR U7753 ( .A(n6334), .B(n6335), .Z(n5814) );
  NOR U7754 ( .A(n1127), .B(n6004), .Z(n6332) );
  XOR U7755 ( .A(n6336), .B(n5772), .Z(out[1106]) );
  XOR U7756 ( .A(n6337), .B(n2431), .Z(n5772) );
  XNOR U7757 ( .A(n6338), .B(n6339), .Z(n2431) );
  XOR U7758 ( .A(n6340), .B(n5774), .Z(out[1105]) );
  XOR U7759 ( .A(n6341), .B(n2438), .Z(n5774) );
  XOR U7760 ( .A(n6342), .B(n6343), .Z(n2438) );
  NOR U7761 ( .A(n1135), .B(n6019), .Z(n6340) );
  XOR U7762 ( .A(n6344), .B(n5777), .Z(out[1104]) );
  XOR U7763 ( .A(n6345), .B(n2445), .Z(n5777) );
  XOR U7764 ( .A(n6346), .B(n6347), .Z(n2445) );
  ANDN U7765 ( .B(n6024), .A(n1139), .Z(n6344) );
  IV U7766 ( .A(n6348), .Z(n1139) );
  XOR U7767 ( .A(n6349), .B(n5779), .Z(out[1103]) );
  XNOR U7768 ( .A(n6350), .B(n3683), .Z(n5779) );
  XOR U7769 ( .A(n6351), .B(n6352), .Z(n3683) );
  NOR U7770 ( .A(n1143), .B(n6029), .Z(n6349) );
  XOR U7771 ( .A(n6353), .B(n5781), .Z(out[1102]) );
  XNOR U7772 ( .A(n6354), .B(n2463), .Z(n5781) );
  XNOR U7773 ( .A(n6355), .B(n6356), .Z(n2463) );
  NOR U7774 ( .A(n6357), .B(n1147), .Z(n6353) );
  XOR U7775 ( .A(n6358), .B(n5788), .Z(out[1101]) );
  XOR U7776 ( .A(n6359), .B(n3693), .Z(n5788) );
  IV U7777 ( .A(n2470), .Z(n3693) );
  XOR U7778 ( .A(n6360), .B(n6361), .Z(n2470) );
  NOR U7779 ( .A(n6362), .B(n1151), .Z(n6358) );
  XOR U7780 ( .A(n6363), .B(n5790), .Z(out[1100]) );
  XNOR U7781 ( .A(n6364), .B(n2477), .Z(n5790) );
  IV U7782 ( .A(n5564), .Z(n2477) );
  XOR U7783 ( .A(n6365), .B(n6366), .Z(n5564) );
  XOR U7784 ( .A(n6367), .B(n2038), .Z(out[10]) );
  XOR U7785 ( .A(n6368), .B(n3322), .Z(n2038) );
  IV U7786 ( .A(n2615), .Z(n3322) );
  NOR U7787 ( .A(n4069), .B(n2037), .Z(n6367) );
  XNOR U7788 ( .A(n2545), .B(n6369), .Z(n2037) );
  IV U7789 ( .A(n3517), .Z(n2545) );
  XNOR U7790 ( .A(n6370), .B(n1758), .Z(n4069) );
  XOR U7791 ( .A(n6371), .B(n4171), .Z(out[109]) );
  XOR U7792 ( .A(n6372), .B(n2512), .Z(n4171) );
  ANDN U7793 ( .B(n3348), .A(n3350), .Z(n6371) );
  XNOR U7794 ( .A(n6373), .B(n2285), .Z(n3350) );
  XOR U7795 ( .A(n6374), .B(n2352), .Z(n3348) );
  XNOR U7796 ( .A(n6375), .B(n5793), .Z(out[1099]) );
  IV U7797 ( .A(n6050), .Z(n5793) );
  XNOR U7798 ( .A(n6376), .B(n2484), .Z(n6050) );
  XNOR U7799 ( .A(n6377), .B(n6378), .Z(n2484) );
  ANDN U7800 ( .B(n1159), .A(n6049), .Z(n6375) );
  XOR U7801 ( .A(n6379), .B(n5795), .Z(out[1098]) );
  XOR U7802 ( .A(n6380), .B(n2491), .Z(n5795) );
  XNOR U7803 ( .A(n6381), .B(n6382), .Z(n2491) );
  ANDN U7804 ( .B(n6055), .A(n1163), .Z(n6379) );
  XOR U7805 ( .A(n6383), .B(n5797), .Z(out[1097]) );
  XNOR U7806 ( .A(n6384), .B(n2498), .Z(n5797) );
  XOR U7807 ( .A(n6385), .B(n6386), .Z(n2498) );
  NOR U7808 ( .A(n6060), .B(n1171), .Z(n6383) );
  XNOR U7809 ( .A(n6387), .B(n5799), .Z(out[1096]) );
  IV U7810 ( .A(n6066), .Z(n5799) );
  XNOR U7811 ( .A(n6388), .B(n2505), .Z(n6066) );
  XNOR U7812 ( .A(n6389), .B(n6390), .Z(n2505) );
  ANDN U7813 ( .B(n1175), .A(n6065), .Z(n6387) );
  XOR U7814 ( .A(n6391), .B(n5801), .Z(out[1095]) );
  XOR U7815 ( .A(n6392), .B(n2512), .Z(n5801) );
  XNOR U7816 ( .A(n6393), .B(n6394), .Z(n2512) );
  NOR U7817 ( .A(n1179), .B(n6075), .Z(n6391) );
  XOR U7818 ( .A(n6395), .B(n5804), .Z(out[1094]) );
  XNOR U7819 ( .A(n6396), .B(n3731), .Z(n5804) );
  IV U7820 ( .A(n2519), .Z(n3731) );
  NOR U7821 ( .A(n6397), .B(n1183), .Z(n6395) );
  XOR U7822 ( .A(n6398), .B(n5807), .Z(out[1093]) );
  XOR U7823 ( .A(n6399), .B(n2526), .Z(n5807) );
  IV U7824 ( .A(n6400), .Z(n2526) );
  ANDN U7825 ( .B(n6085), .A(n6401), .Z(n6398) );
  XOR U7826 ( .A(n6402), .B(n5810), .Z(out[1092]) );
  XNOR U7827 ( .A(n6403), .B(n2537), .Z(n5810) );
  NOR U7828 ( .A(n1191), .B(n6090), .Z(n6402) );
  IV U7829 ( .A(n6404), .Z(n1191) );
  XOR U7830 ( .A(n6405), .B(n5818), .Z(out[1091]) );
  XOR U7831 ( .A(n6406), .B(n2544), .Z(n5818) );
  NOR U7832 ( .A(n6407), .B(n6095), .Z(n6405) );
  XOR U7833 ( .A(n6408), .B(n5821), .Z(out[1090]) );
  XNOR U7834 ( .A(n6409), .B(n2551), .Z(n5821) );
  NOR U7835 ( .A(n6100), .B(n1199), .Z(n6408) );
  XOR U7836 ( .A(n6410), .B(n4174), .Z(out[108]) );
  XOR U7837 ( .A(n6411), .B(n2519), .Z(n4174) );
  XOR U7838 ( .A(n6412), .B(n6413), .Z(n2519) );
  ANDN U7839 ( .B(n3392), .A(n3393), .Z(n6410) );
  XNOR U7840 ( .A(n6414), .B(n2292), .Z(n3393) );
  XOR U7841 ( .A(n6415), .B(n2359), .Z(n3392) );
  XOR U7842 ( .A(n6416), .B(n5823), .Z(out[1089]) );
  XOR U7843 ( .A(n6417), .B(n2558), .Z(n5823) );
  NOR U7844 ( .A(n6418), .B(n1203), .Z(n6416) );
  XOR U7845 ( .A(n6419), .B(n5825), .Z(out[1088]) );
  XNOR U7846 ( .A(n6420), .B(n3757), .Z(n5825) );
  IV U7847 ( .A(n2565), .Z(n3757) );
  NOR U7848 ( .A(n1207), .B(n6110), .Z(n6419) );
  IV U7849 ( .A(n6421), .Z(n1207) );
  XOR U7850 ( .A(n6422), .B(n5827), .Z(out[1087]) );
  XOR U7851 ( .A(n6423), .B(n2539), .Z(n5827) );
  XNOR U7852 ( .A(n5891), .B(n6424), .Z(n2539) );
  XOR U7853 ( .A(n6425), .B(n6426), .Z(n5891) );
  XOR U7854 ( .A(n6324), .B(n2409), .Z(n6426) );
  XNOR U7855 ( .A(n6427), .B(n6428), .Z(n2409) );
  NOR U7856 ( .A(n6429), .B(n6430), .Z(n6427) );
  XOR U7857 ( .A(n6431), .B(n6432), .Z(n6324) );
  NOR U7858 ( .A(n6433), .B(n6434), .Z(n6431) );
  XOR U7859 ( .A(n3652), .B(n6435), .Z(n6425) );
  XOR U7860 ( .A(n5755), .B(n5523), .Z(n6435) );
  XNOR U7861 ( .A(n6436), .B(n6437), .Z(n5523) );
  NOR U7862 ( .A(n6438), .B(n6439), .Z(n6436) );
  XNOR U7863 ( .A(n6440), .B(n6441), .Z(n5755) );
  XNOR U7864 ( .A(n6444), .B(n6445), .Z(n3652) );
  ANDN U7865 ( .B(n6446), .A(n6447), .Z(n6444) );
  ANDN U7866 ( .B(n5608), .A(n6113), .Z(n6422) );
  XNOR U7867 ( .A(n6448), .B(n5829), .Z(out[1086]) );
  XNOR U7868 ( .A(n6449), .B(n2548), .Z(n5829) );
  XNOR U7869 ( .A(n5896), .B(n6450), .Z(n2548) );
  XOR U7870 ( .A(n6451), .B(n6452), .Z(n5896) );
  XOR U7871 ( .A(n6329), .B(n2416), .Z(n6452) );
  XNOR U7872 ( .A(n6453), .B(n6454), .Z(n2416) );
  XNOR U7873 ( .A(n6457), .B(n6458), .Z(n6329) );
  ANDN U7874 ( .B(n6459), .A(n6460), .Z(n6457) );
  XOR U7875 ( .A(n3656), .B(n6461), .Z(n6451) );
  XNOR U7876 ( .A(n5784), .B(n5526), .Z(n6461) );
  XOR U7877 ( .A(n6462), .B(n6463), .Z(n5526) );
  ANDN U7878 ( .B(n6464), .A(n6465), .Z(n6462) );
  XOR U7879 ( .A(n6466), .B(n6467), .Z(n5784) );
  ANDN U7880 ( .B(n6468), .A(n6469), .Z(n6466) );
  NOR U7881 ( .A(n6472), .B(n6473), .Z(n6470) );
  NOR U7882 ( .A(n6474), .B(n5612), .Z(n6448) );
  XOR U7883 ( .A(n6475), .B(n5831), .Z(out[1085]) );
  XOR U7884 ( .A(n6476), .B(n2553), .Z(n5831) );
  XNOR U7885 ( .A(n5906), .B(n6477), .Z(n2553) );
  XOR U7886 ( .A(n6478), .B(n6479), .Z(n5906) );
  XOR U7887 ( .A(n6333), .B(n2423), .Z(n6479) );
  XNOR U7888 ( .A(n6480), .B(n6481), .Z(n2423) );
  XOR U7889 ( .A(n6484), .B(n6485), .Z(n6333) );
  ANDN U7890 ( .B(n6486), .A(n6487), .Z(n6484) );
  XOR U7891 ( .A(n3660), .B(n6488), .Z(n6478) );
  XNOR U7892 ( .A(n5813), .B(n5531), .Z(n6488) );
  XNOR U7893 ( .A(n6489), .B(n6490), .Z(n5531) );
  ANDN U7894 ( .B(n6491), .A(n6492), .Z(n6489) );
  XNOR U7895 ( .A(n6493), .B(n6494), .Z(n5813) );
  ANDN U7896 ( .B(n6495), .A(n6496), .Z(n6493) );
  XNOR U7897 ( .A(n6497), .B(n6498), .Z(n3660) );
  ANDN U7898 ( .B(n5616), .A(n6125), .Z(n6475) );
  XOR U7899 ( .A(n6501), .B(n5833), .Z(out[1084]) );
  XNOR U7900 ( .A(n6502), .B(n2562), .Z(n5833) );
  IV U7901 ( .A(n4913), .Z(n2562) );
  XNOR U7902 ( .A(n5911), .B(n6503), .Z(n4913) );
  XOR U7903 ( .A(n6504), .B(n6505), .Z(n5911) );
  XOR U7904 ( .A(n6337), .B(n2430), .Z(n6505) );
  XOR U7905 ( .A(n6506), .B(n6507), .Z(n2430) );
  XOR U7906 ( .A(n6510), .B(n6511), .Z(n6337) );
  NOR U7907 ( .A(n6512), .B(n6513), .Z(n6510) );
  XOR U7908 ( .A(n3664), .B(n6514), .Z(n6504) );
  XNOR U7909 ( .A(n5840), .B(n5535), .Z(n6514) );
  XNOR U7910 ( .A(n6515), .B(n6516), .Z(n5535) );
  XOR U7911 ( .A(n6517), .B(n4694), .Z(n6516) );
  NOR U7912 ( .A(n6518), .B(n6519), .Z(n6517) );
  XNOR U7913 ( .A(n6520), .B(n6521), .Z(n5840) );
  ANDN U7914 ( .B(n6522), .A(n6523), .Z(n6520) );
  XOR U7915 ( .A(n6524), .B(n6525), .Z(n3664) );
  ANDN U7916 ( .B(n6526), .A(n6527), .Z(n6524) );
  NOR U7917 ( .A(n6130), .B(n5620), .Z(n6501) );
  XOR U7918 ( .A(n6528), .B(n5836), .Z(out[1083]) );
  XOR U7919 ( .A(n6529), .B(n2569), .Z(n5836) );
  XNOR U7920 ( .A(n5916), .B(n6530), .Z(n2569) );
  XOR U7921 ( .A(n6531), .B(n6532), .Z(n5916) );
  XOR U7922 ( .A(n6341), .B(n2437), .Z(n6532) );
  XNOR U7923 ( .A(n6533), .B(n6534), .Z(n2437) );
  XNOR U7924 ( .A(n6537), .B(n6538), .Z(n6341) );
  ANDN U7925 ( .B(n6539), .A(n6540), .Z(n6537) );
  XOR U7926 ( .A(n3668), .B(n6541), .Z(n6531) );
  XNOR U7927 ( .A(n5870), .B(n5538), .Z(n6541) );
  XNOR U7928 ( .A(n6542), .B(n6543), .Z(n5538) );
  ANDN U7929 ( .B(n6544), .A(n6545), .Z(n6542) );
  XOR U7930 ( .A(n6546), .B(n6547), .Z(n5870) );
  NOR U7931 ( .A(n6548), .B(n6549), .Z(n6546) );
  XNOR U7932 ( .A(n6550), .B(n6551), .Z(n3668) );
  ANDN U7933 ( .B(n6552), .A(n6553), .Z(n6550) );
  ANDN U7934 ( .B(n5624), .A(n6135), .Z(n6528) );
  XNOR U7935 ( .A(n6554), .B(n5838), .Z(out[1082]) );
  XOR U7936 ( .A(n6555), .B(n4988), .Z(n5838) );
  XNOR U7937 ( .A(n5921), .B(n6556), .Z(n4988) );
  XOR U7938 ( .A(n6557), .B(n6558), .Z(n5921) );
  XOR U7939 ( .A(n6345), .B(n2444), .Z(n6558) );
  XOR U7940 ( .A(n6559), .B(n6560), .Z(n2444) );
  NOR U7941 ( .A(n6561), .B(n6562), .Z(n6559) );
  XNOR U7942 ( .A(n6563), .B(n6564), .Z(n6345) );
  NOR U7943 ( .A(n6565), .B(n6566), .Z(n6563) );
  XOR U7944 ( .A(n3678), .B(n6567), .Z(n6557) );
  XNOR U7945 ( .A(n5900), .B(n5544), .Z(n6567) );
  XNOR U7946 ( .A(n6568), .B(n6569), .Z(n5544) );
  ANDN U7947 ( .B(n6570), .A(n6571), .Z(n6568) );
  XNOR U7948 ( .A(n6572), .B(n6573), .Z(n5900) );
  NOR U7949 ( .A(n6574), .B(n6575), .Z(n6572) );
  XOR U7950 ( .A(n6576), .B(n6577), .Z(n3678) );
  ANDN U7951 ( .B(n6578), .A(n6579), .Z(n6576) );
  ANDN U7952 ( .B(n5628), .A(n6140), .Z(n6554) );
  XOR U7953 ( .A(n6580), .B(n5844), .Z(out[1081]) );
  XNOR U7954 ( .A(n6581), .B(n5335), .Z(n5844) );
  XNOR U7955 ( .A(n6582), .B(n5927), .Z(n5335) );
  XNOR U7956 ( .A(n6583), .B(n6584), .Z(n5927) );
  XNOR U7957 ( .A(n5548), .B(n3682), .Z(n6584) );
  XOR U7958 ( .A(n6585), .B(n6586), .Z(n3682) );
  NOR U7959 ( .A(n6587), .B(n6588), .Z(n6585) );
  XNOR U7960 ( .A(n6589), .B(n6590), .Z(n5548) );
  ANDN U7961 ( .B(n6591), .A(n6592), .Z(n6589) );
  XNOR U7962 ( .A(n6350), .B(n6593), .Z(n6583) );
  XOR U7963 ( .A(n2451), .B(n5956), .Z(n6593) );
  XNOR U7964 ( .A(n6594), .B(n6595), .Z(n5956) );
  XNOR U7965 ( .A(n6598), .B(n6599), .Z(n2451) );
  ANDN U7966 ( .B(n6600), .A(n6601), .Z(n6598) );
  XOR U7967 ( .A(n6602), .B(n6603), .Z(n6350) );
  NOR U7968 ( .A(n6604), .B(n6605), .Z(n6602) );
  ANDN U7969 ( .B(n5632), .A(n6145), .Z(n6580) );
  XOR U7970 ( .A(n6606), .B(n5846), .Z(out[1080]) );
  XNOR U7971 ( .A(n6607), .B(n2590), .Z(n5846) );
  XNOR U7972 ( .A(n6608), .B(n5933), .Z(n2590) );
  XNOR U7973 ( .A(n6609), .B(n6610), .Z(n5933) );
  XNOR U7974 ( .A(n5552), .B(n3686), .Z(n6610) );
  XNOR U7975 ( .A(n6611), .B(n6612), .Z(n3686) );
  ANDN U7976 ( .B(n6613), .A(n6614), .Z(n6611) );
  XOR U7977 ( .A(n6615), .B(n6616), .Z(n5552) );
  ANDN U7978 ( .B(n6617), .A(n6618), .Z(n6615) );
  XOR U7979 ( .A(n6354), .B(n6619), .Z(n6609) );
  XOR U7980 ( .A(n2462), .B(n6011), .Z(n6619) );
  NOR U7981 ( .A(n6622), .B(n6623), .Z(n6620) );
  XNOR U7982 ( .A(n6624), .B(n6625), .Z(n2462) );
  NOR U7983 ( .A(n6626), .B(n6627), .Z(n6624) );
  XNOR U7984 ( .A(n6628), .B(n6629), .Z(n6354) );
  ANDN U7985 ( .B(n6630), .A(n6631), .Z(n6628) );
  ANDN U7986 ( .B(n5636), .A(n6632), .Z(n6606) );
  XNOR U7987 ( .A(n6633), .B(n4178), .Z(out[107]) );
  XOR U7988 ( .A(n6634), .B(n6400), .Z(n4178) );
  XOR U7989 ( .A(n6635), .B(n6636), .Z(n6400) );
  ANDN U7990 ( .B(n3426), .A(n3428), .Z(n6633) );
  XOR U7991 ( .A(n6637), .B(n2299), .Z(n3428) );
  XOR U7992 ( .A(n6638), .B(n3192), .Z(n3426) );
  XOR U7993 ( .A(n6639), .B(n5849), .Z(out[1079]) );
  XNOR U7994 ( .A(n6640), .B(n2595), .Z(n5849) );
  XNOR U7995 ( .A(n6641), .B(n5938), .Z(n2595) );
  XNOR U7996 ( .A(n6642), .B(n6643), .Z(n5938) );
  XNOR U7997 ( .A(n5556), .B(n3692), .Z(n6643) );
  XNOR U7998 ( .A(n6644), .B(n6645), .Z(n3692) );
  NOR U7999 ( .A(n6646), .B(n6647), .Z(n6644) );
  XOR U8000 ( .A(n6648), .B(n6649), .Z(n5556) );
  ANDN U8001 ( .B(n6650), .A(n6651), .Z(n6648) );
  XOR U8002 ( .A(n6359), .B(n6652), .Z(n6642) );
  XNOR U8003 ( .A(n2469), .B(n6068), .Z(n6652) );
  XNOR U8004 ( .A(n6653), .B(n6654), .Z(n6068) );
  ANDN U8005 ( .B(n6655), .A(n6656), .Z(n6653) );
  XNOR U8006 ( .A(n6657), .B(n6658), .Z(n2469) );
  ANDN U8007 ( .B(n6659), .A(n6660), .Z(n6657) );
  XNOR U8008 ( .A(n6661), .B(n6662), .Z(n6359) );
  ANDN U8009 ( .B(n6663), .A(n6664), .Z(n6661) );
  ANDN U8010 ( .B(n5640), .A(n6155), .Z(n6639) );
  XOR U8011 ( .A(n6665), .B(n5851), .Z(out[1078]) );
  XOR U8012 ( .A(n6666), .B(n2604), .Z(n5851) );
  IV U8013 ( .A(n5348), .Z(n2604) );
  XNOR U8014 ( .A(n6667), .B(n5943), .Z(n5348) );
  XNOR U8015 ( .A(n6668), .B(n6669), .Z(n5943) );
  XNOR U8016 ( .A(n5563), .B(n3698), .Z(n6669) );
  XOR U8017 ( .A(n6670), .B(n6671), .Z(n3698) );
  ANDN U8018 ( .B(n6672), .A(n6673), .Z(n6670) );
  XNOR U8019 ( .A(n6674), .B(n6675), .Z(n5563) );
  ANDN U8020 ( .B(n6676), .A(n6677), .Z(n6674) );
  XNOR U8021 ( .A(n6364), .B(n6678), .Z(n6668) );
  XNOR U8022 ( .A(n2476), .B(n6118), .Z(n6678) );
  XNOR U8023 ( .A(n6679), .B(n6680), .Z(n6118) );
  ANDN U8024 ( .B(n6681), .A(n6682), .Z(n6679) );
  XOR U8025 ( .A(n6683), .B(n6684), .Z(n2476) );
  ANDN U8026 ( .B(n6685), .A(n6686), .Z(n6683) );
  XNOR U8027 ( .A(n6687), .B(n6688), .Z(n6364) );
  ANDN U8028 ( .B(n6689), .A(n6690), .Z(n6687) );
  NOR U8029 ( .A(n6160), .B(n5644), .Z(n6665) );
  XOR U8030 ( .A(n6691), .B(n5853), .Z(out[1077]) );
  XNOR U8031 ( .A(n6692), .B(n2615), .Z(n5853) );
  XNOR U8032 ( .A(n6693), .B(n5948), .Z(n2615) );
  XNOR U8033 ( .A(n6694), .B(n6695), .Z(n5948) );
  XOR U8034 ( .A(n5568), .B(n3701), .Z(n6695) );
  XOR U8035 ( .A(n6696), .B(n6697), .Z(n3701) );
  ANDN U8036 ( .B(n6698), .A(n6699), .Z(n6696) );
  XNOR U8037 ( .A(n6700), .B(n6701), .Z(n5568) );
  XNOR U8038 ( .A(n6376), .B(n6704), .Z(n6694) );
  XOR U8039 ( .A(n2483), .B(n6173), .Z(n6704) );
  ANDN U8040 ( .B(n6707), .A(n6708), .Z(n6705) );
  XNOR U8041 ( .A(n6709), .B(n6710), .Z(n2483) );
  NOR U8042 ( .A(n6711), .B(n6712), .Z(n6709) );
  XOR U8043 ( .A(n6713), .B(n6714), .Z(n6376) );
  ANDN U8044 ( .B(n5652), .A(n6717), .Z(n6691) );
  XNOR U8045 ( .A(n6718), .B(n6171), .Z(out[1076]) );
  XOR U8046 ( .A(n5357), .B(n6719), .Z(n6171) );
  XNOR U8047 ( .A(n5952), .B(n6720), .Z(n5357) );
  XOR U8048 ( .A(n6721), .B(n6722), .Z(n5952) );
  XOR U8049 ( .A(n6380), .B(n2490), .Z(n6722) );
  XNOR U8050 ( .A(n6723), .B(n6724), .Z(n2490) );
  ANDN U8051 ( .B(n6725), .A(n6726), .Z(n6723) );
  ANDN U8052 ( .B(n6729), .A(n6730), .Z(n6727) );
  XOR U8053 ( .A(n3705), .B(n6731), .Z(n6721) );
  XNOR U8054 ( .A(n6228), .B(n5573), .Z(n6731) );
  XOR U8055 ( .A(n6732), .B(n6733), .Z(n5573) );
  XOR U8056 ( .A(n6734), .B(n4694), .Z(n6733) );
  ANDN U8057 ( .B(n6735), .A(n6736), .Z(n6734) );
  XNOR U8058 ( .A(n6737), .B(n6738), .Z(n6228) );
  AND U8059 ( .A(n6739), .B(n6740), .Z(n6737) );
  XNOR U8060 ( .A(n6741), .B(n6742), .Z(n3705) );
  ANDN U8061 ( .B(n6743), .A(n6744), .Z(n6741) );
  NOR U8062 ( .A(n6170), .B(n5656), .Z(n6718) );
  XOR U8063 ( .A(n6745), .B(n5857), .Z(out[1075]) );
  XNOR U8064 ( .A(n6746), .B(n2629), .Z(n5857) );
  XNOR U8065 ( .A(n6747), .B(n5963), .Z(n2629) );
  XNOR U8066 ( .A(n6748), .B(n6749), .Z(n5963) );
  XNOR U8067 ( .A(n5576), .B(n3710), .Z(n6749) );
  XOR U8068 ( .A(n6750), .B(n6751), .Z(n3710) );
  NOR U8069 ( .A(n6752), .B(n6753), .Z(n6750) );
  XOR U8070 ( .A(n6754), .B(n6755), .Z(n5576) );
  AND U8071 ( .A(n6756), .B(n6757), .Z(n6754) );
  XNOR U8072 ( .A(n6384), .B(n6758), .Z(n6748) );
  XOR U8073 ( .A(n2497), .B(n6275), .Z(n6758) );
  XNOR U8074 ( .A(n6759), .B(n6760), .Z(n6275) );
  NOR U8075 ( .A(n6761), .B(n6762), .Z(n6759) );
  XOR U8076 ( .A(n6763), .B(n6764), .Z(n2497) );
  NOR U8077 ( .A(n6765), .B(n6766), .Z(n6763) );
  XNOR U8078 ( .A(n6767), .B(n6768), .Z(n6384) );
  ANDN U8079 ( .B(n5660), .A(n6180), .Z(n6745) );
  XNOR U8080 ( .A(n6771), .B(n5859), .Z(out[1074]) );
  XOR U8081 ( .A(n6772), .B(n2636), .Z(n5859) );
  XNOR U8082 ( .A(n6773), .B(n5968), .Z(n2636) );
  XNOR U8083 ( .A(n6774), .B(n6775), .Z(n5968) );
  XOR U8084 ( .A(n5581), .B(n3716), .Z(n6775) );
  XOR U8085 ( .A(n6776), .B(n6777), .Z(n3716) );
  ANDN U8086 ( .B(n6778), .A(n6779), .Z(n6776) );
  XNOR U8087 ( .A(n6780), .B(n6781), .Z(n5581) );
  ANDN U8088 ( .B(n6782), .A(n6783), .Z(n6780) );
  XNOR U8089 ( .A(n6388), .B(n6784), .Z(n6774) );
  XNOR U8090 ( .A(n2504), .B(n6320), .Z(n6784) );
  XNOR U8091 ( .A(n6785), .B(n6786), .Z(n6320) );
  NOR U8092 ( .A(n6787), .B(n6788), .Z(n6785) );
  XOR U8093 ( .A(n6789), .B(n6790), .Z(n2504) );
  NOR U8094 ( .A(n6791), .B(n6792), .Z(n6789) );
  XNOR U8095 ( .A(n6793), .B(n6794), .Z(n6388) );
  NOR U8096 ( .A(n6795), .B(n6796), .Z(n6793) );
  NOR U8097 ( .A(n6185), .B(n5664), .Z(n6771) );
  XOR U8098 ( .A(n6797), .B(n5861), .Z(out[1073]) );
  XOR U8099 ( .A(n6798), .B(n3338), .Z(n5861) );
  XNOR U8100 ( .A(n6799), .B(n5973), .Z(n3338) );
  XNOR U8101 ( .A(n6800), .B(n6801), .Z(n5973) );
  XNOR U8102 ( .A(n5585), .B(n3721), .Z(n6801) );
  XNOR U8103 ( .A(n6802), .B(n6803), .Z(n3721) );
  XNOR U8104 ( .A(n6806), .B(n6807), .Z(n5585) );
  ANDN U8105 ( .B(n6808), .A(n6809), .Z(n6806) );
  XOR U8106 ( .A(n6392), .B(n6810), .Z(n6800) );
  XNOR U8107 ( .A(n2511), .B(n6372), .Z(n6810) );
  XOR U8108 ( .A(n6811), .B(n6812), .Z(n6372) );
  NOR U8109 ( .A(n6813), .B(n6814), .Z(n6811) );
  XNOR U8110 ( .A(n6815), .B(n6816), .Z(n2511) );
  XNOR U8111 ( .A(n6819), .B(n6820), .Z(n6392) );
  ANDN U8112 ( .B(n6821), .A(n6822), .Z(n6819) );
  ANDN U8113 ( .B(n5668), .A(n6823), .Z(n6797) );
  XOR U8114 ( .A(n6824), .B(n5863), .Z(out[1072]) );
  XOR U8115 ( .A(n6825), .B(n5315), .Z(n5863) );
  XNOR U8116 ( .A(n6826), .B(n5978), .Z(n5315) );
  XNOR U8117 ( .A(n6827), .B(n6828), .Z(n5978) );
  XOR U8118 ( .A(n5590), .B(n3730), .Z(n6828) );
  XOR U8119 ( .A(n6829), .B(n6830), .Z(n3730) );
  AND U8120 ( .A(n6831), .B(n6832), .Z(n6829) );
  XNOR U8121 ( .A(n6833), .B(n6834), .Z(n5590) );
  XNOR U8122 ( .A(n4687), .B(n6835), .Z(n6834) );
  NANDN U8123 ( .A(n6836), .B(n6837), .Z(n6835) );
  XNOR U8124 ( .A(n6396), .B(n6838), .Z(n6827) );
  XOR U8125 ( .A(n2518), .B(n6411), .Z(n6838) );
  XNOR U8126 ( .A(n6839), .B(n6840), .Z(n6411) );
  ANDN U8127 ( .B(n6841), .A(n6842), .Z(n6839) );
  XNOR U8128 ( .A(n6843), .B(n6844), .Z(n2518) );
  XOR U8129 ( .A(n6847), .B(n6848), .Z(n6396) );
  AND U8130 ( .A(n6849), .B(n6850), .Z(n6847) );
  ANDN U8131 ( .B(n5672), .A(n6851), .Z(n6824) );
  XOR U8132 ( .A(n6852), .B(n5874), .Z(out[1071]) );
  XOR U8133 ( .A(n6853), .B(n5382), .Z(n5874) );
  XNOR U8134 ( .A(n6854), .B(n5983), .Z(n5382) );
  XNOR U8135 ( .A(n6855), .B(n6856), .Z(n5983) );
  XNOR U8136 ( .A(n5593), .B(n3736), .Z(n6856) );
  XOR U8137 ( .A(n6857), .B(n6858), .Z(n3736) );
  XOR U8138 ( .A(n6861), .B(n6862), .Z(n5593) );
  AND U8139 ( .A(n6863), .B(n6864), .Z(n6861) );
  XOR U8140 ( .A(n6399), .B(n6865), .Z(n6855) );
  XOR U8141 ( .A(n2525), .B(n6634), .Z(n6865) );
  XNOR U8142 ( .A(n6866), .B(n6867), .Z(n6634) );
  NOR U8143 ( .A(n6868), .B(n6869), .Z(n6866) );
  XNOR U8144 ( .A(n6870), .B(n6871), .Z(n2525) );
  NOR U8145 ( .A(n6872), .B(n6873), .Z(n6870) );
  XNOR U8146 ( .A(n6874), .B(n6875), .Z(n6399) );
  NOR U8147 ( .A(n6876), .B(n6877), .Z(n6874) );
  ANDN U8148 ( .B(n5676), .A(n6878), .Z(n6852) );
  XOR U8149 ( .A(n6879), .B(n5876), .Z(out[1070]) );
  XNOR U8150 ( .A(n6880), .B(n5414), .Z(n5876) );
  XNOR U8151 ( .A(n6881), .B(n5988), .Z(n5414) );
  XNOR U8152 ( .A(n6882), .B(n6883), .Z(n5988) );
  XOR U8153 ( .A(n5597), .B(n3739), .Z(n6883) );
  XOR U8154 ( .A(n6884), .B(n6885), .Z(n3739) );
  XNOR U8155 ( .A(n6888), .B(n6889), .Z(n5597) );
  NOR U8156 ( .A(n6890), .B(n6891), .Z(n6888) );
  XOR U8157 ( .A(n6403), .B(n6892), .Z(n6882) );
  XNOR U8158 ( .A(n2536), .B(n6893), .Z(n6892) );
  XOR U8159 ( .A(n6894), .B(n6895), .Z(n2536) );
  XNOR U8160 ( .A(n6898), .B(n6899), .Z(n6403) );
  NOR U8161 ( .A(n6902), .B(n5680), .Z(n6879) );
  XOR U8162 ( .A(n6903), .B(n4183), .Z(out[106]) );
  XNOR U8163 ( .A(n6893), .B(n2537), .Z(n4183) );
  XNOR U8164 ( .A(n6904), .B(n6905), .Z(n2537) );
  XNOR U8165 ( .A(n6906), .B(n6907), .Z(n6893) );
  ANDN U8166 ( .B(n6908), .A(n6909), .Z(n6906) );
  ANDN U8167 ( .B(n3458), .A(n3460), .Z(n6903) );
  XOR U8168 ( .A(n6910), .B(n2306), .Z(n3460) );
  XNOR U8169 ( .A(n6911), .B(n3196), .Z(n3458) );
  XOR U8170 ( .A(n6912), .B(n5878), .Z(out[1069]) );
  XOR U8171 ( .A(n6913), .B(n2671), .Z(n5878) );
  XNOR U8172 ( .A(n6914), .B(n5993), .Z(n2671) );
  XNOR U8173 ( .A(n6915), .B(n6916), .Z(n5993) );
  XOR U8174 ( .A(n5601), .B(n3744), .Z(n6916) );
  XOR U8175 ( .A(n6917), .B(n6918), .Z(n3744) );
  XOR U8176 ( .A(n6921), .B(n6922), .Z(n5601) );
  XOR U8177 ( .A(n6923), .B(n4407), .Z(n6922) );
  ANDN U8178 ( .B(n6924), .A(n6925), .Z(n6923) );
  XOR U8179 ( .A(n6406), .B(n6926), .Z(n6915) );
  XOR U8180 ( .A(n2543), .B(n6927), .Z(n6926) );
  XOR U8181 ( .A(n6928), .B(n6929), .Z(n2543) );
  NOR U8182 ( .A(n6930), .B(n6931), .Z(n6928) );
  XNOR U8183 ( .A(n6932), .B(n6933), .Z(n6406) );
  NOR U8184 ( .A(n6934), .B(n6935), .Z(n6932) );
  ANDN U8185 ( .B(n5684), .A(n6936), .Z(n6912) );
  XOR U8186 ( .A(n6937), .B(n5880), .Z(out[1068]) );
  XOR U8187 ( .A(n6938), .B(n5515), .Z(n5880) );
  XNOR U8188 ( .A(n6939), .B(n5998), .Z(n5515) );
  XNOR U8189 ( .A(n6940), .B(n6941), .Z(n5998) );
  XOR U8190 ( .A(n5297), .B(n3747), .Z(n6941) );
  XOR U8191 ( .A(n6942), .B(n6943), .Z(n3747) );
  XOR U8192 ( .A(n6946), .B(n6947), .Z(n5297) );
  XOR U8193 ( .A(n6948), .B(n4694), .Z(n6947) );
  NOR U8194 ( .A(n6949), .B(n6950), .Z(n6948) );
  XOR U8195 ( .A(n6409), .B(n6951), .Z(n6940) );
  XOR U8196 ( .A(n2550), .B(n6952), .Z(n6951) );
  XOR U8197 ( .A(n6953), .B(n6954), .Z(n2550) );
  ANDN U8198 ( .B(n6955), .A(n6956), .Z(n6953) );
  XOR U8199 ( .A(n6957), .B(n6958), .Z(n6409) );
  ANDN U8200 ( .B(n6959), .A(n6960), .Z(n6957) );
  NOR U8201 ( .A(n6961), .B(n5688), .Z(n6937) );
  XOR U8202 ( .A(n6962), .B(n5882), .Z(out[1067]) );
  XOR U8203 ( .A(n3363), .B(n6963), .Z(n5882) );
  NOR U8204 ( .A(n5697), .B(n6220), .Z(n6962) );
  XNOR U8205 ( .A(n6964), .B(n5884), .Z(out[1066]) );
  IV U8206 ( .A(n6226), .Z(n5884) );
  XNOR U8207 ( .A(n2217), .B(n6965), .Z(n6226) );
  XOR U8208 ( .A(n6966), .B(n6008), .Z(n2217) );
  XNOR U8209 ( .A(n6967), .B(n6968), .Z(n6008) );
  XNOR U8210 ( .A(n5306), .B(n3756), .Z(n6968) );
  XNOR U8211 ( .A(n6969), .B(n6970), .Z(n3756) );
  NOR U8212 ( .A(n6971), .B(n6972), .Z(n6969) );
  XNOR U8213 ( .A(n6973), .B(n6974), .Z(n5306) );
  ANDN U8214 ( .B(n6975), .A(n6976), .Z(n6973) );
  XNOR U8215 ( .A(n6420), .B(n6977), .Z(n6967) );
  XNOR U8216 ( .A(n2564), .B(n6978), .Z(n6977) );
  XNOR U8217 ( .A(n6979), .B(n6980), .Z(n2564) );
  ANDN U8218 ( .B(n6981), .A(n6982), .Z(n6979) );
  XOR U8219 ( .A(n6983), .B(n6984), .Z(n6420) );
  NOR U8220 ( .A(n6985), .B(n6986), .Z(n6983) );
  NOR U8221 ( .A(n6225), .B(n5701), .Z(n6964) );
  XOR U8222 ( .A(n6987), .B(n5886), .Z(out[1065]) );
  XOR U8223 ( .A(n3371), .B(n6988), .Z(n5886) );
  XOR U8224 ( .A(n6989), .B(n6018), .Z(n3371) );
  XNOR U8225 ( .A(n6990), .B(n6991), .Z(n6018) );
  XOR U8226 ( .A(n5309), .B(n3761), .Z(n6991) );
  XOR U8227 ( .A(n6992), .B(n6993), .Z(n3761) );
  NOR U8228 ( .A(n6994), .B(n6995), .Z(n6992) );
  XNOR U8229 ( .A(n6996), .B(n6997), .Z(n5309) );
  NOR U8230 ( .A(n6998), .B(n6999), .Z(n6996) );
  XNOR U8231 ( .A(n6112), .B(n7000), .Z(n6990) );
  XOR U8232 ( .A(n2571), .B(n7001), .Z(n7000) );
  XNOR U8233 ( .A(n7002), .B(n7003), .Z(n2571) );
  AND U8234 ( .A(n7004), .B(n7005), .Z(n7002) );
  XOR U8235 ( .A(n7006), .B(n7007), .Z(n6112) );
  ANDN U8236 ( .B(n7008), .A(n7009), .Z(n7006) );
  NOR U8237 ( .A(n6235), .B(n5705), .Z(n6987) );
  XNOR U8238 ( .A(n7010), .B(n5888), .Z(out[1064]) );
  XOR U8239 ( .A(n5694), .B(n7011), .Z(n5888) );
  XOR U8240 ( .A(n7012), .B(n6023), .Z(n5694) );
  XNOR U8241 ( .A(n7013), .B(n7014), .Z(n6023) );
  XNOR U8242 ( .A(n5319), .B(n3765), .Z(n7014) );
  XNOR U8243 ( .A(n7015), .B(n7016), .Z(n3765) );
  ANDN U8244 ( .B(n7017), .A(n7018), .Z(n7015) );
  XNOR U8245 ( .A(n7019), .B(n7020), .Z(n5319) );
  NOR U8246 ( .A(n7021), .B(n7022), .Z(n7019) );
  XOR U8247 ( .A(n6115), .B(n7023), .Z(n7013) );
  XNOR U8248 ( .A(n2578), .B(n7024), .Z(n7023) );
  XNOR U8249 ( .A(n7025), .B(n7026), .Z(n2578) );
  ANDN U8250 ( .B(n7027), .A(n7028), .Z(n7025) );
  XNOR U8251 ( .A(n7029), .B(n7030), .Z(n6115) );
  ANDN U8252 ( .B(n7031), .A(n7032), .Z(n7029) );
  ANDN U8253 ( .B(n5709), .A(n6240), .Z(n7010) );
  XOR U8254 ( .A(n7033), .B(n5893), .Z(out[1063]) );
  XOR U8255 ( .A(n2244), .B(n7034), .Z(n5893) );
  IV U8256 ( .A(n5728), .Z(n2244) );
  XNOR U8257 ( .A(n7035), .B(n6028), .Z(n5728) );
  XNOR U8258 ( .A(n7036), .B(n7037), .Z(n6028) );
  XOR U8259 ( .A(n5323), .B(n3769), .Z(n7037) );
  XNOR U8260 ( .A(n7038), .B(n7039), .Z(n3769) );
  ANDN U8261 ( .B(n7040), .A(n7041), .Z(n7038) );
  XNOR U8262 ( .A(n7042), .B(n7043), .Z(n5323) );
  ANDN U8263 ( .B(n7044), .A(n7045), .Z(n7042) );
  XNOR U8264 ( .A(n6122), .B(n7046), .Z(n7036) );
  XNOR U8265 ( .A(n4383), .B(n2586), .Z(n7046) );
  XOR U8266 ( .A(n7047), .B(n7048), .Z(n2586) );
  XOR U8267 ( .A(n7051), .B(n7052), .Z(n4383) );
  AND U8268 ( .A(n7053), .B(n7054), .Z(n7051) );
  XOR U8269 ( .A(n7055), .B(n7056), .Z(n6122) );
  ANDN U8270 ( .B(n7057), .A(n7058), .Z(n7055) );
  AND U8271 ( .A(n1041), .B(n1039), .Z(n7033) );
  XOR U8272 ( .A(n2325), .B(n7059), .Z(n1039) );
  XOR U8273 ( .A(n1798), .B(n7060), .Z(n1041) );
  IV U8274 ( .A(n5195), .Z(n1798) );
  XNOR U8275 ( .A(n6582), .B(n6360), .Z(n5195) );
  XOR U8276 ( .A(n7061), .B(n7062), .Z(n6360) );
  XNOR U8277 ( .A(n5941), .B(n2138), .Z(n7062) );
  XOR U8278 ( .A(n7063), .B(n7064), .Z(n2138) );
  ANDN U8279 ( .B(n6654), .A(n6655), .Z(n7063) );
  XOR U8280 ( .A(n7065), .B(n7066), .Z(n5941) );
  ANDN U8281 ( .B(n6647), .A(n7067), .Z(n7065) );
  XOR U8282 ( .A(n5488), .B(n7068), .Z(n7061) );
  XNOR U8283 ( .A(n4346), .B(n3740), .Z(n7068) );
  XOR U8284 ( .A(n7069), .B(n7070), .Z(n3740) );
  XOR U8285 ( .A(n7072), .B(n7073), .Z(n4346) );
  ANDN U8286 ( .B(n6662), .A(n6663), .Z(n7072) );
  XNOR U8287 ( .A(n7074), .B(n7075), .Z(n5488) );
  ANDN U8288 ( .B(n6658), .A(n6659), .Z(n7074) );
  XOR U8289 ( .A(n7076), .B(n7077), .Z(n6582) );
  XOR U8290 ( .A(n3522), .B(n4900), .Z(n7077) );
  XNOR U8291 ( .A(n7078), .B(n6630), .Z(n4900) );
  AND U8292 ( .A(n7079), .B(n7080), .Z(n7078) );
  XNOR U8293 ( .A(n7081), .B(n7082), .Z(n3522) );
  XNOR U8294 ( .A(n7085), .B(n7086), .Z(n7076) );
  XNOR U8295 ( .A(n4072), .B(n2555), .Z(n7086) );
  XNOR U8296 ( .A(n7087), .B(n6613), .Z(n2555) );
  AND U8297 ( .A(n7088), .B(n7089), .Z(n7087) );
  XNOR U8298 ( .A(n7090), .B(n7091), .Z(n4072) );
  XOR U8299 ( .A(n7094), .B(n6249), .Z(out[1062]) );
  XOR U8300 ( .A(n7095), .B(n2252), .Z(n6249) );
  XNOR U8301 ( .A(n7096), .B(n6033), .Z(n2252) );
  XNOR U8302 ( .A(n7097), .B(n7098), .Z(n6033) );
  XNOR U8303 ( .A(n5328), .B(n3775), .Z(n7098) );
  XOR U8304 ( .A(n7099), .B(n7100), .Z(n3775) );
  ANDN U8305 ( .B(n7101), .A(n7102), .Z(n7099) );
  XNOR U8306 ( .A(n7103), .B(n7104), .Z(n5328) );
  ANDN U8307 ( .B(n7105), .A(n7106), .Z(n7103) );
  XOR U8308 ( .A(n6127), .B(n7107), .Z(n7097) );
  XNOR U8309 ( .A(n4388), .B(n2593), .Z(n7107) );
  XOR U8310 ( .A(n7108), .B(n7109), .Z(n2593) );
  ANDN U8311 ( .B(n7110), .A(n7111), .Z(n7108) );
  XOR U8312 ( .A(n7112), .B(n7113), .Z(n4388) );
  ANDN U8313 ( .B(n7114), .A(n7115), .Z(n7112) );
  XNOR U8314 ( .A(n7116), .B(n7117), .Z(n6127) );
  AND U8315 ( .A(n7118), .B(n7119), .Z(n7116) );
  ANDN U8316 ( .B(n1045), .A(n1043), .Z(n7094) );
  XOR U8317 ( .A(n7121), .B(n1804), .Z(n1045) );
  XOR U8318 ( .A(n6608), .B(n6365), .Z(n1804) );
  XOR U8319 ( .A(n7122), .B(n7123), .Z(n6365) );
  XOR U8320 ( .A(n5492), .B(n4348), .Z(n7123) );
  XNOR U8321 ( .A(n7124), .B(n7125), .Z(n4348) );
  XNOR U8322 ( .A(n7126), .B(n7127), .Z(n5492) );
  ANDN U8323 ( .B(n6684), .A(n6685), .Z(n7126) );
  XNOR U8324 ( .A(n3743), .B(n7128), .Z(n7122) );
  XNOR U8325 ( .A(n5946), .B(n2141), .Z(n7128) );
  XOR U8326 ( .A(n7129), .B(n7130), .Z(n2141) );
  NOR U8327 ( .A(n6681), .B(n6680), .Z(n7129) );
  XOR U8328 ( .A(n7131), .B(n7132), .Z(n5946) );
  NOR U8329 ( .A(n6672), .B(n6671), .Z(n7131) );
  IV U8330 ( .A(n7133), .Z(n6672) );
  ANDN U8331 ( .B(n6675), .A(n6676), .Z(n7134) );
  XOR U8332 ( .A(n7136), .B(n7137), .Z(n6608) );
  XNOR U8333 ( .A(n4903), .B(n4075), .Z(n7137) );
  XOR U8334 ( .A(n7138), .B(n6650), .Z(n4075) );
  NOR U8335 ( .A(n7139), .B(n7070), .Z(n7138) );
  XNOR U8336 ( .A(n7140), .B(n7141), .Z(n4903) );
  NOR U8337 ( .A(n7142), .B(n7073), .Z(n7140) );
  XOR U8338 ( .A(n2559), .B(n7143), .Z(n7136) );
  XNOR U8339 ( .A(n3528), .B(n7144), .Z(n7143) );
  XOR U8340 ( .A(n7145), .B(n7146), .Z(n3528) );
  ANDN U8341 ( .B(n7064), .A(n7147), .Z(n7145) );
  XNOR U8342 ( .A(n7148), .B(n6646), .Z(n2559) );
  IV U8343 ( .A(n7149), .Z(n6646) );
  ANDN U8344 ( .B(n7150), .A(n7066), .Z(n7148) );
  XNOR U8345 ( .A(n7151), .B(n5908), .Z(out[1061]) );
  XOR U8346 ( .A(n7152), .B(n2259), .Z(n5908) );
  XNOR U8347 ( .A(n7153), .B(n6038), .Z(n2259) );
  XNOR U8348 ( .A(n7154), .B(n7155), .Z(n6038) );
  XOR U8349 ( .A(n5332), .B(n3781), .Z(n7155) );
  XOR U8350 ( .A(n7156), .B(n7157), .Z(n3781) );
  NOR U8351 ( .A(n7158), .B(n7159), .Z(n7156) );
  XNOR U8352 ( .A(n7160), .B(n7161), .Z(n5332) );
  ANDN U8353 ( .B(n7162), .A(n7163), .Z(n7160) );
  XNOR U8354 ( .A(n6132), .B(n7164), .Z(n7154) );
  XOR U8355 ( .A(n4392), .B(n2600), .Z(n7164) );
  XNOR U8356 ( .A(n7165), .B(n7166), .Z(n2600) );
  ANDN U8357 ( .B(n7167), .A(n7168), .Z(n7165) );
  XOR U8358 ( .A(n7169), .B(n7170), .Z(n4392) );
  ANDN U8359 ( .B(n7171), .A(n7172), .Z(n7169) );
  XOR U8360 ( .A(n7173), .B(n7174), .Z(n6132) );
  ANDN U8361 ( .B(n7175), .A(n7176), .Z(n7173) );
  AND U8362 ( .A(n1048), .B(n1047), .Z(n7151) );
  XNOR U8363 ( .A(n2339), .B(n7177), .Z(n1047) );
  XOR U8364 ( .A(n1807), .B(n7178), .Z(n1048) );
  XNOR U8365 ( .A(n7179), .B(n5913), .Z(out[1060]) );
  XOR U8366 ( .A(n7180), .B(n3397), .Z(n5913) );
  XNOR U8367 ( .A(n7181), .B(n6042), .Z(n3397) );
  XNOR U8368 ( .A(n7182), .B(n7183), .Z(n6042) );
  XOR U8369 ( .A(n5338), .B(n3785), .Z(n7183) );
  XOR U8370 ( .A(n7184), .B(n7185), .Z(n3785) );
  ANDN U8371 ( .B(n7186), .A(n7187), .Z(n7184) );
  XNOR U8372 ( .A(n7188), .B(n7189), .Z(n5338) );
  ANDN U8373 ( .B(n7190), .A(n7191), .Z(n7188) );
  XOR U8374 ( .A(n6137), .B(n7192), .Z(n7182) );
  XNOR U8375 ( .A(n2610), .B(n4395), .Z(n7192) );
  XNOR U8376 ( .A(n7193), .B(n7194), .Z(n4395) );
  ANDN U8377 ( .B(n7195), .A(n7196), .Z(n7193) );
  XOR U8378 ( .A(n7197), .B(n7198), .Z(n2610) );
  ANDN U8379 ( .B(n7199), .A(n7200), .Z(n7197) );
  XNOR U8380 ( .A(n7201), .B(n7202), .Z(n6137) );
  ANDN U8381 ( .B(n7203), .A(n7204), .Z(n7201) );
  AND U8382 ( .A(n1053), .B(n1051), .Z(n7179) );
  XNOR U8383 ( .A(n2346), .B(n7205), .Z(n1051) );
  XOR U8384 ( .A(n4107), .B(n7206), .Z(n1053) );
  IV U8385 ( .A(n1811), .Z(n4107) );
  XNOR U8386 ( .A(n6667), .B(n6381), .Z(n1811) );
  XOR U8387 ( .A(n7207), .B(n7208), .Z(n6381) );
  XOR U8388 ( .A(n5961), .B(n4352), .Z(n7208) );
  XNOR U8389 ( .A(n7209), .B(n7210), .Z(n4352) );
  ANDN U8390 ( .B(n6730), .A(n6728), .Z(n7209) );
  XNOR U8391 ( .A(n7211), .B(n7212), .Z(n5961) );
  XOR U8392 ( .A(n3752), .B(n7213), .Z(n7207) );
  XNOR U8393 ( .A(n5500), .B(n2151), .Z(n7213) );
  XNOR U8394 ( .A(n7214), .B(n7215), .Z(n2151) );
  NOR U8395 ( .A(n6740), .B(n6738), .Z(n7214) );
  XOR U8396 ( .A(n7216), .B(n7217), .Z(n5500) );
  ANDN U8397 ( .B(n6726), .A(n6724), .Z(n7216) );
  XNOR U8398 ( .A(n7218), .B(n7219), .Z(n3752) );
  NOR U8399 ( .A(n6732), .B(n6735), .Z(n7218) );
  XOR U8400 ( .A(n7220), .B(n7221), .Z(n6667) );
  XNOR U8401 ( .A(n4915), .B(n4082), .Z(n7221) );
  XNOR U8402 ( .A(n7222), .B(n6702), .Z(n4082) );
  ANDN U8403 ( .B(n7223), .A(n7224), .Z(n7222) );
  XNOR U8404 ( .A(n7225), .B(n6715), .Z(n4915) );
  ANDN U8405 ( .B(n7226), .A(n7227), .Z(n7225) );
  XOR U8406 ( .A(n2573), .B(n7228), .Z(n7220) );
  XOR U8407 ( .A(n3534), .B(n7229), .Z(n7228) );
  XNOR U8408 ( .A(n7230), .B(n6708), .Z(n3534) );
  AND U8409 ( .A(n7231), .B(n7232), .Z(n7230) );
  XNOR U8410 ( .A(n7233), .B(n6699), .Z(n2573) );
  IV U8411 ( .A(n7234), .Z(n6699) );
  NOR U8412 ( .A(n7235), .B(n7236), .Z(n7233) );
  XOR U8413 ( .A(n7237), .B(n4186), .Z(out[105]) );
  XOR U8414 ( .A(n6927), .B(n2544), .Z(n4186) );
  XOR U8415 ( .A(n7238), .B(n7239), .Z(n2544) );
  XOR U8416 ( .A(n7240), .B(n7241), .Z(n6927) );
  NOR U8417 ( .A(n7242), .B(n7243), .Z(n7240) );
  ANDN U8418 ( .B(n3495), .A(n3493), .Z(n7237) );
  XNOR U8419 ( .A(n7244), .B(n2380), .Z(n3493) );
  XNOR U8420 ( .A(n7245), .B(n2317), .Z(n3495) );
  XNOR U8421 ( .A(n7246), .B(n5918), .Z(out[1059]) );
  XOR U8422 ( .A(n7247), .B(n2273), .Z(n5918) );
  XNOR U8423 ( .A(n7248), .B(n6047), .Z(n2273) );
  XNOR U8424 ( .A(n7249), .B(n7250), .Z(n6047) );
  XNOR U8425 ( .A(n5342), .B(n3788), .Z(n7250) );
  XOR U8426 ( .A(n7251), .B(n7252), .Z(n3788) );
  XNOR U8427 ( .A(n7255), .B(n7256), .Z(n5342) );
  NOR U8428 ( .A(n7257), .B(n7258), .Z(n7255) );
  XNOR U8429 ( .A(n6142), .B(n7259), .Z(n7249) );
  XNOR U8430 ( .A(n2617), .B(n4403), .Z(n7259) );
  XOR U8431 ( .A(n7260), .B(n7261), .Z(n4403) );
  NOR U8432 ( .A(n7262), .B(n7263), .Z(n7260) );
  XNOR U8433 ( .A(n7264), .B(n7265), .Z(n2617) );
  ANDN U8434 ( .B(n7266), .A(n7267), .Z(n7264) );
  XOR U8435 ( .A(n7268), .B(n7269), .Z(n6142) );
  ANDN U8436 ( .B(n7270), .A(n7271), .Z(n7268) );
  AND U8437 ( .A(n1057), .B(n1055), .Z(n7246) );
  XOR U8438 ( .A(n3435), .B(n7272), .Z(n1055) );
  XOR U8439 ( .A(n1815), .B(n7273), .Z(n1057) );
  IV U8440 ( .A(n5206), .Z(n1815) );
  XNOR U8441 ( .A(n6693), .B(n6385), .Z(n5206) );
  XOR U8442 ( .A(n7274), .B(n7275), .Z(n6385) );
  XNOR U8443 ( .A(n5966), .B(n4354), .Z(n7275) );
  XNOR U8444 ( .A(n7276), .B(n7277), .Z(n4354) );
  NOR U8445 ( .A(n6769), .B(n6768), .Z(n7276) );
  XNOR U8446 ( .A(n7278), .B(n7279), .Z(n5966) );
  AND U8447 ( .A(n6751), .B(n6753), .Z(n7278) );
  XOR U8448 ( .A(n3755), .B(n7280), .Z(n7274) );
  XOR U8449 ( .A(n5504), .B(n2154), .Z(n7280) );
  XOR U8450 ( .A(n7281), .B(n7282), .Z(n2154) );
  NOR U8451 ( .A(n7283), .B(n6760), .Z(n7281) );
  XNOR U8452 ( .A(n7284), .B(n7285), .Z(n5504) );
  AND U8453 ( .A(n6764), .B(n6765), .Z(n7284) );
  XOR U8454 ( .A(n7286), .B(n7287), .Z(n3755) );
  ANDN U8455 ( .B(n7288), .A(n6756), .Z(n7286) );
  XOR U8456 ( .A(n7289), .B(n7290), .Z(n6693) );
  XOR U8457 ( .A(n4918), .B(n4086), .Z(n7290) );
  XOR U8458 ( .A(n7291), .B(n6736), .Z(n4086) );
  ANDN U8459 ( .B(n7292), .A(n7293), .Z(n7291) );
  NOR U8460 ( .A(n7210), .B(n7295), .Z(n7294) );
  IV U8461 ( .A(n7296), .Z(n7210) );
  XOR U8462 ( .A(n2580), .B(n7297), .Z(n7289) );
  XOR U8463 ( .A(n3536), .B(n7298), .Z(n7297) );
  XOR U8464 ( .A(n7299), .B(n6739), .Z(n3536) );
  NOR U8465 ( .A(n7215), .B(n7300), .Z(n7299) );
  XOR U8466 ( .A(n7301), .B(n6743), .Z(n2580) );
  NOR U8467 ( .A(n7302), .B(n7212), .Z(n7301) );
  XOR U8468 ( .A(n7303), .B(n5923), .Z(out[1058]) );
  XOR U8469 ( .A(n7304), .B(n2280), .Z(n5923) );
  XNOR U8470 ( .A(n7305), .B(n6053), .Z(n2280) );
  XNOR U8471 ( .A(n7306), .B(n7307), .Z(n6053) );
  XNOR U8472 ( .A(n5346), .B(n3794), .Z(n7307) );
  XOR U8473 ( .A(n7308), .B(n7309), .Z(n3794) );
  ANDN U8474 ( .B(n7310), .A(n7311), .Z(n7308) );
  XOR U8475 ( .A(n7312), .B(n7313), .Z(n5346) );
  NOR U8476 ( .A(n7314), .B(n7315), .Z(n7312) );
  XNOR U8477 ( .A(n6147), .B(n7316), .Z(n7306) );
  XNOR U8478 ( .A(n2624), .B(n4448), .Z(n7316) );
  XNOR U8479 ( .A(n7317), .B(n7318), .Z(n4448) );
  ANDN U8480 ( .B(n7319), .A(n7320), .Z(n7317) );
  XNOR U8481 ( .A(n7321), .B(n7322), .Z(n2624) );
  ANDN U8482 ( .B(n7323), .A(n7324), .Z(n7321) );
  XOR U8483 ( .A(n7325), .B(n7326), .Z(n6147) );
  AND U8484 ( .A(n1061), .B(n1059), .Z(n7303) );
  XOR U8485 ( .A(n2360), .B(n7329), .Z(n1059) );
  XNOR U8486 ( .A(n6233), .B(n7330), .Z(n2360) );
  XOR U8487 ( .A(n7331), .B(n7332), .Z(n6233) );
  XNOR U8488 ( .A(n3205), .B(n7333), .Z(n7332) );
  XNOR U8489 ( .A(n7334), .B(n7335), .Z(n3205) );
  NOR U8490 ( .A(n7336), .B(n7337), .Z(n7334) );
  XOR U8491 ( .A(n5527), .B(n7338), .Z(n7331) );
  XOR U8492 ( .A(n7339), .B(n2399), .Z(n7338) );
  XNOR U8493 ( .A(n7340), .B(n7341), .Z(n2399) );
  NOR U8494 ( .A(n7342), .B(n7343), .Z(n7340) );
  XNOR U8495 ( .A(n7344), .B(n7345), .Z(n5527) );
  NOR U8496 ( .A(n7346), .B(n7347), .Z(n7344) );
  XOR U8497 ( .A(n1828), .B(n7348), .Z(n1061) );
  IV U8498 ( .A(n5209), .Z(n1828) );
  XNOR U8499 ( .A(n6720), .B(n6389), .Z(n5209) );
  XOR U8500 ( .A(n7349), .B(n7350), .Z(n6389) );
  XNOR U8501 ( .A(n5971), .B(n5517), .Z(n7350) );
  XNOR U8502 ( .A(n7351), .B(n7352), .Z(n5517) );
  AND U8503 ( .A(n6790), .B(n6792), .Z(n7351) );
  XNOR U8504 ( .A(n7353), .B(n7354), .Z(n5971) );
  ANDN U8505 ( .B(n6777), .A(n6778), .Z(n7353) );
  XOR U8506 ( .A(n3760), .B(n7355), .Z(n7349) );
  XNOR U8507 ( .A(n4356), .B(n2157), .Z(n7355) );
  XOR U8508 ( .A(n7356), .B(n7357), .Z(n2157) );
  NOR U8509 ( .A(n7358), .B(n6786), .Z(n7356) );
  XNOR U8510 ( .A(n7359), .B(n7360), .Z(n4356) );
  ANDN U8511 ( .B(n6796), .A(n6794), .Z(n7359) );
  XOR U8512 ( .A(n7361), .B(n7362), .Z(n3760) );
  NOR U8513 ( .A(n6782), .B(n6781), .Z(n7361) );
  XOR U8514 ( .A(n7363), .B(n7364), .Z(n6720) );
  XNOR U8515 ( .A(n4921), .B(n4089), .Z(n7364) );
  XOR U8516 ( .A(n7365), .B(n6757), .Z(n4089) );
  ANDN U8517 ( .B(n7287), .A(n7366), .Z(n7365) );
  XOR U8518 ( .A(n7367), .B(n6770), .Z(n4921) );
  NOR U8519 ( .A(n7277), .B(n7368), .Z(n7367) );
  IV U8520 ( .A(n7369), .Z(n7277) );
  XOR U8521 ( .A(n2587), .B(n7370), .Z(n7363) );
  XNOR U8522 ( .A(n3539), .B(n7371), .Z(n7370) );
  XNOR U8523 ( .A(n7372), .B(n6762), .Z(n3539) );
  AND U8524 ( .A(n7373), .B(n7282), .Z(n7372) );
  XNOR U8525 ( .A(n7374), .B(n6752), .Z(n2587) );
  ANDN U8526 ( .B(n7375), .A(n7279), .Z(n7374) );
  XOR U8527 ( .A(n7376), .B(n5928), .Z(out[1057]) );
  XOR U8528 ( .A(n7377), .B(n3142), .Z(n5928) );
  XNOR U8529 ( .A(n7378), .B(n6058), .Z(n3142) );
  XNOR U8530 ( .A(n7379), .B(n7380), .Z(n6058) );
  XOR U8531 ( .A(n5351), .B(n3800), .Z(n7380) );
  XOR U8532 ( .A(n7381), .B(n7382), .Z(n3800) );
  AND U8533 ( .A(n7383), .B(n7384), .Z(n7381) );
  XNOR U8534 ( .A(n7385), .B(n7386), .Z(n5351) );
  XNOR U8535 ( .A(n6152), .B(n7389), .Z(n7379) );
  XOR U8536 ( .A(n2631), .B(n4494), .Z(n7389) );
  XOR U8537 ( .A(n7390), .B(n7391), .Z(n4494) );
  XOR U8538 ( .A(n7394), .B(n7395), .Z(n2631) );
  ANDN U8539 ( .B(n7396), .A(n7397), .Z(n7394) );
  XOR U8540 ( .A(n7398), .B(n7399), .Z(n6152) );
  ANDN U8541 ( .B(n7400), .A(n7401), .Z(n7398) );
  AND U8542 ( .A(n1065), .B(n1063), .Z(n7376) );
  XOR U8543 ( .A(n3441), .B(n7402), .Z(n1063) );
  IV U8544 ( .A(n2367), .Z(n3441) );
  XNOR U8545 ( .A(n6238), .B(n7403), .Z(n2367) );
  XOR U8546 ( .A(n7404), .B(n7405), .Z(n6238) );
  XNOR U8547 ( .A(n3209), .B(n7406), .Z(n7405) );
  XNOR U8548 ( .A(n7407), .B(n7408), .Z(n3209) );
  ANDN U8549 ( .B(n7409), .A(n7410), .Z(n7407) );
  XNOR U8550 ( .A(n5530), .B(n7411), .Z(n7404) );
  XNOR U8551 ( .A(n7412), .B(n2406), .Z(n7411) );
  XOR U8552 ( .A(n7413), .B(n7414), .Z(n2406) );
  NOR U8553 ( .A(n7415), .B(n7416), .Z(n7413) );
  XOR U8554 ( .A(n7417), .B(n7418), .Z(n5530) );
  NOR U8555 ( .A(n7419), .B(n7420), .Z(n7417) );
  XOR U8556 ( .A(n1832), .B(n7421), .Z(n1065) );
  IV U8557 ( .A(n4117), .Z(n1832) );
  XNOR U8558 ( .A(n6747), .B(n6393), .Z(n4117) );
  XOR U8559 ( .A(n7422), .B(n7423), .Z(n6393) );
  XOR U8560 ( .A(n5976), .B(n5521), .Z(n7423) );
  XOR U8561 ( .A(n7424), .B(n7425), .Z(n5521) );
  NOR U8562 ( .A(n6818), .B(n6816), .Z(n7424) );
  XNOR U8563 ( .A(n7426), .B(n7427), .Z(n5976) );
  NOR U8564 ( .A(n6803), .B(n6804), .Z(n7426) );
  XOR U8565 ( .A(n3766), .B(n7428), .Z(n7422) );
  XOR U8566 ( .A(n4358), .B(n2160), .Z(n7428) );
  XNOR U8567 ( .A(n7429), .B(n7430), .Z(n2160) );
  ANDN U8568 ( .B(n6812), .A(n7431), .Z(n7429) );
  XOR U8569 ( .A(n7432), .B(n7433), .Z(n4358) );
  NOR U8570 ( .A(n7434), .B(n6820), .Z(n7432) );
  XOR U8571 ( .A(n7435), .B(n7436), .Z(n3766) );
  NOR U8572 ( .A(n7437), .B(n6807), .Z(n7435) );
  XOR U8573 ( .A(n7438), .B(n7439), .Z(n6747) );
  XNOR U8574 ( .A(n4924), .B(n4094), .Z(n7439) );
  XNOR U8575 ( .A(n7440), .B(n6783), .Z(n4094) );
  IV U8576 ( .A(n7441), .Z(n6783) );
  ANDN U8577 ( .B(n7362), .A(n7442), .Z(n7440) );
  XNOR U8578 ( .A(n7443), .B(n6795), .Z(n4924) );
  NOR U8579 ( .A(n7360), .B(n7444), .Z(n7443) );
  IV U8580 ( .A(n7445), .Z(n7360) );
  XOR U8581 ( .A(n2596), .B(n7446), .Z(n7438) );
  XNOR U8582 ( .A(n3542), .B(n7447), .Z(n7446) );
  XNOR U8583 ( .A(n7448), .B(n6788), .Z(n3542) );
  ANDN U8584 ( .B(n7449), .A(n7450), .Z(n7448) );
  XNOR U8585 ( .A(n7451), .B(n6779), .Z(n2596) );
  IV U8586 ( .A(n7452), .Z(n6779) );
  NOR U8587 ( .A(n7453), .B(n7354), .Z(n7451) );
  XOR U8588 ( .A(n7454), .B(n5934), .Z(out[1056]) );
  XOR U8589 ( .A(n7455), .B(n2294), .Z(n5934) );
  XNOR U8590 ( .A(n7456), .B(n6064), .Z(n2294) );
  XNOR U8591 ( .A(n7457), .B(n7458), .Z(n6064) );
  XOR U8592 ( .A(n5355), .B(n3806), .Z(n7458) );
  XOR U8593 ( .A(n7459), .B(n7460), .Z(n3806) );
  NOR U8594 ( .A(n7461), .B(n7462), .Z(n7459) );
  XNOR U8595 ( .A(n7463), .B(n7464), .Z(n5355) );
  ANDN U8596 ( .B(n7465), .A(n7466), .Z(n7463) );
  XNOR U8597 ( .A(n6157), .B(n7467), .Z(n7457) );
  XOR U8598 ( .A(n2638), .B(n4538), .Z(n7467) );
  XOR U8599 ( .A(n7468), .B(n7469), .Z(n4538) );
  NOR U8600 ( .A(n7470), .B(n7471), .Z(n7468) );
  XOR U8601 ( .A(n7472), .B(n7473), .Z(n2638) );
  ANDN U8602 ( .B(n7474), .A(n7475), .Z(n7472) );
  XNOR U8603 ( .A(n7476), .B(n7477), .Z(n6157) );
  ANDN U8604 ( .B(n7478), .A(n7479), .Z(n7476) );
  ANDN U8605 ( .B(n1067), .A(n1069), .Z(n7454) );
  XNOR U8606 ( .A(n1837), .B(n7480), .Z(n1069) );
  XNOR U8607 ( .A(n6773), .B(n6412), .Z(n1837) );
  XOR U8608 ( .A(n7481), .B(n7482), .Z(n6412) );
  XNOR U8609 ( .A(n5981), .B(n5525), .Z(n7482) );
  XNOR U8610 ( .A(n7483), .B(n7484), .Z(n5525) );
  NOR U8611 ( .A(n6846), .B(n6844), .Z(n7483) );
  XNOR U8612 ( .A(n7485), .B(n7486), .Z(n5981) );
  NOR U8613 ( .A(n6830), .B(n6832), .Z(n7485) );
  XNOR U8614 ( .A(n3770), .B(n7487), .Z(n7481) );
  XNOR U8615 ( .A(n4360), .B(n2163), .Z(n7487) );
  XNOR U8616 ( .A(n7488), .B(n7489), .Z(n2163) );
  ANDN U8617 ( .B(n6842), .A(n6840), .Z(n7488) );
  IV U8618 ( .A(n7490), .Z(n6840) );
  XNOR U8619 ( .A(n7491), .B(n7492), .Z(n4360) );
  ANDN U8620 ( .B(n6848), .A(n6850), .Z(n7491) );
  XOR U8621 ( .A(n7493), .B(n7494), .Z(n3770) );
  ANDN U8622 ( .B(n6833), .A(n6837), .Z(n7493) );
  XOR U8623 ( .A(n7495), .B(n7496), .Z(n6773) );
  XOR U8624 ( .A(n4928), .B(n4097), .Z(n7496) );
  XOR U8625 ( .A(n7497), .B(n6808), .Z(n4097) );
  AND U8626 ( .A(n7436), .B(n7498), .Z(n7497) );
  NOR U8627 ( .A(n7500), .B(n7501), .Z(n7499) );
  IV U8628 ( .A(n7433), .Z(n7500) );
  XNOR U8629 ( .A(n2601), .B(n7502), .Z(n7495) );
  XNOR U8630 ( .A(n3545), .B(n7503), .Z(n7502) );
  XNOR U8631 ( .A(n7504), .B(n6814), .Z(n3545) );
  ANDN U8632 ( .B(n7505), .A(n7430), .Z(n7504) );
  XOR U8633 ( .A(n7506), .B(n6805), .Z(n2601) );
  NOR U8634 ( .A(n7427), .B(n7507), .Z(n7506) );
  IV U8635 ( .A(n7508), .Z(n7427) );
  XNOR U8636 ( .A(n7509), .B(n3444), .Z(n1067) );
  XOR U8637 ( .A(n7510), .B(n7511), .Z(n6243) );
  XNOR U8638 ( .A(n3213), .B(n7512), .Z(n7511) );
  XNOR U8639 ( .A(n7513), .B(n7514), .Z(n3213) );
  ANDN U8640 ( .B(n7515), .A(n7516), .Z(n7513) );
  XNOR U8641 ( .A(n5534), .B(n7517), .Z(n7510) );
  XOR U8642 ( .A(n7518), .B(n2411), .Z(n7517) );
  XNOR U8643 ( .A(n7519), .B(n7520), .Z(n2411) );
  ANDN U8644 ( .B(n7521), .A(n7522), .Z(n7519) );
  XNOR U8645 ( .A(n7523), .B(n7524), .Z(n5534) );
  NOR U8646 ( .A(n7525), .B(n7526), .Z(n7523) );
  XNOR U8647 ( .A(n7528), .B(n5939), .Z(out[1055]) );
  XOR U8648 ( .A(n7529), .B(n2301), .Z(n5939) );
  XNOR U8649 ( .A(n7530), .B(n6074), .Z(n2301) );
  XNOR U8650 ( .A(n7531), .B(n7532), .Z(n6074) );
  XOR U8651 ( .A(n5360), .B(n3810), .Z(n7532) );
  XOR U8652 ( .A(n7533), .B(n7534), .Z(n3810) );
  NOR U8653 ( .A(n7535), .B(n7536), .Z(n7533) );
  XNOR U8654 ( .A(n7537), .B(n7538), .Z(n5360) );
  XOR U8655 ( .A(n6162), .B(n7541), .Z(n7531) );
  XNOR U8656 ( .A(n2645), .B(n4584), .Z(n7541) );
  XNOR U8657 ( .A(n7542), .B(n7543), .Z(n4584) );
  XNOR U8658 ( .A(n7546), .B(n7547), .Z(n2645) );
  NOR U8659 ( .A(n7548), .B(n7549), .Z(n7546) );
  XNOR U8660 ( .A(n7550), .B(n7551), .Z(n6162) );
  ANDN U8661 ( .B(n7552), .A(n7553), .Z(n7550) );
  ANDN U8662 ( .B(n1071), .A(n1072), .Z(n7528) );
  XOR U8663 ( .A(n3626), .B(n7554), .Z(n1072) );
  IV U8664 ( .A(n1841), .Z(n3626) );
  XNOR U8665 ( .A(n6799), .B(n6635), .Z(n1841) );
  XOR U8666 ( .A(n7555), .B(n7556), .Z(n6635) );
  XOR U8667 ( .A(n5986), .B(n2168), .Z(n7556) );
  NOR U8668 ( .A(n7559), .B(n6867), .Z(n7557) );
  XNOR U8669 ( .A(n7560), .B(n7561), .Z(n5986) );
  ANDN U8670 ( .B(n6858), .A(n6859), .Z(n7560) );
  XOR U8671 ( .A(n3776), .B(n7562), .Z(n7555) );
  XNOR U8672 ( .A(n4365), .B(n5529), .Z(n7562) );
  XOR U8673 ( .A(n7563), .B(n7564), .Z(n5529) );
  NOR U8674 ( .A(n7565), .B(n6871), .Z(n7563) );
  ANDN U8675 ( .B(n6877), .A(n6875), .Z(n7566) );
  XNOR U8676 ( .A(n7568), .B(n7569), .Z(n3776) );
  NOR U8677 ( .A(n6862), .B(n6864), .Z(n7568) );
  IV U8678 ( .A(n7570), .Z(n6862) );
  XOR U8679 ( .A(n7571), .B(n7572), .Z(n6799) );
  XNOR U8680 ( .A(n4932), .B(n4279), .Z(n7572) );
  XNOR U8681 ( .A(n7573), .B(n6836), .Z(n4279) );
  IV U8682 ( .A(n7574), .Z(n6836) );
  NOR U8683 ( .A(n7575), .B(n7576), .Z(n7573) );
  XOR U8684 ( .A(n7577), .B(n6849), .Z(n4932) );
  NOR U8685 ( .A(n7492), .B(n7578), .Z(n7577) );
  IV U8686 ( .A(n7579), .Z(n7492) );
  XOR U8687 ( .A(n2612), .B(n7580), .Z(n7571) );
  XOR U8688 ( .A(n3548), .B(n7581), .Z(n7580) );
  XOR U8689 ( .A(n7582), .B(n6841), .Z(n3548) );
  NOR U8690 ( .A(n7583), .B(n7489), .Z(n7582) );
  XOR U8691 ( .A(n7584), .B(n6831), .Z(n2612) );
  NOR U8692 ( .A(n7486), .B(n7585), .Z(n7584) );
  XOR U8693 ( .A(n3447), .B(n7586), .Z(n1071) );
  IV U8694 ( .A(n2381), .Z(n3447) );
  XNOR U8695 ( .A(n6247), .B(n7587), .Z(n2381) );
  XOR U8696 ( .A(n7588), .B(n7589), .Z(n6247) );
  XNOR U8697 ( .A(n3216), .B(n7590), .Z(n7589) );
  XOR U8698 ( .A(n7591), .B(n7592), .Z(n3216) );
  ANDN U8699 ( .B(n7593), .A(n7594), .Z(n7591) );
  XOR U8700 ( .A(n5539), .B(n7595), .Z(n7588) );
  XNOR U8701 ( .A(n7596), .B(n2420), .Z(n7595) );
  XNOR U8702 ( .A(n7597), .B(n7598), .Z(n2420) );
  XNOR U8703 ( .A(n7601), .B(n7602), .Z(n5539) );
  ANDN U8704 ( .B(n7603), .A(n7604), .Z(n7601) );
  XOR U8705 ( .A(n7605), .B(n5944), .Z(out[1054]) );
  XOR U8706 ( .A(n7606), .B(n2308), .Z(n5944) );
  XNOR U8707 ( .A(n7607), .B(n6079), .Z(n2308) );
  XNOR U8708 ( .A(n7608), .B(n7609), .Z(n6079) );
  XOR U8709 ( .A(n5369), .B(n3815), .Z(n7609) );
  XOR U8710 ( .A(n7610), .B(n7611), .Z(n3815) );
  XNOR U8711 ( .A(n7614), .B(n7615), .Z(n5369) );
  ANDN U8712 ( .B(n7616), .A(n7617), .Z(n7614) );
  XNOR U8713 ( .A(n6167), .B(n7618), .Z(n7608) );
  XOR U8714 ( .A(n2652), .B(n4629), .Z(n7618) );
  XOR U8715 ( .A(n7619), .B(n7620), .Z(n4629) );
  AND U8716 ( .A(n7621), .B(n7622), .Z(n7619) );
  XNOR U8717 ( .A(n7623), .B(n7624), .Z(n2652) );
  ANDN U8718 ( .B(n7625), .A(n7626), .Z(n7623) );
  XOR U8719 ( .A(n7627), .B(n7628), .Z(n6167) );
  AND U8720 ( .A(n1076), .B(n1075), .Z(n7605) );
  XOR U8721 ( .A(n2392), .B(n7631), .Z(n1075) );
  XNOR U8722 ( .A(n6252), .B(n7632), .Z(n2392) );
  XOR U8723 ( .A(n7633), .B(n7634), .Z(n6252) );
  XOR U8724 ( .A(n7635), .B(n3220), .Z(n7634) );
  XNOR U8725 ( .A(n7636), .B(n7637), .Z(n3220) );
  ANDN U8726 ( .B(n7638), .A(n7639), .Z(n7636) );
  XNOR U8727 ( .A(n2426), .B(n7640), .Z(n7633) );
  XOR U8728 ( .A(n4382), .B(n5542), .Z(n7640) );
  XNOR U8729 ( .A(n7641), .B(n7642), .Z(n5542) );
  XOR U8730 ( .A(n7645), .B(n7646), .Z(n4382) );
  ANDN U8731 ( .B(n7647), .A(n7648), .Z(n7645) );
  XNOR U8732 ( .A(n7649), .B(n7650), .Z(n2426) );
  ANDN U8733 ( .B(n7651), .A(n7652), .Z(n7649) );
  XOR U8734 ( .A(n1846), .B(n7653), .Z(n1076) );
  IV U8735 ( .A(n5223), .Z(n1846) );
  XNOR U8736 ( .A(n6826), .B(n6904), .Z(n5223) );
  XOR U8737 ( .A(n7654), .B(n7655), .Z(n6904) );
  XNOR U8738 ( .A(n5991), .B(n2171), .Z(n7655) );
  XNOR U8739 ( .A(n7656), .B(n7657), .Z(n2171) );
  NOR U8740 ( .A(n6908), .B(n6907), .Z(n7656) );
  XNOR U8741 ( .A(n7658), .B(n7659), .Z(n5991) );
  ANDN U8742 ( .B(n6885), .A(n6887), .Z(n7658) );
  XOR U8743 ( .A(n3779), .B(n7660), .Z(n7654) );
  XOR U8744 ( .A(n4367), .B(n5533), .Z(n7660) );
  XNOR U8745 ( .A(n7661), .B(n7662), .Z(n5533) );
  ANDN U8746 ( .B(n6895), .A(n6897), .Z(n7661) );
  XNOR U8747 ( .A(n7663), .B(n7664), .Z(n4367) );
  NOR U8748 ( .A(n6901), .B(n6899), .Z(n7663) );
  XNOR U8749 ( .A(n7665), .B(n7666), .Z(n3779) );
  AND U8750 ( .A(n6890), .B(n6889), .Z(n7665) );
  XOR U8751 ( .A(n7667), .B(n7668), .Z(n6826) );
  XNOR U8752 ( .A(n4935), .B(n7669), .Z(n7668) );
  XNOR U8753 ( .A(n7670), .B(n6876), .Z(n4935) );
  IV U8754 ( .A(n7671), .Z(n6876) );
  ANDN U8755 ( .B(n7567), .A(n7672), .Z(n7670) );
  XOR U8756 ( .A(n2621), .B(n7673), .Z(n7667) );
  XNOR U8757 ( .A(n3551), .B(n7674), .Z(n7673) );
  XNOR U8758 ( .A(n7675), .B(n6869), .Z(n3551) );
  ANDN U8759 ( .B(n7558), .A(n7676), .Z(n7675) );
  XNOR U8760 ( .A(n7677), .B(n6860), .Z(n2621) );
  NOR U8761 ( .A(n7678), .B(n7561), .Z(n7677) );
  XNOR U8762 ( .A(n7679), .B(n5949), .Z(out[1053]) );
  IV U8763 ( .A(n6290), .Z(n5949) );
  XOR U8764 ( .A(n7680), .B(n2319), .Z(n6290) );
  XNOR U8765 ( .A(n7681), .B(n6084), .Z(n2319) );
  XNOR U8766 ( .A(n7682), .B(n7683), .Z(n6084) );
  XNOR U8767 ( .A(n5372), .B(n3821), .Z(n7683) );
  XOR U8768 ( .A(n7684), .B(n7685), .Z(n3821) );
  XOR U8769 ( .A(n7688), .B(n7689), .Z(n5372) );
  NOR U8770 ( .A(n7690), .B(n7691), .Z(n7688) );
  XNOR U8771 ( .A(n6177), .B(n7692), .Z(n7682) );
  XOR U8772 ( .A(n2659), .B(n4674), .Z(n7692) );
  XOR U8773 ( .A(n7693), .B(n7694), .Z(n4674) );
  NOR U8774 ( .A(n7695), .B(n7696), .Z(n7693) );
  XNOR U8775 ( .A(n7697), .B(n7698), .Z(n2659) );
  NOR U8776 ( .A(n7699), .B(n7700), .Z(n7697) );
  XOR U8777 ( .A(n7701), .B(n7702), .Z(n6177) );
  NOR U8778 ( .A(n7703), .B(n7704), .Z(n7701) );
  ANDN U8779 ( .B(n1083), .A(n1085), .Z(n7679) );
  XOR U8780 ( .A(n1850), .B(n7705), .Z(n1085) );
  IV U8781 ( .A(n5227), .Z(n1850) );
  XNOR U8782 ( .A(n6854), .B(n7238), .Z(n5227) );
  XOR U8783 ( .A(n7706), .B(n7707), .Z(n7238) );
  XOR U8784 ( .A(n5996), .B(n2174), .Z(n7707) );
  XNOR U8785 ( .A(n7708), .B(n7709), .Z(n2174) );
  ANDN U8786 ( .B(n7241), .A(n7710), .Z(n7708) );
  XOR U8787 ( .A(n7711), .B(n7712), .Z(n5996) );
  NOR U8788 ( .A(n6920), .B(n6918), .Z(n7711) );
  XNOR U8789 ( .A(n5537), .B(n7713), .Z(n7706) );
  XOR U8790 ( .A(n4370), .B(n3784), .Z(n7713) );
  XNOR U8791 ( .A(n7714), .B(n7715), .Z(n3784) );
  NOR U8792 ( .A(n6921), .B(n6924), .Z(n7714) );
  XOR U8793 ( .A(n7716), .B(n7717), .Z(n4370) );
  ANDN U8794 ( .B(n6935), .A(n6933), .Z(n7716) );
  XNOR U8795 ( .A(n7718), .B(n7719), .Z(n5537) );
  XOR U8796 ( .A(n7720), .B(n7721), .Z(n6854) );
  XNOR U8797 ( .A(n4938), .B(n5606), .Z(n7721) );
  XOR U8798 ( .A(n7722), .B(n6891), .Z(n5606) );
  NOR U8799 ( .A(n7723), .B(n7666), .Z(n7722) );
  XNOR U8800 ( .A(n7724), .B(n6900), .Z(n4938) );
  ANDN U8801 ( .B(n7725), .A(n7664), .Z(n7724) );
  IV U8802 ( .A(n7726), .Z(n7664) );
  XOR U8803 ( .A(n2626), .B(n7727), .Z(n7720) );
  XNOR U8804 ( .A(n3554), .B(n7728), .Z(n7727) );
  XNOR U8805 ( .A(n7729), .B(n6909), .Z(n3554) );
  IV U8806 ( .A(n7730), .Z(n6909) );
  ANDN U8807 ( .B(n7731), .A(n7657), .Z(n7729) );
  IV U8808 ( .A(n7732), .Z(n7657) );
  XOR U8809 ( .A(n7733), .B(n6886), .Z(n2626) );
  XNOR U8810 ( .A(n7735), .B(n2398), .Z(n1083) );
  XOR U8811 ( .A(n6256), .B(n7736), .Z(n2398) );
  XOR U8812 ( .A(n7737), .B(n7738), .Z(n6256) );
  XNOR U8813 ( .A(n7739), .B(n3223), .Z(n7738) );
  XNOR U8814 ( .A(n7740), .B(n7741), .Z(n3223) );
  ANDN U8815 ( .B(n7742), .A(n7743), .Z(n7740) );
  XOR U8816 ( .A(n2433), .B(n7744), .Z(n7737) );
  XNOR U8817 ( .A(n4386), .B(n5547), .Z(n7744) );
  XNOR U8818 ( .A(n7745), .B(n7746), .Z(n5547) );
  ANDN U8819 ( .B(n7747), .A(n7748), .Z(n7745) );
  XNOR U8820 ( .A(n7749), .B(n7750), .Z(n4386) );
  AND U8821 ( .A(n7751), .B(n7752), .Z(n7749) );
  XNOR U8822 ( .A(n7753), .B(n7754), .Z(n2433) );
  ANDN U8823 ( .B(n7755), .A(n7756), .Z(n7753) );
  XOR U8824 ( .A(n7757), .B(n5954), .Z(out[1052]) );
  XNOR U8825 ( .A(n7758), .B(n5476), .Z(n5954) );
  XNOR U8826 ( .A(n7759), .B(n6089), .Z(n5476) );
  XNOR U8827 ( .A(n7760), .B(n7761), .Z(n6089) );
  XOR U8828 ( .A(n5376), .B(n3827), .Z(n7761) );
  XOR U8829 ( .A(n7762), .B(n7763), .Z(n3827) );
  ANDN U8830 ( .B(n7764), .A(n7765), .Z(n7762) );
  XOR U8831 ( .A(n7766), .B(n7767), .Z(n5376) );
  ANDN U8832 ( .B(n7768), .A(n7769), .Z(n7766) );
  XOR U8833 ( .A(n6182), .B(n7770), .Z(n7760) );
  XOR U8834 ( .A(n2666), .B(n4713), .Z(n7770) );
  XOR U8835 ( .A(n7771), .B(n7772), .Z(n4713) );
  NOR U8836 ( .A(n7773), .B(n7774), .Z(n7771) );
  XOR U8837 ( .A(n7775), .B(n7776), .Z(n2666) );
  NOR U8838 ( .A(n7777), .B(n7778), .Z(n7775) );
  XNOR U8839 ( .A(n7779), .B(n7780), .Z(n6182) );
  ANDN U8840 ( .B(n7781), .A(n7782), .Z(n7779) );
  NOR U8841 ( .A(n1089), .B(n1087), .Z(n7757) );
  XNOR U8842 ( .A(n7783), .B(n2405), .Z(n1087) );
  XOR U8843 ( .A(n6260), .B(n7784), .Z(n2405) );
  XOR U8844 ( .A(n7785), .B(n7786), .Z(n6260) );
  XOR U8845 ( .A(n3230), .B(n4391), .Z(n7786) );
  XNOR U8846 ( .A(n7787), .B(n7788), .Z(n4391) );
  ANDN U8847 ( .B(n7789), .A(n7790), .Z(n7787) );
  XOR U8848 ( .A(n7791), .B(n7792), .Z(n3230) );
  ANDN U8849 ( .B(n7793), .A(n7794), .Z(n7791) );
  XNOR U8850 ( .A(n5551), .B(n7795), .Z(n7785) );
  XOR U8851 ( .A(n7796), .B(n2439), .Z(n7795) );
  XNOR U8852 ( .A(n7797), .B(n7798), .Z(n2439) );
  ANDN U8853 ( .B(n7799), .A(n7800), .Z(n7797) );
  XNOR U8854 ( .A(n7801), .B(n7802), .Z(n5551) );
  NOR U8855 ( .A(n7803), .B(n7804), .Z(n7801) );
  XOR U8856 ( .A(n1854), .B(n7805), .Z(n1089) );
  IV U8857 ( .A(n3641), .Z(n1854) );
  XNOR U8858 ( .A(n6881), .B(n7806), .Z(n3641) );
  XOR U8859 ( .A(n7807), .B(n7808), .Z(n6881) );
  XNOR U8860 ( .A(n4942), .B(n5649), .Z(n7808) );
  XNOR U8861 ( .A(n7809), .B(n6925), .Z(n5649) );
  IV U8862 ( .A(n7810), .Z(n6925) );
  NOR U8863 ( .A(n7811), .B(n7715), .Z(n7809) );
  XNOR U8864 ( .A(n7812), .B(n6934), .Z(n4942) );
  XNOR U8865 ( .A(n2633), .B(n7814), .Z(n7807) );
  XOR U8866 ( .A(n3562), .B(n7815), .Z(n7814) );
  XNOR U8867 ( .A(n7816), .B(n7243), .Z(n3562) );
  ANDN U8868 ( .B(n7817), .A(n7709), .Z(n7816) );
  XNOR U8869 ( .A(n7818), .B(n6919), .Z(n2633) );
  ANDN U8870 ( .B(n7819), .A(n7820), .Z(n7818) );
  XOR U8871 ( .A(n7821), .B(n5964), .Z(out[1051]) );
  XOR U8872 ( .A(n7822), .B(n5481), .Z(n5964) );
  XNOR U8873 ( .A(n7823), .B(n6094), .Z(n5481) );
  XNOR U8874 ( .A(n7824), .B(n7825), .Z(n6094) );
  XOR U8875 ( .A(n5383), .B(n3832), .Z(n7825) );
  XOR U8876 ( .A(n7826), .B(n7827), .Z(n3832) );
  AND U8877 ( .A(n7828), .B(n7829), .Z(n7826) );
  XOR U8878 ( .A(n7830), .B(n7831), .Z(n5383) );
  ANDN U8879 ( .B(n7832), .A(n7833), .Z(n7830) );
  XNOR U8880 ( .A(n6187), .B(n7834), .Z(n7824) );
  XOR U8881 ( .A(n2673), .B(n4737), .Z(n7834) );
  XOR U8882 ( .A(n7835), .B(n7836), .Z(n4737) );
  ANDN U8883 ( .B(n7837), .A(n7838), .Z(n7835) );
  XOR U8884 ( .A(n7839), .B(n7840), .Z(n2673) );
  ANDN U8885 ( .B(n7841), .A(n7842), .Z(n7839) );
  XOR U8886 ( .A(n7843), .B(n7844), .Z(n6187) );
  NOR U8887 ( .A(n7845), .B(n7846), .Z(n7843) );
  ANDN U8888 ( .B(n1091), .A(n1093), .Z(n7821) );
  XOR U8889 ( .A(n1858), .B(n7847), .Z(n1093) );
  IV U8890 ( .A(n5232), .Z(n1858) );
  XNOR U8891 ( .A(n6914), .B(n7848), .Z(n5232) );
  XOR U8892 ( .A(n7849), .B(n7850), .Z(n6914) );
  XNOR U8893 ( .A(n4945), .B(n7851), .Z(n7850) );
  XNOR U8894 ( .A(n7852), .B(n6960), .Z(n4945) );
  AND U8895 ( .A(n7853), .B(n7854), .Z(n7852) );
  XNOR U8896 ( .A(n2640), .B(n7855), .Z(n7849) );
  XNOR U8897 ( .A(n3565), .B(n5695), .Z(n7855) );
  XNOR U8898 ( .A(n7856), .B(n6950), .Z(n5695) );
  AND U8899 ( .A(n7857), .B(n7858), .Z(n7856) );
  XNOR U8900 ( .A(n7859), .B(n7860), .Z(n3565) );
  NOR U8901 ( .A(n7861), .B(n7862), .Z(n7859) );
  XOR U8902 ( .A(n7863), .B(n6945), .Z(n2640) );
  ANDN U8903 ( .B(n7864), .A(n7865), .Z(n7863) );
  XNOR U8904 ( .A(n2413), .B(n7866), .Z(n1091) );
  XNOR U8905 ( .A(n6264), .B(n7867), .Z(n2413) );
  XOR U8906 ( .A(n7868), .B(n7869), .Z(n6264) );
  XNOR U8907 ( .A(n3233), .B(n4396), .Z(n7869) );
  XNOR U8908 ( .A(n7870), .B(n7871), .Z(n4396) );
  NOR U8909 ( .A(n7872), .B(n7873), .Z(n7870) );
  XOR U8910 ( .A(n7874), .B(n7875), .Z(n3233) );
  XNOR U8911 ( .A(n5555), .B(n7878), .Z(n7868) );
  XNOR U8912 ( .A(n7879), .B(n2446), .Z(n7878) );
  XNOR U8913 ( .A(n7880), .B(n7881), .Z(n2446) );
  ANDN U8914 ( .B(n7882), .A(n7883), .Z(n7880) );
  XNOR U8915 ( .A(n7884), .B(n7885), .Z(n5555) );
  ANDN U8916 ( .B(n7886), .A(n7887), .Z(n7884) );
  XOR U8917 ( .A(n7888), .B(n5969), .Z(out[1050]) );
  XOR U8918 ( .A(n7889), .B(n2338), .Z(n5969) );
  IV U8919 ( .A(n3173), .Z(n2338) );
  XOR U8920 ( .A(n7890), .B(n6099), .Z(n3173) );
  XNOR U8921 ( .A(n7891), .B(n7892), .Z(n6099) );
  XNOR U8922 ( .A(n5387), .B(n3837), .Z(n7892) );
  XOR U8923 ( .A(n7893), .B(n7894), .Z(n3837) );
  XOR U8924 ( .A(n7897), .B(n7898), .Z(n5387) );
  NOR U8925 ( .A(n7899), .B(n7900), .Z(n7897) );
  XNOR U8926 ( .A(n6192), .B(n7901), .Z(n7891) );
  XOR U8927 ( .A(n2206), .B(n4761), .Z(n7901) );
  XOR U8928 ( .A(n7902), .B(n7903), .Z(n4761) );
  XOR U8929 ( .A(n7906), .B(n7907), .Z(n2206) );
  AND U8930 ( .A(n7908), .B(n7909), .Z(n7906) );
  XNOR U8931 ( .A(n7910), .B(n7911), .Z(n6192) );
  ANDN U8932 ( .B(n7912), .A(n7913), .Z(n7910) );
  ANDN U8933 ( .B(n1095), .A(n1096), .Z(n7888) );
  XNOR U8934 ( .A(n1862), .B(n7914), .Z(n1096) );
  XNOR U8935 ( .A(n6939), .B(n7915), .Z(n1862) );
  XOR U8936 ( .A(n7916), .B(n7917), .Z(n6939) );
  XNOR U8937 ( .A(n4952), .B(n7918), .Z(n7917) );
  NOR U8938 ( .A(n7921), .B(n7922), .Z(n7919) );
  XNOR U8939 ( .A(n2647), .B(n7923), .Z(n7916) );
  XNOR U8940 ( .A(n3567), .B(n5730), .Z(n7923) );
  XOR U8941 ( .A(n7924), .B(n7925), .Z(n5730) );
  ANDN U8942 ( .B(n7926), .A(n7927), .Z(n7924) );
  XNOR U8943 ( .A(n7928), .B(n7929), .Z(n3567) );
  ANDN U8944 ( .B(n7930), .A(n7931), .Z(n7928) );
  XNOR U8945 ( .A(n7932), .B(n7933), .Z(n2647) );
  ANDN U8946 ( .B(n7934), .A(n7935), .Z(n7932) );
  XOR U8947 ( .A(n2418), .B(n7936), .Z(n1095) );
  IV U8948 ( .A(n5070), .Z(n2418) );
  XNOR U8949 ( .A(n6268), .B(n7937), .Z(n5070) );
  XOR U8950 ( .A(n7938), .B(n7939), .Z(n6268) );
  XOR U8951 ( .A(n3237), .B(n4402), .Z(n7939) );
  XOR U8952 ( .A(n7940), .B(n7941), .Z(n4402) );
  ANDN U8953 ( .B(n7942), .A(n7943), .Z(n7940) );
  XOR U8954 ( .A(n7944), .B(n7945), .Z(n3237) );
  ANDN U8955 ( .B(n7946), .A(n7947), .Z(n7944) );
  XOR U8956 ( .A(n5565), .B(n7948), .Z(n7938) );
  XNOR U8957 ( .A(n7949), .B(n2453), .Z(n7948) );
  XNOR U8958 ( .A(n7950), .B(n7951), .Z(n2453) );
  ANDN U8959 ( .B(n7952), .A(n7953), .Z(n7950) );
  XOR U8960 ( .A(n7954), .B(n7955), .Z(n5565) );
  AND U8961 ( .A(n7956), .B(n7957), .Z(n7954) );
  XNOR U8962 ( .A(n7958), .B(n4189), .Z(out[104]) );
  IV U8963 ( .A(n4368), .Z(n4189) );
  XNOR U8964 ( .A(n6952), .B(n2551), .Z(n4368) );
  XNOR U8965 ( .A(n7806), .B(n7959), .Z(n2551) );
  XOR U8966 ( .A(n7960), .B(n7961), .Z(n7806) );
  XNOR U8967 ( .A(n4372), .B(n2177), .Z(n7961) );
  XOR U8968 ( .A(n7962), .B(n7862), .Z(n2177) );
  ANDN U8969 ( .B(n7963), .A(n7964), .Z(n7962) );
  XOR U8970 ( .A(n7965), .B(n7854), .Z(n4372) );
  ANDN U8971 ( .B(n6958), .A(n6959), .Z(n7965) );
  XOR U8972 ( .A(n6001), .B(n7966), .Z(n7960) );
  XOR U8973 ( .A(n5541), .B(n3790), .Z(n7966) );
  XOR U8974 ( .A(n7967), .B(n7857), .Z(n3790) );
  ANDN U8975 ( .B(n6949), .A(n6946), .Z(n7967) );
  XOR U8976 ( .A(n7968), .B(n7969), .Z(n5541) );
  ANDN U8977 ( .B(n6954), .A(n6955), .Z(n7968) );
  XOR U8978 ( .A(n7970), .B(n7864), .Z(n6001) );
  ANDN U8979 ( .B(n6943), .A(n6944), .Z(n7970) );
  XOR U8980 ( .A(n7971), .B(n7963), .Z(n6952) );
  ANDN U8981 ( .B(n7964), .A(n7860), .Z(n7971) );
  IV U8982 ( .A(n7972), .Z(n7860) );
  AND U8983 ( .A(n3526), .B(n3524), .Z(n7958) );
  XNOR U8984 ( .A(n7973), .B(n2391), .Z(n3524) );
  XOR U8985 ( .A(n3420), .B(n7974), .Z(n3526) );
  IV U8986 ( .A(n2325), .Z(n3420) );
  XNOR U8987 ( .A(n6203), .B(n7975), .Z(n2325) );
  XOR U8988 ( .A(n7976), .B(n7977), .Z(n6203) );
  XNOR U8989 ( .A(n3182), .B(n6415), .Z(n7977) );
  XNOR U8990 ( .A(n7978), .B(n7979), .Z(n6415) );
  ANDN U8991 ( .B(n7980), .A(n7981), .Z(n7978) );
  XNOR U8992 ( .A(n7982), .B(n7983), .Z(n3182) );
  ANDN U8993 ( .B(n7984), .A(n7985), .Z(n7982) );
  XNOR U8994 ( .A(n5498), .B(n7986), .Z(n7976) );
  XOR U8995 ( .A(n7987), .B(n2358), .Z(n7986) );
  XNOR U8996 ( .A(n7988), .B(n7989), .Z(n2358) );
  NOR U8997 ( .A(n7990), .B(n7991), .Z(n7988) );
  XNOR U8998 ( .A(n7992), .B(n7993), .Z(n5498) );
  ANDN U8999 ( .B(n7994), .A(n7995), .Z(n7992) );
  XNOR U9000 ( .A(n7996), .B(n5974), .Z(out[1049]) );
  XNOR U9001 ( .A(n7997), .B(n2345), .Z(n5974) );
  XNOR U9002 ( .A(n7998), .B(n6104), .Z(n2345) );
  XNOR U9003 ( .A(n7999), .B(n8000), .Z(n6104) );
  XNOR U9004 ( .A(n5391), .B(n3841), .Z(n8000) );
  XNOR U9005 ( .A(n8001), .B(n8002), .Z(n3841) );
  XNOR U9006 ( .A(n8005), .B(n8006), .Z(n5391) );
  XNOR U9007 ( .A(n6197), .B(n8009), .Z(n7999) );
  XOR U9008 ( .A(n2213), .B(n4790), .Z(n8009) );
  XNOR U9009 ( .A(n8010), .B(n8011), .Z(n4790) );
  ANDN U9010 ( .B(n8012), .A(n8013), .Z(n8010) );
  XNOR U9011 ( .A(n8014), .B(n8015), .Z(n2213) );
  ANDN U9012 ( .B(n8016), .A(n8017), .Z(n8014) );
  XOR U9013 ( .A(n8018), .B(n8019), .Z(n6197) );
  ANDN U9014 ( .B(n8020), .A(n8021), .Z(n8018) );
  AND U9015 ( .A(n1100), .B(n1099), .Z(n7996) );
  XOR U9016 ( .A(n2427), .B(n8022), .Z(n1099) );
  XNOR U9017 ( .A(n6272), .B(n8023), .Z(n2427) );
  XOR U9018 ( .A(n8024), .B(n8025), .Z(n6272) );
  XNOR U9019 ( .A(n3241), .B(n4449), .Z(n8025) );
  XNOR U9020 ( .A(n8026), .B(n8027), .Z(n4449) );
  ANDN U9021 ( .B(n8028), .A(n8029), .Z(n8026) );
  XOR U9022 ( .A(n8030), .B(n8031), .Z(n3241) );
  XOR U9023 ( .A(n5569), .B(n8034), .Z(n8024) );
  XNOR U9024 ( .A(n8035), .B(n2464), .Z(n8034) );
  XNOR U9025 ( .A(n8036), .B(n8037), .Z(n2464) );
  AND U9026 ( .A(n8038), .B(n8039), .Z(n8036) );
  XNOR U9027 ( .A(n8040), .B(n8041), .Z(n5569) );
  AND U9028 ( .A(n8042), .B(n8043), .Z(n8040) );
  XOR U9029 ( .A(n1866), .B(n8044), .Z(n1100) );
  IV U9030 ( .A(n5239), .Z(n1866) );
  XNOR U9031 ( .A(n8045), .B(n8046), .Z(n5239) );
  XNOR U9032 ( .A(n8047), .B(n5979), .Z(out[1048]) );
  XNOR U9033 ( .A(n8048), .B(n2352), .Z(n5979) );
  XNOR U9034 ( .A(n8049), .B(n6109), .Z(n2352) );
  XNOR U9035 ( .A(n8050), .B(n8051), .Z(n6109) );
  XOR U9036 ( .A(n5395), .B(n3847), .Z(n8051) );
  XOR U9037 ( .A(n8052), .B(n8053), .Z(n3847) );
  NOR U9038 ( .A(n8054), .B(n8055), .Z(n8052) );
  XNOR U9039 ( .A(n8056), .B(n8057), .Z(n5395) );
  ANDN U9040 ( .B(n8058), .A(n8059), .Z(n8056) );
  XNOR U9041 ( .A(n6202), .B(n8060), .Z(n8050) );
  XOR U9042 ( .A(n2220), .B(n4817), .Z(n8060) );
  XOR U9043 ( .A(n8061), .B(n8062), .Z(n4817) );
  ANDN U9044 ( .B(n8063), .A(n8064), .Z(n8061) );
  XOR U9045 ( .A(n8065), .B(n8066), .Z(n2220) );
  NOR U9046 ( .A(n8067), .B(n8068), .Z(n8065) );
  XOR U9047 ( .A(n8069), .B(n8070), .Z(n6202) );
  AND U9048 ( .A(n1105), .B(n1103), .Z(n8047) );
  XOR U9049 ( .A(n2434), .B(n8073), .Z(n1103) );
  XNOR U9050 ( .A(n6280), .B(n8074), .Z(n2434) );
  XOR U9051 ( .A(n8075), .B(n8076), .Z(n6280) );
  XOR U9052 ( .A(n3244), .B(n4493), .Z(n8076) );
  XOR U9053 ( .A(n8077), .B(n8078), .Z(n4493) );
  NOR U9054 ( .A(n8079), .B(n8080), .Z(n8077) );
  XOR U9055 ( .A(n8081), .B(n8082), .Z(n3244) );
  NOR U9056 ( .A(n8083), .B(n8084), .Z(n8081) );
  XNOR U9057 ( .A(n5572), .B(n8085), .Z(n8075) );
  XOR U9058 ( .A(n8086), .B(n2471), .Z(n8085) );
  XNOR U9059 ( .A(n8087), .B(n8088), .Z(n2471) );
  NOR U9060 ( .A(n8089), .B(n8090), .Z(n8087) );
  XNOR U9061 ( .A(n8091), .B(n8092), .Z(n5572) );
  ANDN U9062 ( .B(n8093), .A(n8094), .Z(n8091) );
  XOR U9063 ( .A(n1874), .B(n8095), .Z(n1105) );
  IV U9064 ( .A(n5242), .Z(n1874) );
  XNOR U9065 ( .A(n6966), .B(n8096), .Z(n5242) );
  XOR U9066 ( .A(n8097), .B(n8098), .Z(n6966) );
  XNOR U9067 ( .A(n4958), .B(n8099), .Z(n8098) );
  ANDN U9068 ( .B(n8101), .A(n8102), .Z(n8100) );
  XOR U9069 ( .A(n2661), .B(n8103), .Z(n8097) );
  XNOR U9070 ( .A(n3571), .B(n5786), .Z(n8103) );
  XNOR U9071 ( .A(n8104), .B(n8105), .Z(n5786) );
  NOR U9072 ( .A(n8106), .B(n8107), .Z(n8104) );
  XOR U9073 ( .A(n8108), .B(n8109), .Z(n3571) );
  NOR U9074 ( .A(n8110), .B(n8111), .Z(n8108) );
  XOR U9075 ( .A(n8112), .B(n6995), .Z(n2661) );
  XNOR U9076 ( .A(n8115), .B(n5984), .Z(out[1047]) );
  XNOR U9077 ( .A(n7987), .B(n2359), .Z(n5984) );
  XNOR U9078 ( .A(n8116), .B(n8117), .Z(n2359) );
  XNOR U9079 ( .A(n8118), .B(n8119), .Z(n7987) );
  NOR U9080 ( .A(n8120), .B(n8121), .Z(n8118) );
  ANDN U9081 ( .B(n1107), .A(n1108), .Z(n8115) );
  XOR U9082 ( .A(n1878), .B(n8122), .Z(n1108) );
  IV U9083 ( .A(n5245), .Z(n1878) );
  XNOR U9084 ( .A(n6124), .B(n6989), .Z(n5245) );
  XOR U9085 ( .A(n8123), .B(n8124), .Z(n6989) );
  XNOR U9086 ( .A(n4961), .B(n8125), .Z(n8124) );
  XNOR U9087 ( .A(n8126), .B(n7032), .Z(n4961) );
  IV U9088 ( .A(n8127), .Z(n7032) );
  AND U9089 ( .A(n8128), .B(n8129), .Z(n8126) );
  XOR U9090 ( .A(n2668), .B(n8130), .Z(n8123) );
  XNOR U9091 ( .A(n3573), .B(n5815), .Z(n8130) );
  XNOR U9092 ( .A(n8131), .B(n7022), .Z(n5815) );
  NOR U9093 ( .A(n8132), .B(n8133), .Z(n8131) );
  XNOR U9094 ( .A(n8134), .B(n8135), .Z(n3573) );
  AND U9095 ( .A(n8136), .B(n8137), .Z(n8134) );
  XNOR U9096 ( .A(n8138), .B(n8139), .Z(n2668) );
  ANDN U9097 ( .B(n8140), .A(n8141), .Z(n8138) );
  XOR U9098 ( .A(n8142), .B(n8143), .Z(n6124) );
  XOR U9099 ( .A(n4390), .B(n2196), .Z(n8143) );
  XNOR U9100 ( .A(n8144), .B(n8145), .Z(n2196) );
  NOR U9101 ( .A(n7054), .B(n7052), .Z(n8144) );
  XNOR U9102 ( .A(n8146), .B(n8147), .Z(n4390) );
  ANDN U9103 ( .B(n7056), .A(n7057), .Z(n8146) );
  XOR U9104 ( .A(n6031), .B(n8148), .Z(n8142) );
  XNOR U9105 ( .A(n5567), .B(n3814), .Z(n8148) );
  XOR U9106 ( .A(n8149), .B(n8150), .Z(n3814) );
  ANDN U9107 ( .B(n7045), .A(n7043), .Z(n8149) );
  XNOR U9108 ( .A(n8151), .B(n8152), .Z(n5567) );
  ANDN U9109 ( .B(n7048), .A(n7050), .Z(n8151) );
  XNOR U9110 ( .A(n8153), .B(n8154), .Z(n6031) );
  NOR U9111 ( .A(n7040), .B(n7039), .Z(n8153) );
  XNOR U9112 ( .A(n2441), .B(n8155), .Z(n1107) );
  XNOR U9113 ( .A(n6284), .B(n8156), .Z(n2441) );
  XOR U9114 ( .A(n8157), .B(n8158), .Z(n6284) );
  XOR U9115 ( .A(n3247), .B(n4537), .Z(n8158) );
  XOR U9116 ( .A(n8159), .B(n8160), .Z(n4537) );
  ANDN U9117 ( .B(n8161), .A(n8162), .Z(n8159) );
  XNOR U9118 ( .A(n8163), .B(n8164), .Z(n3247) );
  XOR U9119 ( .A(n5577), .B(n8167), .Z(n8157) );
  XOR U9120 ( .A(n8168), .B(n2478), .Z(n8167) );
  XNOR U9121 ( .A(n8169), .B(n8170), .Z(n2478) );
  ANDN U9122 ( .B(n8171), .A(n8172), .Z(n8169) );
  XOR U9123 ( .A(n8173), .B(n8174), .Z(n5577) );
  ANDN U9124 ( .B(n8175), .A(n8176), .Z(n8173) );
  XNOR U9125 ( .A(n8177), .B(n5989), .Z(out[1046]) );
  XOR U9126 ( .A(n8178), .B(n2366), .Z(n5989) );
  IV U9127 ( .A(n3192), .Z(n2366) );
  XOR U9128 ( .A(n8179), .B(n8180), .Z(n3192) );
  AND U9129 ( .A(n1112), .B(n1111), .Z(n8177) );
  XOR U9130 ( .A(n2448), .B(n8181), .Z(n1111) );
  IV U9131 ( .A(n3477), .Z(n2448) );
  XNOR U9132 ( .A(n6288), .B(n8182), .Z(n3477) );
  XOR U9133 ( .A(n8183), .B(n8184), .Z(n6288) );
  XOR U9134 ( .A(n3250), .B(n4583), .Z(n8184) );
  NOR U9135 ( .A(n8187), .B(n8188), .Z(n8185) );
  XNOR U9136 ( .A(n8189), .B(n8190), .Z(n3250) );
  NOR U9137 ( .A(n8191), .B(n8192), .Z(n8189) );
  XNOR U9138 ( .A(n5580), .B(n8193), .Z(n8183) );
  XNOR U9139 ( .A(n8194), .B(n2485), .Z(n8193) );
  XNOR U9140 ( .A(n8195), .B(n8196), .Z(n2485) );
  AND U9141 ( .A(n8197), .B(n8198), .Z(n8195) );
  XOR U9142 ( .A(n8199), .B(n8200), .Z(n5580) );
  NOR U9143 ( .A(n8201), .B(n8202), .Z(n8199) );
  XOR U9144 ( .A(n1882), .B(n8203), .Z(n1112) );
  IV U9145 ( .A(n5252), .Z(n1882) );
  XNOR U9146 ( .A(n6129), .B(n7012), .Z(n5252) );
  XOR U9147 ( .A(n8204), .B(n8205), .Z(n7012) );
  XOR U9148 ( .A(n4964), .B(n8206), .Z(n8205) );
  XNOR U9149 ( .A(n8207), .B(n7058), .Z(n4964) );
  IV U9150 ( .A(n8208), .Z(n7058) );
  NOR U9151 ( .A(n8209), .B(n8147), .Z(n8207) );
  XNOR U9152 ( .A(n2675), .B(n8210), .Z(n8204) );
  XOR U9153 ( .A(n3576), .B(n5841), .Z(n8210) );
  XOR U9154 ( .A(n8211), .B(n7044), .Z(n5841) );
  ANDN U9155 ( .B(n8150), .A(n8212), .Z(n8211) );
  XOR U9156 ( .A(n8213), .B(n7053), .Z(n3576) );
  NOR U9157 ( .A(n8145), .B(n8214), .Z(n8213) );
  IV U9158 ( .A(n8215), .Z(n8145) );
  XNOR U9159 ( .A(n8216), .B(n7041), .Z(n2675) );
  ANDN U9160 ( .B(n8217), .A(n8154), .Z(n8216) );
  XOR U9161 ( .A(n8218), .B(n8219), .Z(n6129) );
  XNOR U9162 ( .A(n4394), .B(n2199), .Z(n8219) );
  XNOR U9163 ( .A(n8220), .B(n8221), .Z(n2199) );
  ANDN U9164 ( .B(n7113), .A(n7114), .Z(n8220) );
  XNOR U9165 ( .A(n8222), .B(n8223), .Z(n4394) );
  NOR U9166 ( .A(n7118), .B(n7117), .Z(n8222) );
  XOR U9167 ( .A(n6036), .B(n8224), .Z(n8218) );
  XOR U9168 ( .A(n5571), .B(n3819), .Z(n8224) );
  XOR U9169 ( .A(n8225), .B(n8226), .Z(n3819) );
  ANDN U9170 ( .B(n7104), .A(n7105), .Z(n8225) );
  XNOR U9171 ( .A(n8227), .B(n8228), .Z(n5571) );
  AND U9172 ( .A(n7109), .B(n7111), .Z(n8227) );
  XOR U9173 ( .A(n8229), .B(n8230), .Z(n6036) );
  XNOR U9174 ( .A(n8231), .B(n5994), .Z(out[1045]) );
  IV U9175 ( .A(n6327), .Z(n5994) );
  XOR U9176 ( .A(n8232), .B(n2373), .Z(n6327) );
  IV U9177 ( .A(n3196), .Z(n2373) );
  XOR U9178 ( .A(n8233), .B(n8234), .Z(n3196) );
  AND U9179 ( .A(n1117), .B(n1115), .Z(n8231) );
  XOR U9180 ( .A(n4199), .B(n8235), .Z(n1115) );
  XNOR U9181 ( .A(n6293), .B(n8236), .Z(n4199) );
  XOR U9182 ( .A(n8237), .B(n8238), .Z(n6293) );
  XNOR U9183 ( .A(n3253), .B(n4630), .Z(n8238) );
  XOR U9184 ( .A(n8239), .B(n8240), .Z(n4630) );
  NOR U9185 ( .A(n8241), .B(n8242), .Z(n8239) );
  XNOR U9186 ( .A(n8243), .B(n8244), .Z(n3253) );
  ANDN U9187 ( .B(n8245), .A(n8246), .Z(n8243) );
  XNOR U9188 ( .A(n5586), .B(n8247), .Z(n8237) );
  XOR U9189 ( .A(n8248), .B(n2494), .Z(n8247) );
  XNOR U9190 ( .A(n8249), .B(n8250), .Z(n2494) );
  AND U9191 ( .A(n8251), .B(n8252), .Z(n8249) );
  XOR U9192 ( .A(n8253), .B(n8254), .Z(n5586) );
  NOR U9193 ( .A(n8255), .B(n8256), .Z(n8253) );
  XOR U9194 ( .A(n3675), .B(n8257), .Z(n1117) );
  IV U9195 ( .A(n1886), .Z(n3675) );
  XNOR U9196 ( .A(n7035), .B(n6133), .Z(n1886) );
  XOR U9197 ( .A(n8258), .B(n8259), .Z(n6133) );
  XNOR U9198 ( .A(n4401), .B(n2202), .Z(n8259) );
  XNOR U9199 ( .A(n8260), .B(n8261), .Z(n2202) );
  NOR U9200 ( .A(n7171), .B(n7170), .Z(n8260) );
  XNOR U9201 ( .A(n8262), .B(n8263), .Z(n4401) );
  NOR U9202 ( .A(n8264), .B(n7175), .Z(n8262) );
  XNOR U9203 ( .A(n6041), .B(n8265), .Z(n8258) );
  XOR U9204 ( .A(n5575), .B(n3829), .Z(n8265) );
  XOR U9205 ( .A(n8266), .B(n8267), .Z(n3829) );
  ANDN U9206 ( .B(n7163), .A(n7161), .Z(n8266) );
  XOR U9207 ( .A(n8268), .B(n8269), .Z(n5575) );
  ANDN U9208 ( .B(n7168), .A(n7166), .Z(n8268) );
  XNOR U9209 ( .A(n8270), .B(n8271), .Z(n6041) );
  AND U9210 ( .A(n7157), .B(n7159), .Z(n8270) );
  XOR U9211 ( .A(n8272), .B(n8273), .Z(n7035) );
  XOR U9212 ( .A(n4967), .B(n8274), .Z(n8273) );
  XNOR U9213 ( .A(n8275), .B(n7119), .Z(n4967) );
  ANDN U9214 ( .B(n8276), .A(n8223), .Z(n8275) );
  XNOR U9215 ( .A(n2208), .B(n8277), .Z(n8272) );
  XNOR U9216 ( .A(n3579), .B(n5871), .Z(n8277) );
  XOR U9217 ( .A(n8278), .B(n7106), .Z(n5871) );
  ANDN U9218 ( .B(n8226), .A(n8279), .Z(n8278) );
  XNOR U9219 ( .A(n8280), .B(n7115), .Z(n3579) );
  NOR U9220 ( .A(n8221), .B(n8281), .Z(n8280) );
  IV U9221 ( .A(n8282), .Z(n8221) );
  XOR U9222 ( .A(n8283), .B(n7102), .Z(n2208) );
  AND U9223 ( .A(n8230), .B(n8284), .Z(n8283) );
  XNOR U9224 ( .A(n8285), .B(n5999), .Z(out[1044]) );
  XOR U9225 ( .A(n8286), .B(n2380), .Z(n5999) );
  XNOR U9226 ( .A(n8287), .B(n8288), .Z(n2380) );
  AND U9227 ( .A(n1120), .B(n1119), .Z(n8285) );
  XOR U9228 ( .A(n2466), .B(n8289), .Z(n1119) );
  IV U9229 ( .A(n5090), .Z(n2466) );
  XNOR U9230 ( .A(n6297), .B(n8290), .Z(n5090) );
  XOR U9231 ( .A(n8291), .B(n8292), .Z(n6297) );
  XOR U9232 ( .A(n3257), .B(n4673), .Z(n8292) );
  XNOR U9233 ( .A(n8293), .B(n8294), .Z(n4673) );
  NOR U9234 ( .A(n8295), .B(n8296), .Z(n8293) );
  XNOR U9235 ( .A(n8297), .B(n8298), .Z(n3257) );
  NOR U9236 ( .A(n8299), .B(n8300), .Z(n8297) );
  XOR U9237 ( .A(n5589), .B(n8301), .Z(n8291) );
  XOR U9238 ( .A(n8302), .B(n2499), .Z(n8301) );
  XNOR U9239 ( .A(n8303), .B(n8304), .Z(n2499) );
  ANDN U9240 ( .B(n8305), .A(n8306), .Z(n8303) );
  XOR U9241 ( .A(n8307), .B(n8308), .Z(n5589) );
  NOR U9242 ( .A(n8309), .B(n8310), .Z(n8307) );
  XOR U9243 ( .A(n1891), .B(n8311), .Z(n1120) );
  IV U9244 ( .A(n5258), .Z(n1891) );
  XNOR U9245 ( .A(n7096), .B(n6138), .Z(n5258) );
  XOR U9246 ( .A(n8312), .B(n8313), .Z(n6138) );
  XNOR U9247 ( .A(n4447), .B(n1976), .Z(n8313) );
  XNOR U9248 ( .A(n8314), .B(n8315), .Z(n1976) );
  NOR U9249 ( .A(n7194), .B(n7195), .Z(n8314) );
  XNOR U9250 ( .A(n8316), .B(n8317), .Z(n4447) );
  ANDN U9251 ( .B(n7204), .A(n7202), .Z(n8316) );
  XOR U9252 ( .A(n6046), .B(n8318), .Z(n8312) );
  XNOR U9253 ( .A(n5579), .B(n3833), .Z(n8318) );
  XOR U9254 ( .A(n8319), .B(n8320), .Z(n3833) );
  ANDN U9255 ( .B(n7191), .A(n7189), .Z(n8319) );
  XOR U9256 ( .A(n8321), .B(n8322), .Z(n5579) );
  AND U9257 ( .A(n7200), .B(n7198), .Z(n8321) );
  XNOR U9258 ( .A(n8323), .B(n8324), .Z(n6046) );
  AND U9259 ( .A(n7185), .B(n7187), .Z(n8323) );
  XOR U9260 ( .A(n8325), .B(n8326), .Z(n7096) );
  XNOR U9261 ( .A(n4971), .B(n8327), .Z(n8326) );
  XOR U9262 ( .A(n8328), .B(n7176), .Z(n4971) );
  NOR U9263 ( .A(n8329), .B(n8330), .Z(n8328) );
  XNOR U9264 ( .A(n2215), .B(n8331), .Z(n8325) );
  XNOR U9265 ( .A(n3581), .B(n5901), .Z(n8331) );
  XNOR U9266 ( .A(n8332), .B(n7162), .Z(n5901) );
  AND U9267 ( .A(n8267), .B(n8333), .Z(n8332) );
  XOR U9268 ( .A(n8334), .B(n7172), .Z(n3581) );
  NOR U9269 ( .A(n8261), .B(n8335), .Z(n8334) );
  IV U9270 ( .A(n8336), .Z(n8261) );
  XOR U9271 ( .A(n8337), .B(n7158), .Z(n2215) );
  NOR U9272 ( .A(n8338), .B(n8271), .Z(n8337) );
  XOR U9273 ( .A(n8339), .B(n6004), .Z(out[1043]) );
  XOR U9274 ( .A(n8340), .B(n2391), .Z(n6004) );
  XNOR U9275 ( .A(n8341), .B(n8342), .Z(n2391) );
  AND U9276 ( .A(n1129), .B(n1127), .Z(n8339) );
  XOR U9277 ( .A(n3485), .B(n8343), .Z(n1127) );
  IV U9278 ( .A(n2473), .Z(n3485) );
  XNOR U9279 ( .A(n6301), .B(n8344), .Z(n2473) );
  XOR U9280 ( .A(n8345), .B(n8346), .Z(n6301) );
  XNOR U9281 ( .A(n3260), .B(n4712), .Z(n8346) );
  XNOR U9282 ( .A(n8347), .B(n8348), .Z(n4712) );
  NOR U9283 ( .A(n8349), .B(n8350), .Z(n8347) );
  XOR U9284 ( .A(n8351), .B(n8352), .Z(n3260) );
  ANDN U9285 ( .B(n8353), .A(n8354), .Z(n8351) );
  XOR U9286 ( .A(n5594), .B(n8355), .Z(n8345) );
  XNOR U9287 ( .A(n8356), .B(n2508), .Z(n8355) );
  XNOR U9288 ( .A(n8357), .B(n8358), .Z(n2508) );
  ANDN U9289 ( .B(n8359), .A(n8360), .Z(n8357) );
  XOR U9290 ( .A(n8361), .B(n8362), .Z(n5594) );
  ANDN U9291 ( .B(n8363), .A(n8364), .Z(n8361) );
  XOR U9292 ( .A(n1895), .B(n8365), .Z(n1129) );
  IV U9293 ( .A(n5262), .Z(n1895) );
  XNOR U9294 ( .A(n7153), .B(n6143), .Z(n5262) );
  XOR U9295 ( .A(n8366), .B(n8367), .Z(n6143) );
  XOR U9296 ( .A(n4492), .B(n1979), .Z(n8367) );
  XNOR U9297 ( .A(n8368), .B(n8369), .Z(n1979) );
  AND U9298 ( .A(n7261), .B(n7262), .Z(n8368) );
  XOR U9299 ( .A(n8370), .B(n8371), .Z(n4492) );
  ANDN U9300 ( .B(n7269), .A(n7270), .Z(n8370) );
  IV U9301 ( .A(n8372), .Z(n7270) );
  XOR U9302 ( .A(n6052), .B(n8373), .Z(n8366) );
  XNOR U9303 ( .A(n5583), .B(n3838), .Z(n8373) );
  XNOR U9304 ( .A(n8374), .B(n8375), .Z(n3838) );
  XNOR U9305 ( .A(n8376), .B(n8377), .Z(n5583) );
  NOR U9306 ( .A(n7266), .B(n7265), .Z(n8376) );
  XOR U9307 ( .A(n8378), .B(n8379), .Z(n6052) );
  ANDN U9308 ( .B(n7252), .A(n7254), .Z(n8378) );
  XOR U9309 ( .A(n8380), .B(n8381), .Z(n7153) );
  XOR U9310 ( .A(n4975), .B(n8382), .Z(n8381) );
  XNOR U9311 ( .A(n8383), .B(n7203), .Z(n4975) );
  XOR U9312 ( .A(n2224), .B(n8385), .Z(n8380) );
  XNOR U9313 ( .A(n3583), .B(n5958), .Z(n8385) );
  XNOR U9314 ( .A(n8386), .B(n7190), .Z(n5958) );
  XOR U9315 ( .A(n8388), .B(n7196), .Z(n3583) );
  ANDN U9316 ( .B(n8389), .A(n8315), .Z(n8388) );
  IV U9317 ( .A(n8390), .Z(n8315) );
  XNOR U9318 ( .A(n8391), .B(n7186), .Z(n2224) );
  ANDN U9319 ( .B(n8392), .A(n8324), .Z(n8391) );
  XNOR U9320 ( .A(n8393), .B(n6009), .Z(out[1042]) );
  XOR U9321 ( .A(n7339), .B(n2400), .Z(n6009) );
  IV U9322 ( .A(n3206), .Z(n2400) );
  XNOR U9323 ( .A(n8394), .B(n8395), .Z(n7339) );
  ANDN U9324 ( .B(n8396), .A(n8397), .Z(n8394) );
  AND U9325 ( .A(n1132), .B(n1131), .Z(n8393) );
  XOR U9326 ( .A(n3489), .B(n8398), .Z(n1131) );
  IV U9327 ( .A(n2480), .Z(n3489) );
  XNOR U9328 ( .A(n6305), .B(n8399), .Z(n2480) );
  XOR U9329 ( .A(n8400), .B(n8401), .Z(n6305) );
  XNOR U9330 ( .A(n3269), .B(n4736), .Z(n8401) );
  XNOR U9331 ( .A(n8402), .B(n8403), .Z(n4736) );
  NOR U9332 ( .A(n8404), .B(n8405), .Z(n8402) );
  XOR U9333 ( .A(n8406), .B(n8407), .Z(n3269) );
  NOR U9334 ( .A(n8408), .B(n8409), .Z(n8406) );
  XOR U9335 ( .A(n5598), .B(n8410), .Z(n8400) );
  XNOR U9336 ( .A(n8411), .B(n2515), .Z(n8410) );
  XOR U9337 ( .A(n8412), .B(n8413), .Z(n2515) );
  NOR U9338 ( .A(n8414), .B(n8415), .Z(n8412) );
  XNOR U9339 ( .A(n8416), .B(n8417), .Z(n5598) );
  XOR U9340 ( .A(n1899), .B(n8420), .Z(n1132) );
  IV U9341 ( .A(n5265), .Z(n1899) );
  XNOR U9342 ( .A(n7181), .B(n6148), .Z(n5265) );
  XOR U9343 ( .A(n8421), .B(n8422), .Z(n6148) );
  XNOR U9344 ( .A(n4536), .B(n1982), .Z(n8422) );
  XOR U9345 ( .A(n8423), .B(n8424), .Z(n1982) );
  NOR U9346 ( .A(n7318), .B(n7319), .Z(n8423) );
  XNOR U9347 ( .A(n8425), .B(n8426), .Z(n4536) );
  ANDN U9348 ( .B(n7326), .A(n7327), .Z(n8425) );
  IV U9349 ( .A(n8427), .Z(n7327) );
  XOR U9350 ( .A(n6057), .B(n8428), .Z(n8421) );
  XOR U9351 ( .A(n5588), .B(n3842), .Z(n8428) );
  XNOR U9352 ( .A(n8429), .B(n8430), .Z(n3842) );
  XOR U9353 ( .A(n8431), .B(n8432), .Z(n5588) );
  ANDN U9354 ( .B(n7324), .A(n7322), .Z(n8431) );
  XOR U9355 ( .A(n8433), .B(n8434), .Z(n6057) );
  NOR U9356 ( .A(n8435), .B(n7309), .Z(n8433) );
  XOR U9357 ( .A(n8436), .B(n8437), .Z(n7181) );
  XNOR U9358 ( .A(n4978), .B(n8438), .Z(n8437) );
  XNOR U9359 ( .A(n8439), .B(n7271), .Z(n4978) );
  IV U9360 ( .A(n8440), .Z(n7271) );
  ANDN U9361 ( .B(n8371), .A(n8441), .Z(n8439) );
  XOR U9362 ( .A(n2229), .B(n8442), .Z(n8436) );
  XOR U9363 ( .A(n3589), .B(n6012), .Z(n8442) );
  XNOR U9364 ( .A(n8443), .B(n7258), .Z(n6012) );
  ANDN U9365 ( .B(n8444), .A(n8375), .Z(n8443) );
  XNOR U9366 ( .A(n8445), .B(n7263), .Z(n3589) );
  ANDN U9367 ( .B(n8446), .A(n8369), .Z(n8445) );
  XOR U9368 ( .A(n8447), .B(n7253), .Z(n2229) );
  ANDN U9369 ( .B(n8379), .A(n8448), .Z(n8447) );
  XOR U9370 ( .A(n8449), .B(n6019), .Z(out[1041]) );
  XNOR U9371 ( .A(n7412), .B(n2407), .Z(n6019) );
  IV U9372 ( .A(n3210), .Z(n2407) );
  XNOR U9373 ( .A(n8450), .B(n8451), .Z(n7412) );
  AND U9374 ( .A(n8452), .B(n8453), .Z(n8450) );
  ANDN U9375 ( .B(n1135), .A(n1136), .Z(n8449) );
  XOR U9376 ( .A(n1903), .B(n8454), .Z(n1136) );
  IV U9377 ( .A(n3695), .Z(n1903) );
  XNOR U9378 ( .A(n7248), .B(n6153), .Z(n3695) );
  XOR U9379 ( .A(n8455), .B(n8456), .Z(n6153) );
  XOR U9380 ( .A(n4582), .B(n1985), .Z(n8456) );
  XNOR U9381 ( .A(n8457), .B(n8458), .Z(n1985) );
  ANDN U9382 ( .B(n7391), .A(n7393), .Z(n8457) );
  XNOR U9383 ( .A(n8459), .B(n8460), .Z(n4582) );
  ANDN U9384 ( .B(n7401), .A(n8461), .Z(n8459) );
  IV U9385 ( .A(n8462), .Z(n7401) );
  XOR U9386 ( .A(n6062), .B(n8463), .Z(n8455) );
  XOR U9387 ( .A(n5592), .B(n3846), .Z(n8463) );
  XNOR U9388 ( .A(n8464), .B(n8465), .Z(n3846) );
  NOR U9389 ( .A(n7388), .B(n7386), .Z(n8464) );
  XNOR U9390 ( .A(n8466), .B(n8467), .Z(n5592) );
  ANDN U9391 ( .B(n7397), .A(n8468), .Z(n8466) );
  XNOR U9392 ( .A(n8469), .B(n8470), .Z(n6062) );
  ANDN U9393 ( .B(n7382), .A(n7384), .Z(n8469) );
  XOR U9394 ( .A(n8471), .B(n8472), .Z(n7248) );
  XOR U9395 ( .A(n4982), .B(n8473), .Z(n8472) );
  XOR U9396 ( .A(n8474), .B(n7328), .Z(n4982) );
  ANDN U9397 ( .B(n8475), .A(n8426), .Z(n8474) );
  XOR U9398 ( .A(n2242), .B(n8476), .Z(n8471) );
  XOR U9399 ( .A(n3591), .B(n6070), .Z(n8476) );
  XOR U9400 ( .A(n8477), .B(n7315), .Z(n6070) );
  ANDN U9401 ( .B(n8478), .A(n8430), .Z(n8477) );
  XNOR U9402 ( .A(n8479), .B(n7320), .Z(n3591) );
  IV U9403 ( .A(n8480), .Z(n7320) );
  ANDN U9404 ( .B(n8424), .A(n8481), .Z(n8479) );
  XOR U9405 ( .A(n8482), .B(n7310), .Z(n2242) );
  ANDN U9406 ( .B(n8434), .A(n8483), .Z(n8482) );
  XOR U9407 ( .A(n2487), .B(n8484), .Z(n1135) );
  IV U9408 ( .A(n4862), .Z(n2487) );
  XNOR U9409 ( .A(n5892), .B(n6309), .Z(n4862) );
  XOR U9410 ( .A(n8485), .B(n8486), .Z(n6309) );
  XNOR U9411 ( .A(n3273), .B(n4760), .Z(n8486) );
  XNOR U9412 ( .A(n8487), .B(n8488), .Z(n4760) );
  NOR U9413 ( .A(n8489), .B(n8490), .Z(n8487) );
  XNOR U9414 ( .A(n8491), .B(n8492), .Z(n3273) );
  NOR U9415 ( .A(n8493), .B(n8494), .Z(n8491) );
  XOR U9416 ( .A(n5602), .B(n8495), .Z(n8485) );
  XOR U9417 ( .A(n8496), .B(n2522), .Z(n8495) );
  XOR U9418 ( .A(n8497), .B(n8498), .Z(n2522) );
  ANDN U9419 ( .B(n8499), .A(n8500), .Z(n8497) );
  XNOR U9420 ( .A(n8501), .B(n8502), .Z(n5602) );
  NOR U9421 ( .A(n8503), .B(n8504), .Z(n8501) );
  XOR U9422 ( .A(n8505), .B(n8506), .Z(n5892) );
  XNOR U9423 ( .A(n3861), .B(n5167), .Z(n8506) );
  XNOR U9424 ( .A(n8507), .B(n8508), .Z(n5167) );
  ANDN U9425 ( .B(n8509), .A(n8510), .Z(n8507) );
  XNOR U9426 ( .A(n8511), .B(n8512), .Z(n3861) );
  ANDN U9427 ( .B(n8513), .A(n8514), .Z(n8511) );
  XNOR U9428 ( .A(n6370), .B(n8515), .Z(n8505) );
  XNOR U9429 ( .A(n1757), .B(n8516), .Z(n8515) );
  XNOR U9430 ( .A(n8517), .B(n8518), .Z(n1757) );
  NOR U9431 ( .A(n8519), .B(n8520), .Z(n8517) );
  XNOR U9432 ( .A(n8521), .B(n8522), .Z(n6370) );
  AND U9433 ( .A(n8523), .B(n8524), .Z(n8521) );
  XNOR U9434 ( .A(n8525), .B(n6024), .Z(out[1040]) );
  XOR U9435 ( .A(n7518), .B(n2412), .Z(n6024) );
  XNOR U9436 ( .A(n8526), .B(n8527), .Z(n7518) );
  NOR U9437 ( .A(n8528), .B(n8529), .Z(n8526) );
  NOR U9438 ( .A(n6348), .B(n1140), .Z(n8525) );
  XOR U9439 ( .A(n1907), .B(n8530), .Z(n1140) );
  IV U9440 ( .A(n4176), .Z(n1907) );
  XNOR U9441 ( .A(n7305), .B(n6158), .Z(n4176) );
  XOR U9442 ( .A(n8531), .B(n8532), .Z(n6158) );
  XNOR U9443 ( .A(n4628), .B(n1988), .Z(n8532) );
  XOR U9444 ( .A(n8533), .B(n8534), .Z(n1988) );
  AND U9445 ( .A(n7469), .B(n7470), .Z(n8533) );
  XOR U9446 ( .A(n8535), .B(n8536), .Z(n4628) );
  NOR U9447 ( .A(n7478), .B(n7477), .Z(n8535) );
  XNOR U9448 ( .A(n6072), .B(n8537), .Z(n8531) );
  XNOR U9449 ( .A(n5596), .B(n3851), .Z(n8537) );
  XOR U9450 ( .A(n8538), .B(n8539), .Z(n3851) );
  NOR U9451 ( .A(n8540), .B(n7464), .Z(n8538) );
  XNOR U9452 ( .A(n8541), .B(n8542), .Z(n5596) );
  AND U9453 ( .A(n7473), .B(n7475), .Z(n8541) );
  XNOR U9454 ( .A(n8543), .B(n8544), .Z(n6072) );
  ANDN U9455 ( .B(n7460), .A(n8545), .Z(n8543) );
  XOR U9456 ( .A(n8546), .B(n8547), .Z(n7305) );
  XNOR U9457 ( .A(n4990), .B(n8548), .Z(n8547) );
  XOR U9458 ( .A(n8549), .B(n7400), .Z(n4990) );
  NOR U9459 ( .A(n8460), .B(n8550), .Z(n8549) );
  IV U9460 ( .A(n8551), .Z(n8460) );
  XOR U9461 ( .A(n2249), .B(n8552), .Z(n8546) );
  XNOR U9462 ( .A(n3594), .B(n6119), .Z(n8552) );
  XOR U9463 ( .A(n8553), .B(n7387), .Z(n6119) );
  ANDN U9464 ( .B(n8554), .A(n8465), .Z(n8553) );
  IV U9465 ( .A(n8555), .Z(n8465) );
  XNOR U9466 ( .A(n8556), .B(n7392), .Z(n3594) );
  XOR U9467 ( .A(n8558), .B(n7383), .Z(n2249) );
  NOR U9468 ( .A(n8470), .B(n8559), .Z(n8558) );
  XOR U9469 ( .A(n2492), .B(n8560), .Z(n6348) );
  XNOR U9470 ( .A(n5897), .B(n6313), .Z(n2492) );
  XOR U9471 ( .A(n8561), .B(n8562), .Z(n6313) );
  XOR U9472 ( .A(n3276), .B(n4792), .Z(n8562) );
  XNOR U9473 ( .A(n8563), .B(n8564), .Z(n4792) );
  ANDN U9474 ( .B(n8565), .A(n8512), .Z(n8563) );
  XNOR U9475 ( .A(n8566), .B(n8567), .Z(n3276) );
  NOR U9476 ( .A(n8518), .B(n8568), .Z(n8566) );
  IV U9477 ( .A(n8569), .Z(n8518) );
  XNOR U9478 ( .A(n5298), .B(n8570), .Z(n8561) );
  XNOR U9479 ( .A(n8571), .B(n2529), .Z(n8570) );
  XNOR U9480 ( .A(n8572), .B(n8573), .Z(n2529) );
  XNOR U9481 ( .A(n8576), .B(n8577), .Z(n5298) );
  XOR U9482 ( .A(n8579), .B(n8580), .Z(n5897) );
  XOR U9483 ( .A(n3867), .B(n5170), .Z(n8580) );
  XNOR U9484 ( .A(n8581), .B(n8582), .Z(n5170) );
  XOR U9485 ( .A(n8584), .B(n8585), .Z(n3867) );
  ANDN U9486 ( .B(n8586), .A(n6428), .Z(n8584) );
  IV U9487 ( .A(n8587), .Z(n6428) );
  XNOR U9488 ( .A(n8588), .B(n8589), .Z(n8579) );
  XNOR U9489 ( .A(n4275), .B(n1763), .Z(n8589) );
  XNOR U9490 ( .A(n8590), .B(n8591), .Z(n1763) );
  ANDN U9491 ( .B(n8592), .A(n8593), .Z(n8590) );
  XNOR U9492 ( .A(n8594), .B(n8595), .Z(n4275) );
  NOR U9493 ( .A(n8596), .B(n6445), .Z(n8594) );
  XOR U9494 ( .A(n8597), .B(n4192), .Z(out[103]) );
  XOR U9495 ( .A(n8598), .B(n2558), .Z(n4192) );
  XNOR U9496 ( .A(n7848), .B(n8599), .Z(n2558) );
  XOR U9497 ( .A(n8600), .B(n8601), .Z(n7848) );
  XNOR U9498 ( .A(n4375), .B(n2180), .Z(n8601) );
  XNOR U9499 ( .A(n8602), .B(n7931), .Z(n2180) );
  IV U9500 ( .A(n8603), .Z(n7931) );
  ANDN U9501 ( .B(n8604), .A(n8605), .Z(n8602) );
  XNOR U9502 ( .A(n8606), .B(n7921), .Z(n4375) );
  IV U9503 ( .A(n8607), .Z(n7921) );
  XOR U9504 ( .A(n6006), .B(n8610), .Z(n8600) );
  XOR U9505 ( .A(n5546), .B(n3796), .Z(n8610) );
  XOR U9506 ( .A(n8611), .B(n7926), .Z(n3796) );
  ANDN U9507 ( .B(n8612), .A(n8613), .Z(n8611) );
  XNOR U9508 ( .A(n8614), .B(n8615), .Z(n5546) );
  NOR U9509 ( .A(n8616), .B(n8617), .Z(n8614) );
  XOR U9510 ( .A(n8618), .B(n7935), .Z(n6006) );
  ANDN U9511 ( .B(n8619), .A(n8620), .Z(n8618) );
  AND U9512 ( .A(n3558), .B(n3560), .Z(n8597) );
  XOR U9513 ( .A(n2332), .B(n8621), .Z(n3560) );
  XNOR U9514 ( .A(n6208), .B(n8622), .Z(n2332) );
  XOR U9515 ( .A(n8623), .B(n8624), .Z(n6208) );
  XOR U9516 ( .A(n3191), .B(n6638), .Z(n8624) );
  XOR U9517 ( .A(n8625), .B(n8626), .Z(n6638) );
  NOR U9518 ( .A(n8627), .B(n8628), .Z(n8625) );
  XOR U9519 ( .A(n8629), .B(n8630), .Z(n3191) );
  NOR U9520 ( .A(n8631), .B(n8632), .Z(n8629) );
  XOR U9521 ( .A(n5502), .B(n8633), .Z(n8623) );
  XOR U9522 ( .A(n8178), .B(n2365), .Z(n8633) );
  XNOR U9523 ( .A(n8634), .B(n8635), .Z(n2365) );
  NOR U9524 ( .A(n8636), .B(n8637), .Z(n8634) );
  XNOR U9525 ( .A(n8638), .B(n8639), .Z(n8178) );
  NOR U9526 ( .A(n8640), .B(n8641), .Z(n8638) );
  XNOR U9527 ( .A(n8642), .B(n8643), .Z(n5502) );
  ANDN U9528 ( .B(n8644), .A(n8645), .Z(n8642) );
  XOR U9529 ( .A(n7333), .B(n3206), .Z(n3558) );
  XOR U9530 ( .A(n8646), .B(n8647), .Z(n3206) );
  XNOR U9531 ( .A(n8648), .B(n8649), .Z(n7333) );
  NOR U9532 ( .A(n8650), .B(n8651), .Z(n8648) );
  XOR U9533 ( .A(n8652), .B(n6029), .Z(out[1039]) );
  XOR U9534 ( .A(n7596), .B(n2421), .Z(n6029) );
  IV U9535 ( .A(n3217), .Z(n2421) );
  XNOR U9536 ( .A(n8653), .B(n8654), .Z(n7596) );
  ANDN U9537 ( .B(n8655), .A(n8656), .Z(n8653) );
  AND U9538 ( .A(n1144), .B(n1143), .Z(n8652) );
  XOR U9539 ( .A(n8657), .B(n2502), .Z(n1143) );
  XOR U9540 ( .A(n5907), .B(n6317), .Z(n2502) );
  XOR U9541 ( .A(n8658), .B(n8659), .Z(n6317) );
  XNOR U9542 ( .A(n3280), .B(n4816), .Z(n8659) );
  XNOR U9543 ( .A(n8660), .B(n6429), .Z(n4816) );
  ANDN U9544 ( .B(n6430), .A(n8585), .Z(n8660) );
  XNOR U9545 ( .A(n8661), .B(n6434), .Z(n3280) );
  ANDN U9546 ( .B(n8591), .A(n8662), .Z(n8661) );
  XNOR U9547 ( .A(n5301), .B(n8663), .Z(n8658) );
  XOR U9548 ( .A(n6423), .B(n2538), .Z(n8663) );
  XNOR U9549 ( .A(n8664), .B(n6438), .Z(n2538) );
  ANDN U9550 ( .B(n6439), .A(n8665), .Z(n8664) );
  XNOR U9551 ( .A(n8666), .B(n6442), .Z(n6423) );
  ANDN U9552 ( .B(n8582), .A(n6443), .Z(n8666) );
  XOR U9553 ( .A(n8667), .B(n6446), .Z(n5301) );
  AND U9554 ( .A(n6447), .B(n8595), .Z(n8667) );
  XOR U9555 ( .A(n8668), .B(n8669), .Z(n5907) );
  XOR U9556 ( .A(n3875), .B(n5172), .Z(n8669) );
  XNOR U9557 ( .A(n8670), .B(n8671), .Z(n5172) );
  NOR U9558 ( .A(n8672), .B(n6467), .Z(n8670) );
  XOR U9559 ( .A(n8673), .B(n8674), .Z(n3875) );
  ANDN U9560 ( .B(n6454), .A(n8675), .Z(n8673) );
  XOR U9561 ( .A(n4277), .B(n8676), .Z(n8668) );
  XNOR U9562 ( .A(n1766), .B(n8677), .Z(n8676) );
  XOR U9563 ( .A(n8678), .B(n8679), .Z(n1766) );
  ANDN U9564 ( .B(n6458), .A(n8680), .Z(n8678) );
  XNOR U9565 ( .A(n8681), .B(n8682), .Z(n4277) );
  NOR U9566 ( .A(n6471), .B(n8683), .Z(n8681) );
  XOR U9567 ( .A(n1911), .B(n8684), .Z(n1144) );
  IV U9568 ( .A(n4181), .Z(n1911) );
  XNOR U9569 ( .A(n7378), .B(n6163), .Z(n4181) );
  XOR U9570 ( .A(n8685), .B(n8686), .Z(n6163) );
  XNOR U9571 ( .A(n4672), .B(n1991), .Z(n8686) );
  XOR U9572 ( .A(n8687), .B(n8688), .Z(n1991) );
  NOR U9573 ( .A(n7544), .B(n7543), .Z(n8687) );
  XNOR U9574 ( .A(n8689), .B(n8690), .Z(n4672) );
  NOR U9575 ( .A(n7552), .B(n7551), .Z(n8689) );
  XNOR U9576 ( .A(n6077), .B(n8691), .Z(n8685) );
  XOR U9577 ( .A(n5600), .B(n3854), .Z(n8691) );
  XOR U9578 ( .A(n8692), .B(n8693), .Z(n3854) );
  NOR U9579 ( .A(n7540), .B(n7538), .Z(n8692) );
  XNOR U9580 ( .A(n8694), .B(n8695), .Z(n5600) );
  ANDN U9581 ( .B(n7548), .A(n7547), .Z(n8694) );
  XNOR U9582 ( .A(n8696), .B(n8697), .Z(n6077) );
  ANDN U9583 ( .B(n7534), .A(n8698), .Z(n8696) );
  XOR U9584 ( .A(n8699), .B(n8700), .Z(n7378) );
  XOR U9585 ( .A(n4993), .B(n8701), .Z(n8700) );
  XOR U9586 ( .A(n8702), .B(n8703), .Z(n4993) );
  ANDN U9587 ( .B(n8536), .A(n8704), .Z(n8702) );
  XNOR U9588 ( .A(n2256), .B(n8705), .Z(n8699) );
  XNOR U9589 ( .A(n3596), .B(n6174), .Z(n8705) );
  XOR U9590 ( .A(n8706), .B(n7465), .Z(n6174) );
  ANDN U9591 ( .B(n8539), .A(n8707), .Z(n8706) );
  XNOR U9592 ( .A(n8708), .B(n7471), .Z(n3596) );
  ANDN U9593 ( .B(n8534), .A(n8709), .Z(n8708) );
  XNOR U9594 ( .A(n8710), .B(n7462), .Z(n2256) );
  ANDN U9595 ( .B(n8711), .A(n8544), .Z(n8710) );
  XNOR U9596 ( .A(n8712), .B(n6034), .Z(out[1038]) );
  IV U9597 ( .A(n6357), .Z(n6034) );
  XOR U9598 ( .A(n5543), .B(n7635), .Z(n6357) );
  XOR U9599 ( .A(n8713), .B(n8714), .Z(n7635) );
  ANDN U9600 ( .B(n8715), .A(n8716), .Z(n8713) );
  XNOR U9601 ( .A(n8717), .B(n8718), .Z(n5543) );
  ANDN U9602 ( .B(n1147), .A(n1148), .Z(n8712) );
  XOR U9603 ( .A(n3708), .B(n8719), .Z(n1148) );
  IV U9604 ( .A(n1919), .Z(n3708) );
  XNOR U9605 ( .A(n7456), .B(n6168), .Z(n1919) );
  XOR U9606 ( .A(n8720), .B(n8721), .Z(n6168) );
  XNOR U9607 ( .A(n4711), .B(n1994), .Z(n8721) );
  XOR U9608 ( .A(n8722), .B(n8723), .Z(n1994) );
  ANDN U9609 ( .B(n7620), .A(n7622), .Z(n8722) );
  XOR U9610 ( .A(n8724), .B(n8725), .Z(n4711) );
  ANDN U9611 ( .B(n7628), .A(n7629), .Z(n8724) );
  XOR U9612 ( .A(n6082), .B(n8726), .Z(n8720) );
  XOR U9613 ( .A(n5296), .B(n3858), .Z(n8726) );
  XNOR U9614 ( .A(n8727), .B(n8728), .Z(n3858) );
  XOR U9615 ( .A(n8729), .B(n8730), .Z(n5296) );
  ANDN U9616 ( .B(n7626), .A(n7624), .Z(n8729) );
  XOR U9617 ( .A(n8731), .B(n8732), .Z(n6082) );
  ANDN U9618 ( .B(n7611), .A(n7612), .Z(n8731) );
  XOR U9619 ( .A(n8733), .B(n8734), .Z(n7456) );
  XNOR U9620 ( .A(n4996), .B(n8735), .Z(n8734) );
  XNOR U9621 ( .A(n8736), .B(n8737), .Z(n4996) );
  NOR U9622 ( .A(n8738), .B(n8739), .Z(n8736) );
  XNOR U9623 ( .A(n2265), .B(n8740), .Z(n8733) );
  XOR U9624 ( .A(n3598), .B(n6229), .Z(n8740) );
  XOR U9625 ( .A(n8741), .B(n7539), .Z(n6229) );
  AND U9626 ( .A(n8693), .B(n8742), .Z(n8741) );
  XNOR U9627 ( .A(n8743), .B(n7545), .Z(n3598) );
  ANDN U9628 ( .B(n8688), .A(n8744), .Z(n8743) );
  XNOR U9629 ( .A(n8745), .B(n7536), .Z(n2265) );
  ANDN U9630 ( .B(n8746), .A(n8697), .Z(n8745) );
  XOR U9631 ( .A(n2506), .B(n8747), .Z(n1147) );
  IV U9632 ( .A(n4878), .Z(n2506) );
  XNOR U9633 ( .A(n5912), .B(n6325), .Z(n4878) );
  XOR U9634 ( .A(n8748), .B(n8749), .Z(n6325) );
  XNOR U9635 ( .A(n3285), .B(n4841), .Z(n8749) );
  XOR U9636 ( .A(n8750), .B(n6455), .Z(n4841) );
  NOR U9637 ( .A(n6456), .B(n8674), .Z(n8750) );
  XNOR U9638 ( .A(n8751), .B(n6459), .Z(n3285) );
  ANDN U9639 ( .B(n8679), .A(n8752), .Z(n8751) );
  XNOR U9640 ( .A(n5305), .B(n8753), .Z(n8748) );
  XNOR U9641 ( .A(n6449), .B(n2547), .Z(n8753) );
  XNOR U9642 ( .A(n8754), .B(n6464), .Z(n2547) );
  IV U9643 ( .A(n8756), .Z(n6465) );
  XOR U9644 ( .A(n8757), .B(n8758), .Z(n6449) );
  NOR U9645 ( .A(n6468), .B(n8671), .Z(n8757) );
  XOR U9646 ( .A(n8759), .B(n6472), .Z(n5305) );
  ANDN U9647 ( .B(n6473), .A(n8682), .Z(n8759) );
  IV U9648 ( .A(n8760), .Z(n8682) );
  XOR U9649 ( .A(n8761), .B(n8762), .Z(n5912) );
  XNOR U9650 ( .A(n3879), .B(n5175), .Z(n8762) );
  XNOR U9651 ( .A(n8763), .B(n8764), .Z(n5175) );
  ANDN U9652 ( .B(n8765), .A(n6494), .Z(n8763) );
  XOR U9653 ( .A(n8766), .B(n8767), .Z(n3879) );
  ANDN U9654 ( .B(n8768), .A(n6481), .Z(n8766) );
  XOR U9655 ( .A(n4285), .B(n8769), .Z(n8761) );
  XOR U9656 ( .A(n1774), .B(n8770), .Z(n8769) );
  XNOR U9657 ( .A(n8771), .B(n8772), .Z(n1774) );
  NOR U9658 ( .A(n8773), .B(n6485), .Z(n8771) );
  XOR U9659 ( .A(n8774), .B(n8775), .Z(n4285) );
  ANDN U9660 ( .B(n8776), .A(n8777), .Z(n8774) );
  XNOR U9661 ( .A(n8778), .B(n6039), .Z(out[1037]) );
  IV U9662 ( .A(n6362), .Z(n6039) );
  XNOR U9663 ( .A(n2432), .B(n7739), .Z(n6362) );
  XOR U9664 ( .A(n8779), .B(n8780), .Z(n7739) );
  ANDN U9665 ( .B(n8781), .A(n8782), .Z(n8779) );
  AND U9666 ( .A(n1153), .B(n1151), .Z(n8778) );
  XNOR U9667 ( .A(n2513), .B(n8785), .Z(n1151) );
  XOR U9668 ( .A(n5917), .B(n6331), .Z(n2513) );
  XNOR U9669 ( .A(n8786), .B(n8787), .Z(n6331) );
  XOR U9670 ( .A(n2552), .B(n5310), .Z(n8787) );
  XOR U9671 ( .A(n8788), .B(n6499), .Z(n5310) );
  NOR U9672 ( .A(n6500), .B(n8775), .Z(n8788) );
  NOR U9673 ( .A(n8790), .B(n8791), .Z(n8789) );
  XOR U9674 ( .A(n3288), .B(n8792), .Z(n8786) );
  XOR U9675 ( .A(n4873), .B(n6476), .Z(n8792) );
  XOR U9676 ( .A(n8793), .B(n6495), .Z(n6476) );
  ANDN U9677 ( .B(n6496), .A(n8764), .Z(n8793) );
  XOR U9678 ( .A(n8794), .B(n6483), .Z(n4873) );
  ANDN U9679 ( .B(n8767), .A(n6482), .Z(n8794) );
  XOR U9680 ( .A(n8795), .B(n6486), .Z(n3288) );
  XOR U9681 ( .A(n8796), .B(n8797), .Z(n5917) );
  XNOR U9682 ( .A(n3884), .B(n5178), .Z(n8797) );
  XNOR U9683 ( .A(n8798), .B(n8799), .Z(n5178) );
  ANDN U9684 ( .B(n8800), .A(n6521), .Z(n8798) );
  XOR U9685 ( .A(n8801), .B(n8802), .Z(n3884) );
  ANDN U9686 ( .B(n8803), .A(n6507), .Z(n8801) );
  XNOR U9687 ( .A(n4287), .B(n8804), .Z(n8796) );
  XOR U9688 ( .A(n1779), .B(n8805), .Z(n8804) );
  XNOR U9689 ( .A(n8806), .B(n8807), .Z(n1779) );
  ANDN U9690 ( .B(n8808), .A(n8809), .Z(n8806) );
  XOR U9691 ( .A(n8810), .B(n8811), .Z(n4287) );
  NOR U9692 ( .A(n6525), .B(n8812), .Z(n8810) );
  XOR U9693 ( .A(n3714), .B(n8813), .Z(n1153) );
  IV U9694 ( .A(n1923), .Z(n3714) );
  XNOR U9695 ( .A(n7530), .B(n6178), .Z(n1923) );
  XOR U9696 ( .A(n8814), .B(n8815), .Z(n6178) );
  XNOR U9697 ( .A(n4735), .B(n1997), .Z(n8815) );
  XNOR U9698 ( .A(n8816), .B(n8817), .Z(n1997) );
  AND U9699 ( .A(n7696), .B(n7694), .Z(n8816) );
  XNOR U9700 ( .A(n8818), .B(n8819), .Z(n4735) );
  ANDN U9701 ( .B(n7702), .A(n8820), .Z(n8818) );
  XOR U9702 ( .A(n6087), .B(n8821), .Z(n8814) );
  XOR U9703 ( .A(n5300), .B(n3864), .Z(n8821) );
  XOR U9704 ( .A(n8822), .B(n8823), .Z(n3864) );
  IV U9705 ( .A(n8824), .Z(n7690) );
  ANDN U9706 ( .B(n7699), .A(n7698), .Z(n8825) );
  XNOR U9707 ( .A(n8827), .B(n8828), .Z(n6087) );
  NOR U9708 ( .A(n7687), .B(n7685), .Z(n8827) );
  XOR U9709 ( .A(n8829), .B(n8830), .Z(n7530) );
  XOR U9710 ( .A(n4999), .B(n8831), .Z(n8830) );
  XOR U9711 ( .A(n8832), .B(n7630), .Z(n4999) );
  NOR U9712 ( .A(n8833), .B(n8725), .Z(n8832) );
  XNOR U9713 ( .A(n2270), .B(n8834), .Z(n8829) );
  XOR U9714 ( .A(n3601), .B(n6276), .Z(n8834) );
  XOR U9715 ( .A(n8835), .B(n7616), .Z(n6276) );
  ANDN U9716 ( .B(n8836), .A(n8728), .Z(n8835) );
  IV U9717 ( .A(n8837), .Z(n8728) );
  XOR U9718 ( .A(n8838), .B(n7621), .Z(n3601) );
  ANDN U9719 ( .B(n8723), .A(n8839), .Z(n8838) );
  XOR U9720 ( .A(n8840), .B(n7613), .Z(n2270) );
  ANDN U9721 ( .B(n8732), .A(n8841), .Z(n8840) );
  XOR U9722 ( .A(n8842), .B(n6044), .Z(out[1036]) );
  XNOR U9723 ( .A(n7796), .B(n2440), .Z(n6044) );
  XNOR U9724 ( .A(n8845), .B(n8846), .Z(n7796) );
  ANDN U9725 ( .B(n8847), .A(n8848), .Z(n8845) );
  ANDN U9726 ( .B(n1157), .A(n1155), .Z(n8842) );
  XOR U9727 ( .A(n2520), .B(n8849), .Z(n1155) );
  IV U9728 ( .A(n4885), .Z(n2520) );
  XNOR U9729 ( .A(n5922), .B(n6334), .Z(n4885) );
  XOR U9730 ( .A(n8850), .B(n8851), .Z(n6334) );
  XOR U9731 ( .A(n3292), .B(n4912), .Z(n8851) );
  XOR U9732 ( .A(n8852), .B(n6508), .Z(n4912) );
  NOR U9733 ( .A(n6509), .B(n8802), .Z(n8852) );
  XNOR U9734 ( .A(n8853), .B(n6513), .Z(n3292) );
  ANDN U9735 ( .B(n6512), .A(n8807), .Z(n8853) );
  IV U9736 ( .A(n8854), .Z(n8807) );
  XNOR U9737 ( .A(n5318), .B(n8855), .Z(n8850) );
  XNOR U9738 ( .A(n6502), .B(n2561), .Z(n8855) );
  XNOR U9739 ( .A(n8856), .B(n6519), .Z(n2561) );
  ANDN U9740 ( .B(n6518), .A(n8857), .Z(n8856) );
  XOR U9741 ( .A(n8858), .B(n6522), .Z(n6502) );
  ANDN U9742 ( .B(n6523), .A(n8799), .Z(n8858) );
  IV U9743 ( .A(n8859), .Z(n8799) );
  XNOR U9744 ( .A(n8860), .B(n6526), .Z(n5318) );
  ANDN U9745 ( .B(n6527), .A(n8861), .Z(n8860) );
  XOR U9746 ( .A(n8862), .B(n8863), .Z(n5922) );
  XNOR U9747 ( .A(n3888), .B(n5186), .Z(n8863) );
  XOR U9748 ( .A(n8864), .B(n8865), .Z(n5186) );
  AND U9749 ( .A(n8866), .B(n6547), .Z(n8864) );
  XNOR U9750 ( .A(n8867), .B(n8868), .Z(n3888) );
  ANDN U9751 ( .B(n8869), .A(n6534), .Z(n8867) );
  XNOR U9752 ( .A(n4289), .B(n8870), .Z(n8862) );
  XOR U9753 ( .A(n1784), .B(n8871), .Z(n8870) );
  XOR U9754 ( .A(n8872), .B(n8873), .Z(n1784) );
  ANDN U9755 ( .B(n8874), .A(n6538), .Z(n8872) );
  IV U9756 ( .A(n8875), .Z(n6538) );
  XNOR U9757 ( .A(n8876), .B(n8877), .Z(n4289) );
  ANDN U9758 ( .B(n8878), .A(n8879), .Z(n8876) );
  XOR U9759 ( .A(n1928), .B(n8880), .Z(n1157) );
  IV U9760 ( .A(n3719), .Z(n1928) );
  XNOR U9761 ( .A(n7607), .B(n6183), .Z(n3719) );
  XOR U9762 ( .A(n8881), .B(n8882), .Z(n6183) );
  XNOR U9763 ( .A(n4759), .B(n2004), .Z(n8882) );
  XNOR U9764 ( .A(n8883), .B(n8884), .Z(n2004) );
  AND U9765 ( .A(n7774), .B(n7772), .Z(n8883) );
  XNOR U9766 ( .A(n8885), .B(n8886), .Z(n4759) );
  NOR U9767 ( .A(n7781), .B(n7780), .Z(n8885) );
  XOR U9768 ( .A(n6092), .B(n8887), .Z(n8881) );
  XOR U9769 ( .A(n5304), .B(n3868), .Z(n8887) );
  XOR U9770 ( .A(n8888), .B(n8889), .Z(n3868) );
  ANDN U9771 ( .B(n7767), .A(n7768), .Z(n8888) );
  XOR U9772 ( .A(n8890), .B(n8891), .Z(n5304) );
  ANDN U9773 ( .B(n7776), .A(n8892), .Z(n8890) );
  XOR U9774 ( .A(n8893), .B(n8894), .Z(n6092) );
  ANDN U9775 ( .B(n7763), .A(n8895), .Z(n8893) );
  XOR U9776 ( .A(n8896), .B(n8897), .Z(n7607) );
  XNOR U9777 ( .A(n5002), .B(n8898), .Z(n8897) );
  XNOR U9778 ( .A(n8899), .B(n7704), .Z(n5002) );
  ANDN U9779 ( .B(n8900), .A(n8819), .Z(n8899) );
  XOR U9780 ( .A(n2277), .B(n8901), .Z(n8896) );
  XOR U9781 ( .A(n3404), .B(n6321), .Z(n8901) );
  XOR U9782 ( .A(n8902), .B(n7691), .Z(n6321) );
  ANDN U9783 ( .B(n8823), .A(n8903), .Z(n8902) );
  XNOR U9784 ( .A(n8904), .B(n7695), .Z(n3404) );
  ANDN U9785 ( .B(n8905), .A(n8817), .Z(n8904) );
  XOR U9786 ( .A(n8906), .B(n7686), .Z(n2277) );
  XOR U9787 ( .A(n8908), .B(n6049), .Z(out[1035]) );
  XOR U9788 ( .A(n7879), .B(n2447), .Z(n6049) );
  IV U9789 ( .A(n3234), .Z(n2447) );
  XOR U9790 ( .A(n8911), .B(n8912), .Z(n7879) );
  AND U9791 ( .A(n8913), .B(n8914), .Z(n8911) );
  ANDN U9792 ( .B(n1161), .A(n1159), .Z(n8908) );
  XOR U9793 ( .A(n2527), .B(n8915), .Z(n1159) );
  IV U9794 ( .A(n4889), .Z(n2527) );
  XNOR U9795 ( .A(n5926), .B(n6338), .Z(n4889) );
  XOR U9796 ( .A(n8916), .B(n8917), .Z(n6338) );
  XNOR U9797 ( .A(n3295), .B(n4950), .Z(n8917) );
  XOR U9798 ( .A(n8918), .B(n6535), .Z(n4950) );
  NOR U9799 ( .A(n6536), .B(n8868), .Z(n8918) );
  XOR U9800 ( .A(n8919), .B(n6539), .Z(n3295) );
  XNOR U9801 ( .A(n5322), .B(n8920), .Z(n8916) );
  XNOR U9802 ( .A(n6529), .B(n2568), .Z(n8920) );
  XOR U9803 ( .A(n8921), .B(n6544), .Z(n2568) );
  XNOR U9804 ( .A(n8923), .B(n6548), .Z(n6529) );
  ANDN U9805 ( .B(n6549), .A(n8865), .Z(n8923) );
  XOR U9806 ( .A(n8924), .B(n6553), .Z(n5322) );
  IV U9807 ( .A(n8925), .Z(n6553) );
  NOR U9808 ( .A(n6552), .B(n8877), .Z(n8924) );
  XOR U9809 ( .A(n8926), .B(n8927), .Z(n5926) );
  XNOR U9810 ( .A(n3892), .B(n5189), .Z(n8927) );
  XOR U9811 ( .A(n8928), .B(n8929), .Z(n5189) );
  NOR U9812 ( .A(n6573), .B(n8930), .Z(n8928) );
  IV U9813 ( .A(n8931), .Z(n6573) );
  XOR U9814 ( .A(n8932), .B(n8933), .Z(n3892) );
  ANDN U9815 ( .B(n6560), .A(n8934), .Z(n8932) );
  XOR U9816 ( .A(n4292), .B(n8935), .Z(n8926) );
  XNOR U9817 ( .A(n1789), .B(n8936), .Z(n8935) );
  XOR U9818 ( .A(n8937), .B(n8938), .Z(n1789) );
  NOR U9819 ( .A(n6564), .B(n8939), .Z(n8937) );
  IV U9820 ( .A(n8940), .Z(n6564) );
  XNOR U9821 ( .A(n8941), .B(n8942), .Z(n4292) );
  ANDN U9822 ( .B(n6577), .A(n8943), .Z(n8941) );
  XOR U9823 ( .A(n1932), .B(n8944), .Z(n1161) );
  IV U9824 ( .A(n3726), .Z(n1932) );
  XNOR U9825 ( .A(n7681), .B(n6188), .Z(n3726) );
  XOR U9826 ( .A(n8945), .B(n8946), .Z(n6188) );
  XNOR U9827 ( .A(n4789), .B(n2008), .Z(n8946) );
  XOR U9828 ( .A(n8947), .B(n8948), .Z(n2008) );
  ANDN U9829 ( .B(n7836), .A(n7837), .Z(n8947) );
  XNOR U9830 ( .A(n8949), .B(n8950), .Z(n4789) );
  XNOR U9831 ( .A(n6097), .B(n8951), .Z(n8945) );
  XOR U9832 ( .A(n5308), .B(n3877), .Z(n8951) );
  XNOR U9833 ( .A(n8952), .B(n8953), .Z(n3877) );
  ANDN U9834 ( .B(n7833), .A(n7831), .Z(n8952) );
  XNOR U9835 ( .A(n8954), .B(n8955), .Z(n5308) );
  XOR U9836 ( .A(n8956), .B(n8957), .Z(n6097) );
  NOR U9837 ( .A(n7829), .B(n7827), .Z(n8956) );
  XOR U9838 ( .A(n8958), .B(n8959), .Z(n7681) );
  XNOR U9839 ( .A(n5005), .B(n8960), .Z(n8959) );
  XNOR U9840 ( .A(n8961), .B(n7782), .Z(n5005) );
  ANDN U9841 ( .B(n8962), .A(n8886), .Z(n8961) );
  XOR U9842 ( .A(n2284), .B(n8963), .Z(n8958) );
  XOR U9843 ( .A(n3407), .B(n6373), .Z(n8963) );
  XNOR U9844 ( .A(n8964), .B(n7769), .Z(n6373) );
  NOR U9845 ( .A(n8965), .B(n8889), .Z(n8964) );
  XNOR U9846 ( .A(n8966), .B(n7773), .Z(n3407) );
  IV U9847 ( .A(n8967), .Z(n7773) );
  NOR U9848 ( .A(n8884), .B(n8968), .Z(n8966) );
  XOR U9849 ( .A(n8969), .B(n7764), .Z(n2284) );
  XNOR U9850 ( .A(n8971), .B(n6055), .Z(out[1034]) );
  XOR U9851 ( .A(n7949), .B(n2454), .Z(n6055) );
  IV U9852 ( .A(n3238), .Z(n2454) );
  XOR U9853 ( .A(n8974), .B(n8975), .Z(n7949) );
  ANDN U9854 ( .B(n8976), .A(n8977), .Z(n8974) );
  ANDN U9855 ( .B(n1163), .A(n1165), .Z(n8971) );
  XOR U9856 ( .A(n1937), .B(n8978), .Z(n1165) );
  IV U9857 ( .A(n3733), .Z(n1937) );
  XNOR U9858 ( .A(n7759), .B(n6193), .Z(n3733) );
  XOR U9859 ( .A(n8979), .B(n8980), .Z(n6193) );
  XOR U9860 ( .A(n4815), .B(n2011), .Z(n8980) );
  XOR U9861 ( .A(n8981), .B(n8982), .Z(n2011) );
  XOR U9862 ( .A(n8983), .B(n8984), .Z(n4815) );
  XNOR U9863 ( .A(n6102), .B(n8985), .Z(n8979) );
  XNOR U9864 ( .A(n5317), .B(n3882), .Z(n8985) );
  XNOR U9865 ( .A(n8986), .B(n8987), .Z(n3882) );
  IV U9866 ( .A(n8988), .Z(n7899) );
  XNOR U9867 ( .A(n8989), .B(n8990), .Z(n5317) );
  ANDN U9868 ( .B(n7907), .A(n7909), .Z(n8989) );
  XOR U9869 ( .A(n8991), .B(n8992), .Z(n6102) );
  NOR U9870 ( .A(n7896), .B(n7894), .Z(n8991) );
  XOR U9871 ( .A(n8993), .B(n8994), .Z(n7759) );
  XNOR U9872 ( .A(n5008), .B(n8995), .Z(n8994) );
  XOR U9873 ( .A(n8996), .B(n7846), .Z(n5008) );
  ANDN U9874 ( .B(n8997), .A(n8950), .Z(n8996) );
  XOR U9875 ( .A(n2291), .B(n8998), .Z(n8993) );
  XOR U9876 ( .A(n3409), .B(n6414), .Z(n8998) );
  XOR U9877 ( .A(n8999), .B(n7832), .Z(n6414) );
  ANDN U9878 ( .B(n9000), .A(n8953), .Z(n8999) );
  XNOR U9879 ( .A(n9001), .B(n9002), .Z(n3409) );
  ANDN U9880 ( .B(n8948), .A(n9003), .Z(n9001) );
  XOR U9881 ( .A(n9004), .B(n7828), .Z(n2291) );
  XNOR U9882 ( .A(n3514), .B(n9006), .Z(n1163) );
  XNOR U9883 ( .A(n5932), .B(n6342), .Z(n3514) );
  XOR U9884 ( .A(n9007), .B(n9008), .Z(n6342) );
  XNOR U9885 ( .A(n3300), .B(n4987), .Z(n9008) );
  XOR U9886 ( .A(n9009), .B(n6562), .Z(n4987) );
  XNOR U9887 ( .A(n9010), .B(n6565), .Z(n3300) );
  AND U9888 ( .A(n8938), .B(n6566), .Z(n9010) );
  XOR U9889 ( .A(n5327), .B(n9011), .Z(n9007) );
  XNOR U9890 ( .A(n6555), .B(n2575), .Z(n9011) );
  XOR U9891 ( .A(n9012), .B(n6570), .Z(n2575) );
  XNOR U9892 ( .A(n9014), .B(n6575), .Z(n6555) );
  XNOR U9893 ( .A(n9015), .B(n6578), .Z(n5327) );
  ANDN U9894 ( .B(n6579), .A(n8942), .Z(n9015) );
  IV U9895 ( .A(n9016), .Z(n8942) );
  XOR U9896 ( .A(n9017), .B(n9018), .Z(n5932) );
  XNOR U9897 ( .A(n3896), .B(n5191), .Z(n9018) );
  XOR U9898 ( .A(n9019), .B(n9020), .Z(n5191) );
  XNOR U9899 ( .A(n9022), .B(n9023), .Z(n3896) );
  ANDN U9900 ( .B(n9024), .A(n6599), .Z(n9022) );
  XOR U9901 ( .A(n4295), .B(n9025), .Z(n9017) );
  XNOR U9902 ( .A(n1793), .B(n9026), .Z(n9025) );
  XOR U9903 ( .A(n9027), .B(n9028), .Z(n1793) );
  XOR U9904 ( .A(n9030), .B(n9031), .Z(n4295) );
  AND U9905 ( .A(n9032), .B(n6586), .Z(n9030) );
  XOR U9906 ( .A(n9033), .B(n6060), .Z(out[1033]) );
  XOR U9907 ( .A(n8035), .B(n2465), .Z(n6060) );
  XOR U9908 ( .A(n9034), .B(n9035), .Z(n2465) );
  XNOR U9909 ( .A(n9036), .B(n9037), .Z(n8035) );
  NOR U9910 ( .A(n9038), .B(n9039), .Z(n9036) );
  ANDN U9911 ( .B(n1171), .A(n1172), .Z(n9033) );
  XNOR U9912 ( .A(n1941), .B(n9040), .Z(n1172) );
  XNOR U9913 ( .A(n7823), .B(n6198), .Z(n1941) );
  XOR U9914 ( .A(n9041), .B(n9042), .Z(n6198) );
  XOR U9915 ( .A(n4840), .B(n2014), .Z(n9042) );
  XNOR U9916 ( .A(n9043), .B(n9044), .Z(n2014) );
  ANDN U9917 ( .B(n8013), .A(n8011), .Z(n9043) );
  XOR U9918 ( .A(n9045), .B(n9046), .Z(n4840) );
  ANDN U9919 ( .B(n8019), .A(n8020), .Z(n9045) );
  XOR U9920 ( .A(n6107), .B(n9047), .Z(n9041) );
  XOR U9921 ( .A(n5321), .B(n3886), .Z(n9047) );
  XOR U9922 ( .A(n9048), .B(n9049), .Z(n3886) );
  NOR U9923 ( .A(n8007), .B(n8006), .Z(n9048) );
  IV U9924 ( .A(n9050), .Z(n8007) );
  XNOR U9925 ( .A(n9051), .B(n9052), .Z(n5321) );
  NOR U9926 ( .A(n8016), .B(n8015), .Z(n9051) );
  XOR U9927 ( .A(n9053), .B(n9054), .Z(n6107) );
  ANDN U9928 ( .B(n8003), .A(n8002), .Z(n9053) );
  XOR U9929 ( .A(n9055), .B(n9056), .Z(n7823) );
  XNOR U9930 ( .A(n5011), .B(n9057), .Z(n9056) );
  XNOR U9931 ( .A(n9058), .B(n7913), .Z(n5011) );
  XNOR U9932 ( .A(n2298), .B(n9060), .Z(n9055) );
  XOR U9933 ( .A(n3411), .B(n6637), .Z(n9060) );
  XOR U9934 ( .A(n9061), .B(n7900), .Z(n6637) );
  ANDN U9935 ( .B(n9062), .A(n8987), .Z(n9061) );
  XNOR U9936 ( .A(n9063), .B(n7905), .Z(n3411) );
  NOR U9937 ( .A(n9064), .B(n8982), .Z(n9063) );
  XNOR U9938 ( .A(n9065), .B(n7895), .Z(n2298) );
  ANDN U9939 ( .B(n9066), .A(n9067), .Z(n9065) );
  XOR U9940 ( .A(n3517), .B(n9068), .Z(n1171) );
  XNOR U9941 ( .A(n5937), .B(n6346), .Z(n3517) );
  XOR U9942 ( .A(n9069), .B(n9070), .Z(n6346) );
  XOR U9943 ( .A(n3303), .B(n5021), .Z(n9070) );
  XOR U9944 ( .A(n9071), .B(n6600), .Z(n5021) );
  ANDN U9945 ( .B(n6601), .A(n9023), .Z(n9071) );
  XNOR U9946 ( .A(n9072), .B(n6605), .Z(n3303) );
  XOR U9947 ( .A(n5334), .B(n9073), .Z(n9069) );
  XOR U9948 ( .A(n6581), .B(n2582), .Z(n9073) );
  XOR U9949 ( .A(n9074), .B(n6591), .Z(n2582) );
  ANDN U9950 ( .B(n6592), .A(n9075), .Z(n9074) );
  XOR U9951 ( .A(n9076), .B(n6597), .Z(n6581) );
  AND U9952 ( .A(n9020), .B(n6596), .Z(n9076) );
  XNOR U9953 ( .A(n9077), .B(n6588), .Z(n5334) );
  AND U9954 ( .A(n6587), .B(n9031), .Z(n9077) );
  XOR U9955 ( .A(n9078), .B(n9079), .Z(n5937) );
  XNOR U9956 ( .A(n3901), .B(n5196), .Z(n9079) );
  XNOR U9957 ( .A(n9080), .B(n7083), .Z(n5196) );
  ANDN U9958 ( .B(n6621), .A(n7084), .Z(n9080) );
  XNOR U9959 ( .A(n9081), .B(n9082), .Z(n3901) );
  NOR U9960 ( .A(n9083), .B(n6625), .Z(n9081) );
  XOR U9961 ( .A(n4297), .B(n9084), .Z(n9078) );
  XNOR U9962 ( .A(n7060), .B(n1799), .Z(n9084) );
  XNOR U9963 ( .A(n9085), .B(n7080), .Z(n1799) );
  NOR U9964 ( .A(n6629), .B(n7079), .Z(n9085) );
  IV U9965 ( .A(n9086), .Z(n6629) );
  XNOR U9966 ( .A(n9087), .B(n7093), .Z(n7060) );
  ANDN U9967 ( .B(n6616), .A(n7092), .Z(n9087) );
  XNOR U9968 ( .A(n9088), .B(n7088), .Z(n4297) );
  NOR U9969 ( .A(n7089), .B(n6612), .Z(n9088) );
  XOR U9970 ( .A(n9089), .B(n6065), .Z(out[1032]) );
  XOR U9971 ( .A(n8086), .B(n2472), .Z(n6065) );
  XNOR U9972 ( .A(n9090), .B(n9091), .Z(n2472) );
  XNOR U9973 ( .A(n9092), .B(n9093), .Z(n8086) );
  ANDN U9974 ( .B(n9094), .A(n9095), .Z(n9092) );
  NOR U9975 ( .A(n1176), .B(n1175), .Z(n9089) );
  XNOR U9976 ( .A(n3521), .B(n7085), .Z(n1175) );
  XOR U9977 ( .A(n9096), .B(n6627), .Z(n7085) );
  IV U9978 ( .A(n2554), .Z(n3521) );
  XNOR U9979 ( .A(n6351), .B(n5942), .Z(n2554) );
  XOR U9980 ( .A(n9097), .B(n9098), .Z(n5942) );
  XOR U9981 ( .A(n3905), .B(n5199), .Z(n9098) );
  XOR U9982 ( .A(n9099), .B(n7147), .Z(n5199) );
  NOR U9983 ( .A(n7064), .B(n6654), .Z(n9099) );
  XOR U9984 ( .A(n9100), .B(n9101), .Z(n6654) );
  XOR U9985 ( .A(n9102), .B(n9103), .Z(n7064) );
  XOR U9986 ( .A(n9104), .B(n9105), .Z(n3905) );
  ANDN U9987 ( .B(n9106), .A(n6658), .Z(n9104) );
  XOR U9988 ( .A(n9107), .B(n9108), .Z(n6658) );
  XOR U9989 ( .A(n4300), .B(n9109), .Z(n9097) );
  XNOR U9990 ( .A(n1803), .B(n7121), .Z(n9109) );
  XOR U9991 ( .A(n9110), .B(n9111), .Z(n7121) );
  ANDN U9992 ( .B(n7070), .A(n7071), .Z(n9110) );
  IV U9993 ( .A(n6649), .Z(n7071) );
  XOR U9994 ( .A(n9114), .B(n9115), .Z(n7070) );
  XNOR U9995 ( .A(n9116), .B(n7142), .Z(n1803) );
  ANDN U9996 ( .B(n7073), .A(n6662), .Z(n9116) );
  XOR U9997 ( .A(n9117), .B(n9118), .Z(n6662) );
  XOR U9998 ( .A(n9119), .B(n9120), .Z(n7073) );
  XOR U9999 ( .A(n9121), .B(n7150), .Z(n4300) );
  ANDN U10000 ( .B(n7066), .A(n6645), .Z(n9121) );
  IV U10001 ( .A(n7067), .Z(n6645) );
  XOR U10002 ( .A(n9122), .B(n9123), .Z(n7067) );
  XOR U10003 ( .A(n9124), .B(n9125), .Z(n7066) );
  XOR U10004 ( .A(n9126), .B(n9127), .Z(n6351) );
  XNOR U10005 ( .A(n3311), .B(n5121), .Z(n9127) );
  XNOR U10006 ( .A(n9128), .B(n9129), .Z(n5121) );
  ANDN U10007 ( .B(n6627), .A(n9082), .Z(n9128) );
  XOR U10008 ( .A(n9130), .B(n9131), .Z(n9082) );
  XOR U10009 ( .A(n9132), .B(n9133), .Z(n6627) );
  NOR U10010 ( .A(n6630), .B(n7080), .Z(n9134) );
  XNOR U10011 ( .A(n9135), .B(n9136), .Z(n7080) );
  XOR U10012 ( .A(n9137), .B(n9138), .Z(n6630) );
  XOR U10013 ( .A(n5339), .B(n9139), .Z(n9126) );
  XNOR U10014 ( .A(n6607), .B(n2589), .Z(n9139) );
  XNOR U10015 ( .A(n9140), .B(n6618), .Z(n2589) );
  ANDN U10016 ( .B(n7091), .A(n7093), .Z(n9140) );
  XOR U10017 ( .A(n9141), .B(n9142), .Z(n7093) );
  IV U10018 ( .A(n6617), .Z(n7091) );
  XOR U10019 ( .A(n9143), .B(n9144), .Z(n6617) );
  XNOR U10020 ( .A(n9145), .B(n6623), .Z(n6607) );
  NOR U10021 ( .A(n7082), .B(n7083), .Z(n9145) );
  XNOR U10022 ( .A(n9146), .B(n9147), .Z(n7083) );
  IV U10023 ( .A(n6622), .Z(n7082) );
  XNOR U10024 ( .A(n9148), .B(n9149), .Z(n6622) );
  XNOR U10025 ( .A(n9150), .B(n6614), .Z(n5339) );
  NOR U10026 ( .A(n6613), .B(n7088), .Z(n9150) );
  XOR U10027 ( .A(n9151), .B(n9152), .Z(n7088) );
  XOR U10028 ( .A(n9153), .B(n9154), .Z(n6613) );
  XOR U10029 ( .A(n9155), .B(n1946), .Z(n1176) );
  XOR U10030 ( .A(n9156), .B(n9157), .Z(n7890) );
  XNOR U10031 ( .A(n5014), .B(n9158), .Z(n9157) );
  XOR U10032 ( .A(n9159), .B(n8021), .Z(n5014) );
  AND U10033 ( .A(n9160), .B(n9046), .Z(n9159) );
  XOR U10034 ( .A(n2305), .B(n9161), .Z(n9156) );
  XOR U10035 ( .A(n3414), .B(n6910), .Z(n9161) );
  XNOR U10036 ( .A(n9162), .B(n8008), .Z(n6910) );
  NOR U10037 ( .A(n9163), .B(n9049), .Z(n9162) );
  XOR U10038 ( .A(n9164), .B(n8012), .Z(n3414) );
  ANDN U10039 ( .B(n9165), .A(n9044), .Z(n9164) );
  IV U10040 ( .A(n9166), .Z(n9044) );
  XNOR U10041 ( .A(n9167), .B(n8004), .Z(n2305) );
  ANDN U10042 ( .B(n9054), .A(n9168), .Z(n9167) );
  XOR U10043 ( .A(n9169), .B(n9170), .Z(n6204) );
  XNOR U10044 ( .A(n9171), .B(n3890), .Z(n9170) );
  ANDN U10045 ( .B(n8057), .A(n8058), .Z(n9172) );
  IV U10046 ( .A(n9174), .Z(n8058) );
  XOR U10047 ( .A(n4870), .B(n9175), .Z(n9169) );
  XOR U10048 ( .A(n2018), .B(n5326), .Z(n9175) );
  XOR U10049 ( .A(n9176), .B(n9177), .Z(n5326) );
  AND U10050 ( .A(n8066), .B(n8068), .Z(n9176) );
  XOR U10051 ( .A(n9178), .B(n9179), .Z(n2018) );
  ANDN U10052 ( .B(n8062), .A(n8063), .Z(n9178) );
  XOR U10053 ( .A(n9180), .B(n9181), .Z(n4870) );
  XOR U10054 ( .A(n9182), .B(n6075), .Z(out[1031]) );
  XOR U10055 ( .A(n8168), .B(n2479), .Z(n6075) );
  XNOR U10056 ( .A(n9183), .B(n9184), .Z(n2479) );
  XNOR U10057 ( .A(n9185), .B(n9186), .Z(n8168) );
  NOR U10058 ( .A(n9187), .B(n9188), .Z(n9185) );
  ANDN U10059 ( .B(n1179), .A(n1180), .Z(n9182) );
  XOR U10060 ( .A(n9189), .B(n1951), .Z(n1180) );
  XOR U10061 ( .A(n9190), .B(n9191), .Z(n7998) );
  XOR U10062 ( .A(n5017), .B(n9192), .Z(n9191) );
  XOR U10063 ( .A(n9193), .B(n8072), .Z(n5017) );
  ANDN U10064 ( .B(n9181), .A(n9194), .Z(n9193) );
  XNOR U10065 ( .A(n2316), .B(n9195), .Z(n9190) );
  XOR U10066 ( .A(n3417), .B(n7245), .Z(n9195) );
  XNOR U10067 ( .A(n9196), .B(n8059), .Z(n7245) );
  IV U10068 ( .A(n9197), .Z(n8059) );
  ANDN U10069 ( .B(n9173), .A(n9198), .Z(n9196) );
  XNOR U10070 ( .A(n9199), .B(n8064), .Z(n3417) );
  AND U10071 ( .A(n9200), .B(n9179), .Z(n9199) );
  XNOR U10072 ( .A(n9201), .B(n8055), .Z(n2316) );
  ANDN U10073 ( .B(n9202), .A(n9203), .Z(n9201) );
  XOR U10074 ( .A(n9204), .B(n9205), .Z(n6209) );
  XOR U10075 ( .A(n9206), .B(n3894), .Z(n9205) );
  XOR U10076 ( .A(n9207), .B(n9208), .Z(n3894) );
  ANDN U10077 ( .B(n9209), .A(n7989), .Z(n9207) );
  XOR U10078 ( .A(n4910), .B(n9210), .Z(n9204) );
  XOR U10079 ( .A(n2021), .B(n5330), .Z(n9210) );
  XNOR U10080 ( .A(n9211), .B(n9212), .Z(n5330) );
  XNOR U10081 ( .A(n9214), .B(n9215), .Z(n2021) );
  ANDN U10082 ( .B(n8119), .A(n9216), .Z(n9214) );
  XOR U10083 ( .A(n9217), .B(n9218), .Z(n4910) );
  XNOR U10084 ( .A(n7144), .B(n2560), .Z(n1179) );
  XOR U10085 ( .A(n5947), .B(n6355), .Z(n2560) );
  XOR U10086 ( .A(n9220), .B(n9221), .Z(n6355) );
  XOR U10087 ( .A(n3315), .B(n5508), .Z(n9221) );
  XOR U10088 ( .A(n9222), .B(n6659), .Z(n5508) );
  XOR U10089 ( .A(n9223), .B(n9224), .Z(n6659) );
  NOR U10090 ( .A(n9225), .B(n9105), .Z(n9222) );
  XNOR U10091 ( .A(n9226), .B(n6663), .Z(n3315) );
  XOR U10092 ( .A(n9227), .B(n9228), .Z(n6663) );
  ANDN U10093 ( .B(n7142), .A(n7141), .Z(n9226) );
  IV U10094 ( .A(n6664), .Z(n7141) );
  XOR U10095 ( .A(n9229), .B(n9230), .Z(n6664) );
  XOR U10096 ( .A(n9231), .B(n9232), .Z(n7142) );
  XOR U10097 ( .A(n5343), .B(n9233), .Z(n9220) );
  XNOR U10098 ( .A(n6640), .B(n2594), .Z(n9233) );
  XOR U10099 ( .A(n9234), .B(n6651), .Z(n2594) );
  XOR U10100 ( .A(n9151), .B(n9235), .Z(n6651) );
  NOR U10101 ( .A(n9111), .B(n6650), .Z(n9234) );
  XOR U10102 ( .A(n9236), .B(n9237), .Z(n6650) );
  IV U10103 ( .A(n7139), .Z(n9111) );
  XOR U10104 ( .A(n9238), .B(n9239), .Z(n7139) );
  XOR U10105 ( .A(n9240), .B(n6655), .Z(n6640) );
  XOR U10106 ( .A(n9241), .B(n9242), .Z(n6655) );
  ANDN U10107 ( .B(n7147), .A(n7146), .Z(n9240) );
  IV U10108 ( .A(n6656), .Z(n7146) );
  XOR U10109 ( .A(n9243), .B(n9244), .Z(n6656) );
  XOR U10110 ( .A(n9245), .B(n9246), .Z(n7147) );
  XNOR U10111 ( .A(n9247), .B(n6647), .Z(n5343) );
  XOR U10112 ( .A(n9248), .B(n9249), .Z(n6647) );
  NOR U10113 ( .A(n7149), .B(n7150), .Z(n9247) );
  XNOR U10114 ( .A(n9250), .B(n9251), .Z(n7150) );
  XOR U10115 ( .A(n9252), .B(n9253), .Z(n7149) );
  XOR U10116 ( .A(n9254), .B(n9255), .Z(n5947) );
  XOR U10117 ( .A(n3910), .B(n5202), .Z(n9255) );
  XNOR U10118 ( .A(n9256), .B(n9257), .Z(n5202) );
  ANDN U10119 ( .B(n6680), .A(n7130), .Z(n9256) );
  IV U10120 ( .A(n9258), .Z(n7130) );
  XNOR U10121 ( .A(n9259), .B(n9260), .Z(n6680) );
  XNOR U10122 ( .A(n9261), .B(n9262), .Z(n3910) );
  ANDN U10123 ( .B(n7127), .A(n6684), .Z(n9261) );
  XOR U10124 ( .A(n9263), .B(n9264), .Z(n6684) );
  XOR U10125 ( .A(n9265), .B(n9266), .Z(n9254) );
  XNOR U10126 ( .A(n7178), .B(n1808), .Z(n9266) );
  XNOR U10127 ( .A(n9267), .B(n9268), .Z(n1808) );
  AND U10128 ( .A(n6688), .B(n7125), .Z(n9267) );
  XOR U10129 ( .A(n9269), .B(n9270), .Z(n6688) );
  XOR U10130 ( .A(n9271), .B(n9272), .Z(n7178) );
  ANDN U10131 ( .B(n7135), .A(n6675), .Z(n9271) );
  XNOR U10132 ( .A(n9273), .B(n9274), .Z(n6675) );
  XNOR U10133 ( .A(n9275), .B(n6660), .Z(n7144) );
  IV U10134 ( .A(n9225), .Z(n6660) );
  XNOR U10135 ( .A(n9276), .B(n9277), .Z(n9225) );
  ANDN U10136 ( .B(n9105), .A(n9106), .Z(n9275) );
  IV U10137 ( .A(n7075), .Z(n9106) );
  XOR U10138 ( .A(n9269), .B(n9278), .Z(n7075) );
  XNOR U10139 ( .A(n9279), .B(n9280), .Z(n9105) );
  XNOR U10140 ( .A(n9281), .B(n6080), .Z(out[1030]) );
  IV U10141 ( .A(n6397), .Z(n6080) );
  XNOR U10142 ( .A(n8194), .B(n2486), .Z(n6397) );
  XNOR U10143 ( .A(n9282), .B(n9283), .Z(n2486) );
  XNOR U10144 ( .A(n9284), .B(n9285), .Z(n8194) );
  ANDN U10145 ( .B(n1183), .A(n1184), .Z(n9281) );
  XNOR U10146 ( .A(n9288), .B(n1955), .Z(n1184) );
  XOR U10147 ( .A(n9289), .B(n9290), .Z(n8049) );
  XNOR U10148 ( .A(n3421), .B(n5025), .Z(n9290) );
  XOR U10149 ( .A(n9291), .B(n7984), .Z(n5025) );
  AND U10150 ( .A(n7985), .B(n9218), .Z(n9291) );
  XNOR U10151 ( .A(n9292), .B(n8121), .Z(n3421) );
  ANDN U10152 ( .B(n8120), .A(n9215), .Z(n9292) );
  XOR U10153 ( .A(n7974), .B(n9293), .Z(n9289) );
  XOR U10154 ( .A(n7059), .B(n2326), .Z(n9293) );
  XOR U10155 ( .A(n9294), .B(n7994), .Z(n2326) );
  AND U10156 ( .A(n9295), .B(n7995), .Z(n9294) );
  XOR U10157 ( .A(n9296), .B(n7980), .Z(n7059) );
  ANDN U10158 ( .B(n7981), .A(n9212), .Z(n9296) );
  XNOR U10159 ( .A(n9297), .B(n7991), .Z(n7974) );
  ANDN U10160 ( .B(n7990), .A(n9208), .Z(n9297) );
  XOR U10161 ( .A(n9298), .B(n9299), .Z(n6214) );
  XOR U10162 ( .A(n9300), .B(n3897), .Z(n9299) );
  XNOR U10163 ( .A(n9301), .B(n9302), .Z(n3897) );
  ANDN U10164 ( .B(n9303), .A(n8635), .Z(n9301) );
  IV U10165 ( .A(n9304), .Z(n8635) );
  XOR U10166 ( .A(n4948), .B(n9305), .Z(n9298) );
  XOR U10167 ( .A(n2024), .B(n5337), .Z(n9305) );
  XNOR U10168 ( .A(n9306), .B(n9307), .Z(n5337) );
  XNOR U10169 ( .A(n9309), .B(n9310), .Z(n2024) );
  NOR U10170 ( .A(n9311), .B(n9312), .Z(n9309) );
  ANDN U10171 ( .B(n9315), .A(n9316), .Z(n9313) );
  IV U10172 ( .A(n8630), .Z(n9316) );
  XNOR U10173 ( .A(n9317), .B(n2567), .Z(n1183) );
  XNOR U10174 ( .A(n5953), .B(n6361), .Z(n2567) );
  XNOR U10175 ( .A(n9318), .B(n9319), .Z(n6361) );
  XNOR U10176 ( .A(n2603), .B(n5347), .Z(n9319) );
  XNOR U10177 ( .A(n9320), .B(n7133), .Z(n5347) );
  XNOR U10178 ( .A(n9321), .B(n9322), .Z(n7133) );
  AND U10179 ( .A(n6673), .B(n9323), .Z(n9320) );
  XNOR U10180 ( .A(n9324), .B(n6676), .Z(n2603) );
  XOR U10181 ( .A(n9325), .B(n9251), .Z(n6676) );
  ANDN U10182 ( .B(n6677), .A(n9272), .Z(n9324) );
  XOR U10183 ( .A(n3318), .B(n9326), .Z(n9318) );
  XOR U10184 ( .A(n5866), .B(n6666), .Z(n9326) );
  XNOR U10185 ( .A(n9327), .B(n6681), .Z(n6666) );
  XNOR U10186 ( .A(n9328), .B(n9329), .Z(n6681) );
  ANDN U10187 ( .B(n9257), .A(n9330), .Z(n9327) );
  XNOR U10188 ( .A(n9331), .B(n6685), .Z(n5866) );
  XNOR U10189 ( .A(n9102), .B(n9332), .Z(n6685) );
  ANDN U10190 ( .B(n9262), .A(n9333), .Z(n9331) );
  XNOR U10191 ( .A(n9334), .B(n6689), .Z(n3318) );
  XOR U10192 ( .A(n9335), .B(n9336), .Z(n6689) );
  ANDN U10193 ( .B(n9268), .A(n9337), .Z(n9334) );
  XOR U10194 ( .A(n9338), .B(n9339), .Z(n5953) );
  XNOR U10195 ( .A(n3914), .B(n5204), .Z(n9339) );
  XOR U10196 ( .A(n9340), .B(n7231), .Z(n5204) );
  NOR U10197 ( .A(n6706), .B(n7232), .Z(n9340) );
  XOR U10198 ( .A(n9341), .B(n9342), .Z(n3914) );
  ANDN U10199 ( .B(n6710), .A(n9343), .Z(n9341) );
  XOR U10200 ( .A(n4108), .B(n9344), .Z(n9338) );
  XOR U10201 ( .A(n7206), .B(n1812), .Z(n9344) );
  XOR U10202 ( .A(n9345), .B(n7226), .Z(n1812) );
  ANDN U10203 ( .B(n7227), .A(n6714), .Z(n9345) );
  XOR U10204 ( .A(n9346), .B(n7223), .Z(n7206) );
  NOR U10205 ( .A(n9347), .B(n6701), .Z(n9346) );
  XNOR U10206 ( .A(n9348), .B(n7235), .Z(n4108) );
  ANDN U10207 ( .B(n7236), .A(n6697), .Z(n9348) );
  XNOR U10208 ( .A(n9349), .B(n4196), .Z(out[102]) );
  IV U10209 ( .A(n4373), .Z(n4196) );
  XOR U10210 ( .A(n6978), .B(n2565), .Z(n4373) );
  XOR U10211 ( .A(n7915), .B(n9350), .Z(n2565) );
  XOR U10212 ( .A(n9351), .B(n9352), .Z(n7915) );
  XNOR U10213 ( .A(n4378), .B(n2187), .Z(n9352) );
  XOR U10214 ( .A(n9353), .B(n9354), .Z(n2187) );
  ANDN U10215 ( .B(n9355), .A(n9356), .Z(n9353) );
  XNOR U10216 ( .A(n9357), .B(n9358), .Z(n4378) );
  AND U10217 ( .A(n6984), .B(n6986), .Z(n9357) );
  XOR U10218 ( .A(n6016), .B(n9359), .Z(n9351) );
  XOR U10219 ( .A(n5550), .B(n3799), .Z(n9359) );
  XOR U10220 ( .A(n9360), .B(n9361), .Z(n3799) );
  NOR U10221 ( .A(n6975), .B(n6974), .Z(n9360) );
  IV U10222 ( .A(n9362), .Z(n6975) );
  XOR U10223 ( .A(n9363), .B(n9364), .Z(n5550) );
  NOR U10224 ( .A(n9365), .B(n6980), .Z(n9363) );
  XOR U10225 ( .A(n9366), .B(n9367), .Z(n6016) );
  ANDN U10226 ( .B(n6971), .A(n6970), .Z(n9366) );
  IV U10227 ( .A(n9368), .Z(n6970) );
  XOR U10228 ( .A(n9369), .B(n9355), .Z(n6978) );
  ANDN U10229 ( .B(n9356), .A(n9370), .Z(n9369) );
  ANDN U10230 ( .B(n3585), .A(n3587), .Z(n9349) );
  XNOR U10231 ( .A(n6213), .B(n9372), .Z(n2339) );
  XOR U10232 ( .A(n9373), .B(n9374), .Z(n6213) );
  XNOR U10233 ( .A(n3195), .B(n6911), .Z(n9374) );
  XOR U10234 ( .A(n9375), .B(n9376), .Z(n6911) );
  NOR U10235 ( .A(n9377), .B(n9378), .Z(n9375) );
  XNOR U10236 ( .A(n9379), .B(n9380), .Z(n3195) );
  ANDN U10237 ( .B(n9381), .A(n9382), .Z(n9379) );
  XOR U10238 ( .A(n5506), .B(n9383), .Z(n9373) );
  XOR U10239 ( .A(n8232), .B(n2372), .Z(n9383) );
  XNOR U10240 ( .A(n9384), .B(n9385), .Z(n2372) );
  ANDN U10241 ( .B(n9386), .A(n9387), .Z(n9384) );
  XOR U10242 ( .A(n9388), .B(n9389), .Z(n8232) );
  NOR U10243 ( .A(n9390), .B(n9391), .Z(n9388) );
  XNOR U10244 ( .A(n9392), .B(n9393), .Z(n5506) );
  NOR U10245 ( .A(n9394), .B(n9395), .Z(n9392) );
  XOR U10246 ( .A(n7406), .B(n3210), .Z(n3585) );
  XOR U10247 ( .A(n9396), .B(n9397), .Z(n3210) );
  XOR U10248 ( .A(n9398), .B(n9399), .Z(n7406) );
  ANDN U10249 ( .B(n9400), .A(n9401), .Z(n9398) );
  XNOR U10250 ( .A(n9402), .B(n6085), .Z(out[1029]) );
  XOR U10251 ( .A(n8248), .B(n2495), .Z(n6085) );
  IV U10252 ( .A(n3254), .Z(n2495) );
  XOR U10253 ( .A(n9403), .B(n9404), .Z(n3254) );
  NOR U10254 ( .A(n9407), .B(n9408), .Z(n9405) );
  ANDN U10255 ( .B(n1189), .A(n1187), .Z(n9402) );
  IV U10256 ( .A(n6401), .Z(n1187) );
  XNOR U10257 ( .A(n7229), .B(n2574), .Z(n6401) );
  XNOR U10258 ( .A(n5962), .B(n6366), .Z(n2574) );
  XNOR U10259 ( .A(n9409), .B(n9410), .Z(n6366) );
  XOR U10260 ( .A(n2614), .B(n5352), .Z(n9410) );
  XOR U10261 ( .A(n9411), .B(n6698), .Z(n5352) );
  ANDN U10262 ( .B(n7235), .A(n7234), .Z(n9411) );
  XOR U10263 ( .A(n9412), .B(n9413), .Z(n7234) );
  XNOR U10264 ( .A(n9414), .B(n9415), .Z(n7235) );
  XNOR U10265 ( .A(n9416), .B(n6703), .Z(n2614) );
  ANDN U10266 ( .B(n6702), .A(n7223), .Z(n9416) );
  XOR U10267 ( .A(n9417), .B(n9418), .Z(n7223) );
  XNOR U10268 ( .A(n9419), .B(n9420), .Z(n6702) );
  XOR U10269 ( .A(n3321), .B(n9421), .Z(n9409) );
  XNOR U10270 ( .A(n6368), .B(n6692), .Z(n9421) );
  XNOR U10271 ( .A(n9422), .B(n6707), .Z(n6692) );
  ANDN U10272 ( .B(n6708), .A(n7231), .Z(n9422) );
  XOR U10273 ( .A(n9423), .B(n9424), .Z(n7231) );
  XNOR U10274 ( .A(n9425), .B(n9426), .Z(n6708) );
  XNOR U10275 ( .A(n9427), .B(n9428), .Z(n6368) );
  ANDN U10276 ( .B(n6712), .A(n9342), .Z(n9427) );
  XNOR U10277 ( .A(n9429), .B(n6716), .Z(n3321) );
  ANDN U10278 ( .B(n6715), .A(n7226), .Z(n9429) );
  XNOR U10279 ( .A(n9430), .B(n9431), .Z(n7226) );
  XOR U10280 ( .A(n9432), .B(n9433), .Z(n6715) );
  XOR U10281 ( .A(n9434), .B(n9435), .Z(n5962) );
  XNOR U10282 ( .A(n3603), .B(n5207), .Z(n9435) );
  XNOR U10283 ( .A(n9436), .B(n7300), .Z(n5207) );
  AND U10284 ( .A(n7215), .B(n6738), .Z(n9436) );
  XOR U10285 ( .A(n9437), .B(n9438), .Z(n6738) );
  XOR U10286 ( .A(n9439), .B(n9440), .Z(n7215) );
  XOR U10287 ( .A(n9441), .B(n9442), .Z(n3603) );
  ANDN U10288 ( .B(n6724), .A(n7217), .Z(n9441) );
  XOR U10289 ( .A(n9443), .B(n9444), .Z(n6724) );
  XOR U10290 ( .A(n4111), .B(n9445), .Z(n9434) );
  XNOR U10291 ( .A(n7273), .B(n1816), .Z(n9445) );
  XNOR U10292 ( .A(n9446), .B(n7295), .Z(n1816) );
  ANDN U10293 ( .B(n6728), .A(n7296), .Z(n9446) );
  XOR U10294 ( .A(n9447), .B(n9448), .Z(n7296) );
  XOR U10295 ( .A(n9449), .B(n9450), .Z(n6728) );
  ANDN U10296 ( .B(n6732), .A(n7219), .Z(n9451) );
  IV U10297 ( .A(n7293), .Z(n7219) );
  XOR U10298 ( .A(n9452), .B(n9453), .Z(n7293) );
  XNOR U10299 ( .A(n9454), .B(n9252), .Z(n6732) );
  XNOR U10300 ( .A(n9455), .B(n7302), .Z(n4111) );
  IV U10301 ( .A(n9456), .Z(n7302) );
  ANDN U10302 ( .B(n7212), .A(n6742), .Z(n9455) );
  XOR U10303 ( .A(n9457), .B(n9458), .Z(n6742) );
  XOR U10304 ( .A(n9459), .B(n9460), .Z(n7212) );
  XNOR U10305 ( .A(n9461), .B(n6712), .Z(n7229) );
  XNOR U10306 ( .A(n9462), .B(n9463), .Z(n6712) );
  ANDN U10307 ( .B(n9342), .A(n9464), .Z(n9461) );
  XNOR U10308 ( .A(n9465), .B(n9466), .Z(n9342) );
  XNOR U10309 ( .A(n9467), .B(n4215), .Z(n1189) );
  IV U10310 ( .A(n1961), .Z(n4215) );
  XOR U10311 ( .A(n9468), .B(n9469), .Z(n8116) );
  XNOR U10312 ( .A(n3424), .B(n5028), .Z(n9469) );
  XNOR U10313 ( .A(n9470), .B(n8631), .Z(n5028) );
  ANDN U10314 ( .B(n8632), .A(n9314), .Z(n9470) );
  XNOR U10315 ( .A(n9471), .B(n8641), .Z(n3424) );
  ANDN U10316 ( .B(n9310), .A(n9472), .Z(n9471) );
  XOR U10317 ( .A(n8621), .B(n9473), .Z(n9468) );
  XNOR U10318 ( .A(n7120), .B(n2333), .Z(n9473) );
  XNOR U10319 ( .A(n9474), .B(n8645), .Z(n2333) );
  ANDN U10320 ( .B(n9475), .A(n8644), .Z(n9474) );
  XOR U10321 ( .A(n9476), .B(n8627), .Z(n7120) );
  ANDN U10322 ( .B(n8628), .A(n9307), .Z(n9476) );
  XNOR U10323 ( .A(n9477), .B(n8637), .Z(n8621) );
  ANDN U10324 ( .B(n9302), .A(n9478), .Z(n9477) );
  XOR U10325 ( .A(n9479), .B(n9480), .Z(n6219) );
  XOR U10326 ( .A(n9481), .B(n3902), .Z(n9480) );
  XOR U10327 ( .A(n9482), .B(n9483), .Z(n3902) );
  NOR U10328 ( .A(n9484), .B(n9385), .Z(n9482) );
  XNOR U10329 ( .A(n4985), .B(n9485), .Z(n9479) );
  XOR U10330 ( .A(n2027), .B(n5341), .Z(n9485) );
  XNOR U10331 ( .A(n9486), .B(n9487), .Z(n5341) );
  ANDN U10332 ( .B(n9488), .A(n9376), .Z(n9486) );
  XNOR U10333 ( .A(n9489), .B(n9490), .Z(n2027) );
  ANDN U10334 ( .B(n9491), .A(n9492), .Z(n9489) );
  XNOR U10335 ( .A(n9493), .B(n9494), .Z(n4985) );
  NOR U10336 ( .A(n9495), .B(n9380), .Z(n9493) );
  XOR U10337 ( .A(n9496), .B(n6090), .Z(out[1028]) );
  XOR U10338 ( .A(n8302), .B(n2500), .Z(n6090) );
  XNOR U10339 ( .A(n9497), .B(n9498), .Z(n2500) );
  XNOR U10340 ( .A(n9499), .B(n9500), .Z(n8302) );
  ANDN U10341 ( .B(n9501), .A(n9502), .Z(n9499) );
  ANDN U10342 ( .B(n1193), .A(n6404), .Z(n9496) );
  XNOR U10343 ( .A(n7298), .B(n2581), .Z(n6404) );
  XNOR U10344 ( .A(n5967), .B(n6378), .Z(n2581) );
  XNOR U10345 ( .A(n9503), .B(n9504), .Z(n6378) );
  XNOR U10346 ( .A(n2620), .B(n5356), .Z(n9504) );
  XNOR U10347 ( .A(n9505), .B(n6744), .Z(n5356) );
  XOR U10348 ( .A(n9506), .B(n9507), .Z(n6744) );
  NOR U10349 ( .A(n9456), .B(n6743), .Z(n9505) );
  XNOR U10350 ( .A(n9508), .B(n9509), .Z(n6743) );
  XNOR U10351 ( .A(n9510), .B(n9511), .Z(n9456) );
  XNOR U10352 ( .A(n9512), .B(n6735), .Z(n2620) );
  XOR U10353 ( .A(n9414), .B(n9513), .Z(n6735) );
  ANDN U10354 ( .B(n6736), .A(n7292), .Z(n9512) );
  XNOR U10355 ( .A(n9138), .B(n9514), .Z(n7292) );
  XNOR U10356 ( .A(n9515), .B(n9516), .Z(n6736) );
  XOR U10357 ( .A(n6719), .B(n9517), .Z(n9503) );
  XNOR U10358 ( .A(n5183), .B(n3325), .Z(n9517) );
  XNOR U10359 ( .A(n9518), .B(n6730), .Z(n3325) );
  XOR U10360 ( .A(n9519), .B(n9520), .Z(n6730) );
  ANDN U10361 ( .B(n7295), .A(n6729), .Z(n9518) );
  XOR U10362 ( .A(n9521), .B(n9522), .Z(n6729) );
  XOR U10363 ( .A(n9523), .B(n9524), .Z(n7295) );
  XNOR U10364 ( .A(n9525), .B(n6726), .Z(n5183) );
  ANDN U10365 ( .B(n9442), .A(n6725), .Z(n9525) );
  IV U10366 ( .A(n9528), .Z(n6725) );
  XNOR U10367 ( .A(n9529), .B(n6740), .Z(n6719) );
  XNOR U10368 ( .A(n9530), .B(n9531), .Z(n6740) );
  ANDN U10369 ( .B(n7300), .A(n6739), .Z(n9529) );
  XOR U10370 ( .A(n9532), .B(n9533), .Z(n6739) );
  XOR U10371 ( .A(n9534), .B(n9535), .Z(n7300) );
  XOR U10372 ( .A(n9536), .B(n9537), .Z(n5967) );
  XOR U10373 ( .A(n1829), .B(n5210), .Z(n9537) );
  XOR U10374 ( .A(n9538), .B(n7373), .Z(n5210) );
  ANDN U10375 ( .B(n6760), .A(n7282), .Z(n9538) );
  XNOR U10376 ( .A(n9539), .B(n9540), .Z(n7282) );
  XNOR U10377 ( .A(n9541), .B(n9542), .Z(n6760) );
  XNOR U10378 ( .A(n9543), .B(n7368), .Z(n1829) );
  ANDN U10379 ( .B(n6768), .A(n7369), .Z(n9543) );
  XOR U10380 ( .A(n9544), .B(n9545), .Z(n7369) );
  XOR U10381 ( .A(n9546), .B(n9547), .Z(n6768) );
  XNOR U10382 ( .A(n4114), .B(n9548), .Z(n9536) );
  XOR U10383 ( .A(n7348), .B(n3608), .Z(n9548) );
  XNOR U10384 ( .A(n9549), .B(n9550), .Z(n3608) );
  ANDN U10385 ( .B(n7285), .A(n6764), .Z(n9549) );
  XOR U10386 ( .A(n9551), .B(n9552), .Z(n6764) );
  XOR U10387 ( .A(n9553), .B(n7366), .Z(n7348) );
  NOR U10388 ( .A(n7288), .B(n7287), .Z(n9553) );
  XOR U10389 ( .A(n9554), .B(n9555), .Z(n7287) );
  IV U10390 ( .A(n6755), .Z(n7288) );
  XOR U10391 ( .A(n9556), .B(n9557), .Z(n6755) );
  XOR U10392 ( .A(n9558), .B(n7375), .Z(n4114) );
  ANDN U10393 ( .B(n7279), .A(n6751), .Z(n9558) );
  XNOR U10394 ( .A(n9559), .B(n9560), .Z(n6751) );
  XOR U10395 ( .A(n9443), .B(n9561), .Z(n7279) );
  XOR U10396 ( .A(n9562), .B(n9528), .Z(n7298) );
  XOR U10397 ( .A(n9563), .B(n9564), .Z(n9528) );
  ANDN U10398 ( .B(n7217), .A(n9442), .Z(n9562) );
  XOR U10399 ( .A(n9565), .B(n9566), .Z(n9442) );
  XOR U10400 ( .A(n9567), .B(n9547), .Z(n7217) );
  XNOR U10401 ( .A(n9568), .B(n4219), .Z(n1193) );
  IV U10402 ( .A(n1969), .Z(n4219) );
  XOR U10403 ( .A(n9569), .B(n9570), .Z(n8179) );
  XOR U10404 ( .A(n3430), .B(n5031), .Z(n9570) );
  XOR U10405 ( .A(n9571), .B(n9381), .Z(n5031) );
  AND U10406 ( .A(n9494), .B(n9382), .Z(n9571) );
  XNOR U10407 ( .A(n9572), .B(n9391), .Z(n3430) );
  ANDN U10408 ( .B(n9490), .A(n9573), .Z(n9572) );
  XNOR U10409 ( .A(n9371), .B(n9574), .Z(n9569) );
  XOR U10410 ( .A(n7177), .B(n2340), .Z(n9574) );
  XNOR U10411 ( .A(n9575), .B(n9395), .Z(n2340) );
  ANDN U10412 ( .B(n9576), .A(n9577), .Z(n9575) );
  XNOR U10413 ( .A(n9578), .B(n9377), .Z(n7177) );
  IV U10414 ( .A(n9579), .Z(n9377) );
  ANDN U10415 ( .B(n9378), .A(n9487), .Z(n9578) );
  XOR U10416 ( .A(n9580), .B(n9386), .Z(n9371) );
  NOR U10417 ( .A(n9581), .B(n9483), .Z(n9580) );
  XOR U10418 ( .A(n9582), .B(n9583), .Z(n6224) );
  XNOR U10419 ( .A(n2030), .B(n3906), .Z(n9583) );
  XNOR U10420 ( .A(n9584), .B(n9585), .Z(n3906) );
  ANDN U10421 ( .B(n9586), .A(n9587), .Z(n9584) );
  XNOR U10422 ( .A(n9588), .B(n9589), .Z(n2030) );
  ANDN U10423 ( .B(n9590), .A(n9591), .Z(n9588) );
  XNOR U10424 ( .A(n9592), .B(n9593), .Z(n9582) );
  XOR U10425 ( .A(n5345), .B(n5020), .Z(n9593) );
  XNOR U10426 ( .A(n9594), .B(n9595), .Z(n5020) );
  ANDN U10427 ( .B(n9596), .A(n9597), .Z(n9594) );
  XNOR U10428 ( .A(n9598), .B(n9599), .Z(n5345) );
  ANDN U10429 ( .B(n9600), .A(n9601), .Z(n9598) );
  XOR U10430 ( .A(n9602), .B(n6095), .Z(out[1027]) );
  XOR U10431 ( .A(n8356), .B(n3261), .Z(n6095) );
  XOR U10432 ( .A(n9603), .B(n9604), .Z(n3261) );
  XNOR U10433 ( .A(n9605), .B(n9606), .Z(n8356) );
  ANDN U10434 ( .B(n9607), .A(n9608), .Z(n9605) );
  ANDN U10435 ( .B(n1197), .A(n1195), .Z(n9602) );
  IV U10436 ( .A(n6407), .Z(n1195) );
  XNOR U10437 ( .A(n7371), .B(n2588), .Z(n6407) );
  XNOR U10438 ( .A(n5972), .B(n6382), .Z(n2588) );
  XNOR U10439 ( .A(n9609), .B(n9610), .Z(n6382) );
  XNOR U10440 ( .A(n2628), .B(n5361), .Z(n9610) );
  XOR U10441 ( .A(n9611), .B(n6753), .Z(n5361) );
  XNOR U10442 ( .A(n9612), .B(n9613), .Z(n6753) );
  ANDN U10443 ( .B(n6752), .A(n7375), .Z(n9611) );
  XOR U10444 ( .A(n9614), .B(n9615), .Z(n7375) );
  XNOR U10445 ( .A(n9616), .B(n9617), .Z(n6752) );
  XNOR U10446 ( .A(n9618), .B(n6756), .Z(n2628) );
  XNOR U10447 ( .A(n9619), .B(n9511), .Z(n6756) );
  ANDN U10448 ( .B(n7366), .A(n6757), .Z(n9618) );
  XNOR U10449 ( .A(n9620), .B(n9621), .Z(n6757) );
  XOR U10450 ( .A(n9229), .B(n9622), .Z(n7366) );
  IV U10451 ( .A(n9623), .Z(n9229) );
  XNOR U10452 ( .A(n3329), .B(n9624), .Z(n9609) );
  XNOR U10453 ( .A(n5217), .B(n6746), .Z(n9624) );
  XOR U10454 ( .A(n9625), .B(n7283), .Z(n6746) );
  IV U10455 ( .A(n6761), .Z(n7283) );
  XOR U10456 ( .A(n9131), .B(n9626), .Z(n6761) );
  ANDN U10457 ( .B(n6762), .A(n7373), .Z(n9625) );
  XOR U10458 ( .A(n9627), .B(n9628), .Z(n7373) );
  XOR U10459 ( .A(n9629), .B(n9630), .Z(n6762) );
  XNOR U10460 ( .A(n9631), .B(n6765), .Z(n5217) );
  XOR U10461 ( .A(n9632), .B(n9633), .Z(n6765) );
  AND U10462 ( .A(n9550), .B(n6766), .Z(n9631) );
  XNOR U10463 ( .A(n9634), .B(n6769), .Z(n3329) );
  XOR U10464 ( .A(n9635), .B(n9636), .Z(n6769) );
  ANDN U10465 ( .B(n7368), .A(n6770), .Z(n9634) );
  XOR U10466 ( .A(n9637), .B(n9638), .Z(n6770) );
  XOR U10467 ( .A(n9639), .B(n9640), .Z(n7368) );
  XOR U10468 ( .A(n9641), .B(n9642), .Z(n5972) );
  XOR U10469 ( .A(n1833), .B(n5212), .Z(n9642) );
  XOR U10470 ( .A(n9643), .B(n7449), .Z(n5212) );
  ANDN U10471 ( .B(n6786), .A(n7357), .Z(n9643) );
  IV U10472 ( .A(n7450), .Z(n7357) );
  XOR U10473 ( .A(n9644), .B(n9645), .Z(n7450) );
  XNOR U10474 ( .A(n9646), .B(n9647), .Z(n6786) );
  XNOR U10475 ( .A(n9648), .B(n7444), .Z(n1833) );
  ANDN U10476 ( .B(n6794), .A(n7445), .Z(n9648) );
  XOR U10477 ( .A(n9649), .B(n9650), .Z(n7445) );
  XOR U10478 ( .A(n4118), .B(n9653), .Z(n9641) );
  XNOR U10479 ( .A(n7421), .B(n3612), .Z(n9653) );
  XNOR U10480 ( .A(n9654), .B(n9655), .Z(n3612) );
  ANDN U10481 ( .B(n7352), .A(n6790), .Z(n9654) );
  XNOR U10482 ( .A(n9656), .B(n9657), .Z(n6790) );
  XOR U10483 ( .A(n9658), .B(n7442), .Z(n7421) );
  ANDN U10484 ( .B(n6781), .A(n7362), .Z(n9658) );
  XOR U10485 ( .A(n9659), .B(n9660), .Z(n7362) );
  XNOR U10486 ( .A(n9661), .B(n9413), .Z(n6781) );
  XNOR U10487 ( .A(n9662), .B(n7453), .Z(n4118) );
  ANDN U10488 ( .B(n7354), .A(n6777), .Z(n9662) );
  XOR U10489 ( .A(n9663), .B(n9664), .Z(n6777) );
  XOR U10490 ( .A(n9665), .B(n9552), .Z(n7354) );
  XNOR U10491 ( .A(n9666), .B(n6766), .Z(n7371) );
  XOR U10492 ( .A(n9667), .B(n9668), .Z(n6766) );
  NOR U10493 ( .A(n9550), .B(n7285), .Z(n9666) );
  XOR U10494 ( .A(n9669), .B(n9652), .Z(n7285) );
  XOR U10495 ( .A(n9670), .B(n9671), .Z(n9550) );
  XOR U10496 ( .A(n9672), .B(n4222), .Z(n1197) );
  IV U10497 ( .A(n1973), .Z(n4222) );
  XOR U10498 ( .A(n9673), .B(n9674), .Z(n8233) );
  XNOR U10499 ( .A(n3432), .B(n5034), .Z(n9674) );
  XNOR U10500 ( .A(n9675), .B(n9676), .Z(n5034) );
  AND U10501 ( .A(n9595), .B(n9677), .Z(n9675) );
  XNOR U10502 ( .A(n9678), .B(n9679), .Z(n3432) );
  ANDN U10503 ( .B(n9589), .A(n9680), .Z(n9678) );
  XNOR U10504 ( .A(n9681), .B(n9682), .Z(n9673) );
  XOR U10505 ( .A(n7205), .B(n2347), .Z(n9682) );
  XOR U10506 ( .A(n9683), .B(n9684), .Z(n2347) );
  ANDN U10507 ( .B(n9685), .A(n9686), .Z(n9683) );
  XOR U10508 ( .A(n9687), .B(n9688), .Z(n7205) );
  ANDN U10509 ( .B(n9689), .A(n9599), .Z(n9687) );
  XOR U10510 ( .A(n9690), .B(n9691), .Z(n6234) );
  XNOR U10511 ( .A(n2033), .B(n3912), .Z(n9691) );
  XNOR U10512 ( .A(n9692), .B(n9693), .Z(n3912) );
  ANDN U10513 ( .B(n9694), .A(n9695), .Z(n9692) );
  XNOR U10514 ( .A(n9696), .B(n9697), .Z(n2033) );
  ANDN U10515 ( .B(n9698), .A(n9699), .Z(n9696) );
  XNOR U10516 ( .A(n9700), .B(n9701), .Z(n9690) );
  XNOR U10517 ( .A(n5350), .B(n5057), .Z(n9701) );
  XOR U10518 ( .A(n9702), .B(n9703), .Z(n5057) );
  ANDN U10519 ( .B(n9704), .A(n9705), .Z(n9702) );
  XNOR U10520 ( .A(n9706), .B(n9707), .Z(n5350) );
  NOR U10521 ( .A(n9708), .B(n9709), .Z(n9706) );
  XOR U10522 ( .A(n9710), .B(n6100), .Z(out[1026]) );
  XNOR U10523 ( .A(n8411), .B(n2516), .Z(n6100) );
  XNOR U10524 ( .A(n9711), .B(n9712), .Z(n2516) );
  XNOR U10525 ( .A(n9713), .B(n9714), .Z(n8411) );
  ANDN U10526 ( .B(n9715), .A(n9716), .Z(n9713) );
  ANDN U10527 ( .B(n1199), .A(n1201), .Z(n9710) );
  XNOR U10528 ( .A(n9717), .B(n1662), .Z(n1201) );
  XOR U10529 ( .A(n9718), .B(n9719), .Z(n8287) );
  XOR U10530 ( .A(n3436), .B(n5037), .Z(n9719) );
  XOR U10531 ( .A(n9720), .B(n9721), .Z(n5037) );
  ANDN U10532 ( .B(n9722), .A(n9703), .Z(n9720) );
  XOR U10533 ( .A(n9723), .B(n9724), .Z(n3436) );
  ANDN U10534 ( .B(n9697), .A(n9725), .Z(n9723) );
  XNOR U10535 ( .A(n9726), .B(n9727), .Z(n9718) );
  XNOR U10536 ( .A(n7272), .B(n2354), .Z(n9727) );
  XNOR U10537 ( .A(n9728), .B(n9729), .Z(n2354) );
  NOR U10538 ( .A(n9730), .B(n9731), .Z(n9728) );
  XOR U10539 ( .A(n9732), .B(n9733), .Z(n7272) );
  ANDN U10540 ( .B(n9734), .A(n9707), .Z(n9732) );
  XOR U10541 ( .A(n9735), .B(n9736), .Z(n6239) );
  XOR U10542 ( .A(n2040), .B(n3915), .Z(n9736) );
  XOR U10543 ( .A(n9737), .B(n9738), .Z(n3915) );
  XNOR U10544 ( .A(n9740), .B(n9741), .Z(n2040) );
  XOR U10545 ( .A(n9743), .B(n9744), .Z(n9735) );
  XOR U10546 ( .A(n5354), .B(n5094), .Z(n9744) );
  XNOR U10547 ( .A(n9745), .B(n9746), .Z(n5094) );
  NOR U10548 ( .A(n7335), .B(n9747), .Z(n9745) );
  XNOR U10549 ( .A(n9748), .B(n9749), .Z(n5354) );
  ANDN U10550 ( .B(n9750), .A(n8649), .Z(n9748) );
  XOR U10551 ( .A(n7447), .B(n3543), .Z(n1199) );
  IV U10552 ( .A(n2597), .Z(n3543) );
  XOR U10553 ( .A(n5977), .B(n6386), .Z(n2597) );
  XNOR U10554 ( .A(n9751), .B(n9752), .Z(n6386) );
  XOR U10555 ( .A(n2635), .B(n5368), .Z(n9752) );
  XNOR U10556 ( .A(n9753), .B(n6778), .Z(n5368) );
  XNOR U10557 ( .A(n9754), .B(n9755), .Z(n6778) );
  ANDN U10558 ( .B(n7453), .A(n7452), .Z(n9753) );
  XNOR U10559 ( .A(n9756), .B(n9757), .Z(n7452) );
  XNOR U10560 ( .A(n9758), .B(n9759), .Z(n7453) );
  XNOR U10561 ( .A(n9760), .B(n6782), .Z(n2635) );
  XOR U10562 ( .A(n9761), .B(n9762), .Z(n6782) );
  ANDN U10563 ( .B(n7442), .A(n7441), .Z(n9760) );
  XOR U10564 ( .A(n9763), .B(n9764), .Z(n7441) );
  XNOR U10565 ( .A(n9765), .B(n9766), .Z(n7442) );
  XOR U10566 ( .A(n3333), .B(n9767), .Z(n9751) );
  XOR U10567 ( .A(n5249), .B(n6772), .Z(n9767) );
  XNOR U10568 ( .A(n9768), .B(n7358), .Z(n6772) );
  IV U10569 ( .A(n6787), .Z(n7358) );
  XOR U10570 ( .A(n9280), .B(n9769), .Z(n6787) );
  ANDN U10571 ( .B(n6788), .A(n7449), .Z(n9768) );
  XNOR U10572 ( .A(n9770), .B(n9771), .Z(n7449) );
  XOR U10573 ( .A(n9772), .B(n9773), .Z(n6788) );
  XNOR U10574 ( .A(n9774), .B(n6792), .Z(n5249) );
  XOR U10575 ( .A(n9539), .B(n9775), .Z(n6792) );
  ANDN U10576 ( .B(n6791), .A(n9776), .Z(n9774) );
  XNOR U10577 ( .A(n9777), .B(n6796), .Z(n3333) );
  XNOR U10578 ( .A(n9778), .B(n9779), .Z(n6796) );
  AND U10579 ( .A(n6795), .B(n7444), .Z(n9777) );
  XNOR U10580 ( .A(n9780), .B(n9781), .Z(n7444) );
  XOR U10581 ( .A(n9782), .B(n9783), .Z(n6795) );
  XOR U10582 ( .A(n9784), .B(n9785), .Z(n5977) );
  XOR U10583 ( .A(n1838), .B(n5219), .Z(n9785) );
  XOR U10584 ( .A(n9786), .B(n7505), .Z(n5219) );
  ANDN U10585 ( .B(n7430), .A(n6812), .Z(n9786) );
  XOR U10586 ( .A(n9787), .B(n9788), .Z(n6812) );
  XNOR U10587 ( .A(n9789), .B(n9790), .Z(n7430) );
  XNOR U10588 ( .A(n9791), .B(n7501), .Z(n1838) );
  ANDN U10589 ( .B(n6820), .A(n7433), .Z(n9791) );
  XOR U10590 ( .A(n9792), .B(n9793), .Z(n7433) );
  XNOR U10591 ( .A(n9794), .B(n9795), .Z(n6820) );
  XOR U10592 ( .A(n4122), .B(n9796), .Z(n9784) );
  XNOR U10593 ( .A(n7480), .B(n3617), .Z(n9796) );
  XNOR U10594 ( .A(n9797), .B(n9798), .Z(n3617) );
  ANDN U10595 ( .B(n6816), .A(n7425), .Z(n9797) );
  XOR U10596 ( .A(n9799), .B(n9800), .Z(n6816) );
  XNOR U10597 ( .A(n9801), .B(n7498), .Z(n7480) );
  ANDN U10598 ( .B(n6807), .A(n7436), .Z(n9801) );
  XNOR U10599 ( .A(n9802), .B(n9803), .Z(n7436) );
  XNOR U10600 ( .A(n9804), .B(n9805), .Z(n6807) );
  XNOR U10601 ( .A(n9806), .B(n7507), .Z(n4122) );
  ANDN U10602 ( .B(n6803), .A(n7508), .Z(n9806) );
  XOR U10603 ( .A(n9807), .B(n9657), .Z(n7508) );
  IV U10604 ( .A(n9808), .Z(n9657) );
  XNOR U10605 ( .A(n9809), .B(n9810), .Z(n6803) );
  XNOR U10606 ( .A(n9811), .B(n6791), .Z(n7447) );
  XOR U10607 ( .A(n9812), .B(n9813), .Z(n6791) );
  NOR U10608 ( .A(n9655), .B(n7352), .Z(n9811) );
  XNOR U10609 ( .A(n9814), .B(n9815), .Z(n7352) );
  IV U10610 ( .A(n9776), .Z(n9655) );
  XNOR U10611 ( .A(n9816), .B(n9817), .Z(n9776) );
  XNOR U10612 ( .A(n9818), .B(n6105), .Z(out[1025]) );
  IV U10613 ( .A(n6418), .Z(n6105) );
  XNOR U10614 ( .A(n8496), .B(n2523), .Z(n6418) );
  XNOR U10615 ( .A(n9819), .B(n9820), .Z(n2523) );
  XOR U10616 ( .A(n9821), .B(n9822), .Z(n8496) );
  NOR U10617 ( .A(n9823), .B(n9824), .Z(n9821) );
  ANDN U10618 ( .B(n1203), .A(n1205), .Z(n9818) );
  XNOR U10619 ( .A(n9825), .B(n1667), .Z(n1205) );
  XOR U10620 ( .A(n9826), .B(n9827), .Z(n8341) );
  XNOR U10621 ( .A(n3439), .B(n5040), .Z(n9827) );
  XNOR U10622 ( .A(n9828), .B(n7336), .Z(n5040) );
  AND U10623 ( .A(n9746), .B(n7337), .Z(n9828) );
  XNOR U10624 ( .A(n9829), .B(n8397), .Z(n3439) );
  ANDN U10625 ( .B(n9741), .A(n8396), .Z(n9829) );
  XNOR U10626 ( .A(n2361), .B(n9830), .Z(n9826) );
  XOR U10627 ( .A(n3985), .B(n7329), .Z(n9830) );
  XNOR U10628 ( .A(n9831), .B(n8650), .Z(n7329) );
  AND U10629 ( .A(n9749), .B(n8651), .Z(n9831) );
  XOR U10630 ( .A(n9832), .B(n7343), .Z(n3985) );
  AND U10631 ( .A(n9738), .B(n7342), .Z(n9832) );
  XNOR U10632 ( .A(n9833), .B(n7347), .Z(n2361) );
  AND U10633 ( .A(n7346), .B(n9834), .Z(n9833) );
  XOR U10634 ( .A(n9835), .B(n9836), .Z(n6244) );
  XNOR U10635 ( .A(n2044), .B(n3604), .Z(n9836) );
  XOR U10636 ( .A(n9837), .B(n9838), .Z(n3604) );
  ANDN U10637 ( .B(n7414), .A(n9839), .Z(n9837) );
  XOR U10638 ( .A(n9840), .B(n9841), .Z(n2044) );
  NOR U10639 ( .A(n9842), .B(n8451), .Z(n9840) );
  XNOR U10640 ( .A(n9843), .B(n9844), .Z(n9835) );
  XNOR U10641 ( .A(n5359), .B(n5125), .Z(n9844) );
  XOR U10642 ( .A(n9845), .B(n9846), .Z(n5125) );
  NOR U10643 ( .A(n7408), .B(n9847), .Z(n9845) );
  IV U10644 ( .A(n9848), .Z(n7408) );
  XNOR U10645 ( .A(n9849), .B(n9850), .Z(n5359) );
  NOR U10646 ( .A(n9851), .B(n9399), .Z(n9849) );
  XOR U10647 ( .A(n7503), .B(n3546), .Z(n1203) );
  IV U10648 ( .A(n2602), .Z(n3546) );
  XOR U10649 ( .A(n5982), .B(n6390), .Z(n2602) );
  XNOR U10650 ( .A(n9852), .B(n9853), .Z(n6390) );
  XOR U10651 ( .A(n2642), .B(n5373), .Z(n9853) );
  XNOR U10652 ( .A(n9854), .B(n6804), .Z(n5373) );
  XOR U10653 ( .A(n9855), .B(n9856), .Z(n6804) );
  ANDN U10654 ( .B(n7507), .A(n6805), .Z(n9854) );
  XOR U10655 ( .A(n9857), .B(n9858), .Z(n6805) );
  XOR U10656 ( .A(n9859), .B(n9860), .Z(n7507) );
  XNOR U10657 ( .A(n9861), .B(n7437), .Z(n2642) );
  IV U10658 ( .A(n6809), .Z(n7437) );
  XNOR U10659 ( .A(n9862), .B(n9759), .Z(n6809) );
  NOR U10660 ( .A(n6808), .B(n7498), .Z(n9861) );
  XOR U10661 ( .A(n9863), .B(n9433), .Z(n7498) );
  IV U10662 ( .A(n9864), .Z(n9433) );
  XOR U10663 ( .A(n9865), .B(n9866), .Z(n6808) );
  XNOR U10664 ( .A(n3337), .B(n9867), .Z(n9852) );
  XOR U10665 ( .A(n5280), .B(n6798), .Z(n9867) );
  XNOR U10666 ( .A(n9868), .B(n7431), .Z(n6798) );
  IV U10667 ( .A(n6813), .Z(n7431) );
  XOR U10668 ( .A(n9869), .B(n9870), .Z(n6813) );
  ANDN U10669 ( .B(n6814), .A(n7505), .Z(n9868) );
  XOR U10670 ( .A(n9871), .B(n9872), .Z(n7505) );
  XOR U10671 ( .A(n9873), .B(n9874), .Z(n6814) );
  XNOR U10672 ( .A(n9875), .B(n6818), .Z(n5280) );
  XOR U10673 ( .A(n9876), .B(n9645), .Z(n6818) );
  ANDN U10674 ( .B(n9798), .A(n6817), .Z(n9875) );
  XOR U10675 ( .A(n9877), .B(n7434), .Z(n3337) );
  IV U10676 ( .A(n6822), .Z(n7434) );
  XOR U10677 ( .A(n9878), .B(n9879), .Z(n6822) );
  ANDN U10678 ( .B(n7501), .A(n6821), .Z(n9877) );
  XNOR U10679 ( .A(n9458), .B(n9880), .Z(n6821) );
  XNOR U10680 ( .A(n9114), .B(n9881), .Z(n7501) );
  XOR U10681 ( .A(n9882), .B(n9883), .Z(n5982) );
  XNOR U10682 ( .A(n1842), .B(n5221), .Z(n9883) );
  XNOR U10683 ( .A(n9884), .B(n7583), .Z(n5221) );
  ANDN U10684 ( .B(n7489), .A(n7490), .Z(n9884) );
  XOR U10685 ( .A(n9885), .B(n9886), .Z(n7490) );
  XOR U10686 ( .A(n9887), .B(n9888), .Z(n7489) );
  XNOR U10687 ( .A(n9889), .B(n7578), .Z(n1842) );
  NOR U10688 ( .A(n7579), .B(n6848), .Z(n9889) );
  XNOR U10689 ( .A(n9890), .B(n9891), .Z(n6848) );
  XNOR U10690 ( .A(n9892), .B(n9893), .Z(n7579) );
  XOR U10691 ( .A(n4125), .B(n9894), .Z(n9882) );
  XNOR U10692 ( .A(n7554), .B(n3627), .Z(n9894) );
  XNOR U10693 ( .A(n9895), .B(n9896), .Z(n3627) );
  ANDN U10694 ( .B(n6844), .A(n9897), .Z(n9895) );
  XOR U10695 ( .A(n9898), .B(n9899), .Z(n6844) );
  XNOR U10696 ( .A(n9900), .B(n7576), .Z(n7554) );
  NOR U10697 ( .A(n7494), .B(n6833), .Z(n9900) );
  XNOR U10698 ( .A(n9617), .B(n9901), .Z(n6833) );
  IV U10699 ( .A(n7575), .Z(n7494) );
  XOR U10700 ( .A(n9902), .B(n9322), .Z(n7575) );
  XNOR U10701 ( .A(n9903), .B(n7585), .Z(n4125) );
  AND U10702 ( .A(n7486), .B(n6830), .Z(n9903) );
  XOR U10703 ( .A(n9904), .B(n9905), .Z(n6830) );
  XOR U10704 ( .A(n9906), .B(n9907), .Z(n7486) );
  XNOR U10705 ( .A(n9909), .B(n9910), .Z(n6817) );
  ANDN U10706 ( .B(n7425), .A(n9798), .Z(n9908) );
  XOR U10707 ( .A(n9911), .B(n9912), .Z(n9798) );
  XOR U10708 ( .A(n9913), .B(n9891), .Z(n7425) );
  XOR U10709 ( .A(n9914), .B(n6110), .Z(out[1024]) );
  XOR U10710 ( .A(n8571), .B(n2530), .Z(n6110) );
  IV U10711 ( .A(n3277), .Z(n2530) );
  XOR U10712 ( .A(n9915), .B(n9916), .Z(n3277) );
  XNOR U10713 ( .A(n9917), .B(n9918), .Z(n8571) );
  NOR U10714 ( .A(n9919), .B(n8508), .Z(n9917) );
  ANDN U10715 ( .B(n1209), .A(n6421), .Z(n9914) );
  XOR U10716 ( .A(n7581), .B(n2613), .Z(n6421) );
  XNOR U10717 ( .A(n5987), .B(n6394), .Z(n2613) );
  XNOR U10718 ( .A(n9920), .B(n9921), .Z(n6394) );
  XOR U10719 ( .A(n2649), .B(n5377), .Z(n9921) );
  XOR U10720 ( .A(n9922), .B(n6832), .Z(n5377) );
  ANDN U10721 ( .B(n7585), .A(n6831), .Z(n9922) );
  XNOR U10722 ( .A(n9924), .B(n9925), .Z(n6831) );
  XOR U10723 ( .A(n9926), .B(n9927), .Z(n7585) );
  XOR U10724 ( .A(n9928), .B(n6837), .Z(n2649) );
  XOR U10725 ( .A(n9929), .B(n9930), .Z(n6837) );
  ANDN U10726 ( .B(n7576), .A(n7574), .Z(n9928) );
  XOR U10727 ( .A(n9931), .B(n9932), .Z(n7574) );
  XOR U10728 ( .A(n9522), .B(n9933), .Z(n7576) );
  XOR U10729 ( .A(n3341), .B(n9934), .Z(n9920) );
  XOR U10730 ( .A(n5314), .B(n6825), .Z(n9934) );
  XNOR U10731 ( .A(n9935), .B(n6842), .Z(n6825) );
  XNOR U10732 ( .A(n9936), .B(n9937), .Z(n6842) );
  ANDN U10733 ( .B(n7583), .A(n6841), .Z(n9935) );
  XOR U10734 ( .A(n9938), .B(n9939), .Z(n6841) );
  XNOR U10735 ( .A(n9940), .B(n9941), .Z(n7583) );
  XNOR U10736 ( .A(n9942), .B(n6846), .Z(n5314) );
  XOR U10737 ( .A(n9943), .B(n9790), .Z(n6846) );
  ANDN U10738 ( .B(n9896), .A(n6845), .Z(n9942) );
  XNOR U10739 ( .A(n9944), .B(n6850), .Z(n3341) );
  XOR U10740 ( .A(n9945), .B(n9946), .Z(n6850) );
  ANDN U10741 ( .B(n7578), .A(n6849), .Z(n9944) );
  XOR U10742 ( .A(n9559), .B(n9947), .Z(n6849) );
  XOR U10743 ( .A(n9948), .B(n9949), .Z(n7578) );
  XOR U10744 ( .A(n9950), .B(n9951), .Z(n5987) );
  XNOR U10745 ( .A(n1847), .B(n5224), .Z(n9951) );
  XNOR U10746 ( .A(n9952), .B(n7676), .Z(n5224) );
  ANDN U10747 ( .B(n6867), .A(n7558), .Z(n9952) );
  XOR U10748 ( .A(n9953), .B(n9954), .Z(n7558) );
  XNOR U10749 ( .A(n9955), .B(n9956), .Z(n6867) );
  XNOR U10750 ( .A(n9957), .B(n7672), .Z(n1847) );
  ANDN U10751 ( .B(n6875), .A(n7567), .Z(n9957) );
  XOR U10752 ( .A(n9958), .B(n9959), .Z(n7567) );
  XOR U10753 ( .A(n9960), .B(n9149), .Z(n6875) );
  XOR U10754 ( .A(n4131), .B(n9961), .Z(n9950) );
  XOR U10755 ( .A(n7653), .B(n3631), .Z(n9961) );
  XOR U10756 ( .A(n9962), .B(n9963), .Z(n3631) );
  ANDN U10757 ( .B(n6871), .A(n7564), .Z(n9962) );
  IV U10758 ( .A(n9964), .Z(n7564) );
  XNOR U10759 ( .A(n9227), .B(n9965), .Z(n6871) );
  IV U10760 ( .A(n9966), .Z(n9227) );
  XOR U10761 ( .A(n9967), .B(n9968), .Z(n7653) );
  ANDN U10762 ( .B(n7569), .A(n7570), .Z(n9967) );
  XOR U10763 ( .A(n9969), .B(n9757), .Z(n7570) );
  XNOR U10764 ( .A(n9970), .B(n7678), .Z(n4131) );
  ANDN U10765 ( .B(n7561), .A(n6858), .Z(n9970) );
  XNOR U10766 ( .A(n9971), .B(n9972), .Z(n6858) );
  XOR U10767 ( .A(n9973), .B(n9899), .Z(n7561) );
  XOR U10768 ( .A(n9974), .B(n6845), .Z(n7581) );
  XOR U10769 ( .A(n9975), .B(n9976), .Z(n6845) );
  NOR U10770 ( .A(n7484), .B(n9896), .Z(n9974) );
  XNOR U10771 ( .A(n9977), .B(n9978), .Z(n9896) );
  IV U10772 ( .A(n9897), .Z(n7484) );
  XOR U10773 ( .A(n9979), .B(n9149), .Z(n9897) );
  XNOR U10774 ( .A(n9980), .B(n4234), .Z(n1209) );
  IV U10775 ( .A(n1675), .Z(n4234) );
  XOR U10776 ( .A(n9981), .B(n9982), .Z(n8646) );
  XNOR U10777 ( .A(n3442), .B(n5044), .Z(n9982) );
  XOR U10778 ( .A(n9983), .B(n7409), .Z(n5044) );
  ANDN U10779 ( .B(n7410), .A(n9846), .Z(n9983) );
  XOR U10780 ( .A(n9984), .B(n8452), .Z(n3442) );
  NOR U10781 ( .A(n9841), .B(n8453), .Z(n9984) );
  XOR U10782 ( .A(n2368), .B(n9985), .Z(n9981) );
  XOR U10783 ( .A(n7402), .B(n3988), .Z(n9985) );
  XOR U10784 ( .A(n9986), .B(n7416), .Z(n3988) );
  AND U10785 ( .A(n7415), .B(n9838), .Z(n9986) );
  XNOR U10786 ( .A(n9987), .B(n9401), .Z(n7402) );
  NOR U10787 ( .A(n9400), .B(n9850), .Z(n9987) );
  XNOR U10788 ( .A(n9988), .B(n7420), .Z(n2368) );
  NOR U10789 ( .A(n9989), .B(n9990), .Z(n9988) );
  XOR U10790 ( .A(n9991), .B(n9992), .Z(n6248) );
  XNOR U10791 ( .A(n2048), .B(n3609), .Z(n9992) );
  XNOR U10792 ( .A(n9993), .B(n9994), .Z(n3609) );
  NOR U10793 ( .A(n7520), .B(n9995), .Z(n9993) );
  XOR U10794 ( .A(n9996), .B(n9997), .Z(n2048) );
  NOR U10795 ( .A(n8527), .B(n9998), .Z(n9996) );
  IV U10796 ( .A(n9999), .Z(n8527) );
  XNOR U10797 ( .A(n10000), .B(n10001), .Z(n9991) );
  XOR U10798 ( .A(n5367), .B(n5153), .Z(n10001) );
  NOR U10799 ( .A(n10004), .B(n7514), .Z(n10002) );
  XNOR U10800 ( .A(n10005), .B(n10006), .Z(n5367) );
  NOR U10801 ( .A(n10007), .B(n10008), .Z(n10005) );
  XOR U10802 ( .A(n10009), .B(n6113), .Z(out[1023]) );
  XOR U10803 ( .A(n7674), .B(n2622), .Z(n6113) );
  XOR U10804 ( .A(n10010), .B(n6873), .Z(n7674) );
  ANDN U10805 ( .B(n9963), .A(n9964), .Z(n10010) );
  XOR U10806 ( .A(n10011), .B(n9244), .Z(n9964) );
  ANDN U10807 ( .B(n5610), .A(n5608), .Z(n10009) );
  XNOR U10808 ( .A(n10012), .B(n1680), .Z(n5608) );
  IV U10809 ( .A(n4237), .Z(n1680) );
  XOR U10810 ( .A(n10013), .B(n10014), .Z(n9396) );
  XNOR U10811 ( .A(n3445), .B(n5048), .Z(n10014) );
  XOR U10812 ( .A(n10015), .B(n7515), .Z(n5048) );
  ANDN U10813 ( .B(n7516), .A(n10003), .Z(n10015) );
  XNOR U10814 ( .A(n10016), .B(n8528), .Z(n3445) );
  ANDN U10815 ( .B(n8529), .A(n9997), .Z(n10016) );
  XOR U10816 ( .A(n2375), .B(n10017), .Z(n10013) );
  XNOR U10817 ( .A(n7509), .B(n3993), .Z(n10017) );
  XOR U10818 ( .A(n10018), .B(n7521), .Z(n3993) );
  XNOR U10819 ( .A(n10019), .B(n10020), .Z(n7509) );
  ANDN U10820 ( .B(n10021), .A(n10006), .Z(n10019) );
  XNOR U10821 ( .A(n10022), .B(n7525), .Z(n2375) );
  ANDN U10822 ( .B(n7526), .A(n10023), .Z(n10022) );
  XOR U10823 ( .A(n10024), .B(n10025), .Z(n6253) );
  XOR U10824 ( .A(n5371), .B(n3615), .Z(n10025) );
  XOR U10825 ( .A(n10026), .B(n10027), .Z(n3615) );
  XNOR U10826 ( .A(n10029), .B(n10030), .Z(n5371) );
  ANDN U10827 ( .B(n10031), .A(n10032), .Z(n10029) );
  XOR U10828 ( .A(n10033), .B(n10034), .Z(n10024) );
  XOR U10829 ( .A(n2052), .B(n5181), .Z(n10034) );
  XNOR U10830 ( .A(n10035), .B(n10036), .Z(n5181) );
  ANDN U10831 ( .B(n7592), .A(n10037), .Z(n10035) );
  XNOR U10832 ( .A(n10038), .B(n10039), .Z(n2052) );
  ANDN U10833 ( .B(n10040), .A(n8654), .Z(n10038) );
  IV U10834 ( .A(n10041), .Z(n8654) );
  XOR U10835 ( .A(n9171), .B(n4871), .Z(n5610) );
  XNOR U10836 ( .A(n10042), .B(n8117), .Z(n4871) );
  XNOR U10837 ( .A(n10043), .B(n10044), .Z(n8117) );
  XNOR U10838 ( .A(n5399), .B(n3850), .Z(n10044) );
  XNOR U10839 ( .A(n10045), .B(n10046), .Z(n3850) );
  ANDN U10840 ( .B(n7993), .A(n7994), .Z(n10045) );
  XOR U10841 ( .A(n10047), .B(n10048), .Z(n7994) );
  XNOR U10842 ( .A(n10049), .B(n9209), .Z(n5399) );
  AND U10843 ( .A(n7989), .B(n7991), .Z(n10049) );
  XOR U10844 ( .A(n10050), .B(n10051), .Z(n7991) );
  XOR U10845 ( .A(n6207), .B(n10053), .Z(n10043) );
  XOR U10846 ( .A(n2227), .B(n4842), .Z(n10053) );
  XOR U10847 ( .A(n10054), .B(n9216), .Z(n4842) );
  ANDN U10848 ( .B(n8121), .A(n8119), .Z(n10054) );
  XOR U10849 ( .A(n10055), .B(n9557), .Z(n8119) );
  XNOR U10850 ( .A(n10056), .B(n10057), .Z(n8121) );
  XNOR U10851 ( .A(n10058), .B(n9213), .Z(n2227) );
  ANDN U10852 ( .B(n7979), .A(n7980), .Z(n10058) );
  XOR U10853 ( .A(n10059), .B(n10060), .Z(n7980) );
  XOR U10854 ( .A(n10061), .B(n10062), .Z(n7979) );
  XNOR U10855 ( .A(n10063), .B(n9219), .Z(n6207) );
  ANDN U10856 ( .B(n7983), .A(n7984), .Z(n10063) );
  XOR U10857 ( .A(n10064), .B(n10065), .Z(n7984) );
  XOR U10858 ( .A(n10066), .B(n10067), .Z(n7983) );
  XOR U10859 ( .A(n10068), .B(n9202), .Z(n9171) );
  NOR U10860 ( .A(n10069), .B(n8053), .Z(n10068) );
  XNOR U10861 ( .A(n10070), .B(n6116), .Z(out[1022]) );
  IV U10862 ( .A(n6474), .Z(n6116) );
  XOR U10863 ( .A(n7728), .B(n4939), .Z(n6474) );
  IV U10864 ( .A(n2627), .Z(n4939) );
  XOR U10865 ( .A(n5997), .B(n6636), .Z(n2627) );
  XNOR U10866 ( .A(n10071), .B(n10072), .Z(n6636) );
  XOR U10867 ( .A(n2663), .B(n5386), .Z(n10072) );
  XNOR U10868 ( .A(n10073), .B(n6887), .Z(n5386) );
  XOR U10869 ( .A(n10074), .B(n10075), .Z(n6887) );
  NOR U10870 ( .A(n7734), .B(n6886), .Z(n10073) );
  XOR U10871 ( .A(n10076), .B(n10077), .Z(n6886) );
  XNOR U10872 ( .A(n10078), .B(n6890), .Z(n2663) );
  XOR U10873 ( .A(n10079), .B(n10080), .Z(n6890) );
  ANDN U10874 ( .B(n6891), .A(n10081), .Z(n10078) );
  XOR U10875 ( .A(n10082), .B(n10083), .Z(n6891) );
  XNOR U10876 ( .A(n3352), .B(n10084), .Z(n10071) );
  XNOR U10877 ( .A(n5413), .B(n6880), .Z(n10084) );
  XNOR U10878 ( .A(n10085), .B(n6908), .Z(n6880) );
  XOR U10879 ( .A(n9671), .B(n10086), .Z(n6908) );
  NOR U10880 ( .A(n7730), .B(n7731), .Z(n10085) );
  XOR U10881 ( .A(n10087), .B(n10088), .Z(n7730) );
  XNOR U10882 ( .A(n10089), .B(n6897), .Z(n5413) );
  XNOR U10883 ( .A(n10090), .B(n9954), .Z(n6897) );
  ANDN U10884 ( .B(n6896), .A(n10091), .Z(n10089) );
  XOR U10885 ( .A(n10092), .B(n6901), .Z(n3352) );
  XOR U10886 ( .A(n10093), .B(n10094), .Z(n6901) );
  ANDN U10887 ( .B(n6900), .A(n7725), .Z(n10092) );
  XOR U10888 ( .A(n10095), .B(n10096), .Z(n6900) );
  XOR U10889 ( .A(n10097), .B(n10098), .Z(n5997) );
  XNOR U10890 ( .A(n1855), .B(n5230), .Z(n10098) );
  XOR U10891 ( .A(n10099), .B(n7817), .Z(n5230) );
  ANDN U10892 ( .B(n7709), .A(n7241), .Z(n10099) );
  XNOR U10893 ( .A(n10100), .B(n10101), .Z(n7241) );
  XOR U10894 ( .A(n10102), .B(n10103), .Z(n7709) );
  XOR U10895 ( .A(n10104), .B(n7813), .Z(n1855) );
  ANDN U10896 ( .B(n6933), .A(n7717), .Z(n10104) );
  XOR U10897 ( .A(n10105), .B(n10106), .Z(n7717) );
  XOR U10898 ( .A(n10107), .B(n10108), .Z(n6933) );
  XNOR U10899 ( .A(n4137), .B(n10109), .Z(n10097) );
  XOR U10900 ( .A(n7805), .B(n3642), .Z(n10109) );
  XOR U10901 ( .A(n10110), .B(n10111), .Z(n3642) );
  ANDN U10902 ( .B(n7719), .A(n6929), .Z(n10110) );
  XOR U10903 ( .A(n10112), .B(n10113), .Z(n6929) );
  XOR U10904 ( .A(n10114), .B(n7811), .Z(n7805) );
  AND U10905 ( .A(n6921), .B(n7715), .Z(n10114) );
  XOR U10906 ( .A(n10115), .B(n9613), .Z(n7715) );
  XOR U10907 ( .A(n10116), .B(n10117), .Z(n6921) );
  XOR U10908 ( .A(n10118), .B(n7819), .Z(n4137) );
  ANDN U10909 ( .B(n6918), .A(n7712), .Z(n10118) );
  IV U10910 ( .A(n7820), .Z(n7712) );
  XOR U10911 ( .A(n10119), .B(n10120), .Z(n7820) );
  XOR U10912 ( .A(n10121), .B(n10122), .Z(n6918) );
  XNOR U10913 ( .A(n10123), .B(n6896), .Z(n7728) );
  XOR U10914 ( .A(n10124), .B(n10125), .Z(n6896) );
  ANDN U10915 ( .B(n10091), .A(n7662), .Z(n10123) );
  IV U10916 ( .A(n10126), .Z(n7662) );
  AND U10917 ( .A(n5614), .B(n5612), .Z(n10070) );
  XOR U10918 ( .A(n10127), .B(n1685), .Z(n5612) );
  XNOR U10919 ( .A(n10128), .B(n6257), .Z(n1685) );
  XNOR U10920 ( .A(n10129), .B(n10130), .Z(n6257) );
  XNOR U10921 ( .A(n5375), .B(n3618), .Z(n10130) );
  XNOR U10922 ( .A(n10131), .B(n10132), .Z(n3618) );
  AND U10923 ( .A(n10133), .B(n7650), .Z(n10131) );
  XNOR U10924 ( .A(n10134), .B(n10135), .Z(n5375) );
  ANDN U10925 ( .B(n10136), .A(n7646), .Z(n10134) );
  XOR U10926 ( .A(n10137), .B(n10138), .Z(n10129) );
  XNOR U10927 ( .A(n2055), .B(n5214), .Z(n10138) );
  XNOR U10928 ( .A(n10139), .B(n10140), .Z(n5214) );
  AND U10929 ( .A(n10141), .B(n7637), .Z(n10139) );
  XNOR U10930 ( .A(n10142), .B(n10143), .Z(n2055) );
  NOR U10931 ( .A(n10144), .B(n8714), .Z(n10142) );
  XOR U10932 ( .A(n9206), .B(n5331), .Z(n5614) );
  XNOR U10933 ( .A(n10145), .B(n8180), .Z(n5331) );
  XNOR U10934 ( .A(n10146), .B(n10147), .Z(n8180) );
  XOR U10935 ( .A(n5403), .B(n3855), .Z(n10147) );
  XNOR U10936 ( .A(n10148), .B(n10149), .Z(n3855) );
  ANDN U10937 ( .B(n8645), .A(n10150), .Z(n10148) );
  XNOR U10938 ( .A(n10151), .B(n10152), .Z(n8645) );
  XNOR U10939 ( .A(n10153), .B(n9303), .Z(n5403) );
  ANDN U10940 ( .B(n8637), .A(n9304), .Z(n10153) );
  XOR U10941 ( .A(n9532), .B(n10154), .Z(n9304) );
  XOR U10942 ( .A(n10155), .B(n9879), .Z(n8637) );
  XNOR U10943 ( .A(n6212), .B(n10156), .Z(n10146) );
  XNOR U10944 ( .A(n2240), .B(n4872), .Z(n10156) );
  XNOR U10945 ( .A(n10157), .B(n9312), .Z(n4872) );
  ANDN U10946 ( .B(n8641), .A(n8639), .Z(n10157) );
  IV U10947 ( .A(n9311), .Z(n8639) );
  XOR U10948 ( .A(n10158), .B(n9413), .Z(n9311) );
  XOR U10949 ( .A(n10159), .B(n10160), .Z(n8641) );
  XOR U10950 ( .A(n10161), .B(n9308), .Z(n2240) );
  ANDN U10951 ( .B(n8627), .A(n8626), .Z(n10161) );
  XOR U10952 ( .A(n9138), .B(n10162), .Z(n8626) );
  XOR U10953 ( .A(n10163), .B(n10164), .Z(n8627) );
  XOR U10954 ( .A(n10165), .B(n10166), .Z(n6212) );
  ANDN U10955 ( .B(n8631), .A(n8630), .Z(n10165) );
  XOR U10956 ( .A(n10167), .B(n10168), .Z(n8630) );
  XOR U10957 ( .A(n9527), .B(n10169), .Z(n8631) );
  XOR U10958 ( .A(n10170), .B(n9295), .Z(n9206) );
  XOR U10959 ( .A(n10171), .B(n10172), .Z(n7993) );
  XOR U10960 ( .A(n10173), .B(n6125), .Z(out[1021]) );
  XOR U10961 ( .A(n7815), .B(n2634), .Z(n6125) );
  XNOR U10962 ( .A(n6002), .B(n6905), .Z(n2634) );
  XNOR U10963 ( .A(n10174), .B(n10175), .Z(n6905) );
  XOR U10964 ( .A(n2670), .B(n5392), .Z(n10175) );
  XNOR U10965 ( .A(n10176), .B(n6920), .Z(n5392) );
  XOR U10966 ( .A(n10177), .B(n10178), .Z(n6920) );
  ANDN U10967 ( .B(n6919), .A(n7819), .Z(n10176) );
  XNOR U10968 ( .A(n10179), .B(n10180), .Z(n7819) );
  XOR U10969 ( .A(n10181), .B(n10182), .Z(n6919) );
  XNOR U10970 ( .A(n10183), .B(n6924), .Z(n2670) );
  XOR U10971 ( .A(n10184), .B(n10185), .Z(n6924) );
  ANDN U10972 ( .B(n7811), .A(n7810), .Z(n10183) );
  XOR U10973 ( .A(n10186), .B(n10187), .Z(n7810) );
  XNOR U10974 ( .A(n9458), .B(n10188), .Z(n7811) );
  XOR U10975 ( .A(n3355), .B(n10189), .Z(n10174) );
  XNOR U10976 ( .A(n5461), .B(n6913), .Z(n10189) );
  XNOR U10977 ( .A(n10190), .B(n7710), .Z(n6913) );
  IV U10978 ( .A(n7242), .Z(n7710) );
  XOR U10979 ( .A(n10191), .B(n9817), .Z(n7242) );
  ANDN U10980 ( .B(n7243), .A(n7817), .Z(n10190) );
  XOR U10981 ( .A(n10192), .B(n10193), .Z(n7817) );
  XOR U10982 ( .A(n10194), .B(n10195), .Z(n7243) );
  XOR U10983 ( .A(n10196), .B(n6930), .Z(n5461) );
  XNOR U10984 ( .A(n10197), .B(n10198), .Z(n6930) );
  ANDN U10985 ( .B(n6931), .A(n10111), .Z(n10196) );
  XNOR U10986 ( .A(n10199), .B(n6935), .Z(n3355) );
  XOR U10987 ( .A(n10200), .B(n10201), .Z(n6935) );
  ANDN U10988 ( .B(n6934), .A(n7813), .Z(n10199) );
  XOR U10989 ( .A(n10202), .B(n10203), .Z(n7813) );
  XOR U10990 ( .A(n10204), .B(n10205), .Z(n6934) );
  XOR U10991 ( .A(n10206), .B(n10207), .Z(n6002) );
  XNOR U10992 ( .A(n5233), .B(n1859), .Z(n10207) );
  XOR U10993 ( .A(n10208), .B(n7853), .Z(n1859) );
  NOR U10994 ( .A(n6958), .B(n7854), .Z(n10208) );
  XNOR U10995 ( .A(n10209), .B(n10210), .Z(n7854) );
  XOR U10996 ( .A(n10211), .B(n9426), .Z(n6958) );
  XNOR U10997 ( .A(n10212), .B(n7861), .Z(n5233) );
  ANDN U10998 ( .B(n7862), .A(n7963), .Z(n10212) );
  XNOR U10999 ( .A(n9132), .B(n10213), .Z(n7963) );
  XNOR U11000 ( .A(n10214), .B(n10215), .Z(n7862) );
  XNOR U11001 ( .A(n3646), .B(n10216), .Z(n10206) );
  XNOR U11002 ( .A(n7847), .B(n4140), .Z(n10216) );
  XNOR U11003 ( .A(n10217), .B(n7865), .Z(n4140) );
  NOR U11004 ( .A(n6943), .B(n7864), .Z(n10217) );
  XOR U11005 ( .A(n10218), .B(n10219), .Z(n7864) );
  XNOR U11006 ( .A(n10220), .B(n10221), .Z(n6943) );
  XOR U11007 ( .A(n10222), .B(n7858), .Z(n7847) );
  ANDN U11008 ( .B(n6946), .A(n7857), .Z(n10222) );
  XNOR U11009 ( .A(n10223), .B(n9755), .Z(n7857) );
  XOR U11010 ( .A(n10224), .B(n10225), .Z(n6946) );
  XOR U11011 ( .A(n10226), .B(n10227), .Z(n3646) );
  ANDN U11012 ( .B(n7969), .A(n6954), .Z(n10226) );
  XNOR U11013 ( .A(n9520), .B(n10228), .Z(n6954) );
  XNOR U11014 ( .A(n10229), .B(n6931), .Z(n7815) );
  XOR U11015 ( .A(n10230), .B(n10231), .Z(n6931) );
  ANDN U11016 ( .B(n10111), .A(n7719), .Z(n10229) );
  XOR U11017 ( .A(n10232), .B(n9426), .Z(n7719) );
  XNOR U11018 ( .A(n10233), .B(n10234), .Z(n10111) );
  NOR U11019 ( .A(n5618), .B(n5616), .Z(n10173) );
  XOR U11020 ( .A(n10235), .B(n1689), .Z(n5616) );
  XNOR U11021 ( .A(n10236), .B(n6261), .Z(n1689) );
  XNOR U11022 ( .A(n10237), .B(n10238), .Z(n6261) );
  XOR U11023 ( .A(n5379), .B(n3628), .Z(n10238) );
  XOR U11024 ( .A(n10239), .B(n10240), .Z(n3628) );
  AND U11025 ( .A(n10241), .B(n7754), .Z(n10239) );
  XNOR U11026 ( .A(n10242), .B(n10243), .Z(n5379) );
  NOR U11027 ( .A(n10244), .B(n7750), .Z(n10242) );
  XOR U11028 ( .A(n10245), .B(n10246), .Z(n10237) );
  XOR U11029 ( .A(n2058), .B(n5248), .Z(n10246) );
  XNOR U11030 ( .A(n10247), .B(n10248), .Z(n5248) );
  ANDN U11031 ( .B(n7741), .A(n10249), .Z(n10247) );
  XNOR U11032 ( .A(n10250), .B(n10251), .Z(n2058) );
  ANDN U11033 ( .B(n10252), .A(n8780), .Z(n10250) );
  XNOR U11034 ( .A(n9300), .B(n2025), .Z(n5618) );
  XNOR U11035 ( .A(n7975), .B(n8234), .Z(n2025) );
  XNOR U11036 ( .A(n10253), .B(n10254), .Z(n8234) );
  XOR U11037 ( .A(n5408), .B(n3859), .Z(n10254) );
  XNOR U11038 ( .A(n10255), .B(n10256), .Z(n3859) );
  ANDN U11039 ( .B(n9395), .A(n10257), .Z(n10255) );
  XNOR U11040 ( .A(n10258), .B(n9329), .Z(n9395) );
  XNOR U11041 ( .A(n10259), .B(n9484), .Z(n5408) );
  ANDN U11042 ( .B(n9385), .A(n9386), .Z(n10259) );
  XOR U11043 ( .A(n10260), .B(n9946), .Z(n9386) );
  XNOR U11044 ( .A(n9630), .B(n10261), .Z(n9385) );
  XOR U11045 ( .A(n6217), .B(n10262), .Z(n10253) );
  XOR U11046 ( .A(n2247), .B(n4911), .Z(n10262) );
  XNOR U11047 ( .A(n10263), .B(n9491), .Z(n4911) );
  ANDN U11048 ( .B(n9391), .A(n9389), .Z(n10263) );
  IV U11049 ( .A(n9492), .Z(n9389) );
  XOR U11050 ( .A(n9509), .B(n10264), .Z(n9492) );
  XNOR U11051 ( .A(n10265), .B(n10266), .Z(n9391) );
  XNOR U11052 ( .A(n10267), .B(n9488), .Z(n2247) );
  ANDN U11053 ( .B(n9376), .A(n9579), .Z(n10267) );
  XOR U11054 ( .A(n10268), .B(n10269), .Z(n9579) );
  XNOR U11055 ( .A(n9623), .B(n10270), .Z(n9376) );
  XOR U11056 ( .A(n10271), .B(n9495), .Z(n6217) );
  ANDN U11057 ( .B(n9380), .A(n9381), .Z(n10271) );
  XOR U11058 ( .A(n9439), .B(n10272), .Z(n9381) );
  XOR U11059 ( .A(n10273), .B(n10274), .Z(n9380) );
  XOR U11060 ( .A(n10275), .B(n10276), .Z(n7975) );
  XOR U11061 ( .A(n1960), .B(n9467), .Z(n10276) );
  XNOR U11062 ( .A(n10277), .B(n8636), .Z(n9467) );
  IV U11063 ( .A(n9478), .Z(n8636) );
  XOR U11064 ( .A(n10278), .B(n10279), .Z(n9478) );
  NOR U11065 ( .A(n9302), .B(n9303), .Z(n10277) );
  XOR U11066 ( .A(n10280), .B(n10281), .Z(n9303) );
  XOR U11067 ( .A(n10282), .B(n10283), .Z(n9302) );
  XNOR U11068 ( .A(n10284), .B(n8632), .Z(n1960) );
  XNOR U11069 ( .A(n10285), .B(n9463), .Z(n8632) );
  ANDN U11070 ( .B(n9314), .A(n9315), .Z(n10284) );
  IV U11071 ( .A(n10166), .Z(n9315) );
  XOR U11072 ( .A(n10286), .B(n10287), .Z(n10166) );
  XOR U11073 ( .A(n10288), .B(n10234), .Z(n9314) );
  XNOR U11074 ( .A(n3754), .B(n10289), .Z(n10275) );
  XNOR U11075 ( .A(n5106), .B(n4214), .Z(n10289) );
  XOR U11076 ( .A(n10290), .B(n8644), .Z(n4214) );
  NOR U11077 ( .A(n10149), .B(n9475), .Z(n10290) );
  XOR U11078 ( .A(n10292), .B(n9472), .Z(n5106) );
  IV U11079 ( .A(n8640), .Z(n9472) );
  XOR U11080 ( .A(n10293), .B(n9764), .Z(n8640) );
  ANDN U11081 ( .B(n9312), .A(n9310), .Z(n10292) );
  XOR U11082 ( .A(n9623), .B(n10294), .Z(n9310) );
  XOR U11083 ( .A(n10295), .B(n10296), .Z(n9312) );
  XNOR U11084 ( .A(n10297), .B(n8628), .Z(n3754) );
  XOR U11085 ( .A(n10116), .B(n10298), .Z(n8628) );
  ANDN U11086 ( .B(n9307), .A(n9308), .Z(n10297) );
  XOR U11087 ( .A(n10299), .B(n10300), .Z(n9308) );
  XNOR U11088 ( .A(n10301), .B(n10302), .Z(n9307) );
  XNOR U11089 ( .A(n10303), .B(n9475), .Z(n9300) );
  XOR U11090 ( .A(n10304), .B(n10305), .Z(n9475) );
  ANDN U11091 ( .B(n10149), .A(n8643), .Z(n10303) );
  IV U11092 ( .A(n10150), .Z(n8643) );
  XNOR U11093 ( .A(n10306), .B(n10307), .Z(n10150) );
  XOR U11094 ( .A(n10308), .B(n9645), .Z(n10149) );
  XOR U11095 ( .A(n10309), .B(n6130), .Z(out[1020]) );
  XNOR U11096 ( .A(n7851), .B(n2641), .Z(n6130) );
  XNOR U11097 ( .A(n6007), .B(n7239), .Z(n2641) );
  XNOR U11098 ( .A(n10310), .B(n10311), .Z(n7239) );
  XNOR U11099 ( .A(n2677), .B(n5396), .Z(n10311) );
  XNOR U11100 ( .A(n10312), .B(n6944), .Z(n5396) );
  XOR U11101 ( .A(n10313), .B(n10314), .Z(n6944) );
  ANDN U11102 ( .B(n7865), .A(n6945), .Z(n10312) );
  XOR U11103 ( .A(n10315), .B(n10316), .Z(n6945) );
  XOR U11104 ( .A(n10317), .B(n10318), .Z(n7865) );
  XOR U11105 ( .A(n10319), .B(n6949), .Z(n2677) );
  XNOR U11106 ( .A(n10320), .B(n10180), .Z(n6949) );
  ANDN U11107 ( .B(n6950), .A(n7858), .Z(n10319) );
  XOR U11108 ( .A(n10321), .B(n10322), .Z(n7858) );
  XNOR U11109 ( .A(n10323), .B(n10324), .Z(n6950) );
  XNOR U11110 ( .A(n3359), .B(n10325), .Z(n10310) );
  XNOR U11111 ( .A(n5514), .B(n6938), .Z(n10325) );
  XNOR U11112 ( .A(n10326), .B(n7964), .Z(n6938) );
  XOR U11113 ( .A(n10327), .B(n9912), .Z(n7964) );
  ANDN U11114 ( .B(n7861), .A(n7972), .Z(n10326) );
  XNOR U11115 ( .A(n10328), .B(n10329), .Z(n7972) );
  XNOR U11116 ( .A(n10330), .B(n10331), .Z(n7861) );
  XNOR U11117 ( .A(n10332), .B(n6955), .Z(n5514) );
  XOR U11118 ( .A(n10333), .B(n10103), .Z(n6955) );
  ANDN U11119 ( .B(n6956), .A(n10227), .Z(n10332) );
  XNOR U11120 ( .A(n10334), .B(n6959), .Z(n3359) );
  XOR U11121 ( .A(n10335), .B(n9424), .Z(n6959) );
  ANDN U11122 ( .B(n6960), .A(n7853), .Z(n10334) );
  XNOR U11123 ( .A(n9659), .B(n10336), .Z(n7853) );
  XOR U11124 ( .A(n10337), .B(n10338), .Z(n6960) );
  XOR U11125 ( .A(n10339), .B(n10340), .Z(n6007) );
  XOR U11126 ( .A(n5236), .B(n1863), .Z(n10340) );
  XNOR U11127 ( .A(n10341), .B(n7922), .Z(n1863) );
  ANDN U11128 ( .B(n8608), .A(n8607), .Z(n10341) );
  XOR U11129 ( .A(n10342), .B(n10343), .Z(n8607) );
  XOR U11130 ( .A(n10344), .B(n7930), .Z(n5236) );
  NOR U11131 ( .A(n8603), .B(n8604), .Z(n10344) );
  XNOR U11132 ( .A(n10345), .B(n10346), .Z(n8603) );
  XNOR U11133 ( .A(n3650), .B(n10347), .Z(n10339) );
  XOR U11134 ( .A(n7914), .B(n4143), .Z(n10347) );
  XOR U11135 ( .A(n10348), .B(n7934), .Z(n4143) );
  ANDN U11136 ( .B(n7935), .A(n8619), .Z(n10348) );
  XOR U11137 ( .A(n9520), .B(n10349), .Z(n7935) );
  XNOR U11138 ( .A(n10350), .B(n7927), .Z(n7914) );
  IV U11139 ( .A(n10351), .Z(n7927) );
  NOR U11140 ( .A(n8612), .B(n7926), .Z(n10350) );
  XNOR U11141 ( .A(n10352), .B(n9856), .Z(n7926) );
  XNOR U11142 ( .A(n10353), .B(n10354), .Z(n3650) );
  ANDN U11143 ( .B(n8617), .A(n8615), .Z(n10353) );
  XNOR U11144 ( .A(n10355), .B(n6956), .Z(n7851) );
  XNOR U11145 ( .A(n10356), .B(n10357), .Z(n6956) );
  XOR U11146 ( .A(n9532), .B(n10358), .Z(n7969) );
  IV U11147 ( .A(n10359), .Z(n9532) );
  XOR U11148 ( .A(n10360), .B(n10361), .Z(n10227) );
  ANDN U11149 ( .B(n5620), .A(n5622), .Z(n10309) );
  XNOR U11150 ( .A(n9481), .B(n2028), .Z(n5622) );
  XNOR U11151 ( .A(n8622), .B(n8288), .Z(n2028) );
  XNOR U11152 ( .A(n10362), .B(n10363), .Z(n8288) );
  XOR U11153 ( .A(n5418), .B(n3863), .Z(n10363) );
  XNOR U11154 ( .A(n10364), .B(n10365), .Z(n3863) );
  NOR U11155 ( .A(n10366), .B(n9684), .Z(n10364) );
  XNOR U11156 ( .A(n10367), .B(n9586), .Z(n5418) );
  ANDN U11157 ( .B(n9587), .A(n10368), .Z(n10367) );
  XOR U11158 ( .A(n6222), .B(n10369), .Z(n10362) );
  XNOR U11159 ( .A(n2254), .B(n4949), .Z(n10369) );
  XNOR U11160 ( .A(n10370), .B(n9590), .Z(n4949) );
  ANDN U11161 ( .B(n9679), .A(n10371), .Z(n10370) );
  XNOR U11162 ( .A(n10372), .B(n9600), .Z(n2254) );
  NOR U11163 ( .A(n10373), .B(n9688), .Z(n10372) );
  XOR U11164 ( .A(n10374), .B(n9596), .Z(n6222) );
  ANDN U11165 ( .B(n9676), .A(n10375), .Z(n10374) );
  XOR U11166 ( .A(n10376), .B(n10377), .Z(n8622) );
  XNOR U11167 ( .A(n1968), .B(n9568), .Z(n10377) );
  XNOR U11168 ( .A(n10378), .B(n9581), .Z(n9568) );
  IV U11169 ( .A(n9387), .Z(n9581) );
  XNOR U11170 ( .A(n10379), .B(n9224), .Z(n9387) );
  AND U11171 ( .A(n9483), .B(n9484), .Z(n10378) );
  XNOR U11172 ( .A(n10380), .B(n10381), .Z(n9484) );
  XNOR U11173 ( .A(n10382), .B(n10125), .Z(n9483) );
  XNOR U11174 ( .A(n10383), .B(n9382), .Z(n1968) );
  XOR U11175 ( .A(n9563), .B(n10384), .Z(n9382) );
  ANDN U11176 ( .B(n9495), .A(n9494), .Z(n10383) );
  XOR U11177 ( .A(n10360), .B(n10385), .Z(n9494) );
  IV U11178 ( .A(n10386), .Z(n10360) );
  XOR U11179 ( .A(n10387), .B(n10388), .Z(n9495) );
  XNOR U11180 ( .A(n3759), .B(n10389), .Z(n10376) );
  XOR U11181 ( .A(n5109), .B(n4218), .Z(n10389) );
  XOR U11182 ( .A(n10390), .B(n9577), .Z(n4218) );
  IV U11183 ( .A(n9394), .Z(n9577) );
  XOR U11184 ( .A(n10391), .B(n9773), .Z(n9394) );
  NOR U11185 ( .A(n10256), .B(n9576), .Z(n10390) );
  XOR U11186 ( .A(n10392), .B(n9573), .Z(n5109) );
  IV U11187 ( .A(n9390), .Z(n9573) );
  XOR U11188 ( .A(n10393), .B(n9866), .Z(n9390) );
  NOR U11189 ( .A(n9491), .B(n9490), .Z(n10392) );
  XNOR U11190 ( .A(n9765), .B(n10394), .Z(n9490) );
  XOR U11191 ( .A(n10395), .B(n10396), .Z(n9491) );
  XNOR U11192 ( .A(n10397), .B(n9378), .Z(n3759) );
  XOR U11193 ( .A(n10224), .B(n10398), .Z(n9378) );
  ANDN U11194 ( .B(n9487), .A(n9488), .Z(n10397) );
  XNOR U11195 ( .A(n10399), .B(n10400), .Z(n9488) );
  XNOR U11196 ( .A(n10401), .B(n10402), .Z(n9487) );
  XNOR U11197 ( .A(n10403), .B(n9576), .Z(n9481) );
  XOR U11198 ( .A(n10404), .B(n10300), .Z(n9576) );
  ANDN U11199 ( .B(n10256), .A(n9393), .Z(n10403) );
  IV U11200 ( .A(n10257), .Z(n9393) );
  XOR U11201 ( .A(n10405), .B(n10406), .Z(n10257) );
  XNOR U11202 ( .A(n10407), .B(n9790), .Z(n10256) );
  XOR U11203 ( .A(n10408), .B(n1693), .Z(n5620) );
  XNOR U11204 ( .A(n8718), .B(n6265), .Z(n1693) );
  XNOR U11205 ( .A(n10409), .B(n10410), .Z(n6265) );
  XNOR U11206 ( .A(n5385), .B(n3632), .Z(n10410) );
  XNOR U11207 ( .A(n10411), .B(n10412), .Z(n3632) );
  ANDN U11208 ( .B(n10413), .A(n7798), .Z(n10411) );
  IV U11209 ( .A(n10414), .Z(n7798) );
  XOR U11210 ( .A(n10415), .B(n10416), .Z(n5385) );
  AND U11211 ( .A(n7788), .B(n10417), .Z(n10415) );
  XOR U11212 ( .A(n10418), .B(n10419), .Z(n10409) );
  XOR U11213 ( .A(n2062), .B(n5278), .Z(n10419) );
  XNOR U11214 ( .A(n10420), .B(n10421), .Z(n5278) );
  ANDN U11215 ( .B(n10422), .A(n7792), .Z(n10420) );
  IV U11216 ( .A(n10423), .Z(n7792) );
  XNOR U11217 ( .A(n10424), .B(n10425), .Z(n2062) );
  ANDN U11218 ( .B(n10426), .A(n10427), .Z(n10424) );
  XOR U11219 ( .A(n10428), .B(n10429), .Z(n8718) );
  XOR U11220 ( .A(n5060), .B(n7735), .Z(n10429) );
  XNOR U11221 ( .A(n10430), .B(n7751), .Z(n7735) );
  ANDN U11222 ( .B(n10243), .A(n7752), .Z(n10430) );
  XNOR U11223 ( .A(n10431), .B(n7742), .Z(n5060) );
  XOR U11224 ( .A(n2397), .B(n10432), .Z(n10428) );
  XNOR U11225 ( .A(n3454), .B(n4002), .Z(n10432) );
  XOR U11226 ( .A(n10433), .B(n7756), .Z(n4002) );
  IV U11227 ( .A(n10434), .Z(n7756) );
  ANDN U11228 ( .B(n10240), .A(n7755), .Z(n10433) );
  XNOR U11229 ( .A(n10435), .B(n8781), .Z(n3454) );
  ANDN U11230 ( .B(n10251), .A(n10436), .Z(n10435) );
  XOR U11231 ( .A(n10437), .B(n7747), .Z(n2397) );
  ANDN U11232 ( .B(n7748), .A(n10438), .Z(n10437) );
  XOR U11233 ( .A(n10439), .B(n4202), .Z(out[101]) );
  XOR U11234 ( .A(n7001), .B(n2572), .Z(n4202) );
  XOR U11235 ( .A(n8046), .B(n10440), .Z(n2572) );
  XOR U11236 ( .A(n10441), .B(n10442), .Z(n8046) );
  XOR U11237 ( .A(n4381), .B(n2190), .Z(n10442) );
  XNOR U11238 ( .A(n10443), .B(n8110), .Z(n2190) );
  IV U11239 ( .A(n10444), .Z(n8110) );
  NOR U11240 ( .A(n10445), .B(n10446), .Z(n10443) );
  XNOR U11241 ( .A(n10447), .B(n8102), .Z(n4381) );
  XOR U11242 ( .A(n6021), .B(n10448), .Z(n10441) );
  XOR U11243 ( .A(n5554), .B(n3804), .Z(n10448) );
  XNOR U11244 ( .A(n10449), .B(n8106), .Z(n3804) );
  IV U11245 ( .A(n10450), .Z(n8106) );
  AND U11246 ( .A(n6999), .B(n6997), .Z(n10449) );
  XOR U11247 ( .A(n10451), .B(n10452), .Z(n5554) );
  NOR U11248 ( .A(n7005), .B(n7003), .Z(n10451) );
  XNOR U11249 ( .A(n10453), .B(n8114), .Z(n6021) );
  XNOR U11250 ( .A(n10454), .B(n10446), .Z(n7001) );
  ANDN U11251 ( .B(n3624), .A(n4376), .Z(n10439) );
  XNOR U11252 ( .A(n7512), .B(n2412), .Z(n4376) );
  XNOR U11253 ( .A(n10128), .B(n10455), .Z(n2412) );
  XOR U11254 ( .A(n10456), .B(n10457), .Z(n10128) );
  XOR U11255 ( .A(n3448), .B(n5051), .Z(n10457) );
  XOR U11256 ( .A(n10458), .B(n7593), .Z(n5051) );
  ANDN U11257 ( .B(n10036), .A(n10459), .Z(n10458) );
  XNOR U11258 ( .A(n10460), .B(n8656), .Z(n3448) );
  ANDN U11259 ( .B(n10039), .A(n8655), .Z(n10460) );
  XNOR U11260 ( .A(n2382), .B(n10461), .Z(n10456) );
  XOR U11261 ( .A(n7586), .B(n3996), .Z(n10461) );
  XOR U11262 ( .A(n10462), .B(n7599), .Z(n3996) );
  ANDN U11263 ( .B(n10027), .A(n7600), .Z(n10462) );
  XNOR U11264 ( .A(n10463), .B(n10464), .Z(n7586) );
  ANDN U11265 ( .B(n10465), .A(n10030), .Z(n10463) );
  XOR U11266 ( .A(n10466), .B(n7603), .Z(n2382) );
  ANDN U11267 ( .B(n10467), .A(n10468), .Z(n10466) );
  XNOR U11268 ( .A(n10469), .B(n10008), .Z(n7512) );
  NOR U11269 ( .A(n10470), .B(n10021), .Z(n10469) );
  XOR U11270 ( .A(n2346), .B(n9681), .Z(n3624) );
  XOR U11271 ( .A(n10471), .B(n10368), .Z(n9681) );
  ANDN U11272 ( .B(n10472), .A(n10473), .Z(n10471) );
  XOR U11273 ( .A(n6218), .B(n10474), .Z(n2346) );
  XOR U11274 ( .A(n10475), .B(n10476), .Z(n6218) );
  XNOR U11275 ( .A(n3199), .B(n7244), .Z(n10476) );
  XNOR U11276 ( .A(n10477), .B(n9601), .Z(n7244) );
  IV U11277 ( .A(n10373), .Z(n9601) );
  XOR U11278 ( .A(n9765), .B(n10478), .Z(n10373) );
  ANDN U11279 ( .B(n9688), .A(n9689), .Z(n10477) );
  XNOR U11280 ( .A(n10479), .B(n9431), .Z(n9688) );
  XNOR U11281 ( .A(n10480), .B(n9597), .Z(n3199) );
  IV U11282 ( .A(n10375), .Z(n9597) );
  XOR U11283 ( .A(n10481), .B(n10482), .Z(n10375) );
  NOR U11284 ( .A(n9676), .B(n9677), .Z(n10480) );
  XNOR U11285 ( .A(n9539), .B(n10483), .Z(n9676) );
  XOR U11286 ( .A(n5518), .B(n10484), .Z(n10475) );
  XOR U11287 ( .A(n8286), .B(n2379), .Z(n10484) );
  XNOR U11288 ( .A(n10485), .B(n9587), .Z(n2379) );
  XNOR U11289 ( .A(n10486), .B(n9773), .Z(n9587) );
  ANDN U11290 ( .B(n10368), .A(n10472), .Z(n10485) );
  XOR U11291 ( .A(n10487), .B(n10488), .Z(n10368) );
  XNOR U11292 ( .A(n10489), .B(n9591), .Z(n8286) );
  IV U11293 ( .A(n10371), .Z(n9591) );
  XNOR U11294 ( .A(n9617), .B(n10490), .Z(n10371) );
  NOR U11295 ( .A(n10491), .B(n9679), .Z(n10489) );
  XNOR U11296 ( .A(n10492), .B(n9251), .Z(n9679) );
  XNOR U11297 ( .A(n10493), .B(n10494), .Z(n5518) );
  ANDN U11298 ( .B(n9684), .A(n9685), .Z(n10493) );
  XOR U11299 ( .A(n10495), .B(n10496), .Z(n9684) );
  XOR U11300 ( .A(n10497), .B(n6135), .Z(out[1019]) );
  XOR U11301 ( .A(n7918), .B(n2648), .Z(n6135) );
  XNOR U11302 ( .A(n6017), .B(n7959), .Z(n2648) );
  XNOR U11303 ( .A(n10498), .B(n10499), .Z(n7959) );
  XNOR U11304 ( .A(n10500), .B(n5400), .Z(n10499) );
  XOR U11305 ( .A(n10501), .B(n8620), .Z(n5400) );
  ANDN U11306 ( .B(n7933), .A(n7934), .Z(n10501) );
  XOR U11307 ( .A(n10502), .B(n10503), .Z(n7934) );
  XOR U11308 ( .A(n6963), .B(n10504), .Z(n10498) );
  XOR U11309 ( .A(n2211), .B(n3364), .Z(n10504) );
  XNOR U11310 ( .A(n10505), .B(n8609), .Z(n3364) );
  ANDN U11311 ( .B(n7922), .A(n7920), .Z(n10505) );
  XNOR U11312 ( .A(n9802), .B(n10506), .Z(n7922) );
  XNOR U11313 ( .A(n10507), .B(n8613), .Z(n2211) );
  NOR U11314 ( .A(n10351), .B(n7925), .Z(n10507) );
  XNOR U11315 ( .A(n10508), .B(n9664), .Z(n10351) );
  XNOR U11316 ( .A(n10509), .B(n8605), .Z(n6963) );
  IV U11317 ( .A(n10510), .Z(n8605) );
  ANDN U11318 ( .B(n7929), .A(n7930), .Z(n10509) );
  XNOR U11319 ( .A(n10511), .B(n10512), .Z(n7930) );
  XOR U11320 ( .A(n10513), .B(n10514), .Z(n6017) );
  XNOR U11321 ( .A(n5240), .B(n1867), .Z(n10514) );
  XOR U11322 ( .A(n10515), .B(n10516), .Z(n1867) );
  ANDN U11323 ( .B(n9358), .A(n6984), .Z(n10515) );
  XOR U11324 ( .A(n9630), .B(n10517), .Z(n6984) );
  XNOR U11325 ( .A(n10518), .B(n10519), .Z(n5240) );
  ANDN U11326 ( .B(n9354), .A(n9355), .Z(n10518) );
  XNOR U11327 ( .A(n10520), .B(n10521), .Z(n9355) );
  XNOR U11328 ( .A(n3654), .B(n10522), .Z(n10513) );
  XOR U11329 ( .A(n8044), .B(n4146), .Z(n10522) );
  XNOR U11330 ( .A(n10523), .B(n10524), .Z(n4146) );
  NOR U11331 ( .A(n9368), .B(n9367), .Z(n10523) );
  XOR U11332 ( .A(n10525), .B(n10526), .Z(n9368) );
  XOR U11333 ( .A(n10527), .B(n10528), .Z(n8044) );
  ANDN U11334 ( .B(n6974), .A(n9361), .Z(n10527) );
  XNOR U11335 ( .A(n10529), .B(n10182), .Z(n6974) );
  XOR U11336 ( .A(n10530), .B(n10531), .Z(n3654) );
  ANDN U11337 ( .B(n6980), .A(n9364), .Z(n10530) );
  XOR U11338 ( .A(n10050), .B(n10532), .Z(n6980) );
  XOR U11339 ( .A(n10533), .B(n10534), .Z(n7918) );
  ANDN U11340 ( .B(n8615), .A(n10354), .Z(n10533) );
  XOR U11341 ( .A(n9630), .B(n10535), .Z(n8615) );
  XNOR U11342 ( .A(n10536), .B(n10537), .Z(n9630) );
  NOR U11343 ( .A(n5626), .B(n5624), .Z(n10497) );
  XNOR U11344 ( .A(n10538), .B(n1698), .Z(n5624) );
  IV U11345 ( .A(n4249), .Z(n1698) );
  XOR U11346 ( .A(n8783), .B(n6269), .Z(n4249) );
  XNOR U11347 ( .A(n10539), .B(n10540), .Z(n6269) );
  XOR U11348 ( .A(n5389), .B(n3637), .Z(n10540) );
  XNOR U11349 ( .A(n10541), .B(n10542), .Z(n3637) );
  NOR U11350 ( .A(n7881), .B(n10543), .Z(n10541) );
  IV U11351 ( .A(n10544), .Z(n7881) );
  XNOR U11352 ( .A(n10545), .B(n10546), .Z(n5389) );
  ANDN U11353 ( .B(n10547), .A(n10548), .Z(n10545) );
  XOR U11354 ( .A(n10549), .B(n10550), .Z(n10539) );
  XNOR U11355 ( .A(n2065), .B(n5312), .Z(n10550) );
  XNOR U11356 ( .A(n10551), .B(n10552), .Z(n5312) );
  ANDN U11357 ( .B(n10553), .A(n7875), .Z(n10551) );
  IV U11358 ( .A(n10554), .Z(n7875) );
  XOR U11359 ( .A(n10555), .B(n10556), .Z(n2065) );
  NOR U11360 ( .A(n8912), .B(n10557), .Z(n10555) );
  XOR U11361 ( .A(n10558), .B(n10559), .Z(n8783) );
  XOR U11362 ( .A(n5064), .B(n7783), .Z(n10559) );
  XOR U11363 ( .A(n10560), .B(n7789), .Z(n7783) );
  NOR U11364 ( .A(n7793), .B(n10421), .Z(n10561) );
  IV U11365 ( .A(n10562), .Z(n7793) );
  XOR U11366 ( .A(n2404), .B(n10563), .Z(n10558) );
  XNOR U11367 ( .A(n3456), .B(n4006), .Z(n10563) );
  XOR U11368 ( .A(n10564), .B(n7799), .Z(n4006) );
  ANDN U11369 ( .B(n7800), .A(n10412), .Z(n10564) );
  XNOR U11370 ( .A(n10565), .B(n8848), .Z(n3456) );
  NOR U11371 ( .A(n8847), .B(n10425), .Z(n10565) );
  XNOR U11372 ( .A(n10566), .B(n7803), .Z(n2404) );
  IV U11373 ( .A(n10567), .Z(n7803) );
  XOR U11374 ( .A(n9592), .B(n2031), .Z(n5626) );
  XNOR U11375 ( .A(n9372), .B(n8342), .Z(n2031) );
  XNOR U11376 ( .A(n10569), .B(n10570), .Z(n8342) );
  XOR U11377 ( .A(n5422), .B(n3869), .Z(n10570) );
  XNOR U11378 ( .A(n10571), .B(n10572), .Z(n3869) );
  ANDN U11379 ( .B(n9729), .A(n10573), .Z(n10571) );
  XNOR U11380 ( .A(n10574), .B(n9694), .Z(n5422) );
  ANDN U11381 ( .B(n9695), .A(n10575), .Z(n10574) );
  XOR U11382 ( .A(n6232), .B(n10576), .Z(n10569) );
  XNOR U11383 ( .A(n2261), .B(n4986), .Z(n10576) );
  XNOR U11384 ( .A(n10577), .B(n9698), .Z(n4986) );
  NOR U11385 ( .A(n10578), .B(n9724), .Z(n10577) );
  XNOR U11386 ( .A(n10579), .B(n9709), .Z(n2261) );
  ANDN U11387 ( .B(n9708), .A(n9733), .Z(n10579) );
  XNOR U11388 ( .A(n10580), .B(n9704), .Z(n6232) );
  ANDN U11389 ( .B(n9705), .A(n9721), .Z(n10580) );
  XOR U11390 ( .A(n10581), .B(n10582), .Z(n9372) );
  XOR U11391 ( .A(n1972), .B(n9672), .Z(n10582) );
  XNOR U11392 ( .A(n10583), .B(n10472), .Z(n9672) );
  XNOR U11393 ( .A(n9102), .B(n10584), .Z(n10472) );
  NOR U11394 ( .A(n9585), .B(n9586), .Z(n10583) );
  XNOR U11395 ( .A(n10047), .B(n10585), .Z(n9586) );
  IV U11396 ( .A(n10473), .Z(n9585) );
  XOR U11397 ( .A(n10586), .B(n10231), .Z(n10473) );
  XNOR U11398 ( .A(n10587), .B(n9677), .Z(n1972) );
  XOR U11399 ( .A(n9667), .B(n10588), .Z(n9677) );
  NOR U11400 ( .A(n9596), .B(n9595), .Z(n10587) );
  XOR U11401 ( .A(n10589), .B(n10590), .Z(n9595) );
  XOR U11402 ( .A(n10591), .B(n10402), .Z(n9596) );
  XNOR U11403 ( .A(n3764), .B(n10592), .Z(n10581) );
  XNOR U11404 ( .A(n5111), .B(n4221), .Z(n10592) );
  XNOR U11405 ( .A(n10593), .B(n9685), .Z(n4221) );
  XOR U11406 ( .A(n10594), .B(n9874), .Z(n9685) );
  ANDN U11407 ( .B(n9686), .A(n10365), .Z(n10593) );
  XNOR U11408 ( .A(n10595), .B(n10491), .Z(n5111) );
  IV U11409 ( .A(n9680), .Z(n10491) );
  XOR U11410 ( .A(n10596), .B(n9932), .Z(n9680) );
  NOR U11411 ( .A(n9590), .B(n9589), .Z(n10595) );
  XNOR U11412 ( .A(n10597), .B(n9864), .Z(n9589) );
  XOR U11413 ( .A(n10598), .B(n10599), .Z(n9590) );
  XOR U11414 ( .A(n10601), .B(n10077), .Z(n9689) );
  ANDN U11415 ( .B(n9599), .A(n9600), .Z(n10600) );
  XOR U11416 ( .A(n10602), .B(n10603), .Z(n9600) );
  XOR U11417 ( .A(n10604), .B(n10605), .Z(n9599) );
  XOR U11418 ( .A(n10606), .B(n9686), .Z(n9592) );
  ANDN U11419 ( .B(n10365), .A(n10494), .Z(n10606) );
  IV U11420 ( .A(n10366), .Z(n10494) );
  XNOR U11421 ( .A(n10608), .B(n10609), .Z(n10366) );
  XOR U11422 ( .A(n10610), .B(n9888), .Z(n10365) );
  XOR U11423 ( .A(n10611), .B(n6140), .Z(out[1018]) );
  XNOR U11424 ( .A(n10612), .B(n2655), .Z(n6140) );
  XNOR U11425 ( .A(n6022), .B(n8599), .Z(n2655) );
  XNOR U11426 ( .A(n10613), .B(n10614), .Z(n8599) );
  XOR U11427 ( .A(n5605), .B(n5404), .Z(n10614) );
  XNOR U11428 ( .A(n10615), .B(n6971), .Z(n5404) );
  XNOR U11429 ( .A(n10616), .B(n9788), .Z(n6971) );
  AND U11430 ( .A(n10524), .B(n6972), .Z(n10615) );
  XNOR U11431 ( .A(n10617), .B(n9365), .Z(n5605) );
  IV U11432 ( .A(n6982), .Z(n9365) );
  XNOR U11433 ( .A(n10618), .B(n10346), .Z(n6982) );
  NOR U11434 ( .A(n10531), .B(n6981), .Z(n10617) );
  XOR U11435 ( .A(n6965), .B(n10619), .Z(n10613) );
  XNOR U11436 ( .A(n2218), .B(n3368), .Z(n10619) );
  XNOR U11437 ( .A(n10620), .B(n6986), .Z(n3368) );
  XOR U11438 ( .A(n10621), .B(n10622), .Z(n6986) );
  NOR U11439 ( .A(n10623), .B(n10516), .Z(n10620) );
  XNOR U11440 ( .A(n10624), .B(n9362), .Z(n2218) );
  XOR U11441 ( .A(n10625), .B(n10626), .Z(n9362) );
  ANDN U11442 ( .B(n10528), .A(n10627), .Z(n10624) );
  XNOR U11443 ( .A(n10628), .B(n9356), .Z(n6965) );
  XOR U11444 ( .A(n10629), .B(n10630), .Z(n9356) );
  ANDN U11445 ( .B(n10519), .A(n10631), .Z(n10628) );
  XOR U11446 ( .A(n10632), .B(n10633), .Z(n6022) );
  XNOR U11447 ( .A(n5243), .B(n1875), .Z(n10633) );
  XOR U11448 ( .A(n10634), .B(n8101), .Z(n1875) );
  ANDN U11449 ( .B(n8102), .A(n7007), .Z(n10634) );
  XOR U11450 ( .A(n10635), .B(n9773), .Z(n7007) );
  XOR U11451 ( .A(n10636), .B(n10637), .Z(n8102) );
  XNOR U11452 ( .A(n10638), .B(n8111), .Z(n5243) );
  ANDN U11453 ( .B(n10446), .A(n10444), .Z(n10638) );
  XOR U11454 ( .A(n10639), .B(n10640), .Z(n10444) );
  XOR U11455 ( .A(n10641), .B(n9463), .Z(n10446) );
  XOR U11456 ( .A(n3659), .B(n10642), .Z(n10632) );
  XOR U11457 ( .A(n8095), .B(n4149), .Z(n10642) );
  XOR U11458 ( .A(n10643), .B(n8113), .Z(n4149) );
  ANDN U11459 ( .B(n6993), .A(n8114), .Z(n10643) );
  XOR U11460 ( .A(n9778), .B(n10644), .Z(n8114) );
  XNOR U11461 ( .A(n10645), .B(n10646), .Z(n6993) );
  XOR U11462 ( .A(n10647), .B(n8107), .Z(n8095) );
  NOR U11463 ( .A(n10450), .B(n6997), .Z(n10647) );
  XNOR U11464 ( .A(n10648), .B(n10316), .Z(n6997) );
  XNOR U11465 ( .A(n10649), .B(n9260), .Z(n10450) );
  XNOR U11466 ( .A(n10650), .B(n10651), .Z(n3659) );
  ANDN U11467 ( .B(n7003), .A(n10452), .Z(n10650) );
  XOR U11468 ( .A(n10652), .B(n9879), .Z(n7003) );
  ANDN U11469 ( .B(n5630), .A(n5628), .Z(n10611) );
  XOR U11470 ( .A(n10653), .B(n1703), .Z(n5628) );
  XNOR U11471 ( .A(n8843), .B(n6273), .Z(n1703) );
  XNOR U11472 ( .A(n10654), .B(n10655), .Z(n6273) );
  XOR U11473 ( .A(n5394), .B(n3643), .Z(n10655) );
  XOR U11474 ( .A(n10656), .B(n10657), .Z(n3643) );
  ANDN U11475 ( .B(n10658), .A(n10659), .Z(n10656) );
  XNOR U11476 ( .A(n10660), .B(n10661), .Z(n5394) );
  ANDN U11477 ( .B(n10662), .A(n7941), .Z(n10660) );
  XNOR U11478 ( .A(n10663), .B(n10664), .Z(n10654) );
  XOR U11479 ( .A(n2068), .B(n5363), .Z(n10664) );
  XNOR U11480 ( .A(n10665), .B(n10666), .Z(n5363) );
  ANDN U11481 ( .B(n10667), .A(n7945), .Z(n10665) );
  XNOR U11482 ( .A(n10668), .B(n10669), .Z(n2068) );
  ANDN U11483 ( .B(n10670), .A(n8975), .Z(n10668) );
  XOR U11484 ( .A(n10671), .B(n10672), .Z(n8843) );
  XOR U11485 ( .A(n3463), .B(n5067), .Z(n10672) );
  XOR U11486 ( .A(n10673), .B(n7876), .Z(n5067) );
  ANDN U11487 ( .B(n10552), .A(n7877), .Z(n10673) );
  XOR U11488 ( .A(n10674), .B(n8913), .Z(n3463) );
  XOR U11489 ( .A(n4009), .B(n10675), .Z(n10671) );
  XOR U11490 ( .A(n7866), .B(n2414), .Z(n10675) );
  XNOR U11491 ( .A(n10676), .B(n7887), .Z(n2414) );
  ANDN U11492 ( .B(n10677), .A(n10678), .Z(n10676) );
  XNOR U11493 ( .A(n10679), .B(n7873), .Z(n7866) );
  ANDN U11494 ( .B(n7872), .A(n10680), .Z(n10679) );
  XOR U11495 ( .A(n10681), .B(n7882), .Z(n4009) );
  XOR U11496 ( .A(n9700), .B(n2034), .Z(n5630) );
  XNOR U11497 ( .A(n10474), .B(n8647), .Z(n2034) );
  XNOR U11498 ( .A(n10682), .B(n10683), .Z(n8647) );
  XOR U11499 ( .A(n5426), .B(n3876), .Z(n10683) );
  XOR U11500 ( .A(n10684), .B(n10685), .Z(n3876) );
  AND U11501 ( .A(n7345), .B(n7347), .Z(n10684) );
  XOR U11502 ( .A(n10686), .B(n10687), .Z(n7347) );
  XNOR U11503 ( .A(n10688), .B(n9739), .Z(n5426) );
  ANDN U11504 ( .B(n7343), .A(n7341), .Z(n10688) );
  XOR U11505 ( .A(n10689), .B(n9939), .Z(n7341) );
  XOR U11506 ( .A(n10690), .B(n10691), .Z(n7343) );
  XNOR U11507 ( .A(n6237), .B(n10692), .Z(n10682) );
  XOR U11508 ( .A(n2268), .B(n5022), .Z(n10692) );
  XNOR U11509 ( .A(n10693), .B(n9742), .Z(n5022) );
  ANDN U11510 ( .B(n8397), .A(n8395), .Z(n10693) );
  XOR U11511 ( .A(n10694), .B(n10695), .Z(n8395) );
  XNOR U11512 ( .A(n9414), .B(n10696), .Z(n8397) );
  XNOR U11513 ( .A(n10697), .B(n9750), .Z(n2268) );
  AND U11514 ( .A(n8649), .B(n8650), .Z(n10697) );
  XOR U11515 ( .A(n10698), .B(n10699), .Z(n8650) );
  XOR U11516 ( .A(n9122), .B(n10700), .Z(n8649) );
  XNOR U11517 ( .A(n10701), .B(n9747), .Z(n6237) );
  AND U11518 ( .A(n7336), .B(n7335), .Z(n10701) );
  XOR U11519 ( .A(n10702), .B(n10703), .Z(n7335) );
  XOR U11520 ( .A(n10704), .B(n9790), .Z(n7336) );
  XOR U11521 ( .A(n10705), .B(n10706), .Z(n10474) );
  XNOR U11522 ( .A(n1661), .B(n9717), .Z(n10706) );
  XNOR U11523 ( .A(n10707), .B(n10708), .Z(n9717) );
  NOR U11524 ( .A(n9693), .B(n9694), .Z(n10707) );
  XNOR U11525 ( .A(n9242), .B(n10709), .Z(n9694) );
  IV U11526 ( .A(n10710), .Z(n9693) );
  XNOR U11527 ( .A(n10711), .B(n9722), .Z(n1661) );
  ANDN U11528 ( .B(n9703), .A(n9704), .Z(n10711) );
  XOR U11529 ( .A(n10604), .B(n10712), .Z(n9704) );
  XOR U11530 ( .A(n10713), .B(n10714), .Z(n9703) );
  XNOR U11531 ( .A(n3768), .B(n10715), .Z(n10705) );
  XOR U11532 ( .A(n5113), .B(n4226), .Z(n10715) );
  XNOR U11533 ( .A(n10716), .B(n10717), .Z(n4226) );
  ANDN U11534 ( .B(n9731), .A(n10572), .Z(n10716) );
  XNOR U11535 ( .A(n10718), .B(n10719), .Z(n5113) );
  NOR U11536 ( .A(n9698), .B(n9697), .Z(n10718) );
  XOR U11537 ( .A(n9522), .B(n10720), .Z(n9697) );
  IV U11538 ( .A(n9122), .Z(n9522) );
  XNOR U11539 ( .A(n10721), .B(n10722), .Z(n9122) );
  XOR U11540 ( .A(n10723), .B(n10724), .Z(n9698) );
  XNOR U11541 ( .A(n10725), .B(n9734), .Z(n3768) );
  AND U11542 ( .A(n9709), .B(n9707), .Z(n10725) );
  XNOR U11543 ( .A(n10726), .B(n10727), .Z(n9707) );
  XOR U11544 ( .A(n10728), .B(n10729), .Z(n9709) );
  XOR U11545 ( .A(n10730), .B(n9731), .Z(n9700) );
  XNOR U11546 ( .A(n10602), .B(n10731), .Z(n9731) );
  XNOR U11547 ( .A(n10732), .B(n9954), .Z(n10572) );
  XOR U11548 ( .A(n10733), .B(n6145), .Z(out[1017]) );
  XOR U11549 ( .A(n8099), .B(n2662), .Z(n6145) );
  XNOR U11550 ( .A(n6027), .B(n9350), .Z(n2662) );
  XNOR U11551 ( .A(n10734), .B(n10735), .Z(n9350) );
  XNOR U11552 ( .A(n5650), .B(n5407), .Z(n10735) );
  XOR U11553 ( .A(n10736), .B(n6994), .Z(n5407) );
  XNOR U11554 ( .A(n10737), .B(n9886), .Z(n6994) );
  ANDN U11555 ( .B(n6995), .A(n8113), .Z(n10736) );
  XOR U11556 ( .A(n10738), .B(n10739), .Z(n8113) );
  XOR U11557 ( .A(n10740), .B(n10741), .Z(n6995) );
  XNOR U11558 ( .A(n10742), .B(n7005), .Z(n5650) );
  XOR U11559 ( .A(n10743), .B(n10744), .Z(n7005) );
  ANDN U11560 ( .B(n10651), .A(n7004), .Z(n10742) );
  XOR U11561 ( .A(n6988), .B(n10745), .Z(n10734) );
  XOR U11562 ( .A(n2223), .B(n3372), .Z(n10745) );
  XNOR U11563 ( .A(n10746), .B(n7009), .Z(n3372) );
  XOR U11564 ( .A(n10747), .B(n9771), .Z(n7009) );
  NOR U11565 ( .A(n7008), .B(n8101), .Z(n10746) );
  XNOR U11566 ( .A(n10748), .B(n10749), .Z(n8101) );
  XNOR U11567 ( .A(n10750), .B(n10221), .Z(n7008) );
  XOR U11568 ( .A(n10751), .B(n6999), .Z(n2223) );
  XOR U11569 ( .A(n10752), .B(n10753), .Z(n6999) );
  ANDN U11570 ( .B(n8107), .A(n8105), .Z(n10751) );
  IV U11571 ( .A(n6998), .Z(n8105) );
  XOR U11572 ( .A(n10754), .B(n10755), .Z(n6998) );
  XOR U11573 ( .A(n10756), .B(n10205), .Z(n8107) );
  XNOR U11574 ( .A(n10757), .B(n10445), .Z(n6988) );
  XOR U11575 ( .A(n10758), .B(n10759), .Z(n10445) );
  ANDN U11576 ( .B(n8111), .A(n8109), .Z(n10757) );
  XOR U11577 ( .A(n10760), .B(n10761), .Z(n8109) );
  XOR U11578 ( .A(n10762), .B(n10763), .Z(n8111) );
  XOR U11579 ( .A(n10764), .B(n10765), .Z(n6027) );
  XNOR U11580 ( .A(n5246), .B(n1879), .Z(n10765) );
  XOR U11581 ( .A(n10766), .B(n8128), .Z(n1879) );
  ANDN U11582 ( .B(n7030), .A(n8129), .Z(n10766) );
  XOR U11583 ( .A(n10767), .B(n8136), .Z(n5246) );
  NOR U11584 ( .A(n10768), .B(n8137), .Z(n10767) );
  XNOR U11585 ( .A(n3663), .B(n10769), .Z(n10764) );
  XNOR U11586 ( .A(n8122), .B(n4152), .Z(n10769) );
  XOR U11587 ( .A(n10770), .B(n8140), .Z(n4152) );
  ANDN U11588 ( .B(n8141), .A(n10771), .Z(n10770) );
  XNOR U11589 ( .A(n10772), .B(n8132), .Z(n8122) );
  IV U11590 ( .A(n10773), .Z(n8132) );
  ANDN U11591 ( .B(n8133), .A(n7020), .Z(n10772) );
  XNOR U11592 ( .A(n10774), .B(n10775), .Z(n3663) );
  AND U11593 ( .A(n7026), .B(n10776), .Z(n10774) );
  XOR U11594 ( .A(n10777), .B(n7004), .Z(n8099) );
  XOR U11595 ( .A(n10778), .B(n10307), .Z(n7004) );
  ANDN U11596 ( .B(n10452), .A(n10651), .Z(n10777) );
  XOR U11597 ( .A(n10779), .B(n10780), .Z(n10651) );
  XOR U11598 ( .A(n10781), .B(n9874), .Z(n10452) );
  ANDN U11599 ( .B(n5634), .A(n5632), .Z(n10733) );
  XOR U11600 ( .A(n10782), .B(n1708), .Z(n5632) );
  XNOR U11601 ( .A(n8909), .B(n6281), .Z(n1708) );
  XNOR U11602 ( .A(n10783), .B(n10784), .Z(n6281) );
  XNOR U11603 ( .A(n5398), .B(n3647), .Z(n10784) );
  XNOR U11604 ( .A(n10785), .B(n10786), .Z(n3647) );
  NOR U11605 ( .A(n10787), .B(n8037), .Z(n10785) );
  XNOR U11606 ( .A(n10788), .B(n10789), .Z(n5398) );
  ANDN U11607 ( .B(n10790), .A(n8027), .Z(n10788) );
  IV U11608 ( .A(n10791), .Z(n8027) );
  XNOR U11609 ( .A(n10792), .B(n10793), .Z(n10783) );
  XNOR U11610 ( .A(n2071), .B(n5410), .Z(n10793) );
  XNOR U11611 ( .A(n10794), .B(n10795), .Z(n5410) );
  NOR U11612 ( .A(n10796), .B(n8031), .Z(n10794) );
  XOR U11613 ( .A(n10797), .B(n10798), .Z(n2071) );
  ANDN U11614 ( .B(n10799), .A(n9037), .Z(n10797) );
  IV U11615 ( .A(n10800), .Z(n9037) );
  XOR U11616 ( .A(n10801), .B(n10802), .Z(n8909) );
  XNOR U11617 ( .A(n3466), .B(n5071), .Z(n10802) );
  XOR U11618 ( .A(n10803), .B(n7946), .Z(n5071) );
  ANDN U11619 ( .B(n7947), .A(n10666), .Z(n10803) );
  XOR U11620 ( .A(n10804), .B(n8976), .Z(n3466) );
  AND U11621 ( .A(n8977), .B(n10669), .Z(n10804) );
  XOR U11622 ( .A(n4024), .B(n10805), .Z(n10801) );
  XOR U11623 ( .A(n7936), .B(n2419), .Z(n10805) );
  XOR U11624 ( .A(n10806), .B(n7956), .Z(n2419) );
  ANDN U11625 ( .B(n10807), .A(n7957), .Z(n10806) );
  XOR U11626 ( .A(n10808), .B(n7942), .Z(n7936) );
  XNOR U11627 ( .A(n10809), .B(n7953), .Z(n4024) );
  NOR U11628 ( .A(n7952), .B(n10657), .Z(n10809) );
  XNOR U11629 ( .A(n9743), .B(n2041), .Z(n5634) );
  XNOR U11630 ( .A(n10810), .B(n9397), .Z(n2041) );
  XNOR U11631 ( .A(n10811), .B(n10812), .Z(n9397) );
  XNOR U11632 ( .A(n5430), .B(n3880), .Z(n10812) );
  XNOR U11633 ( .A(n10813), .B(n10814), .Z(n3880) );
  ANDN U11634 ( .B(n7420), .A(n7418), .Z(n10813) );
  IV U11635 ( .A(n10815), .Z(n7418) );
  XNOR U11636 ( .A(n10816), .B(n10817), .Z(n7420) );
  XNOR U11637 ( .A(n10818), .B(n9839), .Z(n5430) );
  ANDN U11638 ( .B(n7416), .A(n7414), .Z(n10818) );
  XOR U11639 ( .A(n10819), .B(n10820), .Z(n7414) );
  XNOR U11640 ( .A(n10821), .B(n9424), .Z(n7416) );
  IV U11641 ( .A(n10822), .Z(n9424) );
  XOR U11642 ( .A(n6242), .B(n10823), .Z(n10811) );
  XNOR U11643 ( .A(n2275), .B(n5058), .Z(n10823) );
  XOR U11644 ( .A(n10824), .B(n9842), .Z(n5058) );
  ANDN U11645 ( .B(n8451), .A(n8452), .Z(n10824) );
  XNOR U11646 ( .A(n10825), .B(n9511), .Z(n8452) );
  XNOR U11647 ( .A(n10116), .B(n10826), .Z(n8451) );
  XNOR U11648 ( .A(n10827), .B(n9851), .Z(n2275) );
  AND U11649 ( .A(n9401), .B(n9399), .Z(n10827) );
  XOR U11650 ( .A(n9637), .B(n10828), .Z(n9399) );
  XOR U11651 ( .A(n9780), .B(n10829), .Z(n9401) );
  XNOR U11652 ( .A(n10830), .B(n9847), .Z(n6242) );
  NOR U11653 ( .A(n9848), .B(n7409), .Z(n10830) );
  XOR U11654 ( .A(n10831), .B(n9888), .Z(n7409) );
  XOR U11655 ( .A(n10832), .B(n10833), .Z(n9848) );
  XNOR U11656 ( .A(n10834), .B(n9834), .Z(n9743) );
  ANDN U11657 ( .B(n10685), .A(n7345), .Z(n10834) );
  XOR U11658 ( .A(n10835), .B(n10836), .Z(n7345) );
  XNOR U11659 ( .A(n10837), .B(n6150), .Z(out[1016]) );
  IV U11660 ( .A(n6632), .Z(n6150) );
  XNOR U11661 ( .A(n8125), .B(n2669), .Z(n6632) );
  XNOR U11662 ( .A(n6032), .B(n10440), .Z(n2669) );
  XNOR U11663 ( .A(n10838), .B(n10839), .Z(n10440) );
  XOR U11664 ( .A(n5693), .B(n5417), .Z(n10839) );
  XNOR U11665 ( .A(n10840), .B(n7017), .Z(n5417) );
  NOR U11666 ( .A(n8139), .B(n8140), .Z(n10840) );
  XOR U11667 ( .A(n10841), .B(n10842), .Z(n8140) );
  IV U11668 ( .A(n7018), .Z(n8139) );
  XOR U11669 ( .A(n9119), .B(n10843), .Z(n7018) );
  XNOR U11670 ( .A(n10844), .B(n10845), .Z(n5693) );
  ANDN U11671 ( .B(n10775), .A(n7027), .Z(n10844) );
  XOR U11672 ( .A(n7011), .B(n10846), .Z(n10838) );
  XOR U11673 ( .A(n2232), .B(n3376), .Z(n10846) );
  XNOR U11674 ( .A(n10847), .B(n7031), .Z(n3376) );
  NOR U11675 ( .A(n8127), .B(n8128), .Z(n10847) );
  XNOR U11676 ( .A(n9506), .B(n10848), .Z(n8128) );
  XNOR U11677 ( .A(n10849), .B(n10850), .Z(n8127) );
  XNOR U11678 ( .A(n10851), .B(n10852), .Z(n2232) );
  ANDN U11679 ( .B(n7022), .A(n10773), .Z(n10851) );
  XOR U11680 ( .A(n10853), .B(n10338), .Z(n10773) );
  XNOR U11681 ( .A(n10854), .B(n10855), .Z(n7022) );
  XNOR U11682 ( .A(n10856), .B(n10857), .Z(n7011) );
  NOR U11683 ( .A(n10858), .B(n8136), .Z(n10856) );
  XNOR U11684 ( .A(n10859), .B(n10860), .Z(n8136) );
  XOR U11685 ( .A(n10861), .B(n10862), .Z(n6032) );
  XNOR U11686 ( .A(n5253), .B(n1883), .Z(n10862) );
  XNOR U11687 ( .A(n10863), .B(n8209), .Z(n1883) );
  ANDN U11688 ( .B(n8147), .A(n7056), .Z(n10863) );
  XOR U11689 ( .A(n10864), .B(n9939), .Z(n7056) );
  XNOR U11690 ( .A(n10380), .B(n10865), .Z(n8147) );
  XNOR U11691 ( .A(n10866), .B(n8214), .Z(n5253) );
  ANDN U11692 ( .B(n7052), .A(n8215), .Z(n10866) );
  XOR U11693 ( .A(n10867), .B(n10868), .Z(n8215) );
  XNOR U11694 ( .A(n10869), .B(n10870), .Z(n7052) );
  XNOR U11695 ( .A(n3667), .B(n10871), .Z(n10861) );
  XOR U11696 ( .A(n8203), .B(n4155), .Z(n10871) );
  XOR U11697 ( .A(n10872), .B(n8217), .Z(n4155) );
  AND U11698 ( .A(n8154), .B(n7039), .Z(n10872) );
  XOR U11699 ( .A(n10873), .B(n10874), .Z(n7039) );
  XOR U11700 ( .A(n10875), .B(n9946), .Z(n8154) );
  XOR U11701 ( .A(n10876), .B(n8212), .Z(n8203) );
  XNOR U11702 ( .A(n10177), .B(n10877), .Z(n8150) );
  IV U11703 ( .A(n9438), .Z(n10177) );
  XOR U11704 ( .A(n10878), .B(n10879), .Z(n7043) );
  XOR U11705 ( .A(n10880), .B(n10881), .Z(n3667) );
  ANDN U11706 ( .B(n8152), .A(n7048), .Z(n10880) );
  XNOR U11707 ( .A(n10882), .B(n10488), .Z(n7048) );
  XOR U11708 ( .A(n10883), .B(n7027), .Z(n8125) );
  XOR U11709 ( .A(n10884), .B(n10406), .Z(n7027) );
  NOR U11710 ( .A(n10775), .B(n10776), .Z(n10883) );
  XOR U11711 ( .A(n10885), .B(n10886), .Z(n10775) );
  NOR U11712 ( .A(n5637), .B(n5636), .Z(n10837) );
  XOR U11713 ( .A(n10887), .B(n3818), .Z(n5636) );
  IV U11714 ( .A(n1713), .Z(n3818) );
  XOR U11715 ( .A(n8972), .B(n6285), .Z(n1713) );
  XNOR U11716 ( .A(n10888), .B(n10889), .Z(n6285) );
  XOR U11717 ( .A(n5402), .B(n3651), .Z(n10889) );
  XOR U11718 ( .A(n10890), .B(n10891), .Z(n3651) );
  ANDN U11719 ( .B(n10892), .A(n8088), .Z(n10890) );
  IV U11720 ( .A(n10893), .Z(n8088) );
  XNOR U11721 ( .A(n10894), .B(n10895), .Z(n5402) );
  NOR U11722 ( .A(n10896), .B(n8078), .Z(n10894) );
  XOR U11723 ( .A(n10897), .B(n10898), .Z(n10888) );
  XNOR U11724 ( .A(n2078), .B(n5459), .Z(n10898) );
  XNOR U11725 ( .A(n10899), .B(n10900), .Z(n5459) );
  ANDN U11726 ( .B(n10901), .A(n10902), .Z(n10899) );
  XNOR U11727 ( .A(n10903), .B(n10904), .Z(n2078) );
  ANDN U11728 ( .B(n10905), .A(n10906), .Z(n10903) );
  XOR U11729 ( .A(n10907), .B(n10908), .Z(n8972) );
  XNOR U11730 ( .A(n3470), .B(n5075), .Z(n10908) );
  XOR U11731 ( .A(n10909), .B(n8033), .Z(n5075) );
  ANDN U11732 ( .B(n8032), .A(n10795), .Z(n10909) );
  XNOR U11733 ( .A(n10910), .B(n9039), .Z(n3470) );
  XNOR U11734 ( .A(n4058), .B(n10911), .Z(n10907) );
  XOR U11735 ( .A(n8022), .B(n2428), .Z(n10911) );
  XOR U11736 ( .A(n10912), .B(n8042), .Z(n2428) );
  NOR U11737 ( .A(n10913), .B(n8043), .Z(n10912) );
  XOR U11738 ( .A(n10914), .B(n8028), .Z(n8022) );
  NOR U11739 ( .A(n10915), .B(n10789), .Z(n10914) );
  XOR U11740 ( .A(n10916), .B(n8038), .Z(n4058) );
  NOR U11741 ( .A(n10917), .B(n8039), .Z(n10916) );
  XOR U11742 ( .A(n9843), .B(n2045), .Z(n5637) );
  XNOR U11743 ( .A(n7330), .B(n10455), .Z(n2045) );
  XNOR U11744 ( .A(n10918), .B(n10919), .Z(n10455) );
  XNOR U11745 ( .A(n5436), .B(n3885), .Z(n10919) );
  XNOR U11746 ( .A(n10920), .B(n10921), .Z(n3885) );
  AND U11747 ( .A(n7525), .B(n7524), .Z(n10920) );
  XOR U11748 ( .A(n10922), .B(n9870), .Z(n7525) );
  XNOR U11749 ( .A(n10923), .B(n9995), .Z(n5436) );
  ANDN U11750 ( .B(n7520), .A(n7521), .Z(n10923) );
  XNOR U11751 ( .A(n10924), .B(n9535), .Z(n7521) );
  XOR U11752 ( .A(n10925), .B(n10088), .Z(n7520) );
  XNOR U11753 ( .A(n6246), .B(n10926), .Z(n10918) );
  XOR U11754 ( .A(n2282), .B(n5095), .Z(n10926) );
  XNOR U11755 ( .A(n10927), .B(n9998), .Z(n5095) );
  ANDN U11756 ( .B(n8528), .A(n9999), .Z(n10927) );
  XOR U11757 ( .A(n10928), .B(n10929), .Z(n9999) );
  XOR U11758 ( .A(n9614), .B(n10930), .Z(n8528) );
  XNOR U11759 ( .A(n10931), .B(n10932), .Z(n2282) );
  ANDN U11760 ( .B(n10008), .A(n10020), .Z(n10931) );
  IV U11761 ( .A(n10470), .Z(n10020) );
  XOR U11762 ( .A(n9114), .B(n10933), .Z(n10470) );
  IV U11763 ( .A(n10934), .Z(n9114) );
  XOR U11764 ( .A(n10935), .B(n9783), .Z(n10008) );
  XOR U11765 ( .A(n10936), .B(n10004), .Z(n6246) );
  ANDN U11766 ( .B(n7514), .A(n7515), .Z(n10936) );
  XNOR U11767 ( .A(n10937), .B(n9954), .Z(n7515) );
  XOR U11768 ( .A(n10938), .B(n9420), .Z(n7514) );
  XOR U11769 ( .A(n10939), .B(n10940), .Z(n7330) );
  XOR U11770 ( .A(n1674), .B(n9980), .Z(n10940) );
  XNOR U11771 ( .A(n10941), .B(n7415), .Z(n9980) );
  XOR U11772 ( .A(n9439), .B(n10942), .Z(n7415) );
  ANDN U11773 ( .B(n9839), .A(n9838), .Z(n10941) );
  XNOR U11774 ( .A(n10943), .B(n10172), .Z(n9838) );
  XNOR U11775 ( .A(n10944), .B(n10945), .Z(n9839) );
  XNOR U11776 ( .A(n10946), .B(n7410), .Z(n1674) );
  XNOR U11777 ( .A(n10947), .B(n10948), .Z(n7410) );
  AND U11778 ( .A(n9846), .B(n9847), .Z(n10946) );
  XNOR U11779 ( .A(n10949), .B(n10950), .Z(n9847) );
  XOR U11780 ( .A(n10885), .B(n10951), .Z(n9846) );
  XOR U11781 ( .A(n3778), .B(n10952), .Z(n10939) );
  XOR U11782 ( .A(n5117), .B(n4233), .Z(n10952) );
  XNOR U11783 ( .A(n10953), .B(n7419), .Z(n4233) );
  IV U11784 ( .A(n9989), .Z(n7419) );
  XOR U11785 ( .A(n10954), .B(n10088), .Z(n9989) );
  ANDN U11786 ( .B(n9990), .A(n10814), .Z(n10953) );
  XOR U11787 ( .A(n10955), .B(n8453), .Z(n5117) );
  XOR U11788 ( .A(n10186), .B(n10956), .Z(n8453) );
  XOR U11789 ( .A(n10957), .B(n10958), .Z(n9842) );
  XOR U11790 ( .A(n10959), .B(n9783), .Z(n9841) );
  XNOR U11791 ( .A(n10961), .B(n10962), .Z(n9400) );
  AND U11792 ( .A(n9851), .B(n9850), .Z(n10960) );
  XOR U11793 ( .A(n10963), .B(n10964), .Z(n9850) );
  XNOR U11794 ( .A(n10965), .B(n10966), .Z(n9851) );
  XOR U11795 ( .A(n10967), .B(n9990), .Z(n9843) );
  XOR U11796 ( .A(n10968), .B(n10969), .Z(n9990) );
  ANDN U11797 ( .B(n10814), .A(n10815), .Z(n10967) );
  XOR U11798 ( .A(n10970), .B(n10971), .Z(n10815) );
  XOR U11799 ( .A(n10972), .B(n10103), .Z(n10814) );
  XOR U11800 ( .A(n10973), .B(n6155), .Z(out[1015]) );
  XNOR U11801 ( .A(n8206), .B(n2676), .Z(n6155) );
  XNOR U11802 ( .A(n6037), .B(n10974), .Z(n2676) );
  XOR U11803 ( .A(n10975), .B(n10976), .Z(n6037) );
  XNOR U11804 ( .A(n5256), .B(n1887), .Z(n10976) );
  XNOR U11805 ( .A(n10977), .B(n8276), .Z(n1887) );
  AND U11806 ( .A(n8223), .B(n7117), .Z(n10977) );
  XNOR U11807 ( .A(n10978), .B(n10979), .Z(n7117) );
  XOR U11808 ( .A(n10980), .B(n10981), .Z(n8223) );
  XNOR U11809 ( .A(n10982), .B(n8281), .Z(n5256) );
  NOR U11810 ( .A(n8282), .B(n7113), .Z(n10982) );
  XNOR U11811 ( .A(n10983), .B(n9813), .Z(n7113) );
  XOR U11812 ( .A(n10984), .B(n10985), .Z(n8282) );
  XNOR U11813 ( .A(n3676), .B(n10986), .Z(n10975) );
  XNOR U11814 ( .A(n8257), .B(n4159), .Z(n10986) );
  XNOR U11815 ( .A(n10987), .B(n8284), .Z(n4159) );
  NOR U11816 ( .A(n7100), .B(n8230), .Z(n10987) );
  XNOR U11817 ( .A(n10988), .B(n9147), .Z(n8230) );
  XOR U11818 ( .A(n10989), .B(n10990), .Z(n7100) );
  XNOR U11819 ( .A(n10991), .B(n10992), .Z(n8257) );
  NOR U11820 ( .A(n7104), .B(n8226), .Z(n10991) );
  XOR U11821 ( .A(n9541), .B(n10993), .Z(n8226) );
  IV U11822 ( .A(n10313), .Z(n9541) );
  XOR U11823 ( .A(n10994), .B(n10741), .Z(n7104) );
  XNOR U11824 ( .A(n10995), .B(n10996), .Z(n3676) );
  NOR U11825 ( .A(n10997), .B(n7109), .Z(n10995) );
  XOR U11826 ( .A(n10998), .B(n9246), .Z(n7109) );
  IV U11827 ( .A(n10094), .Z(n9246) );
  XNOR U11828 ( .A(n10999), .B(n7049), .Z(n8206) );
  XOR U11829 ( .A(n10978), .B(n11000), .Z(n8152) );
  ANDN U11830 ( .B(n5642), .A(n5640), .Z(n10973) );
  XOR U11831 ( .A(n11001), .B(n1718), .Z(n5640) );
  XNOR U11832 ( .A(n9035), .B(n6289), .Z(n1718) );
  XNOR U11833 ( .A(n11002), .B(n11003), .Z(n6289) );
  XOR U11834 ( .A(n5406), .B(n3655), .Z(n11003) );
  XOR U11835 ( .A(n11004), .B(n11005), .Z(n3655) );
  ANDN U11836 ( .B(n11006), .A(n11007), .Z(n11004) );
  XNOR U11837 ( .A(n11008), .B(n11009), .Z(n5406) );
  ANDN U11838 ( .B(n11010), .A(n8160), .Z(n11008) );
  XNOR U11839 ( .A(n11011), .B(n11012), .Z(n11002) );
  XNOR U11840 ( .A(n2081), .B(n5512), .Z(n11012) );
  XNOR U11841 ( .A(n11013), .B(n11014), .Z(n5512) );
  ANDN U11842 ( .B(n11015), .A(n11016), .Z(n11013) );
  XOR U11843 ( .A(n11017), .B(n11018), .Z(n2081) );
  ANDN U11844 ( .B(n11019), .A(n9186), .Z(n11017) );
  IV U11845 ( .A(n11020), .Z(n9186) );
  XOR U11846 ( .A(n11021), .B(n11022), .Z(n9035) );
  XOR U11847 ( .A(n3472), .B(n5078), .Z(n11022) );
  XNOR U11848 ( .A(n11023), .B(n8084), .Z(n5078) );
  NOR U11849 ( .A(n11024), .B(n10900), .Z(n11023) );
  XNOR U11850 ( .A(n11025), .B(n9095), .Z(n3472) );
  NOR U11851 ( .A(n9094), .B(n10904), .Z(n11025) );
  XOR U11852 ( .A(n4092), .B(n11026), .Z(n11021) );
  XOR U11853 ( .A(n8073), .B(n2435), .Z(n11026) );
  XOR U11854 ( .A(n11027), .B(n8093), .Z(n2435) );
  ANDN U11855 ( .B(n8094), .A(n11028), .Z(n11027) );
  XNOR U11856 ( .A(n11029), .B(n8079), .Z(n8073) );
  IV U11857 ( .A(n11030), .Z(n8079) );
  ANDN U11858 ( .B(n8080), .A(n10895), .Z(n11029) );
  XNOR U11859 ( .A(n11031), .B(n8089), .Z(n4092) );
  ANDN U11860 ( .B(n8090), .A(n10891), .Z(n11031) );
  XOR U11861 ( .A(n10000), .B(n2049), .Z(n5642) );
  XNOR U11862 ( .A(n7403), .B(n11032), .Z(n2049) );
  XOR U11863 ( .A(n11033), .B(n11034), .Z(n7403) );
  XOR U11864 ( .A(n3783), .B(n5119), .Z(n11034) );
  XNOR U11865 ( .A(n11035), .B(n8529), .Z(n5119) );
  XNOR U11866 ( .A(n11036), .B(n10324), .Z(n8529) );
  XOR U11867 ( .A(n9458), .B(n11037), .Z(n9997) );
  XOR U11868 ( .A(n11038), .B(n11039), .Z(n9998) );
  XOR U11869 ( .A(n11040), .B(n10021), .Z(n3783) );
  XNOR U11870 ( .A(n10878), .B(n11041), .Z(n10021) );
  ANDN U11871 ( .B(n10006), .A(n10932), .Z(n11040) );
  IV U11872 ( .A(n10007), .Z(n10932) );
  XNOR U11873 ( .A(n11042), .B(n11043), .Z(n10007) );
  XNOR U11874 ( .A(n11044), .B(n11045), .Z(n10006) );
  XNOR U11875 ( .A(n4236), .B(n11046), .Z(n11033) );
  XOR U11876 ( .A(n1679), .B(n10012), .Z(n11046) );
  XNOR U11877 ( .A(n11047), .B(n7522), .Z(n10012) );
  XNOR U11878 ( .A(n9539), .B(n11048), .Z(n7522) );
  ANDN U11879 ( .B(n9995), .A(n9994), .Z(n11047) );
  XOR U11880 ( .A(n11049), .B(n10307), .Z(n9994) );
  XNOR U11881 ( .A(n11051), .B(n7516), .Z(n1679) );
  XNOR U11882 ( .A(n10282), .B(n11052), .Z(n7516) );
  XOR U11883 ( .A(n11053), .B(n10964), .Z(n10004) );
  XOR U11884 ( .A(n11054), .B(n11055), .Z(n10003) );
  XNOR U11885 ( .A(n11056), .B(n7526), .Z(n4236) );
  XOR U11886 ( .A(n11057), .B(n10195), .Z(n7526) );
  ANDN U11887 ( .B(n10023), .A(n10921), .Z(n11056) );
  IV U11888 ( .A(n11058), .Z(n10921) );
  XOR U11889 ( .A(n11059), .B(n10023), .Z(n10000) );
  XOR U11890 ( .A(n10965), .B(n11060), .Z(n10023) );
  NOR U11891 ( .A(n11058), .B(n7524), .Z(n11059) );
  XOR U11892 ( .A(n11061), .B(n11062), .Z(n7524) );
  XOR U11893 ( .A(n10214), .B(n11063), .Z(n11058) );
  XOR U11894 ( .A(n11064), .B(n6160), .Z(out[1014]) );
  XOR U11895 ( .A(n8274), .B(n2209), .Z(n6160) );
  IV U11896 ( .A(n4968), .Z(n2209) );
  XOR U11897 ( .A(n6123), .B(n6043), .Z(n4968) );
  XOR U11898 ( .A(n11065), .B(n11066), .Z(n6043) );
  XNOR U11899 ( .A(n3680), .B(n4164), .Z(n11066) );
  XNOR U11900 ( .A(n11067), .B(n8338), .Z(n4164) );
  ANDN U11901 ( .B(n8271), .A(n7157), .Z(n11067) );
  XOR U11902 ( .A(n11068), .B(n11069), .Z(n7157) );
  XOR U11903 ( .A(n11070), .B(n10094), .Z(n8271) );
  XNOR U11904 ( .A(n11071), .B(n11072), .Z(n3680) );
  ANDN U11905 ( .B(n7166), .A(n8269), .Z(n11071) );
  XOR U11906 ( .A(n10690), .B(n11073), .Z(n7166) );
  XOR U11907 ( .A(n5259), .B(n11074), .Z(n11065) );
  XNOR U11908 ( .A(n8311), .B(n1892), .Z(n11074) );
  XNOR U11909 ( .A(n11075), .B(n8330), .Z(n1892) );
  ANDN U11910 ( .B(n8264), .A(n8263), .Z(n11075) );
  IV U11911 ( .A(n8329), .Z(n8263) );
  XOR U11912 ( .A(n10151), .B(n11076), .Z(n8329) );
  IV U11913 ( .A(n9242), .Z(n10151) );
  IV U11914 ( .A(n7174), .Z(n8264) );
  XOR U11915 ( .A(n11077), .B(n11078), .Z(n7174) );
  XOR U11916 ( .A(n11079), .B(n8333), .Z(n8311) );
  ANDN U11917 ( .B(n7161), .A(n8267), .Z(n11079) );
  XNOR U11918 ( .A(n11080), .B(n9647), .Z(n8267) );
  IV U11919 ( .A(n11081), .Z(n9647) );
  XNOR U11920 ( .A(n9119), .B(n11082), .Z(n7161) );
  XNOR U11921 ( .A(n11083), .B(n8335), .Z(n5259) );
  ANDN U11922 ( .B(n7170), .A(n8336), .Z(n11083) );
  XNOR U11923 ( .A(n11084), .B(n11085), .Z(n8336) );
  XNOR U11924 ( .A(n11086), .B(n9910), .Z(n7170) );
  XOR U11925 ( .A(n11087), .B(n11088), .Z(n6123) );
  XOR U11926 ( .A(n3383), .B(n5756), .Z(n11088) );
  XOR U11927 ( .A(n11089), .B(n7111), .Z(n5756) );
  XNOR U11928 ( .A(n11090), .B(n10868), .Z(n7111) );
  NOR U11929 ( .A(n10996), .B(n7110), .Z(n11089) );
  XNOR U11930 ( .A(n11091), .B(n7118), .Z(n3383) );
  XOR U11931 ( .A(n11092), .B(n11093), .Z(n7118) );
  NOR U11932 ( .A(n8276), .B(n7119), .Z(n11091) );
  XNOR U11933 ( .A(n11094), .B(n10646), .Z(n7119) );
  XOR U11934 ( .A(n11095), .B(n9755), .Z(n8276) );
  XNOR U11935 ( .A(n5427), .B(n11096), .Z(n11087) );
  XNOR U11936 ( .A(n7095), .B(n2251), .Z(n11096) );
  XNOR U11937 ( .A(n11097), .B(n7105), .Z(n2251) );
  XOR U11938 ( .A(n11098), .B(n11099), .Z(n7105) );
  ANDN U11939 ( .B(n7106), .A(n10992), .Z(n11097) );
  IV U11940 ( .A(n8279), .Z(n10992) );
  XOR U11941 ( .A(n11100), .B(n11101), .Z(n8279) );
  XOR U11942 ( .A(n11102), .B(n11103), .Z(n7106) );
  XNOR U11943 ( .A(n11104), .B(n7114), .Z(n7095) );
  XOR U11944 ( .A(n11105), .B(n11106), .Z(n7114) );
  AND U11945 ( .A(n7115), .B(n8281), .Z(n11104) );
  XOR U11946 ( .A(n10399), .B(n11107), .Z(n8281) );
  XOR U11947 ( .A(n11108), .B(n11109), .Z(n7115) );
  XNOR U11948 ( .A(n11110), .B(n7101), .Z(n5427) );
  XOR U11949 ( .A(n11111), .B(n11112), .Z(n7101) );
  ANDN U11950 ( .B(n7102), .A(n8284), .Z(n11110) );
  XOR U11951 ( .A(n11113), .B(n11114), .Z(n8284) );
  XNOR U11952 ( .A(n11115), .B(n11116), .Z(n7102) );
  XOR U11953 ( .A(n11117), .B(n7110), .Z(n8274) );
  XNOR U11954 ( .A(n11118), .B(n11119), .Z(n7110) );
  ANDN U11955 ( .B(n10996), .A(n8228), .Z(n11117) );
  IV U11956 ( .A(n10997), .Z(n8228) );
  XOR U11957 ( .A(n11120), .B(n10088), .Z(n10997) );
  IV U11958 ( .A(n11078), .Z(n10088) );
  XOR U11959 ( .A(n11121), .B(n11122), .Z(n11078) );
  XNOR U11960 ( .A(n11123), .B(n11124), .Z(n10996) );
  AND U11961 ( .A(n5646), .B(n5644), .Z(n11064) );
  XNOR U11962 ( .A(n11125), .B(n1727), .Z(n5644) );
  XOR U11963 ( .A(n11126), .B(n11127), .Z(n9090) );
  XNOR U11964 ( .A(n3474), .B(n5081), .Z(n11127) );
  XOR U11965 ( .A(n11128), .B(n8165), .Z(n5081) );
  ANDN U11966 ( .B(n11014), .A(n8166), .Z(n11128) );
  XNOR U11967 ( .A(n11129), .B(n9188), .Z(n3474) );
  ANDN U11968 ( .B(n9187), .A(n11018), .Z(n11129) );
  XNOR U11969 ( .A(n4129), .B(n11130), .Z(n11126) );
  XOR U11970 ( .A(n8155), .B(n2442), .Z(n11130) );
  XOR U11971 ( .A(n11131), .B(n8175), .Z(n2442) );
  ANDN U11972 ( .B(n8176), .A(n11132), .Z(n11131) );
  XOR U11973 ( .A(n11133), .B(n8161), .Z(n8155) );
  XOR U11974 ( .A(n11134), .B(n8171), .Z(n4129) );
  NOR U11975 ( .A(n11135), .B(n11005), .Z(n11134) );
  XOR U11976 ( .A(n11136), .B(n11137), .Z(n6294) );
  XOR U11977 ( .A(n5416), .B(n3661), .Z(n11137) );
  XOR U11978 ( .A(n11138), .B(n11139), .Z(n3661) );
  ANDN U11979 ( .B(n11140), .A(n11141), .Z(n11138) );
  XNOR U11980 ( .A(n11142), .B(n11143), .Z(n5416) );
  ANDN U11981 ( .B(n8186), .A(n11144), .Z(n11142) );
  XNOR U11982 ( .A(n11145), .B(n11146), .Z(n11136) );
  XOR U11983 ( .A(n2085), .B(n5558), .Z(n11146) );
  XOR U11984 ( .A(n11147), .B(n11148), .Z(n5558) );
  XOR U11985 ( .A(n11150), .B(n11151), .Z(n2085) );
  XOR U11986 ( .A(n10033), .B(n5182), .Z(n5646) );
  XOR U11987 ( .A(n8717), .B(n7527), .Z(n5182) );
  XOR U11988 ( .A(n11153), .B(n11154), .Z(n7527) );
  XOR U11989 ( .A(n10127), .B(n4240), .Z(n11154) );
  XNOR U11990 ( .A(n11155), .B(n7604), .Z(n4240) );
  IV U11991 ( .A(n10468), .Z(n7604) );
  XOR U11992 ( .A(n11156), .B(n10329), .Z(n10468) );
  NOR U11993 ( .A(n11157), .B(n10467), .Z(n11155) );
  XOR U11994 ( .A(n11158), .B(n7600), .Z(n10127) );
  XOR U11995 ( .A(n11159), .B(n9645), .Z(n7600) );
  NOR U11996 ( .A(n10028), .B(n10027), .Z(n11158) );
  XNOR U11997 ( .A(n11160), .B(n10406), .Z(n10027) );
  XOR U11998 ( .A(n3787), .B(n11161), .Z(n11153) );
  XNOR U11999 ( .A(n5129), .B(n1684), .Z(n11161) );
  XOR U12000 ( .A(n11162), .B(n10459), .Z(n1684) );
  IV U12001 ( .A(n7594), .Z(n10459) );
  XOR U12002 ( .A(n11163), .B(n10125), .Z(n7594) );
  XNOR U12003 ( .A(n11164), .B(n11124), .Z(n10036) );
  XOR U12004 ( .A(n11165), .B(n8655), .Z(n5129) );
  XNOR U12005 ( .A(n11166), .B(n11167), .Z(n8655) );
  NOR U12006 ( .A(n10040), .B(n10039), .Z(n11165) );
  XOR U12007 ( .A(n10321), .B(n11168), .Z(n10039) );
  IV U12008 ( .A(n9559), .Z(n10321) );
  XNOR U12009 ( .A(n11169), .B(n10465), .Z(n3787) );
  XNOR U12010 ( .A(n11170), .B(n10057), .Z(n10030) );
  XOR U12011 ( .A(n11171), .B(n11172), .Z(n8717) );
  XOR U12012 ( .A(n6255), .B(n2296), .Z(n11172) );
  XNOR U12013 ( .A(n11173), .B(n10136), .Z(n2296) );
  AND U12014 ( .A(n7646), .B(n7648), .Z(n11173) );
  XOR U12015 ( .A(n11174), .B(n9559), .Z(n7646) );
  XNOR U12016 ( .A(n11175), .B(n11176), .Z(n9559) );
  XNOR U12017 ( .A(n11177), .B(n10141), .Z(n6255) );
  NOR U12018 ( .A(n11178), .B(n7637), .Z(n11177) );
  XNOR U12019 ( .A(n9620), .B(n11179), .Z(n7637) );
  XOR U12020 ( .A(n3893), .B(n11180), .Z(n11171) );
  XOR U12021 ( .A(n5154), .B(n5443), .Z(n11180) );
  XNOR U12022 ( .A(n11181), .B(n10133), .Z(n5443) );
  ANDN U12023 ( .B(n7652), .A(n7650), .Z(n11181) );
  XNOR U12024 ( .A(n11182), .B(n10329), .Z(n7650) );
  XNOR U12025 ( .A(n11183), .B(n11184), .Z(n5154) );
  ANDN U12026 ( .B(n8714), .A(n11185), .Z(n11183) );
  XNOR U12027 ( .A(n11186), .B(n10182), .Z(n8714) );
  XNOR U12028 ( .A(n11187), .B(n11188), .Z(n3893) );
  ANDN U12029 ( .B(n7643), .A(n7642), .Z(n11187) );
  XNOR U12030 ( .A(n11189), .B(n10467), .Z(n10033) );
  XOR U12031 ( .A(n11190), .B(n11043), .Z(n10467) );
  ANDN U12032 ( .B(n11157), .A(n7602), .Z(n11189) );
  XNOR U12033 ( .A(n11191), .B(n6165), .Z(out[1013]) );
  IV U12034 ( .A(n6717), .Z(n6165) );
  XOR U12035 ( .A(n8327), .B(n5902), .Z(n6717) );
  XOR U12036 ( .A(n6128), .B(n6048), .Z(n5902) );
  XOR U12037 ( .A(n11192), .B(n11193), .Z(n6048) );
  XNOR U12038 ( .A(n3685), .B(n4167), .Z(n11193) );
  XNOR U12039 ( .A(n11194), .B(n8392), .Z(n4167) );
  ANDN U12040 ( .B(n8324), .A(n7185), .Z(n11194) );
  XOR U12041 ( .A(n11195), .B(n11196), .Z(n7185) );
  XNOR U12042 ( .A(n10690), .B(n11197), .Z(n8324) );
  XNOR U12043 ( .A(n11198), .B(n11199), .Z(n3685) );
  NOR U12044 ( .A(n8322), .B(n7198), .Z(n11198) );
  XOR U12045 ( .A(n11200), .B(n10822), .Z(n7198) );
  XOR U12046 ( .A(n5263), .B(n11201), .Z(n11192) );
  XOR U12047 ( .A(n8365), .B(n1896), .Z(n11201) );
  XNOR U12048 ( .A(n11202), .B(n8384), .Z(n1896) );
  ANDN U12049 ( .B(n7202), .A(n8317), .Z(n11202) );
  XNOR U12050 ( .A(n11203), .B(n9329), .Z(n8317) );
  XOR U12051 ( .A(n11204), .B(n11205), .Z(n7202) );
  XNOR U12052 ( .A(n11206), .B(n11207), .Z(n8365) );
  ANDN U12053 ( .B(n7189), .A(n8320), .Z(n11206) );
  XNOR U12054 ( .A(n11208), .B(n9788), .Z(n8320) );
  XNOR U12055 ( .A(n11209), .B(n11210), .Z(n7189) );
  XNOR U12056 ( .A(n11211), .B(n8389), .Z(n5263) );
  ANDN U12057 ( .B(n7194), .A(n8390), .Z(n11211) );
  XNOR U12058 ( .A(n11212), .B(n11213), .Z(n8390) );
  XNOR U12059 ( .A(n10947), .B(n11214), .Z(n7194) );
  XOR U12060 ( .A(n11215), .B(n11216), .Z(n6128) );
  XOR U12061 ( .A(n3388), .B(n5785), .Z(n11216) );
  XOR U12062 ( .A(n11218), .B(n10985), .Z(n7168) );
  ANDN U12063 ( .B(n11072), .A(n7167), .Z(n11217) );
  XNOR U12064 ( .A(n11219), .B(n7175), .Z(n3388) );
  XOR U12065 ( .A(n11220), .B(n11221), .Z(n7175) );
  AND U12066 ( .A(n7176), .B(n8330), .Z(n11219) );
  XNOR U12067 ( .A(n11222), .B(n9856), .Z(n8330) );
  XNOR U12068 ( .A(n11223), .B(n11224), .Z(n7176) );
  XOR U12069 ( .A(n5431), .B(n11225), .Z(n11215) );
  XOR U12070 ( .A(n7152), .B(n2258), .Z(n11225) );
  XOR U12071 ( .A(n11226), .B(n7163), .Z(n2258) );
  XOR U12072 ( .A(n11227), .B(n11114), .Z(n7163) );
  NOR U12073 ( .A(n8333), .B(n7162), .Z(n11226) );
  XOR U12074 ( .A(n11228), .B(n11229), .Z(n7162) );
  XOR U12075 ( .A(n11230), .B(n10221), .Z(n8333) );
  XNOR U12076 ( .A(n11231), .B(n7171), .Z(n7152) );
  XOR U12077 ( .A(n11232), .B(n10714), .Z(n7171) );
  AND U12078 ( .A(n7172), .B(n8335), .Z(n11231) );
  XOR U12079 ( .A(n10602), .B(n11233), .Z(n8335) );
  XNOR U12080 ( .A(n11234), .B(n11235), .Z(n7172) );
  XOR U12081 ( .A(n11236), .B(n7159), .Z(n5431) );
  XOR U12082 ( .A(n9132), .B(n11237), .Z(n7159) );
  XOR U12083 ( .A(n11238), .B(n11239), .Z(n8338) );
  XNOR U12084 ( .A(n11240), .B(n9448), .Z(n7158) );
  XNOR U12085 ( .A(n11241), .B(n7167), .Z(n8327) );
  XOR U12086 ( .A(n11242), .B(n11243), .Z(n7167) );
  ANDN U12087 ( .B(n8269), .A(n11072), .Z(n11241) );
  XNOR U12088 ( .A(n11244), .B(n11245), .Z(n11072) );
  XNOR U12089 ( .A(n11246), .B(n10195), .Z(n8269) );
  ANDN U12090 ( .B(n5654), .A(n5652), .Z(n11191) );
  XNOR U12091 ( .A(n11247), .B(n1732), .Z(n5652) );
  XOR U12092 ( .A(n11248), .B(n11249), .Z(n9183) );
  XOR U12093 ( .A(n3478), .B(n5084), .Z(n11249) );
  XNOR U12094 ( .A(n11250), .B(n8192), .Z(n5084) );
  ANDN U12095 ( .B(n8191), .A(n11148), .Z(n11250) );
  XOR U12096 ( .A(n11251), .B(n9287), .Z(n3478) );
  NOR U12097 ( .A(n11151), .B(n9286), .Z(n11251) );
  XNOR U12098 ( .A(n4162), .B(n11252), .Z(n11248) );
  XNOR U12099 ( .A(n8181), .B(n2449), .Z(n11252) );
  XNOR U12100 ( .A(n11253), .B(n8201), .Z(n2449) );
  ANDN U12101 ( .B(n8202), .A(n11254), .Z(n11253) );
  XOR U12102 ( .A(n11255), .B(n8188), .Z(n8181) );
  ANDN U12103 ( .B(n11143), .A(n11256), .Z(n11255) );
  XOR U12104 ( .A(n11257), .B(n8197), .Z(n4162) );
  NOR U12105 ( .A(n11139), .B(n8198), .Z(n11257) );
  XOR U12106 ( .A(n11258), .B(n11259), .Z(n6298) );
  XNOR U12107 ( .A(n5421), .B(n3665), .Z(n11259) );
  XOR U12108 ( .A(n11260), .B(n11261), .Z(n3665) );
  ANDN U12109 ( .B(n11262), .A(n8250), .Z(n11260) );
  IV U12110 ( .A(n11263), .Z(n8250) );
  XNOR U12111 ( .A(n11264), .B(n11265), .Z(n5421) );
  ANDN U12112 ( .B(n8240), .A(n11266), .Z(n11264) );
  XOR U12113 ( .A(n11267), .B(n11268), .Z(n11258) );
  XOR U12114 ( .A(n2088), .B(n4305), .Z(n11268) );
  XNOR U12115 ( .A(n11269), .B(n11270), .Z(n4305) );
  ANDN U12116 ( .B(n11271), .A(n8244), .Z(n11269) );
  XNOR U12117 ( .A(n11272), .B(n11273), .Z(n2088) );
  XOR U12118 ( .A(n10137), .B(n2056), .Z(n5654) );
  IV U12119 ( .A(n5215), .Z(n2056) );
  XOR U12120 ( .A(n7587), .B(n8784), .Z(n5215) );
  XOR U12121 ( .A(n11275), .B(n11276), .Z(n8784) );
  XNOR U12122 ( .A(n5448), .B(n3898), .Z(n11276) );
  XNOR U12123 ( .A(n11277), .B(n11278), .Z(n3898) );
  NOR U12124 ( .A(n7746), .B(n7747), .Z(n11277) );
  XOR U12125 ( .A(n9671), .B(n11279), .Z(n7747) );
  IV U12126 ( .A(n11280), .Z(n9671) );
  XNOR U12127 ( .A(n11281), .B(n10241), .Z(n5448) );
  NOR U12128 ( .A(n10434), .B(n7754), .Z(n11281) );
  XNOR U12129 ( .A(n11282), .B(n11283), .Z(n7754) );
  XOR U12130 ( .A(n11284), .B(n9872), .Z(n10434) );
  XNOR U12131 ( .A(n6259), .B(n11285), .Z(n11275) );
  XNOR U12132 ( .A(n2303), .B(n5184), .Z(n11285) );
  XNOR U12133 ( .A(n11286), .B(n10252), .Z(n5184) );
  ANDN U12134 ( .B(n8780), .A(n8781), .Z(n11286) );
  XOR U12135 ( .A(n11287), .B(n11288), .Z(n8781) );
  XNOR U12136 ( .A(n11289), .B(n10316), .Z(n8780) );
  XOR U12137 ( .A(n11290), .B(n10244), .Z(n2303) );
  ANDN U12138 ( .B(n7750), .A(n7751), .Z(n11290) );
  XOR U12139 ( .A(n9452), .B(n11291), .Z(n7751) );
  XOR U12140 ( .A(n11292), .B(n9664), .Z(n7750) );
  XOR U12141 ( .A(n11293), .B(n10249), .Z(n6259) );
  NOR U12142 ( .A(n7741), .B(n7742), .Z(n11293) );
  XOR U12143 ( .A(n11294), .B(n11295), .Z(n7742) );
  XOR U12144 ( .A(n11296), .B(n9764), .Z(n7741) );
  XOR U12145 ( .A(n11297), .B(n11298), .Z(n7587) );
  XOR U12146 ( .A(n3793), .B(n5132), .Z(n11298) );
  XOR U12147 ( .A(n11299), .B(n8715), .Z(n5132) );
  NOR U12148 ( .A(n11184), .B(n10143), .Z(n11299) );
  IV U12149 ( .A(n10144), .Z(n11184) );
  XOR U12150 ( .A(n11300), .B(n11301), .Z(n10144) );
  XOR U12151 ( .A(n11302), .B(n7647), .Z(n3793) );
  ANDN U12152 ( .B(n10135), .A(n10136), .Z(n11302) );
  XNOR U12153 ( .A(n11303), .B(n11304), .Z(n10136) );
  XNOR U12154 ( .A(n4242), .B(n11305), .Z(n11297) );
  XOR U12155 ( .A(n1688), .B(n10235), .Z(n11305) );
  XOR U12156 ( .A(n11306), .B(n7651), .Z(n10235) );
  ANDN U12157 ( .B(n11307), .A(n10133), .Z(n11306) );
  XOR U12158 ( .A(n9280), .B(n11308), .Z(n10133) );
  IV U12159 ( .A(n10816), .Z(n9280) );
  NOR U12160 ( .A(n10141), .B(n10140), .Z(n11309) );
  XOR U12161 ( .A(n11310), .B(n10057), .Z(n10141) );
  XOR U12162 ( .A(n11311), .B(n7644), .Z(n4242) );
  ANDN U12163 ( .B(n11312), .A(n11188), .Z(n11311) );
  IV U12164 ( .A(n11313), .Z(n11188) );
  XOR U12165 ( .A(n11314), .B(n11312), .Z(n10137) );
  ANDN U12166 ( .B(n7642), .A(n11313), .Z(n11314) );
  XOR U12167 ( .A(n10743), .B(n11315), .Z(n11313) );
  XNOR U12168 ( .A(n11316), .B(n10396), .Z(n7642) );
  XOR U12169 ( .A(n11317), .B(n6170), .Z(out[1012]) );
  XNOR U12170 ( .A(n8382), .B(n5959), .Z(n6170) );
  XOR U12171 ( .A(n6134), .B(n6054), .Z(n5959) );
  XOR U12172 ( .A(n11318), .B(n11319), .Z(n6054) );
  XNOR U12173 ( .A(n3689), .B(n4170), .Z(n11319) );
  XNOR U12174 ( .A(n11320), .B(n8448), .Z(n4170) );
  NOR U12175 ( .A(n7252), .B(n8379), .Z(n11320) );
  XNOR U12176 ( .A(n11321), .B(n10822), .Z(n8379) );
  XOR U12177 ( .A(n11322), .B(n11323), .Z(n10822) );
  XNOR U12178 ( .A(n11324), .B(n11325), .Z(n7252) );
  XOR U12179 ( .A(n11326), .B(n11327), .Z(n3689) );
  AND U12180 ( .A(n8377), .B(n7265), .Z(n11326) );
  XOR U12181 ( .A(n11328), .B(n9535), .Z(n7265) );
  XNOR U12182 ( .A(n5266), .B(n11329), .Z(n11318) );
  XOR U12183 ( .A(n8420), .B(n1900), .Z(n11329) );
  XOR U12184 ( .A(n11330), .B(n11331), .Z(n1900) );
  NOR U12185 ( .A(n7269), .B(n8371), .Z(n11330) );
  XOR U12186 ( .A(n11332), .B(n10945), .Z(n8371) );
  IV U12187 ( .A(n10496), .Z(n10945) );
  XNOR U12188 ( .A(n11333), .B(n10329), .Z(n7269) );
  XNOR U12189 ( .A(n11334), .B(n8444), .Z(n8420) );
  ANDN U12190 ( .B(n8375), .A(n7256), .Z(n11334) );
  XOR U12191 ( .A(n11335), .B(n11116), .Z(n7256) );
  XOR U12192 ( .A(n11336), .B(n9886), .Z(n8375) );
  XOR U12193 ( .A(n11337), .B(n8446), .Z(n5266) );
  ANDN U12194 ( .B(n8369), .A(n7261), .Z(n11337) );
  XNOR U12195 ( .A(n10282), .B(n11338), .Z(n7261) );
  XOR U12196 ( .A(n11339), .B(n11340), .Z(n8369) );
  XOR U12197 ( .A(n11341), .B(n11342), .Z(n6134) );
  XNOR U12198 ( .A(n3396), .B(n5816), .Z(n11342) );
  XOR U12199 ( .A(n11343), .B(n7200), .Z(n5816) );
  XNOR U12200 ( .A(n11344), .B(n11085), .Z(n7200) );
  XOR U12201 ( .A(n11345), .B(n7204), .Z(n3396) );
  XNOR U12202 ( .A(n11346), .B(n10193), .Z(n7204) );
  NOR U12203 ( .A(n8384), .B(n7203), .Z(n11345) );
  XOR U12204 ( .A(n10873), .B(n11347), .Z(n7203) );
  XOR U12205 ( .A(n9101), .B(n11348), .Z(n8384) );
  XNOR U12206 ( .A(n5435), .B(n11349), .Z(n11341) );
  XOR U12207 ( .A(n7180), .B(n2263), .Z(n11349) );
  XOR U12208 ( .A(n11350), .B(n7191), .Z(n2263) );
  XNOR U12209 ( .A(n11351), .B(n11352), .Z(n7191) );
  NOR U12210 ( .A(n8387), .B(n7190), .Z(n11350) );
  XOR U12211 ( .A(n9107), .B(n11353), .Z(n7190) );
  IV U12212 ( .A(n11207), .Z(n8387) );
  XNOR U12213 ( .A(n11354), .B(n10850), .Z(n11207) );
  XNOR U12214 ( .A(n11355), .B(n7195), .Z(n7180) );
  XNOR U12215 ( .A(n11356), .B(n11357), .Z(n7195) );
  ANDN U12216 ( .B(n7196), .A(n8389), .Z(n11355) );
  XNOR U12217 ( .A(n11358), .B(n10729), .Z(n8389) );
  XNOR U12218 ( .A(n11359), .B(n11360), .Z(n7196) );
  XOR U12219 ( .A(n11361), .B(n7187), .Z(n5435) );
  XNOR U12220 ( .A(n11362), .B(n9277), .Z(n7187) );
  NOR U12221 ( .A(n7186), .B(n8392), .Z(n11361) );
  XNOR U12222 ( .A(n11363), .B(n11364), .Z(n8392) );
  XOR U12223 ( .A(n9544), .B(n11365), .Z(n7186) );
  XNOR U12224 ( .A(n11366), .B(n7199), .Z(n8382) );
  XOR U12225 ( .A(n11367), .B(n10971), .Z(n7199) );
  ANDN U12226 ( .B(n8322), .A(n11199), .Z(n11366) );
  XOR U12227 ( .A(n11368), .B(n11369), .Z(n11199) );
  XNOR U12228 ( .A(n11370), .B(n10329), .Z(n8322) );
  XOR U12229 ( .A(n11371), .B(n11372), .Z(n10329) );
  AND U12230 ( .A(n5658), .B(n5656), .Z(n11317) );
  XNOR U12231 ( .A(n11373), .B(n1736), .Z(n5656) );
  XOR U12232 ( .A(n11374), .B(n11375), .Z(n9282) );
  XOR U12233 ( .A(n3480), .B(n5087), .Z(n11375) );
  XOR U12234 ( .A(n11376), .B(n8245), .Z(n5087) );
  ANDN U12235 ( .B(n11270), .A(n11377), .Z(n11376) );
  XNOR U12236 ( .A(n11378), .B(n9408), .Z(n3480) );
  AND U12237 ( .A(n9407), .B(n11273), .Z(n11378) );
  XNOR U12238 ( .A(n4198), .B(n11379), .Z(n11374) );
  XNOR U12239 ( .A(n8235), .B(n2456), .Z(n11379) );
  XNOR U12240 ( .A(n11380), .B(n8256), .Z(n2456) );
  ANDN U12241 ( .B(n11381), .A(n11382), .Z(n11380) );
  XNOR U12242 ( .A(n11383), .B(n8242), .Z(n8235) );
  ANDN U12243 ( .B(n8241), .A(n11384), .Z(n11383) );
  XOR U12244 ( .A(n11385), .B(n8251), .Z(n4198) );
  NOR U12245 ( .A(n11261), .B(n8252), .Z(n11385) );
  XOR U12246 ( .A(n11386), .B(n11387), .Z(n6302) );
  XOR U12247 ( .A(n5425), .B(n3669), .Z(n11387) );
  XOR U12248 ( .A(n11388), .B(n11389), .Z(n3669) );
  NOR U12249 ( .A(n8304), .B(n11390), .Z(n11388) );
  IV U12250 ( .A(n11391), .Z(n8304) );
  XNOR U12251 ( .A(n11392), .B(n11393), .Z(n5425) );
  ANDN U12252 ( .B(n11394), .A(n8294), .Z(n11392) );
  IV U12253 ( .A(n11395), .Z(n8294) );
  XNOR U12254 ( .A(n11396), .B(n11397), .Z(n11386) );
  XOR U12255 ( .A(n2091), .B(n4309), .Z(n11397) );
  XNOR U12256 ( .A(n11398), .B(n11399), .Z(n4309) );
  ANDN U12257 ( .B(n11400), .A(n8298), .Z(n11398) );
  IV U12258 ( .A(n11401), .Z(n8298) );
  XOR U12259 ( .A(n11402), .B(n11403), .Z(n2091) );
  ANDN U12260 ( .B(n11404), .A(n11405), .Z(n11402) );
  XOR U12261 ( .A(n10245), .B(n5380), .Z(n5658) );
  XOR U12262 ( .A(n7632), .B(n8844), .Z(n5380) );
  XOR U12263 ( .A(n11406), .B(n11407), .Z(n8844) );
  XOR U12264 ( .A(n5451), .B(n3903), .Z(n11407) );
  XOR U12265 ( .A(n11408), .B(n11409), .Z(n3903) );
  NOR U12266 ( .A(n10567), .B(n7802), .Z(n11408) );
  XOR U12267 ( .A(n11410), .B(n9817), .Z(n10567) );
  XNOR U12268 ( .A(n10413), .B(n11411), .Z(n5451) );
  XOR U12269 ( .A(n4677), .B(n11412), .Z(n11411) );
  OR U12270 ( .A(n7799), .B(n10414), .Z(n11412) );
  XOR U12271 ( .A(n11413), .B(n11414), .Z(n10414) );
  XNOR U12272 ( .A(n11415), .B(n11416), .Z(n7799) );
  ANDN U12273 ( .B(n11417), .A(rc_i[2]), .Z(n4677) );
  XOR U12274 ( .A(n6263), .B(n11418), .Z(n11406) );
  XOR U12275 ( .A(n2314), .B(n5216), .Z(n11418) );
  XNOR U12276 ( .A(n11419), .B(n10426), .Z(n5216) );
  ANDN U12277 ( .B(n8848), .A(n8846), .Z(n11419) );
  IV U12278 ( .A(n10427), .Z(n8846) );
  XOR U12279 ( .A(n11420), .B(n10962), .Z(n10427) );
  XNOR U12280 ( .A(n11421), .B(n10080), .Z(n8848) );
  XNOR U12281 ( .A(n11422), .B(n10417), .Z(n2314) );
  NOR U12282 ( .A(n7788), .B(n7789), .Z(n11422) );
  XOR U12283 ( .A(n9554), .B(n11423), .Z(n7789) );
  IV U12284 ( .A(n10202), .Z(n9554) );
  XOR U12285 ( .A(n10095), .B(n11424), .Z(n7788) );
  XNOR U12286 ( .A(n11425), .B(n10422), .Z(n6263) );
  ANDN U12287 ( .B(n7794), .A(n10423), .Z(n11425) );
  XOR U12288 ( .A(n11426), .B(n9866), .Z(n10423) );
  XNOR U12289 ( .A(n11427), .B(n10346), .Z(n7794) );
  XOR U12290 ( .A(n11428), .B(n11429), .Z(n7632) );
  XOR U12291 ( .A(n3798), .B(n5135), .Z(n11429) );
  XNOR U12292 ( .A(n11430), .B(n10436), .Z(n5135) );
  IV U12293 ( .A(n8782), .Z(n10436) );
  XOR U12294 ( .A(n10754), .B(n11431), .Z(n8782) );
  NOR U12295 ( .A(n10252), .B(n10251), .Z(n11430) );
  XOR U12296 ( .A(n9809), .B(n11432), .Z(n10251) );
  IV U12297 ( .A(n10095), .Z(n9809) );
  XOR U12298 ( .A(n11433), .B(n11434), .Z(n10252) );
  XNOR U12299 ( .A(n11435), .B(n7752), .Z(n3798) );
  XOR U12300 ( .A(n11436), .B(n11437), .Z(n7752) );
  ANDN U12301 ( .B(n10244), .A(n10243), .Z(n11435) );
  XOR U12302 ( .A(n9151), .B(n11438), .Z(n10243) );
  XOR U12303 ( .A(n11439), .B(n11440), .Z(n10244) );
  XNOR U12304 ( .A(n4245), .B(n11441), .Z(n11428) );
  XOR U12305 ( .A(n1692), .B(n10408), .Z(n11441) );
  XNOR U12306 ( .A(n11442), .B(n7755), .Z(n10408) );
  XOR U12307 ( .A(n11443), .B(n11444), .Z(n7755) );
  NOR U12308 ( .A(n10241), .B(n10240), .Z(n11442) );
  XOR U12309 ( .A(n11445), .B(n11446), .Z(n10240) );
  XOR U12310 ( .A(n11447), .B(n11448), .Z(n10241) );
  XNOR U12311 ( .A(n11450), .B(n10357), .Z(n7743) );
  ANDN U12312 ( .B(n10249), .A(n10248), .Z(n11449) );
  XOR U12313 ( .A(n11451), .B(n11369), .Z(n10248) );
  XOR U12314 ( .A(n10159), .B(n11452), .Z(n10249) );
  XOR U12315 ( .A(n11453), .B(n7748), .Z(n4245) );
  XNOR U12316 ( .A(n11454), .B(n11414), .Z(n7748) );
  ANDN U12317 ( .B(n10438), .A(n11278), .Z(n11453) );
  XNOR U12318 ( .A(n11455), .B(n10438), .Z(n10245) );
  XOR U12319 ( .A(n10167), .B(n11456), .Z(n10438) );
  AND U12320 ( .A(n7746), .B(n11278), .Z(n11455) );
  XOR U12321 ( .A(n11457), .B(n11458), .Z(n11278) );
  XOR U12322 ( .A(n11459), .B(n11460), .Z(n7746) );
  XOR U12323 ( .A(n11461), .B(n6180), .Z(out[1011]) );
  XOR U12324 ( .A(n8438), .B(n6013), .Z(n6180) );
  XOR U12325 ( .A(n6139), .B(n6059), .Z(n6013) );
  XOR U12326 ( .A(n11462), .B(n11463), .Z(n6059) );
  XOR U12327 ( .A(n3696), .B(n4173), .Z(n11463) );
  XNOR U12328 ( .A(n11464), .B(n8483), .Z(n4173) );
  ANDN U12329 ( .B(n7309), .A(n8434), .Z(n11464) );
  XNOR U12330 ( .A(n11465), .B(n11466), .Z(n8434) );
  XOR U12331 ( .A(n11467), .B(n11468), .Z(n7309) );
  XOR U12332 ( .A(n11469), .B(n11470), .Z(n3696) );
  ANDN U12333 ( .B(n7322), .A(n8432), .Z(n11469) );
  XOR U12334 ( .A(n10621), .B(n11471), .Z(n7322) );
  IV U12335 ( .A(n9627), .Z(n10621) );
  XNOR U12336 ( .A(n5268), .B(n11472), .Z(n11462) );
  XNOR U12337 ( .A(n8454), .B(n1904), .Z(n11472) );
  XOR U12338 ( .A(n11473), .B(n8475), .Z(n1904) );
  ANDN U12339 ( .B(n8426), .A(n7326), .Z(n11473) );
  XOR U12340 ( .A(n11474), .B(n11283), .Z(n7326) );
  XOR U12341 ( .A(n9530), .B(n11475), .Z(n8426) );
  XNOR U12342 ( .A(n11476), .B(n8478), .Z(n8454) );
  ANDN U12343 ( .B(n8430), .A(n7313), .Z(n11476) );
  XOR U12344 ( .A(n11477), .B(n9448), .Z(n7313) );
  XNOR U12345 ( .A(n11478), .B(n11479), .Z(n8430) );
  XNOR U12346 ( .A(n11480), .B(n8481), .Z(n5268) );
  ANDN U12347 ( .B(n7318), .A(n8424), .Z(n11480) );
  XNOR U12348 ( .A(n11481), .B(n11482), .Z(n8424) );
  XNOR U12349 ( .A(n11483), .B(n10125), .Z(n7318) );
  XOR U12350 ( .A(n11484), .B(n11485), .Z(n6139) );
  XOR U12351 ( .A(n3400), .B(n5842), .Z(n11485) );
  XNOR U12352 ( .A(n11486), .B(n7266), .Z(n5842) );
  XOR U12353 ( .A(n11487), .B(n11213), .Z(n7266) );
  ANDN U12354 ( .B(n7267), .A(n11327), .Z(n11486) );
  XOR U12355 ( .A(n11488), .B(n8372), .Z(n3400) );
  XOR U12356 ( .A(n11489), .B(n11490), .Z(n8372) );
  ANDN U12357 ( .B(n8441), .A(n8440), .Z(n11488) );
  XOR U12358 ( .A(n11491), .B(n10990), .Z(n8440) );
  IV U12359 ( .A(n11331), .Z(n8441) );
  XOR U12360 ( .A(n11492), .B(n9260), .Z(n11331) );
  XOR U12361 ( .A(n5439), .B(n11493), .Z(n11484) );
  XOR U12362 ( .A(n7247), .B(n2272), .Z(n11493) );
  XNOR U12363 ( .A(n11494), .B(n7257), .Z(n2272) );
  XNOR U12364 ( .A(n11495), .B(n11364), .Z(n7257) );
  ANDN U12365 ( .B(n7258), .A(n8444), .Z(n11494) );
  XNOR U12366 ( .A(n11496), .B(n10526), .Z(n8444) );
  XOR U12367 ( .A(n9263), .B(n11497), .Z(n7258) );
  XNOR U12368 ( .A(n11498), .B(n7262), .Z(n7247) );
  XNOR U12369 ( .A(n10885), .B(n11499), .Z(n7262) );
  ANDN U12370 ( .B(n7263), .A(n8446), .Z(n11498) );
  XNOR U12371 ( .A(n10968), .B(n11500), .Z(n8446) );
  IV U12372 ( .A(n11501), .Z(n10968) );
  XNOR U12373 ( .A(n11502), .B(n11503), .Z(n7263) );
  XNOR U12374 ( .A(n11504), .B(n7254), .Z(n5439) );
  XOR U12375 ( .A(n11505), .B(n10521), .Z(n7254) );
  ANDN U12376 ( .B(n8448), .A(n7253), .Z(n11504) );
  XOR U12377 ( .A(n11506), .B(n9650), .Z(n7253) );
  XOR U12378 ( .A(n11507), .B(n11508), .Z(n8448) );
  XNOR U12379 ( .A(n11509), .B(n7267), .Z(n8438) );
  XOR U12380 ( .A(n11510), .B(n11511), .Z(n7267) );
  ANDN U12381 ( .B(n11327), .A(n8377), .Z(n11509) );
  XOR U12382 ( .A(n11512), .B(n11513), .Z(n8377) );
  XOR U12383 ( .A(n11514), .B(n11515), .Z(n11327) );
  ANDN U12384 ( .B(n5662), .A(n5660), .Z(n11461) );
  XNOR U12385 ( .A(n11516), .B(n1741), .Z(n5660) );
  XOR U12386 ( .A(n11517), .B(n11518), .Z(n9403) );
  XNOR U12387 ( .A(n3482), .B(n5091), .Z(n11518) );
  XNOR U12388 ( .A(n11519), .B(n8300), .Z(n5091) );
  AND U12389 ( .A(n8299), .B(n11399), .Z(n11519) );
  XNOR U12390 ( .A(n11520), .B(n9502), .Z(n3482) );
  NOR U12391 ( .A(n11403), .B(n9501), .Z(n11520) );
  XOR U12392 ( .A(n4231), .B(n11521), .Z(n11517) );
  XNOR U12393 ( .A(n8289), .B(n2467), .Z(n11521) );
  XNOR U12394 ( .A(n11522), .B(n8309), .Z(n2467) );
  IV U12395 ( .A(n11523), .Z(n8309) );
  ANDN U12396 ( .B(n8310), .A(n11524), .Z(n11522) );
  XOR U12397 ( .A(n11525), .B(n8295), .Z(n8289) );
  ANDN U12398 ( .B(n8296), .A(n11393), .Z(n11525) );
  XNOR U12399 ( .A(n11526), .B(n8306), .Z(n4231) );
  ANDN U12400 ( .B(n11389), .A(n8305), .Z(n11526) );
  XOR U12401 ( .A(n11527), .B(n11528), .Z(n6306) );
  XNOR U12402 ( .A(n5429), .B(n3677), .Z(n11528) );
  NOR U12403 ( .A(n11531), .B(n8358), .Z(n11529) );
  XNOR U12404 ( .A(n11532), .B(n11533), .Z(n5429) );
  NOR U12405 ( .A(n8348), .B(n11534), .Z(n11532) );
  XNOR U12406 ( .A(n11535), .B(n11536), .Z(n11527) );
  XNOR U12407 ( .A(n2094), .B(n4314), .Z(n11536) );
  XNOR U12408 ( .A(n11537), .B(n11538), .Z(n4314) );
  AND U12409 ( .A(n8352), .B(n11539), .Z(n11537) );
  XNOR U12410 ( .A(n11540), .B(n11541), .Z(n2094) );
  XOR U12411 ( .A(n10418), .B(n5279), .Z(n5662) );
  XOR U12412 ( .A(n7736), .B(n8910), .Z(n5279) );
  XOR U12413 ( .A(n11543), .B(n11544), .Z(n8910) );
  XNOR U12414 ( .A(n5456), .B(n3907), .Z(n11544) );
  XOR U12415 ( .A(n11545), .B(n11546), .Z(n3907) );
  ANDN U12416 ( .B(n7887), .A(n7885), .Z(n11545) );
  XOR U12417 ( .A(n11547), .B(n11548), .Z(n7887) );
  XOR U12418 ( .A(n11549), .B(n10543), .Z(n5456) );
  NOR U12419 ( .A(n10544), .B(n7882), .Z(n11549) );
  XOR U12420 ( .A(n11092), .B(n11550), .Z(n7882) );
  XOR U12421 ( .A(n11551), .B(n10761), .Z(n10544) );
  XOR U12422 ( .A(n6267), .B(n11552), .Z(n11543) );
  XOR U12423 ( .A(n2321), .B(n5250), .Z(n11552) );
  XOR U12424 ( .A(n11553), .B(n10557), .Z(n5250) );
  XNOR U12425 ( .A(n11554), .B(n10185), .Z(n8913) );
  XOR U12426 ( .A(n10878), .B(n11555), .Z(n8912) );
  XNOR U12427 ( .A(n11556), .B(n10547), .Z(n2321) );
  ANDN U12428 ( .B(n7873), .A(n7871), .Z(n11556) );
  IV U12429 ( .A(n10548), .Z(n7871) );
  XOR U12430 ( .A(n11557), .B(n9905), .Z(n10548) );
  XNOR U12431 ( .A(n11558), .B(n11559), .Z(n7873) );
  XNOR U12432 ( .A(n11560), .B(n10553), .Z(n6267) );
  NOR U12433 ( .A(n10554), .B(n7876), .Z(n11560) );
  XNOR U12434 ( .A(n10743), .B(n11561), .Z(n7876) );
  XOR U12435 ( .A(n11562), .B(n9932), .Z(n10554) );
  XOR U12436 ( .A(n11563), .B(n11564), .Z(n7736) );
  XOR U12437 ( .A(n3803), .B(n5138), .Z(n11564) );
  XNOR U12438 ( .A(n11565), .B(n8847), .Z(n5138) );
  XOR U12439 ( .A(n11566), .B(n10855), .Z(n8847) );
  ANDN U12440 ( .B(n10425), .A(n10426), .Z(n11565) );
  XOR U12441 ( .A(n11567), .B(n11568), .Z(n10426) );
  XOR U12442 ( .A(n11569), .B(n10205), .Z(n10425) );
  IV U12443 ( .A(n9905), .Z(n10205) );
  XOR U12444 ( .A(n11570), .B(n11571), .Z(n9905) );
  XOR U12445 ( .A(n11572), .B(n7790), .Z(n3803) );
  XNOR U12446 ( .A(n11573), .B(n11116), .Z(n7790) );
  NOR U12447 ( .A(n10416), .B(n10417), .Z(n11572) );
  XNOR U12448 ( .A(n11574), .B(n10482), .Z(n10417) );
  XNOR U12449 ( .A(n11575), .B(n9251), .Z(n10416) );
  XNOR U12450 ( .A(n4248), .B(n11576), .Z(n11563) );
  XOR U12451 ( .A(n1697), .B(n10538), .Z(n11576) );
  XOR U12452 ( .A(n11577), .B(n7800), .Z(n10538) );
  XOR U12453 ( .A(n11578), .B(n9954), .Z(n7800) );
  XNOR U12454 ( .A(n11579), .B(n11580), .Z(n9954) );
  ANDN U12455 ( .B(n10412), .A(n10413), .Z(n11577) );
  XOR U12456 ( .A(n11581), .B(n9937), .Z(n10413) );
  XOR U12457 ( .A(n11582), .B(n10836), .Z(n10412) );
  XOR U12458 ( .A(n11583), .B(n10562), .Z(n1697) );
  XOR U12459 ( .A(n11584), .B(n11585), .Z(n10562) );
  ANDN U12460 ( .B(n10421), .A(n10422), .Z(n11583) );
  XNOR U12461 ( .A(n9151), .B(n11586), .Z(n10422) );
  IV U12462 ( .A(n10265), .Z(n9151) );
  XNOR U12463 ( .A(n11587), .B(n11588), .Z(n10265) );
  XOR U12464 ( .A(n11589), .B(n11515), .Z(n10421) );
  XOR U12465 ( .A(n11590), .B(n7804), .Z(n4248) );
  XNOR U12466 ( .A(n11591), .B(n10761), .Z(n7804) );
  ANDN U12467 ( .B(n11409), .A(n10568), .Z(n11590) );
  XNOR U12468 ( .A(n11592), .B(n10568), .Z(n10418) );
  XOR U12469 ( .A(n11593), .B(n10274), .Z(n10568) );
  IV U12470 ( .A(n11440), .Z(n10274) );
  ANDN U12471 ( .B(n7802), .A(n11409), .Z(n11592) );
  XOR U12472 ( .A(n11594), .B(n11595), .Z(n11409) );
  XOR U12473 ( .A(n11596), .B(n10724), .Z(n7802) );
  XOR U12474 ( .A(n11597), .B(n6185), .Z(out[1010]) );
  XOR U12475 ( .A(n8473), .B(n2243), .Z(n6185) );
  XNOR U12476 ( .A(n6063), .B(n6144), .Z(n2243) );
  XNOR U12477 ( .A(n11598), .B(n11599), .Z(n6144) );
  XOR U12478 ( .A(n2279), .B(n5444), .Z(n11599) );
  XNOR U12479 ( .A(n11600), .B(n8435), .Z(n5444) );
  IV U12480 ( .A(n7311), .Z(n8435) );
  XOR U12481 ( .A(n11601), .B(n9463), .Z(n7311) );
  ANDN U12482 ( .B(n8483), .A(n7310), .Z(n11600) );
  XNOR U12483 ( .A(n11602), .B(n11603), .Z(n7310) );
  XOR U12484 ( .A(n11604), .B(n11605), .Z(n8483) );
  XNOR U12485 ( .A(n11606), .B(n7314), .Z(n2279) );
  XNOR U12486 ( .A(n11607), .B(n11508), .Z(n7314) );
  ANDN U12487 ( .B(n7315), .A(n8478), .Z(n11606) );
  XNOR U12488 ( .A(n11608), .B(n10646), .Z(n8478) );
  XNOR U12489 ( .A(n9459), .B(n11609), .Z(n7315) );
  XNOR U12490 ( .A(n3137), .B(n11610), .Z(n11598) );
  XOR U12491 ( .A(n5872), .B(n7304), .Z(n11610) );
  XNOR U12492 ( .A(n11611), .B(n7319), .Z(n7304) );
  XOR U12493 ( .A(n11054), .B(n11612), .Z(n7319) );
  ANDN U12494 ( .B(n8481), .A(n8480), .Z(n11611) );
  XNOR U12495 ( .A(n11613), .B(n11614), .Z(n8480) );
  XNOR U12496 ( .A(n10965), .B(n11615), .Z(n8481) );
  XNOR U12497 ( .A(n11616), .B(n7324), .Z(n5872) );
  XNOR U12498 ( .A(n11617), .B(n11340), .Z(n7324) );
  NOR U12499 ( .A(n11470), .B(n7323), .Z(n11616) );
  XOR U12500 ( .A(n11618), .B(n8427), .Z(n3137) );
  XOR U12501 ( .A(n11619), .B(n10512), .Z(n8427) );
  NOR U12502 ( .A(n7328), .B(n8475), .Z(n11618) );
  XNOR U12503 ( .A(n11620), .B(n10075), .Z(n8475) );
  XOR U12504 ( .A(n11621), .B(n11069), .Z(n7328) );
  XOR U12505 ( .A(n11622), .B(n11623), .Z(n6063) );
  XNOR U12506 ( .A(n5270), .B(n1908), .Z(n11623) );
  XNOR U12507 ( .A(n11624), .B(n8550), .Z(n1908) );
  ANDN U12508 ( .B(n8461), .A(n8551), .Z(n11624) );
  XOR U12509 ( .A(n10686), .B(n11625), .Z(n8551) );
  IV U12510 ( .A(n9131), .Z(n10686) );
  IV U12511 ( .A(n7399), .Z(n8461) );
  XNOR U12512 ( .A(n11626), .B(n11414), .Z(n7399) );
  XOR U12513 ( .A(n11627), .B(n8557), .Z(n5270) );
  ANDN U12514 ( .B(n8458), .A(n7391), .Z(n11627) );
  XNOR U12515 ( .A(n11628), .B(n10231), .Z(n7391) );
  XNOR U12516 ( .A(n11629), .B(n11630), .Z(n8458) );
  XOR U12517 ( .A(n3700), .B(n11631), .Z(n11622) );
  XNOR U12518 ( .A(n8530), .B(n4177), .Z(n11631) );
  XNOR U12519 ( .A(n11632), .B(n8559), .Z(n4177) );
  ANDN U12520 ( .B(n8470), .A(n7382), .Z(n11632) );
  XNOR U12521 ( .A(n11633), .B(n11634), .Z(n7382) );
  XNOR U12522 ( .A(n9627), .B(n11635), .Z(n8470) );
  ANDN U12523 ( .B(n7386), .A(n8555), .Z(n11636) );
  XNOR U12524 ( .A(n11637), .B(n11638), .Z(n8555) );
  XOR U12525 ( .A(n9544), .B(n11639), .Z(n7386) );
  XNOR U12526 ( .A(n11640), .B(n11641), .Z(n3700) );
  ANDN U12527 ( .B(n8468), .A(n11642), .Z(n11640) );
  IV U12528 ( .A(n7395), .Z(n8468) );
  XNOR U12529 ( .A(n11643), .B(n9771), .Z(n7395) );
  XOR U12530 ( .A(n11644), .B(n7323), .Z(n8473) );
  XOR U12531 ( .A(n11645), .B(n10296), .Z(n7323) );
  XNOR U12532 ( .A(n11646), .B(n11414), .Z(n8432) );
  XOR U12533 ( .A(n11647), .B(n11648), .Z(n11470) );
  AND U12534 ( .A(n5666), .B(n5664), .Z(n11597) );
  XOR U12535 ( .A(n11649), .B(n1745), .Z(n5664) );
  XOR U12536 ( .A(n11650), .B(n11651), .Z(n9497) );
  XNOR U12537 ( .A(n3486), .B(n5098), .Z(n11651) );
  XNOR U12538 ( .A(n11652), .B(n8354), .Z(n5098) );
  ANDN U12539 ( .B(n11538), .A(n8353), .Z(n11652) );
  XNOR U12540 ( .A(n11653), .B(n9608), .Z(n3486) );
  ANDN U12541 ( .B(n11541), .A(n9607), .Z(n11653) );
  XOR U12542 ( .A(n4258), .B(n11654), .Z(n11650) );
  XOR U12543 ( .A(n8343), .B(n2474), .Z(n11654) );
  XOR U12544 ( .A(n11655), .B(n8363), .Z(n2474) );
  ANDN U12545 ( .B(n11656), .A(n11657), .Z(n11655) );
  XOR U12546 ( .A(n11658), .B(n8350), .Z(n8343) );
  XOR U12547 ( .A(n11659), .B(n8359), .Z(n4258) );
  ANDN U12548 ( .B(n8360), .A(n11530), .Z(n11659) );
  XOR U12549 ( .A(n11660), .B(n11661), .Z(n6310) );
  XNOR U12550 ( .A(n5434), .B(n3681), .Z(n11661) );
  XOR U12551 ( .A(n11662), .B(n11663), .Z(n3681) );
  ANDN U12552 ( .B(n11664), .A(n11665), .Z(n11662) );
  XNOR U12553 ( .A(n11666), .B(n11667), .Z(n5434) );
  NOR U12554 ( .A(n11668), .B(n11669), .Z(n11666) );
  XNOR U12555 ( .A(n11670), .B(n11671), .Z(n11660) );
  XNOR U12556 ( .A(n2097), .B(n4317), .Z(n11671) );
  XOR U12557 ( .A(n11672), .B(n11673), .Z(n4317) );
  AND U12558 ( .A(n8407), .B(n11674), .Z(n11672) );
  XNOR U12559 ( .A(n11675), .B(n11676), .Z(n2097) );
  ANDN U12560 ( .B(n11677), .A(n9714), .Z(n11675) );
  IV U12561 ( .A(n11678), .Z(n9714) );
  XOR U12562 ( .A(n10549), .B(n5390), .Z(n5666) );
  XOR U12563 ( .A(n7784), .B(n8973), .Z(n5390) );
  XOR U12564 ( .A(n11679), .B(n11680), .Z(n8973) );
  XNOR U12565 ( .A(n5465), .B(n3911), .Z(n11680) );
  NOR U12566 ( .A(n7956), .B(n7955), .Z(n11681) );
  XNOR U12567 ( .A(n11683), .B(n9978), .Z(n7956) );
  XNOR U12568 ( .A(n11684), .B(n10658), .Z(n5465) );
  ANDN U12569 ( .B(n7953), .A(n7951), .Z(n11684) );
  IV U12570 ( .A(n10659), .Z(n7951) );
  XOR U12571 ( .A(n11685), .B(n11686), .Z(n10659) );
  XOR U12572 ( .A(n11687), .B(n11688), .Z(n7953) );
  XOR U12573 ( .A(n6271), .B(n11689), .Z(n11679) );
  XOR U12574 ( .A(n2328), .B(n5281), .Z(n11689) );
  XNOR U12575 ( .A(n11690), .B(n10670), .Z(n5281) );
  XNOR U12576 ( .A(n11691), .B(n10180), .Z(n8976) );
  XOR U12577 ( .A(n11692), .B(n10741), .Z(n8975) );
  XNOR U12578 ( .A(n11693), .B(n10662), .Z(n2328) );
  ANDN U12579 ( .B(n7941), .A(n7942), .Z(n11693) );
  XNOR U12580 ( .A(n9248), .B(n11694), .Z(n7942) );
  XNOR U12581 ( .A(n11695), .B(n9972), .Z(n7941) );
  XNOR U12582 ( .A(n11696), .B(n10667), .Z(n6271) );
  ANDN U12583 ( .B(n7945), .A(n7946), .Z(n11696) );
  XOR U12584 ( .A(n11697), .B(n10640), .Z(n7946) );
  XNOR U12585 ( .A(n11698), .B(n11699), .Z(n7945) );
  XOR U12586 ( .A(n11700), .B(n11701), .Z(n7784) );
  XNOR U12587 ( .A(n3808), .B(n5141), .Z(n11701) );
  XOR U12588 ( .A(n11702), .B(n8914), .Z(n5141) );
  XNOR U12589 ( .A(n11703), .B(n11704), .Z(n8914) );
  ANDN U12590 ( .B(n10557), .A(n10556), .Z(n11702) );
  XOR U12591 ( .A(n11705), .B(n9972), .Z(n10556) );
  IV U12592 ( .A(n10338), .Z(n9972) );
  XNOR U12593 ( .A(n11706), .B(n11707), .Z(n10338) );
  XOR U12594 ( .A(n11708), .B(n9136), .Z(n10557) );
  XOR U12595 ( .A(n11710), .B(n9448), .Z(n7872) );
  NOR U12596 ( .A(n10546), .B(n10547), .Z(n11709) );
  XNOR U12597 ( .A(n11711), .B(n11712), .Z(n10547) );
  IV U12598 ( .A(n10680), .Z(n10546) );
  XOR U12599 ( .A(n11713), .B(n11714), .Z(n10680) );
  XOR U12600 ( .A(n4251), .B(n11715), .Z(n11700) );
  XOR U12601 ( .A(n1702), .B(n10653), .Z(n11715) );
  XNOR U12602 ( .A(n11716), .B(n7883), .Z(n10653) );
  XNOR U12603 ( .A(n11717), .B(n10198), .Z(n7883) );
  ANDN U12604 ( .B(n10543), .A(n10542), .Z(n11716) );
  XOR U12605 ( .A(n11718), .B(n10971), .Z(n10542) );
  XNOR U12606 ( .A(n9565), .B(n11719), .Z(n10543) );
  XOR U12607 ( .A(n11720), .B(n7877), .Z(n1702) );
  XOR U12608 ( .A(n11721), .B(n11722), .Z(n7877) );
  NOR U12609 ( .A(n10553), .B(n10552), .Z(n11720) );
  XNOR U12610 ( .A(n11723), .B(n11648), .Z(n10552) );
  XOR U12611 ( .A(n11724), .B(n9251), .Z(n10553) );
  XOR U12612 ( .A(n11725), .B(n11726), .Z(n9251) );
  XNOR U12613 ( .A(n11727), .B(n10677), .Z(n4251) );
  IV U12614 ( .A(n7886), .Z(n10677) );
  XOR U12615 ( .A(n11728), .B(n11686), .Z(n7886) );
  XNOR U12616 ( .A(n11729), .B(n10678), .Z(n10549) );
  XNOR U12617 ( .A(n11730), .B(n10482), .Z(n10678) );
  ANDN U12618 ( .B(n7885), .A(n11546), .Z(n11729) );
  XNOR U12619 ( .A(n11731), .B(n10868), .Z(n11546) );
  XOR U12620 ( .A(n11732), .B(n11733), .Z(n7885) );
  XNOR U12621 ( .A(n11734), .B(n4205), .Z(out[100]) );
  IV U12622 ( .A(n4379), .Z(n4205) );
  XOR U12623 ( .A(n7024), .B(n2579), .Z(n4379) );
  XNOR U12624 ( .A(n8096), .B(n10974), .Z(n2579) );
  XNOR U12625 ( .A(n11735), .B(n11736), .Z(n10974) );
  XOR U12626 ( .A(n5729), .B(n5423), .Z(n11736) );
  XOR U12627 ( .A(n11737), .B(n7040), .Z(n5423) );
  XOR U12628 ( .A(n11637), .B(n11738), .Z(n7040) );
  ANDN U12629 ( .B(n7041), .A(n8217), .Z(n11737) );
  XNOR U12630 ( .A(n11739), .B(n11099), .Z(n8217) );
  XOR U12631 ( .A(n11740), .B(n11210), .Z(n7041) );
  XNOR U12632 ( .A(n11741), .B(n7050), .Z(n5729) );
  XNOR U12633 ( .A(n11742), .B(n11595), .Z(n7050) );
  ANDN U12634 ( .B(n7049), .A(n10881), .Z(n11741) );
  XOR U12635 ( .A(n11054), .B(n11743), .Z(n10881) );
  XOR U12636 ( .A(n11744), .B(n10609), .Z(n7049) );
  XOR U12637 ( .A(n7034), .B(n11745), .Z(n11735) );
  XOR U12638 ( .A(n2245), .B(n3379), .Z(n11745) );
  XNOR U12639 ( .A(n11746), .B(n7057), .Z(n3379) );
  XOR U12640 ( .A(n11747), .B(n9940), .Z(n7057) );
  ANDN U12641 ( .B(n8209), .A(n8208), .Z(n11746) );
  XOR U12642 ( .A(n11748), .B(n10526), .Z(n8208) );
  XNOR U12643 ( .A(n11749), .B(n9613), .Z(n8209) );
  XOR U12644 ( .A(n11750), .B(n7045), .Z(n2245) );
  XOR U12645 ( .A(n11751), .B(n10842), .Z(n7045) );
  ANDN U12646 ( .B(n8212), .A(n7044), .Z(n11750) );
  XOR U12647 ( .A(n11752), .B(n11704), .Z(n7044) );
  XNOR U12648 ( .A(n11753), .B(n11754), .Z(n8212) );
  XNOR U12649 ( .A(n11755), .B(n7054), .Z(n7034) );
  XNOR U12650 ( .A(n11756), .B(n10386), .Z(n7054) );
  ANDN U12651 ( .B(n8214), .A(n7053), .Z(n11755) );
  XOR U12652 ( .A(n11757), .B(n11758), .Z(n7053) );
  XOR U12653 ( .A(n11759), .B(n10300), .Z(n8214) );
  XOR U12654 ( .A(n11760), .B(n11761), .Z(n8096) );
  XNOR U12655 ( .A(n4385), .B(n2193), .Z(n11761) );
  XOR U12656 ( .A(n11762), .B(n8137), .Z(n2193) );
  XOR U12657 ( .A(n11763), .B(n11595), .Z(n8137) );
  ANDN U12658 ( .B(n10857), .A(n11764), .Z(n11762) );
  XOR U12659 ( .A(n11765), .B(n8129), .Z(n4385) );
  XOR U12660 ( .A(n10280), .B(n11766), .Z(n8129) );
  NOR U12661 ( .A(n7031), .B(n7030), .Z(n11765) );
  XOR U12662 ( .A(n11767), .B(n11768), .Z(n7030) );
  XOR U12663 ( .A(n11769), .B(n9872), .Z(n7031) );
  XNOR U12664 ( .A(n6026), .B(n11770), .Z(n11760) );
  XOR U12665 ( .A(n5562), .B(n3809), .Z(n11770) );
  XNOR U12666 ( .A(n11771), .B(n8133), .Z(n3809) );
  XNOR U12667 ( .A(n11772), .B(n10075), .Z(n8133) );
  ANDN U12668 ( .B(n7020), .A(n10852), .Z(n11771) );
  IV U12669 ( .A(n7021), .Z(n10852) );
  XOR U12670 ( .A(n10738), .B(n11773), .Z(n7021) );
  XOR U12671 ( .A(n11774), .B(n10962), .Z(n7020) );
  XNOR U12672 ( .A(n11775), .B(n10776), .Z(n5562) );
  XOR U12673 ( .A(n11776), .B(n9939), .Z(n10776) );
  ANDN U12674 ( .B(n7028), .A(n7026), .Z(n11775) );
  XOR U12675 ( .A(n11777), .B(n11778), .Z(n7026) );
  IV U12676 ( .A(n10845), .Z(n7028) );
  XOR U12677 ( .A(n11779), .B(n11458), .Z(n10845) );
  XNOR U12678 ( .A(n11780), .B(n8141), .Z(n6026) );
  XNOR U12679 ( .A(n11781), .B(n9879), .Z(n8141) );
  ANDN U12680 ( .B(n10771), .A(n7017), .Z(n11780) );
  XOR U12681 ( .A(n11782), .B(n11479), .Z(n7017) );
  IV U12682 ( .A(n7016), .Z(n10771) );
  XOR U12683 ( .A(n11783), .B(n11224), .Z(n7016) );
  XNOR U12684 ( .A(n11784), .B(n11764), .Z(n7024) );
  IV U12685 ( .A(n10768), .Z(n11764) );
  XOR U12686 ( .A(n9563), .B(n11785), .Z(n10768) );
  NOR U12687 ( .A(n8135), .B(n10857), .Z(n11784) );
  XNOR U12688 ( .A(n11786), .B(n10234), .Z(n10857) );
  IV U12689 ( .A(n10858), .Z(n8135) );
  XOR U12690 ( .A(n11787), .B(n11686), .Z(n10858) );
  ANDN U12691 ( .B(n3671), .A(n3673), .Z(n11734) );
  XOR U12692 ( .A(n3435), .B(n9726), .Z(n3673) );
  XOR U12693 ( .A(n11788), .B(n10575), .Z(n9726) );
  ANDN U12694 ( .B(n10708), .A(n10710), .Z(n11788) );
  XOR U12695 ( .A(n11789), .B(n10357), .Z(n10710) );
  IV U12696 ( .A(n2353), .Z(n3435) );
  XNOR U12697 ( .A(n6223), .B(n10810), .Z(n2353) );
  XOR U12698 ( .A(n11790), .B(n11791), .Z(n10810) );
  XOR U12699 ( .A(n1666), .B(n9825), .Z(n11791) );
  XOR U12700 ( .A(n11792), .B(n7342), .Z(n9825) );
  XOR U12701 ( .A(n9527), .B(n11793), .Z(n7342) );
  NOR U12702 ( .A(n9739), .B(n9738), .Z(n11792) );
  XOR U12703 ( .A(n11584), .B(n11794), .Z(n9738) );
  XNOR U12704 ( .A(n11795), .B(n9329), .Z(n9739) );
  XNOR U12705 ( .A(n11796), .B(n7337), .Z(n1666) );
  XOR U12706 ( .A(n11797), .B(n9910), .Z(n7337) );
  ANDN U12707 ( .B(n9747), .A(n9746), .Z(n11796) );
  XOR U12708 ( .A(n11356), .B(n11798), .Z(n9746) );
  XOR U12709 ( .A(n11799), .B(n10727), .Z(n9747) );
  XOR U12710 ( .A(n3774), .B(n11800), .Z(n11790) );
  XOR U12711 ( .A(n5115), .B(n4228), .Z(n11800) );
  XNOR U12712 ( .A(n11801), .B(n7346), .Z(n4228) );
  XOR U12713 ( .A(n10819), .B(n11802), .Z(n7346) );
  IV U12714 ( .A(n10978), .Z(n10819) );
  NOR U12715 ( .A(n9834), .B(n10685), .Z(n11801) );
  XOR U12716 ( .A(n11803), .B(n10198), .Z(n10685) );
  XOR U12717 ( .A(n11804), .B(n11805), .Z(n9834) );
  XOR U12718 ( .A(n11806), .B(n8396), .Z(n5115) );
  XOR U12719 ( .A(n11807), .B(n10082), .Z(n8396) );
  NOR U12720 ( .A(n9742), .B(n9741), .Z(n11806) );
  XOR U12721 ( .A(n11808), .B(n11809), .Z(n9741) );
  XNOR U12722 ( .A(n11811), .B(n8651), .Z(n3774) );
  XNOR U12723 ( .A(n11812), .B(n10316), .Z(n8651) );
  NOR U12724 ( .A(n9749), .B(n9750), .Z(n11811) );
  XOR U12725 ( .A(n11501), .B(n11813), .Z(n9750) );
  XOR U12726 ( .A(n11814), .B(n11815), .Z(n9749) );
  XOR U12727 ( .A(n11816), .B(n11817), .Z(n6223) );
  XNOR U12728 ( .A(n3202), .B(n7973), .Z(n11817) );
  XNOR U12729 ( .A(n11818), .B(n9708), .Z(n7973) );
  XOR U12730 ( .A(n11819), .B(n9864), .Z(n9708) );
  ANDN U12731 ( .B(n9733), .A(n9734), .Z(n11818) );
  XNOR U12732 ( .A(n11821), .B(n9524), .Z(n9733) );
  XNOR U12733 ( .A(n11822), .B(n9705), .Z(n3202) );
  XNOR U12734 ( .A(n11711), .B(n11823), .Z(n9705) );
  XNOR U12735 ( .A(n11824), .B(n11825), .Z(n9722) );
  XOR U12736 ( .A(n11826), .B(n9645), .Z(n9721) );
  XNOR U12737 ( .A(n11827), .B(n11828), .Z(n9645) );
  XOR U12738 ( .A(n5522), .B(n11829), .Z(n11816) );
  XOR U12739 ( .A(n8340), .B(n2390), .Z(n11829) );
  XNOR U12740 ( .A(n11830), .B(n9695), .Z(n2390) );
  XNOR U12741 ( .A(n11831), .B(n9874), .Z(n9695) );
  IV U12742 ( .A(n11768), .Z(n9874) );
  XOR U12743 ( .A(n11832), .B(n11833), .Z(n11768) );
  ANDN U12744 ( .B(n10575), .A(n10708), .Z(n11830) );
  XOR U12745 ( .A(n11834), .B(n10065), .Z(n10708) );
  XOR U12746 ( .A(n11835), .B(n10094), .Z(n10575) );
  XNOR U12747 ( .A(n11836), .B(n11837), .Z(n10094) );
  XNOR U12748 ( .A(n11838), .B(n9699), .Z(n8340) );
  IV U12749 ( .A(n10578), .Z(n9699) );
  XNOR U12750 ( .A(n11839), .B(n9757), .Z(n10578) );
  ANDN U12751 ( .B(n9724), .A(n10719), .Z(n11838) );
  IV U12752 ( .A(n9725), .Z(n10719) );
  XOR U12753 ( .A(n11698), .B(n11840), .Z(n9725) );
  XNOR U12754 ( .A(n11841), .B(n11842), .Z(n9724) );
  XOR U12755 ( .A(n11843), .B(n10573), .Z(n5522) );
  XOR U12756 ( .A(n11445), .B(n11844), .Z(n10573) );
  NOR U12757 ( .A(n10717), .B(n9729), .Z(n11843) );
  XOR U12758 ( .A(n9530), .B(n11845), .Z(n9729) );
  IV U12759 ( .A(n9730), .Z(n10717) );
  XNOR U12760 ( .A(n11846), .B(n9939), .Z(n9730) );
  XOR U12761 ( .A(n7590), .B(n3217), .Z(n3671) );
  XOR U12762 ( .A(n10236), .B(n11032), .Z(n3217) );
  XNOR U12763 ( .A(n11849), .B(n11850), .Z(n11032) );
  XOR U12764 ( .A(n5440), .B(n3889), .Z(n11850) );
  XNOR U12765 ( .A(n11851), .B(n11157), .Z(n3889) );
  XOR U12766 ( .A(n11852), .B(n10346), .Z(n11157) );
  ANDN U12767 ( .B(n7602), .A(n7603), .Z(n11851) );
  XNOR U12768 ( .A(n11853), .B(n9466), .Z(n7603) );
  XOR U12769 ( .A(n11854), .B(n11855), .Z(n7602) );
  XNOR U12770 ( .A(n11856), .B(n10028), .Z(n5440) );
  XOR U12771 ( .A(n9131), .B(n11857), .Z(n10028) );
  XNOR U12772 ( .A(n11858), .B(n11859), .Z(n9131) );
  ANDN U12773 ( .B(n7598), .A(n7599), .Z(n11856) );
  XNOR U12774 ( .A(n9627), .B(n11860), .Z(n7599) );
  XOR U12775 ( .A(n11861), .B(n11862), .Z(n9627) );
  XOR U12776 ( .A(n11863), .B(n10195), .Z(n7598) );
  IV U12777 ( .A(n11205), .Z(n10195) );
  XOR U12778 ( .A(n11864), .B(n11865), .Z(n11205) );
  XNOR U12779 ( .A(n6251), .B(n11866), .Z(n11849) );
  XNOR U12780 ( .A(n2289), .B(n5126), .Z(n11866) );
  XNOR U12781 ( .A(n11867), .B(n10040), .Z(n5126) );
  XNOR U12782 ( .A(n11868), .B(n11869), .Z(n10040) );
  ANDN U12783 ( .B(n8656), .A(n10041), .Z(n11867) );
  XNOR U12784 ( .A(n11870), .B(n10077), .Z(n10041) );
  XNOR U12785 ( .A(n11871), .B(n9759), .Z(n8656) );
  XNOR U12786 ( .A(n11872), .B(n10032), .Z(n2289) );
  XOR U12787 ( .A(n11873), .B(n11874), .Z(n10032) );
  NOR U12788 ( .A(n10031), .B(n10464), .Z(n11872) );
  XOR U12789 ( .A(n11875), .B(n10037), .Z(n6251) );
  XOR U12790 ( .A(n11876), .B(n11877), .Z(n10037) );
  NOR U12791 ( .A(n7593), .B(n7592), .Z(n11875) );
  XNOR U12792 ( .A(n11878), .B(n11879), .Z(n7592) );
  XOR U12793 ( .A(n11880), .B(n10198), .Z(n7593) );
  XOR U12794 ( .A(n11881), .B(n11882), .Z(n10236) );
  XOR U12795 ( .A(n3452), .B(n5054), .Z(n11882) );
  XNOR U12796 ( .A(n11883), .B(n11178), .Z(n5054) );
  IV U12797 ( .A(n7639), .Z(n11178) );
  XOR U12798 ( .A(n11884), .B(n10103), .Z(n7639) );
  IV U12799 ( .A(n11885), .Z(n10103) );
  ANDN U12800 ( .B(n10140), .A(n7638), .Z(n11883) );
  XOR U12801 ( .A(n11886), .B(n10231), .Z(n7638) );
  XNOR U12802 ( .A(n11244), .B(n11887), .Z(n10140) );
  XNOR U12803 ( .A(n11888), .B(n11185), .Z(n3452) );
  IV U12804 ( .A(n8716), .Z(n11185) );
  XOR U12805 ( .A(n11889), .B(n9929), .Z(n8716) );
  ANDN U12806 ( .B(n10143), .A(n8715), .Z(n11888) );
  XOR U12807 ( .A(n11890), .B(n11891), .Z(n8715) );
  XNOR U12808 ( .A(n11892), .B(n9664), .Z(n10143) );
  XOR U12809 ( .A(n2393), .B(n11893), .Z(n11881) );
  XOR U12810 ( .A(n7631), .B(n3999), .Z(n11893) );
  XOR U12811 ( .A(n11894), .B(n7652), .Z(n3999) );
  XOR U12812 ( .A(n11895), .B(n9771), .Z(n7652) );
  NOR U12813 ( .A(n11307), .B(n7651), .Z(n11894) );
  XOR U12814 ( .A(n11896), .B(n9790), .Z(n7651) );
  IV U12815 ( .A(n10132), .Z(n11307) );
  XNOR U12816 ( .A(n11899), .B(n10609), .Z(n10132) );
  XOR U12817 ( .A(n11900), .B(n7648), .Z(n7631) );
  XOR U12818 ( .A(n11901), .B(n11902), .Z(n7648) );
  NOR U12819 ( .A(n7647), .B(n10135), .Z(n11900) );
  XNOR U12820 ( .A(n10159), .B(n11903), .Z(n10135) );
  IV U12821 ( .A(n11904), .Z(n10159) );
  XOR U12822 ( .A(n9119), .B(n11905), .Z(n7647) );
  XNOR U12823 ( .A(n11906), .B(n7643), .Z(n2393) );
  XNOR U12824 ( .A(n11907), .B(n11908), .Z(n7643) );
  NOR U12825 ( .A(n7644), .B(n11312), .Z(n11906) );
  XOR U12826 ( .A(n11909), .B(n10067), .Z(n11312) );
  XOR U12827 ( .A(n11910), .B(n11513), .Z(n7644) );
  IV U12828 ( .A(n11283), .Z(n11513) );
  XOR U12829 ( .A(n11911), .B(n10031), .Z(n7590) );
  XNOR U12830 ( .A(n9458), .B(n11912), .Z(n10031) );
  XNOR U12831 ( .A(n11913), .B(n11914), .Z(n9458) );
  ANDN U12832 ( .B(n10464), .A(n10465), .Z(n11911) );
  XOR U12833 ( .A(n11915), .B(n10741), .Z(n10465) );
  XNOR U12834 ( .A(n11916), .B(n9949), .Z(n10464) );
  XNOR U12835 ( .A(n11917), .B(n6190), .Z(out[1009]) );
  IV U12836 ( .A(n6823), .Z(n6190) );
  XNOR U12837 ( .A(n8548), .B(n2250), .Z(n6823) );
  XNOR U12838 ( .A(n6073), .B(n6149), .Z(n2250) );
  XNOR U12839 ( .A(n11918), .B(n11919), .Z(n6149) );
  XOR U12840 ( .A(n2286), .B(n5447), .Z(n11919) );
  XOR U12841 ( .A(n11920), .B(n7384), .Z(n5447) );
  XNOR U12842 ( .A(n9563), .B(n11921), .Z(n7384) );
  IV U12843 ( .A(n11922), .Z(n9563) );
  ANDN U12844 ( .B(n8559), .A(n7383), .Z(n11920) );
  XOR U12845 ( .A(n11923), .B(n9893), .Z(n7383) );
  XOR U12846 ( .A(n11924), .B(n11925), .Z(n8559) );
  XNOR U12847 ( .A(n11926), .B(n7388), .Z(n2286) );
  XOR U12848 ( .A(n11604), .B(n11927), .Z(n7388) );
  ANDN U12849 ( .B(n7387), .A(n8554), .Z(n11926) );
  XOR U12850 ( .A(n11928), .B(n11929), .Z(n8554) );
  XNOR U12851 ( .A(n11930), .B(n11931), .Z(n7387) );
  XNOR U12852 ( .A(n3141), .B(n11932), .Z(n11918) );
  XOR U12853 ( .A(n5903), .B(n7377), .Z(n11932) );
  XNOR U12854 ( .A(n11933), .B(n7393), .Z(n7377) );
  XOR U12855 ( .A(n11934), .B(n11124), .Z(n7393) );
  ANDN U12856 ( .B(n7392), .A(n8557), .Z(n11933) );
  XNOR U12857 ( .A(n11935), .B(n11043), .Z(n8557) );
  XNOR U12858 ( .A(n11936), .B(n11937), .Z(n7392) );
  XNOR U12859 ( .A(n11938), .B(n7397), .Z(n5903) );
  XNOR U12860 ( .A(n11939), .B(n11482), .Z(n7397) );
  ANDN U12861 ( .B(n11641), .A(n7396), .Z(n11938) );
  XOR U12862 ( .A(n11940), .B(n8462), .Z(n3141) );
  XOR U12863 ( .A(n11941), .B(n11942), .Z(n8462) );
  ANDN U12864 ( .B(n8550), .A(n7400), .Z(n11940) );
  XNOR U12865 ( .A(n11943), .B(n11196), .Z(n7400) );
  XOR U12866 ( .A(n9438), .B(n11944), .Z(n8550) );
  XOR U12867 ( .A(n11945), .B(n11946), .Z(n6073) );
  XOR U12868 ( .A(n5272), .B(n1912), .Z(n11946) );
  XNOR U12869 ( .A(n11947), .B(n8704), .Z(n1912) );
  ANDN U12870 ( .B(n7477), .A(n8536), .Z(n11947) );
  XNOR U12871 ( .A(n10816), .B(n11948), .Z(n8536) );
  XNOR U12872 ( .A(n11949), .B(n11950), .Z(n10816) );
  XOR U12873 ( .A(n11951), .B(n11952), .Z(n7477) );
  XNOR U12874 ( .A(n11953), .B(n8709), .Z(n5272) );
  NOR U12875 ( .A(n7469), .B(n8534), .Z(n11953) );
  XOR U12876 ( .A(n11954), .B(n11955), .Z(n8534) );
  XOR U12877 ( .A(n11956), .B(n10357), .Z(n7469) );
  XOR U12878 ( .A(n3704), .B(n11957), .Z(n11945) );
  XNOR U12879 ( .A(n8684), .B(n4182), .Z(n11957) );
  XOR U12880 ( .A(n11958), .B(n8711), .Z(n4182) );
  ANDN U12881 ( .B(n8544), .A(n7460), .Z(n11958) );
  XNOR U12882 ( .A(n11959), .B(n11960), .Z(n7460) );
  XNOR U12883 ( .A(n11961), .B(n9771), .Z(n8544) );
  XOR U12884 ( .A(n11962), .B(n11963), .Z(n9771) );
  XOR U12885 ( .A(n11964), .B(n8707), .Z(n8684) );
  ANDN U12886 ( .B(n7464), .A(n8539), .Z(n11964) );
  XOR U12887 ( .A(n10100), .B(n11965), .Z(n8539) );
  IV U12888 ( .A(n11111), .Z(n10100) );
  XOR U12889 ( .A(n11966), .B(n9650), .Z(n7464) );
  XNOR U12890 ( .A(n11967), .B(n11968), .Z(n3704) );
  ANDN U12891 ( .B(n8542), .A(n7473), .Z(n11967) );
  XOR U12892 ( .A(n11970), .B(n7396), .Z(n8548) );
  XOR U12893 ( .A(n11971), .B(n10396), .Z(n7396) );
  NOR U12894 ( .A(n8467), .B(n11641), .Z(n11970) );
  XOR U12895 ( .A(n11972), .B(n11973), .Z(n11641) );
  IV U12896 ( .A(n11642), .Z(n8467) );
  XOR U12897 ( .A(n11974), .B(n10761), .Z(n11642) );
  IV U12898 ( .A(n11952), .Z(n10761) );
  XOR U12899 ( .A(n11975), .B(n11976), .Z(n11952) );
  ANDN U12900 ( .B(n5670), .A(n5668), .Z(n11917) );
  XOR U12901 ( .A(n11977), .B(n1749), .Z(n5668) );
  XOR U12902 ( .A(n11978), .B(n11979), .Z(n9603) );
  XOR U12903 ( .A(n3490), .B(n5101), .Z(n11979) );
  XNOR U12904 ( .A(n11980), .B(n8409), .Z(n5101) );
  ANDN U12905 ( .B(n11981), .A(n11982), .Z(n11980) );
  XNOR U12906 ( .A(n11983), .B(n9716), .Z(n3490) );
  ANDN U12907 ( .B(n11676), .A(n9715), .Z(n11983) );
  XOR U12908 ( .A(n4282), .B(n11984), .Z(n11978) );
  XOR U12909 ( .A(n8398), .B(n2481), .Z(n11984) );
  XOR U12910 ( .A(n11985), .B(n8419), .Z(n2481) );
  ANDN U12911 ( .B(n8418), .A(n11986), .Z(n11985) );
  XOR U12912 ( .A(n11987), .B(n8404), .Z(n8398) );
  ANDN U12913 ( .B(n8405), .A(n11667), .Z(n11987) );
  XNOR U12914 ( .A(n11988), .B(n8414), .Z(n4282) );
  ANDN U12915 ( .B(n8415), .A(n11663), .Z(n11988) );
  XOR U12916 ( .A(n11989), .B(n11990), .Z(n6314) );
  XOR U12917 ( .A(n5438), .B(n3687), .Z(n11990) );
  XNOR U12918 ( .A(n11991), .B(n11992), .Z(n3687) );
  ANDN U12919 ( .B(n8498), .A(n11993), .Z(n11991) );
  XNOR U12920 ( .A(n11994), .B(n11995), .Z(n5438) );
  ANDN U12921 ( .B(n11996), .A(n8488), .Z(n11994) );
  IV U12922 ( .A(n11997), .Z(n8488) );
  XNOR U12923 ( .A(n11998), .B(n11999), .Z(n11989) );
  XNOR U12924 ( .A(n2100), .B(n4319), .Z(n11999) );
  XOR U12925 ( .A(n12000), .B(n12001), .Z(n4319) );
  NOR U12926 ( .A(n12002), .B(n8492), .Z(n12000) );
  XOR U12927 ( .A(n12003), .B(n12004), .Z(n2100) );
  ANDN U12928 ( .B(n12005), .A(n12006), .Z(n12003) );
  XOR U12929 ( .A(n10663), .B(n2069), .Z(n5670) );
  XNOR U12930 ( .A(n7867), .B(n9034), .Z(n2069) );
  XNOR U12931 ( .A(n12007), .B(n12008), .Z(n9034) );
  XOR U12932 ( .A(n5470), .B(n3916), .Z(n12008) );
  XNOR U12933 ( .A(n12009), .B(n12010), .Z(n3916) );
  NOR U12934 ( .A(n12011), .B(n8042), .Z(n12009) );
  XNOR U12935 ( .A(n12012), .B(n12013), .Z(n8042) );
  XNOR U12936 ( .A(n12014), .B(n12015), .Z(n5470) );
  ANDN U12937 ( .B(n8037), .A(n8038), .Z(n12014) );
  XOR U12938 ( .A(n12016), .B(n10193), .Z(n8038) );
  XNOR U12939 ( .A(n12017), .B(n12018), .Z(n8037) );
  XOR U12940 ( .A(n6279), .B(n12019), .Z(n12007) );
  XNOR U12941 ( .A(n2335), .B(n5313), .Z(n12019) );
  XNOR U12942 ( .A(n12020), .B(n10799), .Z(n5313) );
  ANDN U12943 ( .B(n9039), .A(n10800), .Z(n12020) );
  XOR U12944 ( .A(n9119), .B(n12021), .Z(n10800) );
  XOR U12945 ( .A(n12023), .B(n12024), .Z(n11862) );
  XNOR U12946 ( .A(n10087), .B(n11120), .Z(n12024) );
  XNOR U12947 ( .A(n12025), .B(n12026), .Z(n11120) );
  ANDN U12948 ( .B(n12027), .A(n12028), .Z(n12025) );
  XNOR U12949 ( .A(n12029), .B(n12030), .Z(n10087) );
  ANDN U12950 ( .B(n12031), .A(n12032), .Z(n12029) );
  XOR U12951 ( .A(n10925), .B(n12033), .Z(n12023) );
  XOR U12952 ( .A(n10954), .B(n11077), .Z(n12033) );
  XNOR U12953 ( .A(n12034), .B(n12035), .Z(n11077) );
  NOR U12954 ( .A(n12036), .B(n12037), .Z(n12034) );
  XOR U12955 ( .A(n12038), .B(n12039), .Z(n10954) );
  ANDN U12956 ( .B(n12040), .A(n12041), .Z(n12038) );
  XNOR U12957 ( .A(n12042), .B(n12043), .Z(n10925) );
  NOR U12958 ( .A(n12044), .B(n12045), .Z(n12042) );
  XOR U12959 ( .A(n10317), .B(n12046), .Z(n9039) );
  XOR U12960 ( .A(n12047), .B(n12048), .Z(n2335) );
  NOR U12961 ( .A(n10791), .B(n8028), .Z(n12047) );
  XOR U12962 ( .A(n12049), .B(n9322), .Z(n8028) );
  XNOR U12963 ( .A(n12050), .B(n11754), .Z(n10791) );
  XNOR U12964 ( .A(n12051), .B(n10796), .Z(n6279) );
  ANDN U12965 ( .B(n8031), .A(n8033), .Z(n12051) );
  XNOR U12966 ( .A(n12052), .B(n11595), .Z(n8033) );
  XOR U12967 ( .A(n10082), .B(n12053), .Z(n8031) );
  XOR U12968 ( .A(n12054), .B(n12055), .Z(n7867) );
  XNOR U12969 ( .A(n3813), .B(n5143), .Z(n12055) );
  XNOR U12970 ( .A(n12056), .B(n8977), .Z(n5143) );
  XOR U12971 ( .A(n12057), .B(n11103), .Z(n8977) );
  NOR U12972 ( .A(n10670), .B(n10669), .Z(n12056) );
  XNOR U12973 ( .A(n12058), .B(n11754), .Z(n10669) );
  XOR U12974 ( .A(n10163), .B(n12059), .Z(n10670) );
  XOR U12975 ( .A(n12060), .B(n7943), .Z(n3813) );
  XNOR U12976 ( .A(n9544), .B(n12061), .Z(n7943) );
  NOR U12977 ( .A(n10661), .B(n10662), .Z(n12060) );
  XOR U12978 ( .A(n10703), .B(n12062), .Z(n10662) );
  IV U12979 ( .A(n9236), .Z(n10703) );
  XNOR U12980 ( .A(n9414), .B(n12063), .Z(n10661) );
  XOR U12981 ( .A(n4259), .B(n12064), .Z(n12054) );
  XNOR U12982 ( .A(n1707), .B(n10782), .Z(n12064) );
  XOR U12983 ( .A(n12065), .B(n7952), .Z(n10782) );
  XNOR U12984 ( .A(n12066), .B(n11885), .Z(n7952) );
  XOR U12985 ( .A(n12067), .B(n12068), .Z(n11885) );
  ANDN U12986 ( .B(n10657), .A(n10658), .Z(n12065) );
  XOR U12987 ( .A(n11280), .B(n12069), .Z(n10658) );
  XOR U12988 ( .A(n12070), .B(n11511), .Z(n10657) );
  XNOR U12989 ( .A(n12071), .B(n7947), .Z(n1707) );
  XOR U12990 ( .A(n12072), .B(n10307), .Z(n7947) );
  ANDN U12991 ( .B(n10666), .A(n10667), .Z(n12071) );
  XOR U12992 ( .A(n12073), .B(n11842), .Z(n10667) );
  XOR U12993 ( .A(n11972), .B(n12074), .Z(n10666) );
  XOR U12994 ( .A(n12075), .B(n7957), .Z(n4259) );
  XOR U12995 ( .A(n11758), .B(n12076), .Z(n7957) );
  ANDN U12996 ( .B(n11682), .A(n10807), .Z(n12075) );
  XNOR U12997 ( .A(n12077), .B(n10807), .Z(n10663) );
  XOR U12998 ( .A(n9143), .B(n12078), .Z(n10807) );
  IV U12999 ( .A(n11711), .Z(n9143) );
  ANDN U13000 ( .B(n7955), .A(n11682), .Z(n12077) );
  XOR U13001 ( .A(n12079), .B(n10985), .Z(n11682) );
  XNOR U13002 ( .A(n10958), .B(n12080), .Z(n7955) );
  XNOR U13003 ( .A(n12081), .B(n6195), .Z(out[1008]) );
  IV U13004 ( .A(n6851), .Z(n6195) );
  XNOR U13005 ( .A(n8701), .B(n2257), .Z(n6851) );
  XNOR U13006 ( .A(n6078), .B(n6154), .Z(n2257) );
  XNOR U13007 ( .A(n12082), .B(n12083), .Z(n6154) );
  XNOR U13008 ( .A(n2293), .B(n5453), .Z(n12083) );
  XNOR U13009 ( .A(n12084), .B(n8545), .Z(n5453) );
  IV U13010 ( .A(n7461), .Z(n8545) );
  XOR U13011 ( .A(n10869), .B(n12085), .Z(n7461) );
  ANDN U13012 ( .B(n7462), .A(n8711), .Z(n12084) );
  XNOR U13013 ( .A(n12086), .B(n9450), .Z(n8711) );
  XNOR U13014 ( .A(n12087), .B(n9959), .Z(n7462) );
  XNOR U13015 ( .A(n12088), .B(n8540), .Z(n2293) );
  IV U13016 ( .A(n7466), .Z(n8540) );
  XOR U13017 ( .A(n12089), .B(n12090), .Z(n7466) );
  ANDN U13018 ( .B(n8707), .A(n7465), .Z(n12088) );
  XOR U13019 ( .A(n12091), .B(n9552), .Z(n7465) );
  XNOR U13020 ( .A(n12092), .B(n12093), .Z(n8707) );
  XOR U13021 ( .A(n3150), .B(n12094), .Z(n12082) );
  XOR U13022 ( .A(n5957), .B(n7455), .Z(n12094) );
  XNOR U13023 ( .A(n12095), .B(n7470), .Z(n7455) );
  XOR U13024 ( .A(n12096), .B(n12097), .Z(n7470) );
  AND U13025 ( .A(n8709), .B(n7471), .Z(n12095) );
  XNOR U13026 ( .A(n12098), .B(n12099), .Z(n7471) );
  XOR U13027 ( .A(n12100), .B(n10067), .Z(n8709) );
  XNOR U13028 ( .A(n12101), .B(n7475), .Z(n5957) );
  XNOR U13029 ( .A(n12102), .B(n12103), .Z(n7475) );
  ANDN U13030 ( .B(n11968), .A(n7474), .Z(n12101) );
  XNOR U13031 ( .A(n12104), .B(n7478), .Z(n3150) );
  XOR U13032 ( .A(n12105), .B(n10763), .Z(n7478) );
  ANDN U13033 ( .B(n8704), .A(n8703), .Z(n12104) );
  IV U13034 ( .A(n7479), .Z(n8703) );
  XOR U13035 ( .A(n12106), .B(n12107), .Z(n7479) );
  XOR U13036 ( .A(n10313), .B(n12108), .Z(n8704) );
  XOR U13037 ( .A(n12109), .B(n12110), .Z(n6078) );
  XNOR U13038 ( .A(n5274), .B(n1920), .Z(n12110) );
  XNOR U13039 ( .A(n12111), .B(n8739), .Z(n1920) );
  ANDN U13040 ( .B(n7551), .A(n8690), .Z(n12111) );
  IV U13041 ( .A(n8738), .Z(n8690) );
  XOR U13042 ( .A(n12112), .B(n11448), .Z(n8738) );
  XOR U13043 ( .A(n12113), .B(n11686), .Z(n7551) );
  IV U13044 ( .A(n12114), .Z(n11686) );
  XNOR U13045 ( .A(n12115), .B(n8744), .Z(n5274) );
  ANDN U13046 ( .B(n7543), .A(n8688), .Z(n12115) );
  XNOR U13047 ( .A(n12116), .B(n12117), .Z(n8688) );
  XNOR U13048 ( .A(n11584), .B(n12118), .Z(n7543) );
  XOR U13049 ( .A(n3709), .B(n12119), .Z(n12109) );
  XNOR U13050 ( .A(n8719), .B(n4185), .Z(n12119) );
  XOR U13051 ( .A(n12120), .B(n8746), .Z(n4185) );
  ANDN U13052 ( .B(n8697), .A(n7534), .Z(n12120) );
  XOR U13053 ( .A(n12121), .B(n12122), .Z(n7534) );
  XOR U13054 ( .A(n12123), .B(n9872), .Z(n8697) );
  XNOR U13055 ( .A(n12126), .B(n8742), .Z(n8719) );
  ANDN U13056 ( .B(n7538), .A(n8693), .Z(n12126) );
  XOR U13057 ( .A(n9132), .B(n12127), .Z(n8693) );
  IV U13058 ( .A(n12128), .Z(n9132) );
  XOR U13059 ( .A(n12129), .B(n9793), .Z(n7538) );
  XOR U13060 ( .A(n12130), .B(n12131), .Z(n3709) );
  ANDN U13061 ( .B(n7547), .A(n8695), .Z(n12130) );
  XOR U13062 ( .A(n9940), .B(n12132), .Z(n7547) );
  XOR U13063 ( .A(n12133), .B(n7474), .Z(n8701) );
  XNOR U13064 ( .A(n12134), .B(n10599), .Z(n7474) );
  IV U13065 ( .A(n11460), .Z(n10599) );
  NOR U13066 ( .A(n11968), .B(n8542), .Z(n12133) );
  XNOR U13067 ( .A(n12135), .B(n12114), .Z(n8542) );
  XNOR U13068 ( .A(n12136), .B(n12137), .Z(n12114) );
  XNOR U13069 ( .A(n9113), .B(n12138), .Z(n11968) );
  NOR U13070 ( .A(n5673), .B(n5672), .Z(n12081) );
  XNOR U13071 ( .A(n12139), .B(n1754), .Z(n5672) );
  XOR U13072 ( .A(n6318), .B(n9711), .Z(n1754) );
  XOR U13073 ( .A(n12140), .B(n12141), .Z(n9711) );
  XNOR U13074 ( .A(n3497), .B(n4863), .Z(n12141) );
  XNOR U13075 ( .A(n12142), .B(n8493), .Z(n4863) );
  ANDN U13076 ( .B(n8494), .A(n12001), .Z(n12142) );
  XNOR U13077 ( .A(n12143), .B(n9824), .Z(n3497) );
  NOR U13078 ( .A(n12144), .B(n12004), .Z(n12143) );
  XOR U13079 ( .A(n4311), .B(n12145), .Z(n12140) );
  XNOR U13080 ( .A(n8484), .B(n2488), .Z(n12145) );
  XNOR U13081 ( .A(n12146), .B(n8504), .Z(n2488) );
  ANDN U13082 ( .B(n8503), .A(n12147), .Z(n12146) );
  XOR U13083 ( .A(n12148), .B(n8490), .Z(n8484) );
  XOR U13084 ( .A(n12149), .B(n8499), .Z(n4311) );
  ANDN U13085 ( .B(n8500), .A(n12150), .Z(n12149) );
  XNOR U13086 ( .A(n12151), .B(n12152), .Z(n6318) );
  XOR U13087 ( .A(n5442), .B(n3691), .Z(n12152) );
  XOR U13088 ( .A(n12153), .B(n12154), .Z(n3691) );
  NOR U13089 ( .A(n12155), .B(n8573), .Z(n12153) );
  XNOR U13090 ( .A(n12156), .B(n8513), .Z(n5442) );
  NOR U13091 ( .A(n12157), .B(n8564), .Z(n12156) );
  XNOR U13092 ( .A(n4321), .B(n12158), .Z(n12151) );
  XNOR U13093 ( .A(n5890), .B(n2105), .Z(n12158) );
  XNOR U13094 ( .A(n12159), .B(n8510), .Z(n2105) );
  IV U13095 ( .A(n12160), .Z(n8510) );
  NOR U13096 ( .A(n9918), .B(n8509), .Z(n12159) );
  IV U13097 ( .A(n12161), .Z(n9918) );
  XOR U13098 ( .A(n12162), .B(n8523), .Z(n5890) );
  NOR U13099 ( .A(n8577), .B(n8524), .Z(n12162) );
  XNOR U13100 ( .A(n12163), .B(n8520), .Z(n4321) );
  XOR U13101 ( .A(n10792), .B(n2072), .Z(n5673) );
  XNOR U13102 ( .A(n7937), .B(n9091), .Z(n2072) );
  XNOR U13103 ( .A(n12164), .B(n12165), .Z(n9091) );
  XNOR U13104 ( .A(n5477), .B(n3605), .Z(n12165) );
  XOR U13105 ( .A(n12166), .B(n12167), .Z(n3605) );
  ANDN U13106 ( .B(n8092), .A(n8093), .Z(n12166) );
  XOR U13107 ( .A(n12168), .B(n12169), .Z(n8093) );
  XOR U13108 ( .A(n12170), .B(n10892), .Z(n5477) );
  ANDN U13109 ( .B(n8089), .A(n10893), .Z(n12170) );
  XOR U13110 ( .A(n11109), .B(n12171), .Z(n10893) );
  XOR U13111 ( .A(n12172), .B(n10331), .Z(n8089) );
  XOR U13112 ( .A(n6283), .B(n12173), .Z(n12164) );
  XOR U13113 ( .A(n2342), .B(n5365), .Z(n12173) );
  XOR U13114 ( .A(n12174), .B(n12175), .Z(n5365) );
  ANDN U13115 ( .B(n9095), .A(n9093), .Z(n12174) );
  IV U13116 ( .A(n10906), .Z(n9093) );
  XOR U13117 ( .A(n12176), .B(n11210), .Z(n10906) );
  XOR U13118 ( .A(n12177), .B(n10626), .Z(n9095) );
  XOR U13119 ( .A(n12178), .B(n10896), .Z(n2342) );
  ANDN U13120 ( .B(n8078), .A(n11030), .Z(n12178) );
  XNOR U13121 ( .A(n12179), .B(n10749), .Z(n11030) );
  XOR U13122 ( .A(n12180), .B(n10122), .Z(n8078) );
  XNOR U13123 ( .A(n12181), .B(n10901), .Z(n6283) );
  ANDN U13124 ( .B(n8084), .A(n8082), .Z(n12181) );
  IV U13125 ( .A(n10902), .Z(n8082) );
  XOR U13126 ( .A(n12182), .B(n12183), .Z(n10902) );
  XNOR U13127 ( .A(n12184), .B(n10868), .Z(n8084) );
  XOR U13128 ( .A(n12185), .B(n12186), .Z(n7937) );
  XNOR U13129 ( .A(n3817), .B(n5145), .Z(n12186) );
  XOR U13130 ( .A(n9124), .B(n12188), .Z(n9038) );
  IV U13131 ( .A(n11228), .Z(n9124) );
  NOR U13132 ( .A(n10798), .B(n10799), .Z(n12187) );
  XNOR U13133 ( .A(n12189), .B(n10269), .Z(n10799) );
  XOR U13134 ( .A(n12190), .B(n11101), .Z(n10798) );
  XNOR U13135 ( .A(n12191), .B(n8029), .Z(n3817) );
  IV U13136 ( .A(n10915), .Z(n8029) );
  XOR U13137 ( .A(n12192), .B(n9650), .Z(n10915) );
  ANDN U13138 ( .B(n10789), .A(n10790), .Z(n12191) );
  IV U13139 ( .A(n12048), .Z(n10790) );
  XOR U13140 ( .A(n12193), .B(n10833), .Z(n12048) );
  XNOR U13141 ( .A(n12194), .B(n9511), .Z(n10789) );
  XOR U13142 ( .A(n4283), .B(n12195), .Z(n12185) );
  XNOR U13143 ( .A(n1712), .B(n10887), .Z(n12195) );
  XOR U13144 ( .A(n12196), .B(n8039), .Z(n10887) );
  XNOR U13145 ( .A(n11294), .B(n12197), .Z(n8039) );
  ANDN U13146 ( .B(n10787), .A(n10786), .Z(n12196) );
  IV U13147 ( .A(n10917), .Z(n10786) );
  XOR U13148 ( .A(n12198), .B(n11855), .Z(n10917) );
  IV U13149 ( .A(n12015), .Z(n10787) );
  XNOR U13150 ( .A(n12199), .B(n9817), .Z(n12015) );
  XNOR U13151 ( .A(n12200), .B(n8032), .Z(n1712) );
  XNOR U13152 ( .A(n12201), .B(n10406), .Z(n8032) );
  AND U13153 ( .A(n10796), .B(n10795), .Z(n12200) );
  XOR U13154 ( .A(n9113), .B(n12202), .Z(n10795) );
  XNOR U13155 ( .A(n9414), .B(n12203), .Z(n10796) );
  XOR U13156 ( .A(n12204), .B(n12205), .Z(n9414) );
  XOR U13157 ( .A(n12206), .B(n8043), .Z(n4283) );
  XOR U13158 ( .A(n11109), .B(n12207), .Z(n8043) );
  ANDN U13159 ( .B(n10913), .A(n12010), .Z(n12206) );
  IV U13160 ( .A(n12208), .Z(n10913) );
  XOR U13161 ( .A(n12209), .B(n12208), .Z(n10792) );
  XOR U13162 ( .A(n9236), .B(n12210), .Z(n12208) );
  ANDN U13163 ( .B(n12010), .A(n8041), .Z(n12209) );
  IV U13164 ( .A(n12011), .Z(n8041) );
  XOR U13165 ( .A(n12211), .B(n11039), .Z(n12011) );
  XOR U13166 ( .A(n12212), .B(n11085), .Z(n12010) );
  XNOR U13167 ( .A(n12213), .B(n6200), .Z(out[1007]) );
  IV U13168 ( .A(n6878), .Z(n6200) );
  XNOR U13169 ( .A(n8735), .B(n2266), .Z(n6878) );
  XNOR U13170 ( .A(n6083), .B(n6159), .Z(n2266) );
  XNOR U13171 ( .A(n12214), .B(n12215), .Z(n6159) );
  XNOR U13172 ( .A(n2300), .B(n5457), .Z(n12215) );
  XNOR U13173 ( .A(n12216), .B(n8698), .Z(n5457) );
  IV U13174 ( .A(n7535), .Z(n8698) );
  XOR U13175 ( .A(n12217), .B(n11825), .Z(n7535) );
  ANDN U13176 ( .B(n7536), .A(n8746), .Z(n12216) );
  XNOR U13177 ( .A(n12218), .B(n9547), .Z(n8746) );
  XOR U13178 ( .A(n12219), .B(n12220), .Z(n7536) );
  XNOR U13179 ( .A(n12221), .B(n7540), .Z(n2300) );
  XNOR U13180 ( .A(n12222), .B(n9450), .Z(n7540) );
  NOR U13181 ( .A(n7539), .B(n8742), .Z(n12221) );
  XNOR U13182 ( .A(n12223), .B(n10990), .Z(n8742) );
  XNOR U13183 ( .A(n12224), .B(n9808), .Z(n7539) );
  XOR U13184 ( .A(n3153), .B(n12225), .Z(n12214) );
  XOR U13185 ( .A(n6014), .B(n7529), .Z(n12225) );
  XNOR U13186 ( .A(n12226), .B(n7544), .Z(n7529) );
  XNOR U13187 ( .A(n12227), .B(n11369), .Z(n7544) );
  ANDN U13188 ( .B(n8744), .A(n7545), .Z(n12226) );
  XOR U13189 ( .A(n12228), .B(n10287), .Z(n7545) );
  XOR U13190 ( .A(n11303), .B(n12229), .Z(n8744) );
  XNOR U13191 ( .A(n12230), .B(n7548), .Z(n6014) );
  XOR U13192 ( .A(n12231), .B(n12232), .Z(n7548) );
  ANDN U13193 ( .B(n7549), .A(n12131), .Z(n12230) );
  XNOR U13194 ( .A(n12233), .B(n7552), .Z(n3153) );
  XOR U13195 ( .A(n12234), .B(n10305), .Z(n7552) );
  ANDN U13196 ( .B(n8739), .A(n8737), .Z(n12233) );
  IV U13197 ( .A(n7553), .Z(n8737) );
  XOR U13198 ( .A(n12235), .B(n12236), .Z(n7553) );
  XOR U13199 ( .A(n12237), .B(n11081), .Z(n8739) );
  XOR U13200 ( .A(n12238), .B(n12239), .Z(n6083) );
  XNOR U13201 ( .A(n5276), .B(n1924), .Z(n12239) );
  XNOR U13202 ( .A(n12240), .B(n8833), .Z(n1924) );
  ANDN U13203 ( .B(n8725), .A(n7628), .Z(n12240) );
  XOR U13204 ( .A(n12017), .B(n12241), .Z(n7628) );
  XOR U13205 ( .A(n12242), .B(n9937), .Z(n8725) );
  IV U13206 ( .A(n9466), .Z(n9937) );
  XOR U13207 ( .A(n12243), .B(n12244), .Z(n9466) );
  XNOR U13208 ( .A(n12245), .B(n8839), .Z(n5276) );
  NOR U13209 ( .A(n8723), .B(n7620), .Z(n12245) );
  XNOR U13210 ( .A(n12246), .B(n10172), .Z(n7620) );
  XOR U13211 ( .A(n12247), .B(n12248), .Z(n8723) );
  XNOR U13212 ( .A(n3715), .B(n12249), .Z(n12238) );
  XNOR U13213 ( .A(n8813), .B(n4188), .Z(n12249) );
  XNOR U13214 ( .A(n12250), .B(n8841), .Z(n4188) );
  NOR U13215 ( .A(n7611), .B(n8732), .Z(n12250) );
  XOR U13216 ( .A(n9940), .B(n12251), .Z(n8732) );
  IV U13217 ( .A(n11415), .Z(n9940) );
  XNOR U13218 ( .A(n12252), .B(n12253), .Z(n11415) );
  XOR U13219 ( .A(n12254), .B(n12255), .Z(n7611) );
  XOR U13220 ( .A(n12256), .B(n8836), .Z(n8813) );
  NOR U13221 ( .A(n8837), .B(n7615), .Z(n12256) );
  XNOR U13222 ( .A(n12257), .B(n9893), .Z(n7615) );
  XOR U13223 ( .A(n12258), .B(n9277), .Z(n8837) );
  XOR U13224 ( .A(n12259), .B(n12260), .Z(n3715) );
  ANDN U13225 ( .B(n7624), .A(n8730), .Z(n12259) );
  XOR U13226 ( .A(n11092), .B(n12261), .Z(n7624) );
  XOR U13227 ( .A(n12262), .B(n7549), .Z(n8735) );
  XOR U13228 ( .A(n12263), .B(n10724), .Z(n7549) );
  XOR U13229 ( .A(n11758), .B(n12264), .Z(n8695) );
  IV U13230 ( .A(n12017), .Z(n11758) );
  XNOR U13231 ( .A(n12265), .B(n12266), .Z(n12017) );
  XOR U13232 ( .A(n12267), .B(n9274), .Z(n12131) );
  ANDN U13233 ( .B(n5678), .A(n5676), .Z(n12213) );
  XNOR U13234 ( .A(n8516), .B(n3862), .Z(n5676) );
  IV U13235 ( .A(n1758), .Z(n3862) );
  XOR U13236 ( .A(n12268), .B(n12269), .Z(n9819) );
  XOR U13237 ( .A(n3499), .B(n4867), .Z(n12269) );
  XNOR U13238 ( .A(n12270), .B(n8568), .Z(n4867) );
  ANDN U13239 ( .B(n8520), .A(n8569), .Z(n12270) );
  XNOR U13240 ( .A(n12271), .B(n10724), .Z(n8569) );
  XOR U13241 ( .A(n12272), .B(n9858), .Z(n8520) );
  IV U13242 ( .A(n10695), .Z(n9858) );
  XOR U13243 ( .A(n12273), .B(n12274), .Z(n3499) );
  ANDN U13244 ( .B(n8508), .A(n12160), .Z(n12273) );
  XOR U13245 ( .A(n12275), .B(n11196), .Z(n12160) );
  XNOR U13246 ( .A(n9966), .B(n12276), .Z(n8508) );
  XNOR U13247 ( .A(n4340), .B(n12277), .Z(n12268) );
  XOR U13248 ( .A(n8560), .B(n2493), .Z(n12277) );
  XOR U13249 ( .A(n12278), .B(n8578), .Z(n2493) );
  ANDN U13250 ( .B(n8522), .A(n8523), .Z(n12278) );
  XNOR U13251 ( .A(n10082), .B(n12279), .Z(n8523) );
  IV U13252 ( .A(n12280), .Z(n10082) );
  XOR U13253 ( .A(n12281), .B(n10402), .Z(n8522) );
  IV U13254 ( .A(n12282), .Z(n10402) );
  XOR U13255 ( .A(n12283), .B(n8565), .Z(n8560) );
  ANDN U13256 ( .B(n8512), .A(n8513), .Z(n12283) );
  XNOR U13257 ( .A(n12284), .B(n10626), .Z(n8513) );
  IV U13258 ( .A(n10503), .Z(n10626) );
  XOR U13259 ( .A(n12285), .B(n10637), .Z(n8512) );
  XOR U13260 ( .A(n12286), .B(n8575), .Z(n4340) );
  ANDN U13261 ( .B(n8574), .A(n12154), .Z(n12286) );
  XOR U13262 ( .A(n12287), .B(n12288), .Z(n6326) );
  XOR U13263 ( .A(n5446), .B(n3697), .Z(n12288) );
  XNOR U13264 ( .A(n12289), .B(n12290), .Z(n3697) );
  AND U13265 ( .A(n6438), .B(n6437), .Z(n12289) );
  XOR U13266 ( .A(n12291), .B(n12282), .Z(n6438) );
  XNOR U13267 ( .A(n12292), .B(n8586), .Z(n5446) );
  ANDN U13268 ( .B(n6429), .A(n8587), .Z(n12292) );
  XOR U13269 ( .A(n12293), .B(n10324), .Z(n8587) );
  XNOR U13270 ( .A(n12294), .B(n11196), .Z(n6429) );
  XOR U13271 ( .A(n4324), .B(n12295), .Z(n12287) );
  XNOR U13272 ( .A(n5895), .B(n2109), .Z(n12295) );
  XNOR U13273 ( .A(n12296), .B(n8583), .Z(n2109) );
  ANDN U13274 ( .B(n6442), .A(n6441), .Z(n12296) );
  XOR U13275 ( .A(n9659), .B(n12297), .Z(n6441) );
  XOR U13276 ( .A(n12298), .B(n12299), .Z(n6442) );
  XNOR U13277 ( .A(n12300), .B(n12301), .Z(n5895) );
  ANDN U13278 ( .B(n6445), .A(n6446), .Z(n12300) );
  XOR U13279 ( .A(n9639), .B(n12302), .Z(n6446) );
  XOR U13280 ( .A(n12303), .B(n9142), .Z(n6445) );
  XNOR U13281 ( .A(n12304), .B(n8592), .Z(n4324) );
  ANDN U13282 ( .B(n6434), .A(n6432), .Z(n12304) );
  IV U13283 ( .A(n8593), .Z(n6432) );
  XOR U13284 ( .A(n12305), .B(n10503), .Z(n8593) );
  XOR U13285 ( .A(n12306), .B(n12307), .Z(n10503) );
  XOR U13286 ( .A(n9107), .B(n12308), .Z(n6434) );
  XNOR U13287 ( .A(n12309), .B(n8574), .Z(n8516) );
  XOR U13288 ( .A(n12311), .B(n12312), .Z(n12154) );
  XNOR U13289 ( .A(n10897), .B(n2079), .Z(n5678) );
  XNOR U13290 ( .A(n8023), .B(n9184), .Z(n2079) );
  XNOR U13291 ( .A(n12313), .B(n12314), .Z(n9184) );
  XNOR U13292 ( .A(n5482), .B(n3610), .Z(n12314) );
  XOR U13293 ( .A(n12315), .B(n12316), .Z(n3610) );
  ANDN U13294 ( .B(n8174), .A(n8175), .Z(n12315) );
  XOR U13295 ( .A(n12317), .B(n10234), .Z(n8175) );
  XOR U13296 ( .A(n12318), .B(n12319), .Z(n5482) );
  NOR U13297 ( .A(n8170), .B(n8171), .Z(n12318) );
  XOR U13298 ( .A(n12320), .B(n10512), .Z(n8171) );
  IV U13299 ( .A(n11007), .Z(n8170) );
  XNOR U13300 ( .A(n12321), .B(n11235), .Z(n11007) );
  XNOR U13301 ( .A(n6287), .B(n12322), .Z(n12313) );
  XOR U13302 ( .A(n2349), .B(n5411), .Z(n12322) );
  XNOR U13303 ( .A(n12323), .B(n11019), .Z(n5411) );
  ANDN U13304 ( .B(n9188), .A(n11020), .Z(n12323) );
  XOR U13305 ( .A(n12324), .B(n11116), .Z(n11020) );
  IV U13306 ( .A(n12325), .Z(n11116) );
  XNOR U13307 ( .A(n12326), .B(n12327), .Z(n9188) );
  XNOR U13308 ( .A(n12328), .B(n11010), .Z(n2349) );
  ANDN U13309 ( .B(n8160), .A(n8161), .Z(n12328) );
  XNOR U13310 ( .A(n12329), .B(n12330), .Z(n8161) );
  XOR U13311 ( .A(n12331), .B(n10221), .Z(n8160) );
  XOR U13312 ( .A(n12332), .B(n12333), .Z(n6287) );
  NOR U13313 ( .A(n8164), .B(n8165), .Z(n12332) );
  XNOR U13314 ( .A(n12334), .B(n10985), .Z(n8165) );
  IV U13315 ( .A(n11016), .Z(n8164) );
  XNOR U13316 ( .A(n12335), .B(n10324), .Z(n11016) );
  XOR U13317 ( .A(n12336), .B(n12337), .Z(n8023) );
  XOR U13318 ( .A(n3826), .B(n5147), .Z(n12337) );
  XNOR U13319 ( .A(n12338), .B(n9094), .Z(n5147) );
  XOR U13320 ( .A(n9107), .B(n12339), .Z(n9094) );
  ANDN U13321 ( .B(n10904), .A(n10905), .Z(n12338) );
  IV U13322 ( .A(n12175), .Z(n10905) );
  XOR U13323 ( .A(n12340), .B(n9431), .Z(n12175) );
  XOR U13324 ( .A(n12341), .B(n10221), .Z(n10904) );
  XNOR U13325 ( .A(n11858), .B(n12342), .Z(n10221) );
  XOR U13326 ( .A(n12343), .B(n12344), .Z(n11858) );
  XNOR U13327 ( .A(n12345), .B(n10520), .Z(n12344) );
  XOR U13328 ( .A(n12346), .B(n12347), .Z(n10520) );
  ANDN U13329 ( .B(n12348), .A(n12349), .Z(n12346) );
  XNOR U13330 ( .A(n11505), .B(n12350), .Z(n12343) );
  XNOR U13331 ( .A(n12351), .B(n12352), .Z(n12350) );
  XNOR U13332 ( .A(n12353), .B(n12354), .Z(n11505) );
  ANDN U13333 ( .B(n12355), .A(n12356), .Z(n12353) );
  XNOR U13334 ( .A(n12357), .B(n8080), .Z(n3826) );
  XOR U13335 ( .A(n12358), .B(n11603), .Z(n8080) );
  IV U13336 ( .A(n9793), .Z(n11603) );
  XOR U13337 ( .A(n12359), .B(n12360), .Z(n10896) );
  XNOR U13338 ( .A(n9614), .B(n12361), .Z(n10895) );
  IV U13339 ( .A(n9761), .Z(n9614) );
  XOR U13340 ( .A(n4312), .B(n12362), .Z(n12336) );
  XNOR U13341 ( .A(n1717), .B(n11001), .Z(n12362) );
  XNOR U13342 ( .A(n12363), .B(n8090), .Z(n11001) );
  XNOR U13343 ( .A(n12364), .B(n10346), .Z(n8090) );
  XNOR U13344 ( .A(n12365), .B(n12366), .Z(n10346) );
  ANDN U13345 ( .B(n10891), .A(n10892), .Z(n12363) );
  XOR U13346 ( .A(n12367), .B(n9912), .Z(n10892) );
  XOR U13347 ( .A(n12368), .B(n12369), .Z(n10891) );
  XNOR U13348 ( .A(n12370), .B(n8083), .Z(n1717) );
  IV U13349 ( .A(n11024), .Z(n8083) );
  XNOR U13350 ( .A(n12371), .B(n10609), .Z(n11024) );
  ANDN U13351 ( .B(n10900), .A(n10901), .Z(n12370) );
  XNOR U13352 ( .A(n12372), .B(n9511), .Z(n10901) );
  XNOR U13353 ( .A(n12373), .B(n12374), .Z(n9511) );
  XNOR U13354 ( .A(n12375), .B(n9274), .Z(n10900) );
  XNOR U13355 ( .A(n12376), .B(n8094), .Z(n4312) );
  XOR U13356 ( .A(n12377), .B(n11235), .Z(n8094) );
  ANDN U13357 ( .B(n12167), .A(n12378), .Z(n12376) );
  XNOR U13358 ( .A(n12379), .B(n12378), .Z(n10897) );
  IV U13359 ( .A(n11028), .Z(n12378) );
  XOR U13360 ( .A(n12380), .B(n12381), .Z(n11028) );
  NOR U13361 ( .A(n12167), .B(n8092), .Z(n12379) );
  XNOR U13362 ( .A(n12382), .B(n11869), .Z(n8092) );
  XNOR U13363 ( .A(n12383), .B(n11213), .Z(n12167) );
  XNOR U13364 ( .A(n12384), .B(n6205), .Z(out[1006]) );
  IV U13365 ( .A(n6902), .Z(n6205) );
  XNOR U13366 ( .A(n8831), .B(n2271), .Z(n6902) );
  XNOR U13367 ( .A(n6088), .B(n6164), .Z(n2271) );
  XNOR U13368 ( .A(n12385), .B(n12386), .Z(n6164) );
  XOR U13369 ( .A(n2307), .B(n5464), .Z(n12386) );
  XNOR U13370 ( .A(n12387), .B(n7612), .Z(n5464) );
  XOR U13371 ( .A(n12388), .B(n9910), .Z(n7612) );
  ANDN U13372 ( .B(n8841), .A(n7613), .Z(n12387) );
  XOR U13373 ( .A(n12389), .B(n10106), .Z(n7613) );
  IV U13374 ( .A(n12299), .Z(n10106) );
  XOR U13375 ( .A(n9652), .B(n12390), .Z(n8841) );
  XOR U13376 ( .A(n12391), .B(n7617), .Z(n2307) );
  XOR U13377 ( .A(n12392), .B(n9547), .Z(n7617) );
  NOR U13378 ( .A(n8836), .B(n7616), .Z(n12391) );
  XOR U13379 ( .A(n12393), .B(n9800), .Z(n7616) );
  XNOR U13380 ( .A(n12394), .B(n12395), .Z(n8836) );
  XOR U13381 ( .A(n3157), .B(n12396), .Z(n12385) );
  XOR U13382 ( .A(n6069), .B(n7606), .Z(n12396) );
  XNOR U13383 ( .A(n12397), .B(n7622), .Z(n7606) );
  XOR U13384 ( .A(n12398), .B(n12399), .Z(n7622) );
  ANDN U13385 ( .B(n8839), .A(n7621), .Z(n12397) );
  XOR U13386 ( .A(n12400), .B(n10302), .Z(n7621) );
  IV U13387 ( .A(n10388), .Z(n10302) );
  XOR U13388 ( .A(n12401), .B(n11440), .Z(n8839) );
  XNOR U13389 ( .A(n12402), .B(n7626), .Z(n6069) );
  XNOR U13390 ( .A(n12403), .B(n12117), .Z(n7626) );
  NOR U13391 ( .A(n12260), .B(n7625), .Z(n12402) );
  XNOR U13392 ( .A(n12404), .B(n7629), .Z(n3157) );
  XNOR U13393 ( .A(n12405), .B(n10300), .Z(n7629) );
  ANDN U13394 ( .B(n8833), .A(n7630), .Z(n12404) );
  XOR U13395 ( .A(n12406), .B(n11634), .Z(n7630) );
  XNOR U13396 ( .A(n12407), .B(n9788), .Z(n8833) );
  XOR U13397 ( .A(n12408), .B(n12409), .Z(n6088) );
  XNOR U13398 ( .A(n5283), .B(n1929), .Z(n12409) );
  XOR U13399 ( .A(n12410), .B(n8900), .Z(n1929) );
  ANDN U13400 ( .B(n8819), .A(n7702), .Z(n12410) );
  XNOR U13401 ( .A(n12411), .B(n12412), .Z(n7702) );
  XOR U13402 ( .A(n9565), .B(n12413), .Z(n8819) );
  XOR U13403 ( .A(n12414), .B(n8905), .Z(n5283) );
  ANDN U13404 ( .B(n8817), .A(n7694), .Z(n12414) );
  XNOR U13405 ( .A(n12415), .B(n10307), .Z(n7694) );
  XNOR U13406 ( .A(n12416), .B(n12417), .Z(n10307) );
  XOR U13407 ( .A(n12418), .B(n12419), .Z(n8817) );
  XNOR U13408 ( .A(n3720), .B(n12420), .Z(n12408) );
  XNOR U13409 ( .A(n8880), .B(n4191), .Z(n12420) );
  XOR U13410 ( .A(n12421), .B(n8907), .Z(n4191) );
  ANDN U13411 ( .B(n7685), .A(n8828), .Z(n12421) );
  XOR U13412 ( .A(n12422), .B(n12423), .Z(n8828) );
  XOR U13413 ( .A(n12424), .B(n12425), .Z(n7685) );
  XNOR U13414 ( .A(n12426), .B(n8903), .Z(n8880) );
  IV U13415 ( .A(n12427), .Z(n8903) );
  NOR U13416 ( .A(n7689), .B(n8823), .Z(n12426) );
  XOR U13417 ( .A(n12345), .B(n10521), .Z(n8823) );
  XNOR U13418 ( .A(n12428), .B(n12429), .Z(n12345) );
  ANDN U13419 ( .B(n12430), .A(n12431), .Z(n12428) );
  XOR U13420 ( .A(n12432), .B(n9959), .Z(n7689) );
  XOR U13421 ( .A(n12433), .B(n12434), .Z(n3720) );
  ANDN U13422 ( .B(n7698), .A(n8826), .Z(n12433) );
  XOR U13423 ( .A(n12435), .B(n11688), .Z(n7698) );
  XOR U13424 ( .A(n12436), .B(n7625), .Z(n8831) );
  XOR U13425 ( .A(n12437), .B(n11733), .Z(n7625) );
  XNOR U13426 ( .A(n9153), .B(n12438), .Z(n12260) );
  XOR U13427 ( .A(n11109), .B(n12439), .Z(n8730) );
  IV U13428 ( .A(n12411), .Z(n11109) );
  XNOR U13429 ( .A(n10721), .B(n12440), .Z(n12411) );
  XOR U13430 ( .A(n12441), .B(n12442), .Z(n10721) );
  XOR U13431 ( .A(n12443), .B(n12444), .Z(n12442) );
  XOR U13432 ( .A(n11941), .B(n12445), .Z(n12441) );
  XOR U13433 ( .A(n12446), .B(n12447), .Z(n12445) );
  XOR U13434 ( .A(n12448), .B(n12449), .Z(n11941) );
  ANDN U13435 ( .B(n12450), .A(n12451), .Z(n12448) );
  ANDN U13436 ( .B(n5680), .A(n5682), .Z(n12384) );
  XOR U13437 ( .A(n11011), .B(n2082), .Z(n5682) );
  XNOR U13438 ( .A(n8074), .B(n9283), .Z(n2082) );
  XNOR U13439 ( .A(n12452), .B(n12453), .Z(n9283) );
  XOR U13440 ( .A(n5485), .B(n3613), .Z(n12453) );
  XNOR U13441 ( .A(n12454), .B(n12455), .Z(n3613) );
  ANDN U13442 ( .B(n8201), .A(n8200), .Z(n12454) );
  IV U13443 ( .A(n12456), .Z(n8200) );
  XOR U13444 ( .A(n10386), .B(n12457), .Z(n8201) );
  XNOR U13445 ( .A(n12458), .B(n11140), .Z(n5485) );
  NOR U13446 ( .A(n8196), .B(n8197), .Z(n12458) );
  XNOR U13447 ( .A(n12443), .B(n11942), .Z(n8197) );
  XNOR U13448 ( .A(n12459), .B(n12460), .Z(n12443) );
  ANDN U13449 ( .B(n12461), .A(n12462), .Z(n12459) );
  IV U13450 ( .A(n11141), .Z(n8196) );
  XOR U13451 ( .A(n12463), .B(n11360), .Z(n11141) );
  XOR U13452 ( .A(n6292), .B(n12464), .Z(n12452) );
  XOR U13453 ( .A(n2356), .B(n5460), .Z(n12464) );
  XNOR U13454 ( .A(n12465), .B(n11152), .Z(n5460) );
  ANDN U13455 ( .B(n9285), .A(n9287), .Z(n12465) );
  XOR U13456 ( .A(n10738), .B(n12466), .Z(n9287) );
  XNOR U13457 ( .A(n12467), .B(n9448), .Z(n9285) );
  XNOR U13458 ( .A(n12468), .B(n12253), .Z(n9448) );
  XNOR U13459 ( .A(n12469), .B(n12470), .Z(n12253) );
  XOR U13460 ( .A(n11474), .B(n11282), .Z(n12470) );
  XNOR U13461 ( .A(n12471), .B(n12472), .Z(n11282) );
  ANDN U13462 ( .B(n12473), .A(n12474), .Z(n12471) );
  XOR U13463 ( .A(n12475), .B(n12476), .Z(n11474) );
  NOR U13464 ( .A(n12477), .B(n12478), .Z(n12475) );
  XOR U13465 ( .A(n12479), .B(n12480), .Z(n12469) );
  XOR U13466 ( .A(n11512), .B(n11910), .Z(n12480) );
  XOR U13467 ( .A(n12481), .B(n12482), .Z(n11910) );
  ANDN U13468 ( .B(n12483), .A(n12484), .Z(n12481) );
  XNOR U13469 ( .A(n12485), .B(n12486), .Z(n11512) );
  ANDN U13470 ( .B(n12487), .A(n12488), .Z(n12485) );
  XOR U13471 ( .A(n12489), .B(n11144), .Z(n2356) );
  ANDN U13472 ( .B(n8188), .A(n8186), .Z(n12489) );
  XNOR U13473 ( .A(n12490), .B(n10850), .Z(n8186) );
  XNOR U13474 ( .A(n12491), .B(n9613), .Z(n8188) );
  XNOR U13475 ( .A(n12492), .B(n11149), .Z(n6292) );
  ANDN U13476 ( .B(n8192), .A(n8190), .Z(n12492) );
  XOR U13477 ( .A(n12493), .B(n12494), .Z(n8190) );
  XNOR U13478 ( .A(n12495), .B(n11085), .Z(n8192) );
  XOR U13479 ( .A(n12496), .B(n12497), .Z(n8074) );
  XNOR U13480 ( .A(n3831), .B(n5149), .Z(n12497) );
  XOR U13481 ( .A(n12498), .B(n9187), .Z(n5149) );
  XNOR U13482 ( .A(n12499), .B(n12500), .Z(n9187) );
  ANDN U13483 ( .B(n11018), .A(n11019), .Z(n12498) );
  XNOR U13484 ( .A(n12501), .B(n9524), .Z(n11019) );
  XOR U13485 ( .A(n12502), .B(n10850), .Z(n11018) );
  XNOR U13486 ( .A(n12504), .B(n9893), .Z(n8162) );
  NOR U13487 ( .A(n11009), .B(n11010), .Z(n12503) );
  XNOR U13488 ( .A(n9515), .B(n12505), .Z(n11010) );
  XNOR U13489 ( .A(n12506), .B(n9759), .Z(n11009) );
  XNOR U13490 ( .A(n4339), .B(n12507), .Z(n12496) );
  XOR U13491 ( .A(n1726), .B(n11125), .Z(n12507) );
  XNOR U13492 ( .A(n12508), .B(n8172), .Z(n11125) );
  IV U13493 ( .A(n11135), .Z(n8172) );
  XNOR U13494 ( .A(n10743), .B(n12509), .Z(n11135) );
  ANDN U13495 ( .B(n11005), .A(n11006), .Z(n12508) );
  IV U13496 ( .A(n12319), .Z(n11006) );
  XOR U13497 ( .A(n12510), .B(n9978), .Z(n12319) );
  XOR U13498 ( .A(n12511), .B(n11460), .Z(n11005) );
  XNOR U13499 ( .A(n12512), .B(n8166), .Z(n1726) );
  XOR U13500 ( .A(n11118), .B(n12513), .Z(n8166) );
  NOR U13501 ( .A(n11015), .B(n11014), .Z(n12512) );
  XOR U13502 ( .A(n9153), .B(n12514), .Z(n11014) );
  IV U13503 ( .A(n12333), .Z(n11015) );
  XOR U13504 ( .A(n9761), .B(n12515), .Z(n12333) );
  XNOR U13505 ( .A(n12516), .B(n12517), .Z(n9761) );
  XNOR U13506 ( .A(n12518), .B(n8176), .Z(n4339) );
  XOR U13507 ( .A(n12519), .B(n12520), .Z(n8176) );
  AND U13508 ( .A(n12316), .B(n11132), .Z(n12518) );
  XOR U13509 ( .A(n12521), .B(n11132), .Z(n11011) );
  XOR U13510 ( .A(n12522), .B(n12360), .Z(n11132) );
  IV U13511 ( .A(n9420), .Z(n12360) );
  NOR U13512 ( .A(n12316), .B(n8174), .Z(n12521) );
  XOR U13513 ( .A(n11301), .B(n12523), .Z(n8174) );
  XNOR U13514 ( .A(n12524), .B(n11340), .Z(n12316) );
  XNOR U13515 ( .A(n1762), .B(n8588), .Z(n5680) );
  XOR U13516 ( .A(n12525), .B(n8665), .Z(n8588) );
  ANDN U13517 ( .B(n12290), .A(n6437), .Z(n12525) );
  XOR U13518 ( .A(n10885), .B(n12526), .Z(n6437) );
  IV U13519 ( .A(n12527), .Z(n10885) );
  XNOR U13520 ( .A(n9915), .B(n6330), .Z(n1762) );
  XOR U13521 ( .A(n12528), .B(n12529), .Z(n6330) );
  XNOR U13522 ( .A(n5905), .B(n2113), .Z(n12529) );
  XNOR U13523 ( .A(n12530), .B(n8672), .Z(n2113) );
  ANDN U13524 ( .B(n6467), .A(n8758), .Z(n12530) );
  IV U13525 ( .A(n6469), .Z(n8758) );
  XOR U13526 ( .A(n12531), .B(n10209), .Z(n6469) );
  XNOR U13527 ( .A(n12532), .B(n9802), .Z(n6467) );
  IV U13528 ( .A(n9248), .Z(n9802) );
  XNOR U13529 ( .A(n11861), .B(n11371), .Z(n9248) );
  XOR U13530 ( .A(n12533), .B(n12534), .Z(n11371) );
  XNOR U13531 ( .A(n12467), .B(n11477), .Z(n12534) );
  XNOR U13532 ( .A(n12535), .B(n12536), .Z(n11477) );
  NOR U13533 ( .A(n12537), .B(n12538), .Z(n12535) );
  XOR U13534 ( .A(n12539), .B(n12540), .Z(n12467) );
  NOR U13535 ( .A(n12541), .B(n12542), .Z(n12539) );
  XOR U13536 ( .A(n11240), .B(n12543), .Z(n12533) );
  XOR U13537 ( .A(n9447), .B(n11710), .Z(n12543) );
  XNOR U13538 ( .A(n12544), .B(n12545), .Z(n11710) );
  NOR U13539 ( .A(n12546), .B(n12547), .Z(n12544) );
  XNOR U13540 ( .A(n12548), .B(n12549), .Z(n9447) );
  AND U13541 ( .A(n12550), .B(n12551), .Z(n12548) );
  XOR U13542 ( .A(n12552), .B(n12553), .Z(n11240) );
  ANDN U13543 ( .B(n12554), .A(n12555), .Z(n12552) );
  XOR U13544 ( .A(n12556), .B(n12557), .Z(n11861) );
  XNOR U13545 ( .A(n12558), .B(n12559), .Z(n12557) );
  XOR U13546 ( .A(n12560), .B(n12561), .Z(n12556) );
  XNOR U13547 ( .A(n12303), .B(n9141), .Z(n12561) );
  XNOR U13548 ( .A(n12562), .B(n12563), .Z(n9141) );
  XNOR U13549 ( .A(n12566), .B(n12567), .Z(n12303) );
  ANDN U13550 ( .B(n12568), .A(n12569), .Z(n12566) );
  XOR U13551 ( .A(n12570), .B(n8683), .Z(n5905) );
  XOR U13552 ( .A(n9780), .B(n12571), .Z(n6472) );
  XOR U13553 ( .A(n9238), .B(n12572), .Z(n6471) );
  XOR U13554 ( .A(n3702), .B(n12573), .Z(n12528) );
  XNOR U13555 ( .A(n4326), .B(n5450), .Z(n12573) );
  XOR U13556 ( .A(n12574), .B(n12575), .Z(n5450) );
  ANDN U13557 ( .B(n6455), .A(n6454), .Z(n12574) );
  XOR U13558 ( .A(n12576), .B(n11166), .Z(n6454) );
  XNOR U13559 ( .A(n12577), .B(n12107), .Z(n6455) );
  XNOR U13560 ( .A(n12578), .B(n8680), .Z(n4326) );
  NOR U13561 ( .A(n6459), .B(n6458), .Z(n12578) );
  XOR U13562 ( .A(n10752), .B(n12579), .Z(n6458) );
  XNOR U13563 ( .A(n9263), .B(n12580), .Z(n6459) );
  XOR U13564 ( .A(n12581), .B(n12582), .Z(n3702) );
  ANDN U13565 ( .B(n6463), .A(n6464), .Z(n12581) );
  XOR U13566 ( .A(n10604), .B(n12583), .Z(n6464) );
  XOR U13567 ( .A(n12584), .B(n12585), .Z(n9915) );
  XOR U13568 ( .A(n4875), .B(n8657), .Z(n12585) );
  XNOR U13569 ( .A(n12586), .B(n6430), .Z(n8657) );
  XOR U13570 ( .A(n10313), .B(n12587), .Z(n6430) );
  XNOR U13571 ( .A(n12588), .B(n12589), .Z(n10313) );
  ANDN U13572 ( .B(n8585), .A(n8586), .Z(n12586) );
  XOR U13573 ( .A(n12326), .B(n12590), .Z(n8586) );
  XOR U13574 ( .A(n12591), .B(n10280), .Z(n8585) );
  XNOR U13575 ( .A(n12592), .B(n6433), .Z(n4875) );
  IV U13576 ( .A(n8662), .Z(n6433) );
  XOR U13577 ( .A(n12593), .B(n12247), .Z(n8662) );
  NOR U13578 ( .A(n8592), .B(n8591), .Z(n12592) );
  XOR U13579 ( .A(n12594), .B(n11733), .Z(n8591) );
  XOR U13580 ( .A(n9924), .B(n12595), .Z(n8592) );
  IV U13581 ( .A(n10116), .Z(n9924) );
  XOR U13582 ( .A(n2501), .B(n12598), .Z(n12584) );
  XOR U13583 ( .A(n3501), .B(n4362), .Z(n12598) );
  XNOR U13584 ( .A(n12599), .B(n6439), .Z(n4362) );
  XOR U13585 ( .A(n11501), .B(n12600), .Z(n6439) );
  XOR U13586 ( .A(n12601), .B(n11568), .Z(n12290) );
  XNOR U13587 ( .A(n12602), .B(n11482), .Z(n8665) );
  XOR U13588 ( .A(n12603), .B(n6443), .Z(n3501) );
  XOR U13589 ( .A(n9269), .B(n12604), .Z(n6443) );
  IV U13590 ( .A(n11604), .Z(n9269) );
  XNOR U13591 ( .A(n12605), .B(n12606), .Z(n11604) );
  NOR U13592 ( .A(n8583), .B(n8582), .Z(n12603) );
  XOR U13593 ( .A(n12607), .B(n10120), .Z(n8582) );
  XOR U13594 ( .A(n12608), .B(n12107), .Z(n8583) );
  XNOR U13595 ( .A(n12609), .B(n6447), .Z(n2501) );
  XOR U13596 ( .A(n12610), .B(n12096), .Z(n6447) );
  NOR U13597 ( .A(n12301), .B(n8595), .Z(n12609) );
  XOR U13598 ( .A(n12611), .B(n12612), .Z(n8595) );
  IV U13599 ( .A(n8596), .Z(n12301) );
  XOR U13600 ( .A(n10186), .B(n12613), .Z(n8596) );
  XNOR U13601 ( .A(n12614), .B(n6210), .Z(out[1005]) );
  IV U13602 ( .A(n6936), .Z(n6210) );
  XOR U13603 ( .A(n8898), .B(n2278), .Z(n6936) );
  XNOR U13604 ( .A(n6093), .B(n6169), .Z(n2278) );
  XNOR U13605 ( .A(n12615), .B(n12616), .Z(n6169) );
  XNOR U13606 ( .A(n2318), .B(n5472), .Z(n12616) );
  XNOR U13607 ( .A(n12617), .B(n7687), .Z(n5472) );
  XOR U13608 ( .A(n9975), .B(n12618), .Z(n7687) );
  IV U13609 ( .A(n10947), .Z(n9975) );
  ANDN U13610 ( .B(n7686), .A(n8907), .Z(n12617) );
  XNOR U13611 ( .A(n12619), .B(n9795), .Z(n8907) );
  XOR U13612 ( .A(n10209), .B(n12620), .Z(n7686) );
  XNOR U13613 ( .A(n12621), .B(n8824), .Z(n2318) );
  XOR U13614 ( .A(n9652), .B(n12622), .Z(n8824) );
  ANDN U13615 ( .B(n7691), .A(n12427), .Z(n12621) );
  XOR U13616 ( .A(n12623), .B(n11196), .Z(n12427) );
  XOR U13617 ( .A(n12626), .B(n9899), .Z(n7691) );
  XOR U13618 ( .A(n3162), .B(n12627), .Z(n12615) );
  XNOR U13619 ( .A(n6120), .B(n7680), .Z(n12627) );
  XNOR U13620 ( .A(n12628), .B(n7696), .Z(n7680) );
  XNOR U13621 ( .A(n12629), .B(n11648), .Z(n7696) );
  ANDN U13622 ( .B(n7695), .A(n8905), .Z(n12628) );
  XNOR U13623 ( .A(n12630), .B(n10482), .Z(n8905) );
  XOR U13624 ( .A(n12631), .B(n12282), .Z(n7695) );
  XOR U13625 ( .A(n12632), .B(n12633), .Z(n12282) );
  XNOR U13626 ( .A(n12634), .B(n7699), .Z(n6120) );
  XOR U13627 ( .A(n12247), .B(n12635), .Z(n7699) );
  ANDN U13628 ( .B(n7700), .A(n12434), .Z(n12634) );
  XNOR U13629 ( .A(n12636), .B(n8820), .Z(n3162) );
  IV U13630 ( .A(n7703), .Z(n8820) );
  XOR U13631 ( .A(n10399), .B(n12637), .Z(n7703) );
  ANDN U13632 ( .B(n7704), .A(n8900), .Z(n12636) );
  XOR U13633 ( .A(n12638), .B(n9886), .Z(n8900) );
  XNOR U13634 ( .A(n12639), .B(n11960), .Z(n7704) );
  XOR U13635 ( .A(n12640), .B(n12641), .Z(n6093) );
  XOR U13636 ( .A(n5285), .B(n1933), .Z(n12641) );
  AND U13637 ( .A(n8886), .B(n7780), .Z(n12642) );
  XNOR U13638 ( .A(n12643), .B(n11235), .Z(n7780) );
  XOR U13639 ( .A(n11280), .B(n12644), .Z(n8886) );
  XNOR U13640 ( .A(n12645), .B(n12646), .Z(n11280) );
  XNOR U13641 ( .A(n12647), .B(n8968), .Z(n5285) );
  ANDN U13642 ( .B(n8884), .A(n7772), .Z(n12647) );
  XNOR U13643 ( .A(n12648), .B(n10406), .Z(n7772) );
  XNOR U13644 ( .A(n12649), .B(n12650), .Z(n10406) );
  XOR U13645 ( .A(n12651), .B(n12652), .Z(n8884) );
  XNOR U13646 ( .A(n3727), .B(n12653), .Z(n12640) );
  XOR U13647 ( .A(n8944), .B(n4195), .Z(n12653) );
  XOR U13648 ( .A(n12654), .B(n8970), .Z(n4195) );
  NOR U13649 ( .A(n7763), .B(n8894), .Z(n12654) );
  XNOR U13650 ( .A(n12655), .B(n11221), .Z(n8894) );
  XNOR U13651 ( .A(n12656), .B(n9224), .Z(n7763) );
  XNOR U13652 ( .A(n12657), .B(n8965), .Z(n8944) );
  IV U13653 ( .A(n12658), .Z(n8965) );
  ANDN U13654 ( .B(n8889), .A(n7767), .Z(n12657) );
  XOR U13655 ( .A(n12659), .B(n12220), .Z(n7767) );
  XNOR U13656 ( .A(n12660), .B(n9463), .Z(n8889) );
  XOR U13657 ( .A(n12661), .B(n12662), .Z(n9463) );
  XNOR U13658 ( .A(n12663), .B(n12664), .Z(n3727) );
  NOR U13659 ( .A(n8891), .B(n7776), .Z(n12663) );
  XOR U13660 ( .A(n12665), .B(n10193), .Z(n7776) );
  XNOR U13661 ( .A(n12666), .B(n7700), .Z(n8898) );
  XOR U13662 ( .A(n10958), .B(n12667), .Z(n7700) );
  XOR U13663 ( .A(n9252), .B(n12668), .Z(n12434) );
  XOR U13664 ( .A(n12669), .B(n11235), .Z(n8826) );
  XNOR U13665 ( .A(n12670), .B(n12671), .Z(n11235) );
  ANDN U13666 ( .B(n5686), .A(n5684), .Z(n12614) );
  XNOR U13667 ( .A(n8677), .B(n5173), .Z(n5684) );
  XNOR U13668 ( .A(n12672), .B(n12673), .Z(n6424) );
  XNOR U13669 ( .A(n4398), .B(n2507), .Z(n12673) );
  XNOR U13670 ( .A(n12674), .B(n6473), .Z(n2507) );
  XNOR U13671 ( .A(n12675), .B(n11369), .Z(n6473) );
  ANDN U13672 ( .B(n8683), .A(n8760), .Z(n12674) );
  XNOR U13673 ( .A(n12676), .B(n10727), .Z(n8760) );
  XOR U13674 ( .A(n12677), .B(n10324), .Z(n8683) );
  XOR U13675 ( .A(n12678), .B(n12679), .Z(n10324) );
  XNOR U13676 ( .A(n12680), .B(n8756), .Z(n4398) );
  XNOR U13677 ( .A(n10965), .B(n12681), .Z(n8756) );
  NOR U13678 ( .A(n8755), .B(n12582), .Z(n12680) );
  XOR U13679 ( .A(n3504), .B(n12682), .Z(n12672) );
  XOR U13680 ( .A(n8747), .B(n4879), .Z(n12682) );
  XNOR U13681 ( .A(n12683), .B(n6460), .Z(n4879) );
  IV U13682 ( .A(n8752), .Z(n6460) );
  XOR U13683 ( .A(n12684), .B(n12685), .Z(n8752) );
  ANDN U13684 ( .B(n8680), .A(n8679), .Z(n12683) );
  XNOR U13685 ( .A(n10958), .B(n12686), .Z(n8679) );
  IV U13686 ( .A(n12687), .Z(n10958) );
  XOR U13687 ( .A(n10928), .B(n12688), .Z(n8680) );
  XNOR U13688 ( .A(n12689), .B(n6456), .Z(n8747) );
  XOR U13689 ( .A(n12690), .B(n11081), .Z(n6456) );
  ANDN U13690 ( .B(n8674), .A(n12575), .Z(n12689) );
  IV U13691 ( .A(n8675), .Z(n12575) );
  XOR U13692 ( .A(n12691), .B(n10738), .Z(n8675) );
  XNOR U13693 ( .A(n12692), .B(n12693), .Z(n8674) );
  XNOR U13694 ( .A(n12694), .B(n6468), .Z(n3504) );
  XOR U13695 ( .A(n12695), .B(n11925), .Z(n6468) );
  AND U13696 ( .A(n8672), .B(n8671), .Z(n12694) );
  XNOR U13697 ( .A(n12696), .B(n10219), .Z(n8671) );
  XOR U13698 ( .A(n12697), .B(n12235), .Z(n8672) );
  XOR U13699 ( .A(n12698), .B(n12699), .Z(n6335) );
  XOR U13700 ( .A(n5455), .B(n3706), .Z(n12699) );
  XNOR U13701 ( .A(n12700), .B(n12701), .Z(n3706) );
  ANDN U13702 ( .B(n6490), .A(n6491), .Z(n12700) );
  XOR U13703 ( .A(n12702), .B(n10727), .Z(n6491) );
  XNOR U13704 ( .A(n12703), .B(n8768), .Z(n5455) );
  ANDN U13705 ( .B(n6481), .A(n6483), .Z(n12703) );
  XOR U13706 ( .A(n12235), .B(n12704), .Z(n6483) );
  IV U13707 ( .A(n11467), .Z(n12235) );
  XOR U13708 ( .A(n12705), .B(n12706), .Z(n6481) );
  XOR U13709 ( .A(n4329), .B(n12707), .Z(n12698) );
  XOR U13710 ( .A(n5910), .B(n2117), .Z(n12707) );
  XOR U13711 ( .A(n12708), .B(n8765), .Z(n2117) );
  ANDN U13712 ( .B(n6494), .A(n6495), .Z(n12708) );
  XNOR U13713 ( .A(n12709), .B(n10343), .Z(n6495) );
  XNOR U13714 ( .A(n12710), .B(n9322), .Z(n6494) );
  XNOR U13715 ( .A(n12711), .B(n8776), .Z(n5910) );
  ANDN U13716 ( .B(n6499), .A(n6498), .Z(n12711) );
  IV U13717 ( .A(n8777), .Z(n6498) );
  XOR U13718 ( .A(n12712), .B(n12713), .Z(n8777) );
  XOR U13719 ( .A(n10934), .B(n12714), .Z(n6499) );
  XNOR U13720 ( .A(n12715), .B(n8773), .Z(n4329) );
  IV U13721 ( .A(n12716), .Z(n8773) );
  ANDN U13722 ( .B(n6485), .A(n6486), .Z(n12715) );
  XNOR U13723 ( .A(n12717), .B(n12718), .Z(n6486) );
  XOR U13724 ( .A(n10738), .B(n12719), .Z(n6485) );
  XOR U13725 ( .A(n12722), .B(n8755), .Z(n8677) );
  XOR U13726 ( .A(n12723), .B(n12103), .Z(n8755) );
  IV U13727 ( .A(n11630), .Z(n12103) );
  ANDN U13728 ( .B(n12582), .A(n6463), .Z(n12722) );
  XNOR U13729 ( .A(n12724), .B(n11054), .Z(n6463) );
  XOR U13730 ( .A(n12725), .B(n10060), .Z(n12582) );
  XOR U13731 ( .A(n11145), .B(n2086), .Z(n5686) );
  XNOR U13732 ( .A(n8156), .B(n9404), .Z(n2086) );
  XNOR U13733 ( .A(n12726), .B(n12727), .Z(n9404) );
  XNOR U13734 ( .A(n5490), .B(n3619), .Z(n12727) );
  XOR U13735 ( .A(n12728), .B(n12729), .Z(n3619) );
  ANDN U13736 ( .B(n8256), .A(n8254), .Z(n12728) );
  IV U13737 ( .A(n12730), .Z(n8254) );
  XNOR U13738 ( .A(n11106), .B(n12731), .Z(n8256) );
  XNOR U13739 ( .A(n12732), .B(n11262), .Z(n5490) );
  NOR U13740 ( .A(n11263), .B(n8251), .Z(n12732) );
  XNOR U13741 ( .A(n12733), .B(n10763), .Z(n8251) );
  IV U13742 ( .A(n12734), .Z(n10763) );
  XOR U13743 ( .A(n12735), .B(n12736), .Z(n11263) );
  XOR U13744 ( .A(n6296), .B(n12737), .Z(n12726) );
  XOR U13745 ( .A(n2363), .B(n5513), .Z(n12737) );
  XOR U13746 ( .A(n12738), .B(n11274), .Z(n5513) );
  ANDN U13747 ( .B(n9408), .A(n9406), .Z(n12738) );
  XNOR U13748 ( .A(n9544), .B(n12739), .Z(n9406) );
  XNOR U13749 ( .A(n12740), .B(n12741), .Z(n9544) );
  XNOR U13750 ( .A(n12742), .B(n10842), .Z(n9408) );
  XNOR U13751 ( .A(n12743), .B(n11266), .Z(n2363) );
  ANDN U13752 ( .B(n8242), .A(n8240), .Z(n12743) );
  XOR U13753 ( .A(n12744), .B(n10526), .Z(n8240) );
  XNOR U13754 ( .A(n12745), .B(n9755), .Z(n8242) );
  XNOR U13755 ( .A(n12746), .B(n11271), .Z(n6296) );
  ANDN U13756 ( .B(n8244), .A(n8245), .Z(n12746) );
  XOR U13757 ( .A(n12747), .B(n11213), .Z(n8245) );
  XOR U13758 ( .A(n12748), .B(n11891), .Z(n8244) );
  XOR U13759 ( .A(n12749), .B(n12750), .Z(n8156) );
  XNOR U13760 ( .A(n3836), .B(n5151), .Z(n12750) );
  XOR U13761 ( .A(n12751), .B(n9286), .Z(n5151) );
  XOR U13762 ( .A(n12717), .B(n12752), .Z(n9286) );
  ANDN U13763 ( .B(n11151), .A(n11152), .Z(n12751) );
  XOR U13764 ( .A(n10698), .B(n12753), .Z(n11152) );
  XOR U13765 ( .A(n12754), .B(n10526), .Z(n11151) );
  XNOR U13766 ( .A(n12755), .B(n12756), .Z(n10526) );
  XNOR U13767 ( .A(n12757), .B(n8187), .Z(n3836) );
  IV U13768 ( .A(n11256), .Z(n8187) );
  XOR U13769 ( .A(n12758), .B(n9959), .Z(n11256) );
  ANDN U13770 ( .B(n11144), .A(n11143), .Z(n12757) );
  XOR U13771 ( .A(n9929), .B(n12759), .Z(n11143) );
  XNOR U13772 ( .A(n9620), .B(n12760), .Z(n11144) );
  XNOR U13773 ( .A(n4363), .B(n12761), .Z(n12749) );
  XOR U13774 ( .A(n1731), .B(n11247), .Z(n12761) );
  XOR U13775 ( .A(n12762), .B(n8198), .Z(n11247) );
  XNOR U13776 ( .A(n12763), .B(n11458), .Z(n8198) );
  IV U13777 ( .A(n10640), .Z(n11458) );
  XOR U13778 ( .A(n12764), .B(n12765), .Z(n10640) );
  ANDN U13779 ( .B(n11139), .A(n11140), .Z(n12762) );
  XOR U13780 ( .A(n12766), .B(n10630), .Z(n11140) );
  XNOR U13781 ( .A(n12767), .B(n10724), .Z(n11139) );
  XOR U13782 ( .A(n12768), .B(n12769), .Z(n10724) );
  XNOR U13783 ( .A(n12770), .B(n8191), .Z(n1731) );
  XOR U13784 ( .A(n12771), .B(n11243), .Z(n8191) );
  IV U13785 ( .A(n10836), .Z(n11243) );
  ANDN U13786 ( .B(n11148), .A(n11149), .Z(n12770) );
  XOR U13787 ( .A(n12772), .B(n9759), .Z(n11149) );
  XNOR U13788 ( .A(n12773), .B(n12774), .Z(n9759) );
  XOR U13789 ( .A(n9252), .B(n12775), .Z(n11148) );
  XNOR U13790 ( .A(n12776), .B(n8202), .Z(n4363) );
  XNOR U13791 ( .A(n12777), .B(n11503), .Z(n8202) );
  ANDN U13792 ( .B(n11254), .A(n12455), .Z(n12776) );
  XOR U13793 ( .A(n12778), .B(n11254), .Z(n11145) );
  XNOR U13794 ( .A(n11878), .B(n12779), .Z(n11254) );
  IV U13795 ( .A(n9515), .Z(n11878) );
  ANDN U13796 ( .B(n12455), .A(n12456), .Z(n12778) );
  XOR U13797 ( .A(n12311), .B(n12780), .Z(n12456) );
  XOR U13798 ( .A(n12781), .B(n11482), .Z(n12455) );
  XNOR U13799 ( .A(n12782), .B(n6215), .Z(out[1004]) );
  IV U13800 ( .A(n6961), .Z(n6215) );
  XOR U13801 ( .A(n8960), .B(n2285), .Z(n6961) );
  XNOR U13802 ( .A(n6098), .B(n6179), .Z(n2285) );
  XNOR U13803 ( .A(n12783), .B(n12784), .Z(n6179) );
  XOR U13804 ( .A(n2323), .B(n5475), .Z(n12784) );
  XNOR U13805 ( .A(n12785), .B(n8895), .Z(n5475) );
  IV U13806 ( .A(n7765), .Z(n8895) );
  XOR U13807 ( .A(n10282), .B(n12786), .Z(n7765) );
  IV U13808 ( .A(n12787), .Z(n10282) );
  NOR U13809 ( .A(n8970), .B(n7764), .Z(n12785) );
  XOR U13810 ( .A(n12788), .B(n10343), .Z(n7764) );
  XOR U13811 ( .A(n12789), .B(n9891), .Z(n8970) );
  XOR U13812 ( .A(n12790), .B(n7768), .Z(n2323) );
  XOR U13813 ( .A(n12791), .B(n9815), .Z(n7768) );
  ANDN U13814 ( .B(n7769), .A(n12658), .Z(n12790) );
  XOR U13815 ( .A(n12792), .B(n12107), .Z(n12658) );
  IV U13816 ( .A(n11325), .Z(n12107) );
  XOR U13817 ( .A(n12794), .B(n12795), .Z(n12205) );
  XNOR U13818 ( .A(n9763), .B(n12796), .Z(n12795) );
  XNOR U13819 ( .A(n12797), .B(n12798), .Z(n9763) );
  ANDN U13820 ( .B(n12799), .A(n12800), .Z(n12797) );
  XOR U13821 ( .A(n11296), .B(n12801), .Z(n12794) );
  XOR U13822 ( .A(n10293), .B(n12802), .Z(n12801) );
  XNOR U13823 ( .A(n12803), .B(n12804), .Z(n10293) );
  ANDN U13824 ( .B(n12805), .A(n12806), .Z(n12803) );
  XNOR U13825 ( .A(n12807), .B(n12808), .Z(n11296) );
  NOR U13826 ( .A(n12809), .B(n12810), .Z(n12807) );
  XOR U13827 ( .A(n9966), .B(n12811), .Z(n7769) );
  XNOR U13828 ( .A(n3166), .B(n12812), .Z(n12783) );
  XNOR U13829 ( .A(n6175), .B(n7758), .Z(n12812) );
  XNOR U13830 ( .A(n12813), .B(n7774), .Z(n7758) );
  XOR U13831 ( .A(n11972), .B(n12814), .Z(n7774) );
  ANDN U13832 ( .B(n8968), .A(n8967), .Z(n12813) );
  XOR U13833 ( .A(n12611), .B(n12815), .Z(n8967) );
  IV U13834 ( .A(n10604), .Z(n12611) );
  XOR U13835 ( .A(n11711), .B(n12818), .Z(n8968) );
  XOR U13836 ( .A(n12819), .B(n12820), .Z(n11949) );
  XNOR U13837 ( .A(n10056), .B(n11170), .Z(n12820) );
  XNOR U13838 ( .A(n12821), .B(n12822), .Z(n11170) );
  XOR U13839 ( .A(n12825), .B(n12826), .Z(n10056) );
  NOR U13840 ( .A(n12827), .B(n12828), .Z(n12825) );
  XOR U13841 ( .A(n11310), .B(n12829), .Z(n12819) );
  XOR U13842 ( .A(n12830), .B(n12831), .Z(n12829) );
  XNOR U13843 ( .A(n12832), .B(n12833), .Z(n11310) );
  ANDN U13844 ( .B(n12834), .A(n12835), .Z(n12832) );
  XNOR U13845 ( .A(n12837), .B(n8892), .Z(n6175) );
  IV U13846 ( .A(n7777), .Z(n8892) );
  XOR U13847 ( .A(n12838), .B(n12419), .Z(n7777) );
  AND U13848 ( .A(n12664), .B(n7778), .Z(n12837) );
  XNOR U13849 ( .A(n12839), .B(n7781), .Z(n3166) );
  XNOR U13850 ( .A(n10602), .B(n12840), .Z(n7781) );
  ANDN U13851 ( .B(n7782), .A(n8962), .Z(n12839) );
  XOR U13852 ( .A(n12841), .B(n9956), .Z(n8962) );
  IV U13853 ( .A(n11479), .Z(n9956) );
  XOR U13854 ( .A(n12842), .B(n12843), .Z(n7782) );
  XOR U13855 ( .A(n12844), .B(n12845), .Z(n6098) );
  XOR U13856 ( .A(n5287), .B(n1938), .Z(n12845) );
  XOR U13857 ( .A(n12846), .B(n8997), .Z(n1938) );
  ANDN U13858 ( .B(n8950), .A(n7844), .Z(n12846) );
  XOR U13859 ( .A(n12847), .B(n12520), .Z(n7844) );
  XNOR U13860 ( .A(n12848), .B(n9817), .Z(n8950) );
  XNOR U13861 ( .A(n12849), .B(n12850), .Z(n9817) );
  XNOR U13862 ( .A(n12851), .B(n9003), .Z(n5287) );
  NOR U13863 ( .A(n8948), .B(n7836), .Z(n12851) );
  XOR U13864 ( .A(n12852), .B(n10609), .Z(n7836) );
  XNOR U13865 ( .A(n12679), .B(n12853), .Z(n10609) );
  XOR U13866 ( .A(n12854), .B(n12855), .Z(n12679) );
  XNOR U13867 ( .A(n12856), .B(n10379), .Z(n12855) );
  XOR U13868 ( .A(n12857), .B(n12858), .Z(n10379) );
  XNOR U13869 ( .A(n9223), .B(n12861), .Z(n12854) );
  XNOR U13870 ( .A(n12862), .B(n12656), .Z(n12861) );
  XOR U13871 ( .A(n12863), .B(n12864), .Z(n12656) );
  ANDN U13872 ( .B(n12865), .A(n12866), .Z(n12863) );
  XNOR U13873 ( .A(n12867), .B(n12868), .Z(n9223) );
  XOR U13874 ( .A(n12871), .B(n12872), .Z(n12559) );
  ANDN U13875 ( .B(n12873), .A(n12874), .Z(n12871) );
  XNOR U13876 ( .A(n3734), .B(n12875), .Z(n12844) );
  XNOR U13877 ( .A(n8978), .B(n4201), .Z(n12875) );
  XOR U13878 ( .A(n12876), .B(n9005), .Z(n4201) );
  ANDN U13879 ( .B(n7827), .A(n8957), .Z(n12876) );
  XNOR U13880 ( .A(n12877), .B(n10193), .Z(n8957) );
  XNOR U13881 ( .A(n12878), .B(n12879), .Z(n10193) );
  XNOR U13882 ( .A(n12880), .B(n12881), .Z(n7827) );
  XNOR U13883 ( .A(n12882), .B(n9000), .Z(n8978) );
  AND U13884 ( .A(n8953), .B(n7831), .Z(n12882) );
  XOR U13885 ( .A(n12883), .B(n12299), .Z(n7831) );
  XOR U13886 ( .A(n11922), .B(n12884), .Z(n8953) );
  XNOR U13887 ( .A(n12885), .B(n12886), .Z(n11922) );
  XOR U13888 ( .A(n12887), .B(n12888), .Z(n3734) );
  ANDN U13889 ( .B(n8955), .A(n7840), .Z(n12887) );
  XNOR U13890 ( .A(n12889), .B(n11490), .Z(n7840) );
  IV U13891 ( .A(n10331), .Z(n11490) );
  XNOR U13892 ( .A(n12890), .B(n7778), .Z(n8960) );
  XNOR U13893 ( .A(n12891), .B(n11039), .Z(n7778) );
  ANDN U13894 ( .B(n8891), .A(n12664), .Z(n12890) );
  XOR U13895 ( .A(n12892), .B(n12893), .Z(n12664) );
  XNOR U13896 ( .A(n12894), .B(n12520), .Z(n8891) );
  IV U13897 ( .A(n11360), .Z(n12520) );
  XOR U13898 ( .A(n12895), .B(n12896), .Z(n11360) );
  ANDN U13899 ( .B(n5688), .A(n5690), .Z(n12782) );
  XNOR U13900 ( .A(n11267), .B(n2089), .Z(n5690) );
  XNOR U13901 ( .A(n8182), .B(n9498), .Z(n2089) );
  XNOR U13902 ( .A(n12897), .B(n12898), .Z(n9498) );
  XNOR U13903 ( .A(n5494), .B(n3629), .Z(n12898) );
  XNOR U13904 ( .A(n12899), .B(n12900), .Z(n3629) );
  ANDN U13905 ( .B(n8308), .A(n11523), .Z(n12899) );
  XOR U13906 ( .A(n12901), .B(n10714), .Z(n11523) );
  XNOR U13907 ( .A(n12902), .B(n11390), .Z(n5494) );
  ANDN U13908 ( .B(n8306), .A(n11391), .Z(n12902) );
  XNOR U13909 ( .A(n12903), .B(n11614), .Z(n11391) );
  XOR U13910 ( .A(n12904), .B(n10860), .Z(n8306) );
  XOR U13911 ( .A(n6300), .B(n12905), .Z(n12897) );
  XOR U13912 ( .A(n2370), .B(n5559), .Z(n12905) );
  XOR U13913 ( .A(n12906), .B(n12907), .Z(n5559) );
  ANDN U13914 ( .B(n9502), .A(n9500), .Z(n12906) );
  IV U13915 ( .A(n11405), .Z(n9500) );
  XNOR U13916 ( .A(n12908), .B(n9650), .Z(n11405) );
  XNOR U13917 ( .A(n12909), .B(n12910), .Z(n9650) );
  XOR U13918 ( .A(n12911), .B(n11099), .Z(n9502) );
  XOR U13919 ( .A(n12912), .B(n12913), .Z(n2370) );
  ANDN U13920 ( .B(n8295), .A(n11395), .Z(n12912) );
  XNOR U13921 ( .A(n12914), .B(n10646), .Z(n11395) );
  XNOR U13922 ( .A(n12915), .B(n9856), .Z(n8295) );
  XNOR U13923 ( .A(n12916), .B(n11400), .Z(n6300) );
  ANDN U13924 ( .B(n8300), .A(n11401), .Z(n12916) );
  XNOR U13925 ( .A(n10754), .B(n12917), .Z(n11401) );
  XNOR U13926 ( .A(n12918), .B(n11340), .Z(n8300) );
  XNOR U13927 ( .A(n12919), .B(n12920), .Z(n11340) );
  XOR U13928 ( .A(n12921), .B(n12922), .Z(n8182) );
  XNOR U13929 ( .A(n3840), .B(n5156), .Z(n12922) );
  XNOR U13930 ( .A(n12923), .B(n9407), .Z(n5156) );
  XOR U13931 ( .A(n11930), .B(n12924), .Z(n9407) );
  NOR U13932 ( .A(n11274), .B(n11273), .Z(n12923) );
  XNOR U13933 ( .A(n12925), .B(n10646), .Z(n11273) );
  XOR U13934 ( .A(n12926), .B(n12243), .Z(n10646) );
  XOR U13935 ( .A(n12927), .B(n12928), .Z(n12243) );
  XNOR U13936 ( .A(n12929), .B(n10870), .Z(n12928) );
  XNOR U13937 ( .A(n12930), .B(n12931), .Z(n10870) );
  NOR U13938 ( .A(n12932), .B(n12933), .Z(n12930) );
  XOR U13939 ( .A(n12085), .B(n12934), .Z(n12927) );
  XNOR U13940 ( .A(n9668), .B(n10588), .Z(n12934) );
  XNOR U13941 ( .A(n12935), .B(n12936), .Z(n10588) );
  ANDN U13942 ( .B(n12937), .A(n12938), .Z(n12935) );
  XOR U13943 ( .A(n12939), .B(n12940), .Z(n9668) );
  ANDN U13944 ( .B(n12941), .A(n12942), .Z(n12939) );
  XNOR U13945 ( .A(n12943), .B(n12944), .Z(n12085) );
  ANDN U13946 ( .B(n12945), .A(n12946), .Z(n12943) );
  XOR U13947 ( .A(n12947), .B(n12948), .Z(n11274) );
  XNOR U13948 ( .A(n12949), .B(n8241), .Z(n3840) );
  XOR U13949 ( .A(n12950), .B(n12220), .Z(n8241) );
  ANDN U13950 ( .B(n11266), .A(n11265), .Z(n12949) );
  IV U13951 ( .A(n11384), .Z(n11265) );
  XOR U13952 ( .A(n12951), .B(n11288), .Z(n11384) );
  IV U13953 ( .A(n9927), .Z(n11288) );
  XOR U13954 ( .A(n12802), .B(n9764), .Z(n11266) );
  XNOR U13955 ( .A(n12952), .B(n12953), .Z(n12802) );
  NOR U13956 ( .A(n12954), .B(n12955), .Z(n12952) );
  XOR U13957 ( .A(n4399), .B(n12956), .Z(n12921) );
  XOR U13958 ( .A(n1735), .B(n11373), .Z(n12956) );
  XOR U13959 ( .A(n12957), .B(n8252), .Z(n11373) );
  XNOR U13960 ( .A(n12958), .B(n11595), .Z(n8252) );
  XNOR U13961 ( .A(n12959), .B(n12960), .Z(n11595) );
  ANDN U13962 ( .B(n11261), .A(n11262), .Z(n12957) );
  XOR U13963 ( .A(n12961), .B(n12169), .Z(n11262) );
  XNOR U13964 ( .A(n12962), .B(n11733), .Z(n11261) );
  XNOR U13965 ( .A(n12963), .B(n12964), .Z(n11733) );
  XNOR U13966 ( .A(n12965), .B(n8246), .Z(n1735) );
  IV U13967 ( .A(n11377), .Z(n8246) );
  XOR U13968 ( .A(n12966), .B(n10971), .Z(n11377) );
  NOR U13969 ( .A(n11271), .B(n11270), .Z(n12965) );
  XOR U13970 ( .A(n12967), .B(n9557), .Z(n11270) );
  XNOR U13971 ( .A(n9929), .B(n12968), .Z(n11271) );
  IV U13972 ( .A(n9859), .Z(n9929) );
  XNOR U13973 ( .A(n12971), .B(n8255), .Z(n4399) );
  IV U13974 ( .A(n11382), .Z(n8255) );
  XOR U13975 ( .A(n12972), .B(n11614), .Z(n11382) );
  ANDN U13976 ( .B(n12729), .A(n11381), .Z(n12971) );
  XNOR U13977 ( .A(n12973), .B(n11381), .Z(n11267) );
  XOR U13978 ( .A(n9620), .B(n12974), .Z(n11381) );
  NOR U13979 ( .A(n12730), .B(n12729), .Z(n12973) );
  XOR U13980 ( .A(n12975), .B(n11630), .Z(n12729) );
  XOR U13981 ( .A(n12976), .B(n11568), .Z(n12730) );
  XNOR U13982 ( .A(n8770), .B(n5176), .Z(n5688) );
  XOR U13983 ( .A(n6339), .B(n6450), .Z(n5176) );
  XNOR U13984 ( .A(n12977), .B(n12978), .Z(n6450) );
  XNOR U13985 ( .A(n4787), .B(n2514), .Z(n12978) );
  XNOR U13986 ( .A(n12979), .B(n6500), .Z(n2514) );
  XOR U13987 ( .A(n12980), .B(n12399), .Z(n6500) );
  IV U13988 ( .A(n11515), .Z(n12399) );
  ANDN U13989 ( .B(n8775), .A(n8776), .Z(n12979) );
  XOR U13990 ( .A(n11166), .B(n12981), .Z(n8776) );
  XOR U13991 ( .A(n11814), .B(n12982), .Z(n8775) );
  XNOR U13992 ( .A(n12983), .B(n6492), .Z(n4787) );
  IV U13993 ( .A(n8790), .Z(n6492) );
  XNOR U13994 ( .A(n12984), .B(n11043), .Z(n8790) );
  AND U13995 ( .A(n12701), .B(n8791), .Z(n12983) );
  XNOR U13996 ( .A(n3507), .B(n12985), .Z(n12977) );
  XOR U13997 ( .A(n8785), .B(n4882), .Z(n12985) );
  XNOR U13998 ( .A(n12986), .B(n6487), .Z(n4882) );
  XOR U13999 ( .A(n12987), .B(n12652), .Z(n6487) );
  ANDN U14000 ( .B(n8772), .A(n12716), .Z(n12986) );
  XNOR U14001 ( .A(n12988), .B(n10077), .Z(n12716) );
  XNOR U14002 ( .A(n12989), .B(n11039), .Z(n8772) );
  XOR U14003 ( .A(n12990), .B(n6482), .Z(n8785) );
  XNOR U14004 ( .A(n12991), .B(n9788), .Z(n6482) );
  XNOR U14005 ( .A(n12992), .B(n12993), .Z(n9788) );
  NOR U14006 ( .A(n8768), .B(n8767), .Z(n12990) );
  XOR U14007 ( .A(n10047), .B(n12994), .Z(n8767) );
  IV U14008 ( .A(n10980), .Z(n10047) );
  XNOR U14009 ( .A(n12995), .B(n10842), .Z(n8768) );
  XNOR U14010 ( .A(n12996), .B(n6496), .Z(n3507) );
  XNOR U14011 ( .A(n12997), .B(n9450), .Z(n6496) );
  ANDN U14012 ( .B(n8764), .A(n8765), .Z(n12996) );
  XNOR U14013 ( .A(n12998), .B(n11634), .Z(n8765) );
  XOR U14014 ( .A(n9520), .B(n12999), .Z(n8764) );
  IV U14015 ( .A(n13000), .Z(n9520) );
  XNOR U14016 ( .A(n13001), .B(n13002), .Z(n6339) );
  XOR U14017 ( .A(n5463), .B(n3712), .Z(n13002) );
  XOR U14018 ( .A(n13003), .B(n13004), .Z(n3712) );
  ANDN U14019 ( .B(n6519), .A(n6515), .Z(n13003) );
  XNOR U14020 ( .A(n10950), .B(n13005), .Z(n6519) );
  XNOR U14021 ( .A(n13006), .B(n8803), .Z(n5463) );
  ANDN U14022 ( .B(n6507), .A(n6508), .Z(n13006) );
  XNOR U14023 ( .A(n13007), .B(n11634), .Z(n6508) );
  IV U14024 ( .A(n13008), .Z(n11634) );
  XNOR U14025 ( .A(n10754), .B(n13009), .Z(n6507) );
  XOR U14026 ( .A(n4332), .B(n13010), .Z(n13001) );
  XOR U14027 ( .A(n5915), .B(n2121), .Z(n13010) );
  XOR U14028 ( .A(n13011), .B(n8800), .Z(n2121) );
  ANDN U14029 ( .B(n6521), .A(n6522), .Z(n13011) );
  XNOR U14030 ( .A(n13012), .B(n13013), .Z(n6522) );
  XNOR U14031 ( .A(n13014), .B(n10749), .Z(n6521) );
  XOR U14032 ( .A(n13015), .B(n8812), .Z(n5915) );
  ANDN U14033 ( .B(n6525), .A(n6526), .Z(n13015) );
  XOR U14034 ( .A(n13016), .B(n9949), .Z(n6526) );
  XNOR U14035 ( .A(n13017), .B(n9418), .Z(n6525) );
  XOR U14036 ( .A(n13018), .B(n8808), .Z(n4332) );
  ANDN U14037 ( .B(n6513), .A(n6511), .Z(n13018) );
  IV U14038 ( .A(n8809), .Z(n6511) );
  XOR U14039 ( .A(n13019), .B(n10842), .Z(n8809) );
  XOR U14040 ( .A(n13020), .B(n11827), .Z(n10842) );
  XOR U14041 ( .A(n13021), .B(n13022), .Z(n11827) );
  XNOR U14042 ( .A(n13023), .B(n13024), .Z(n13022) );
  XOR U14043 ( .A(n12188), .B(n13025), .Z(n13021) );
  XNOR U14044 ( .A(n9125), .B(n11229), .Z(n13025) );
  XNOR U14045 ( .A(n13026), .B(n13027), .Z(n11229) );
  AND U14046 ( .A(n13028), .B(n13029), .Z(n13026) );
  XNOR U14047 ( .A(n13030), .B(n13031), .Z(n9125) );
  ANDN U14048 ( .B(n13032), .A(n13033), .Z(n13030) );
  XNOR U14049 ( .A(n13034), .B(n13035), .Z(n12188) );
  ANDN U14050 ( .B(n13036), .A(n13037), .Z(n13034) );
  XOR U14051 ( .A(n9443), .B(n13038), .Z(n6513) );
  IV U14052 ( .A(n11930), .Z(n9443) );
  XNOR U14053 ( .A(n13039), .B(n13040), .Z(n11930) );
  XNOR U14054 ( .A(n13041), .B(n8791), .Z(n8770) );
  XOR U14055 ( .A(n13042), .B(n11955), .Z(n8791) );
  IV U14056 ( .A(n12232), .Z(n11955) );
  NOR U14057 ( .A(n12701), .B(n6490), .Z(n13041) );
  XNOR U14058 ( .A(n13043), .B(n11124), .Z(n6490) );
  XOR U14059 ( .A(n9231), .B(n13044), .Z(n12701) );
  IV U14060 ( .A(n10163), .Z(n9231) );
  XOR U14061 ( .A(n13045), .B(n6220), .Z(out[1003]) );
  XOR U14062 ( .A(n8995), .B(n2292), .Z(n6220) );
  XNOR U14063 ( .A(n6103), .B(n6184), .Z(n2292) );
  XNOR U14064 ( .A(n13046), .B(n13047), .Z(n6184) );
  XNOR U14065 ( .A(n2330), .B(n5480), .Z(n13047) );
  XOR U14066 ( .A(n13048), .B(n7829), .Z(n5480) );
  XNOR U14067 ( .A(n13049), .B(n10125), .Z(n7829) );
  XNOR U14068 ( .A(n12517), .B(n13050), .Z(n10125) );
  XOR U14069 ( .A(n13051), .B(n13052), .Z(n12517) );
  XOR U14070 ( .A(n12766), .B(n10629), .Z(n13052) );
  XOR U14071 ( .A(n13053), .B(n13054), .Z(n10629) );
  ANDN U14072 ( .B(n13055), .A(n13056), .Z(n13053) );
  XNOR U14073 ( .A(n13057), .B(n13058), .Z(n12766) );
  XNOR U14074 ( .A(n12012), .B(n13061), .Z(n13051) );
  XNOR U14075 ( .A(n13062), .B(n13063), .Z(n13061) );
  XOR U14076 ( .A(n13064), .B(n13065), .Z(n12012) );
  NOR U14077 ( .A(n13066), .B(n13067), .Z(n13064) );
  NOR U14078 ( .A(n9005), .B(n7828), .Z(n13048) );
  XOR U14079 ( .A(n13068), .B(n13069), .Z(n7828) );
  XNOR U14080 ( .A(n13070), .B(n9149), .Z(n9005) );
  XNOR U14081 ( .A(n13071), .B(n7833), .Z(n2330) );
  XNOR U14082 ( .A(n13072), .B(n9891), .Z(n7833) );
  NOR U14083 ( .A(n7832), .B(n9000), .Z(n13071) );
  XNOR U14084 ( .A(n11467), .B(n13073), .Z(n9000) );
  XNOR U14085 ( .A(n13074), .B(n12373), .Z(n11467) );
  XOR U14086 ( .A(n13075), .B(n13076), .Z(n12373) );
  XOR U14087 ( .A(n9865), .B(n13077), .Z(n13076) );
  XNOR U14088 ( .A(n13078), .B(n13067), .Z(n9865) );
  ANDN U14089 ( .B(n13079), .A(n13080), .Z(n13078) );
  XOR U14090 ( .A(n11426), .B(n13081), .Z(n13075) );
  XOR U14091 ( .A(n10393), .B(n13082), .Z(n13081) );
  XNOR U14092 ( .A(n13083), .B(n13084), .Z(n10393) );
  NOR U14093 ( .A(n13085), .B(n13086), .Z(n13083) );
  XNOR U14094 ( .A(n13087), .B(n13056), .Z(n11426) );
  NOR U14095 ( .A(n13088), .B(n13089), .Z(n13087) );
  XOR U14096 ( .A(n13090), .B(n10120), .Z(n7832) );
  IV U14097 ( .A(n9336), .Z(n10120) );
  XOR U14098 ( .A(n3169), .B(n13091), .Z(n13046) );
  XNOR U14099 ( .A(n6230), .B(n7822), .Z(n13091) );
  XNOR U14100 ( .A(n13092), .B(n7837), .Z(n7822) );
  XOR U14101 ( .A(n9113), .B(n13093), .Z(n7837) );
  ANDN U14102 ( .B(n9003), .A(n9002), .Z(n13092) );
  IV U14103 ( .A(n7838), .Z(n9002) );
  XNOR U14104 ( .A(n13094), .B(n10727), .Z(n7838) );
  XNOR U14105 ( .A(n13095), .B(n12342), .Z(n10727) );
  XNOR U14106 ( .A(n13096), .B(n13097), .Z(n12342) );
  XNOR U14107 ( .A(n12229), .B(n13098), .Z(n13097) );
  XNOR U14108 ( .A(n13099), .B(n13100), .Z(n12229) );
  NOR U14109 ( .A(n13101), .B(n13102), .Z(n13099) );
  XNOR U14110 ( .A(n10168), .B(n13103), .Z(n13096) );
  XNOR U14111 ( .A(n11304), .B(n11456), .Z(n13103) );
  XOR U14112 ( .A(n13104), .B(n13105), .Z(n11456) );
  AND U14113 ( .A(n13106), .B(n13107), .Z(n13104) );
  XOR U14114 ( .A(n13108), .B(n13109), .Z(n11304) );
  NOR U14115 ( .A(n13110), .B(n13111), .Z(n13108) );
  XNOR U14116 ( .A(n13112), .B(n13113), .Z(n10168) );
  NOR U14117 ( .A(n13114), .B(n13115), .Z(n13112) );
  XOR U14118 ( .A(n9236), .B(n13116), .Z(n9003) );
  XNOR U14119 ( .A(n13117), .B(n13118), .Z(n9236) );
  XOR U14120 ( .A(n13119), .B(n7842), .Z(n6230) );
  XOR U14121 ( .A(n13120), .B(n13121), .Z(n7842) );
  NOR U14122 ( .A(n12888), .B(n7841), .Z(n13119) );
  XNOR U14123 ( .A(n13122), .B(n7845), .Z(n3169) );
  XOR U14124 ( .A(n13123), .B(n10729), .Z(n7845) );
  ANDN U14125 ( .B(n7846), .A(n8997), .Z(n13122) );
  XOR U14126 ( .A(n11637), .B(n13124), .Z(n8997) );
  XOR U14127 ( .A(n13125), .B(n12255), .Z(n7846) );
  XOR U14128 ( .A(n13126), .B(n13127), .Z(n6103) );
  XOR U14129 ( .A(n5289), .B(n1942), .Z(n13127) );
  XOR U14130 ( .A(n13128), .B(n9059), .Z(n1942) );
  AND U14131 ( .A(n7911), .B(n8984), .Z(n13128) );
  XOR U14132 ( .A(n13129), .B(n9912), .Z(n8984) );
  IV U14133 ( .A(n11548), .Z(n9912) );
  XOR U14134 ( .A(n13130), .B(n13131), .Z(n11548) );
  XOR U14135 ( .A(n13132), .B(n11503), .Z(n7911) );
  XNOR U14136 ( .A(n13133), .B(n9064), .Z(n5289) );
  ANDN U14137 ( .B(n8982), .A(n7903), .Z(n13133) );
  XOR U14138 ( .A(n11118), .B(n13134), .Z(n7903) );
  IV U14139 ( .A(n11445), .Z(n11118) );
  XNOR U14140 ( .A(n13135), .B(n12307), .Z(n11445) );
  XNOR U14141 ( .A(n13136), .B(n13137), .Z(n12307) );
  XNOR U14142 ( .A(n13138), .B(n11055), .Z(n13137) );
  XNOR U14143 ( .A(n13139), .B(n13140), .Z(n11055) );
  ANDN U14144 ( .B(n13141), .A(n13142), .Z(n13139) );
  XOR U14145 ( .A(n11612), .B(n13143), .Z(n13136) );
  XNOR U14146 ( .A(n12724), .B(n11743), .Z(n13143) );
  XNOR U14147 ( .A(n13144), .B(n13145), .Z(n11743) );
  AND U14148 ( .A(n13146), .B(n13147), .Z(n13144) );
  XNOR U14149 ( .A(n13148), .B(n13149), .Z(n12724) );
  ANDN U14150 ( .B(n13150), .A(n13151), .Z(n13148) );
  XNOR U14151 ( .A(n13152), .B(n13153), .Z(n11612) );
  NOR U14152 ( .A(n13154), .B(n13155), .Z(n13152) );
  XOR U14153 ( .A(n9238), .B(n13156), .Z(n8982) );
  XOR U14154 ( .A(n3738), .B(n13157), .Z(n13126) );
  XOR U14155 ( .A(n9040), .B(n4204), .Z(n13157) );
  XOR U14156 ( .A(n13158), .B(n9066), .Z(n4204) );
  ANDN U14157 ( .B(n7894), .A(n8992), .Z(n13158) );
  IV U14158 ( .A(n9067), .Z(n8992) );
  XOR U14159 ( .A(n13159), .B(n10331), .Z(n9067) );
  XNOR U14160 ( .A(n13160), .B(n13161), .Z(n10331) );
  XNOR U14161 ( .A(n13162), .B(n10065), .Z(n7894) );
  ANDN U14162 ( .B(n8987), .A(n7898), .Z(n13163) );
  XOR U14163 ( .A(n10209), .B(n13164), .Z(n7898) );
  XOR U14164 ( .A(n9667), .B(n12929), .Z(n8987) );
  XNOR U14165 ( .A(n13165), .B(n13166), .Z(n12929) );
  AND U14166 ( .A(n13167), .B(n13168), .Z(n13165) );
  IV U14167 ( .A(n10869), .Z(n9667) );
  XOR U14168 ( .A(n11587), .B(n12836), .Z(n10869) );
  XOR U14169 ( .A(n13169), .B(n13170), .Z(n12836) );
  XNOR U14170 ( .A(n13171), .B(n11928), .Z(n13170) );
  XNOR U14171 ( .A(n13172), .B(n13173), .Z(n11928) );
  ANDN U14172 ( .B(n12938), .A(n12936), .Z(n13172) );
  XOR U14173 ( .A(n11783), .B(n13174), .Z(n13169) );
  XNOR U14174 ( .A(n11223), .B(n13175), .Z(n13174) );
  XOR U14175 ( .A(n13176), .B(n13177), .Z(n11223) );
  AND U14176 ( .A(n12942), .B(n12940), .Z(n13176) );
  XOR U14177 ( .A(n13178), .B(n13179), .Z(n11783) );
  AND U14178 ( .A(n12932), .B(n12931), .Z(n13178) );
  XOR U14179 ( .A(n13180), .B(n13181), .Z(n11587) );
  XNOR U14180 ( .A(n13182), .B(n11719), .Z(n13181) );
  XOR U14181 ( .A(n13183), .B(n13184), .Z(n11719) );
  ANDN U14182 ( .B(n13185), .A(n13186), .Z(n13183) );
  XNOR U14183 ( .A(n11908), .B(n13187), .Z(n13180) );
  XOR U14184 ( .A(n9566), .B(n12413), .Z(n13187) );
  XOR U14185 ( .A(n13188), .B(n13189), .Z(n12413) );
  ANDN U14186 ( .B(n13190), .A(n13191), .Z(n13188) );
  XOR U14187 ( .A(n13192), .B(n13193), .Z(n9566) );
  ANDN U14188 ( .B(n13194), .A(n13195), .Z(n13192) );
  XOR U14189 ( .A(n13196), .B(n13197), .Z(n11908) );
  ANDN U14190 ( .B(n13198), .A(n13199), .Z(n13196) );
  XNOR U14191 ( .A(n13200), .B(n13201), .Z(n3738) );
  ANDN U14192 ( .B(n8990), .A(n7907), .Z(n13200) );
  XNOR U14193 ( .A(n13202), .B(n10512), .Z(n7907) );
  IV U14194 ( .A(n13203), .Z(n10512) );
  XOR U14195 ( .A(n13204), .B(n7841), .Z(n8995) );
  XOR U14196 ( .A(n13205), .B(n11869), .Z(n7841) );
  ANDN U14197 ( .B(n12888), .A(n8955), .Z(n13204) );
  XOR U14198 ( .A(n13206), .B(n12736), .Z(n8955) );
  IV U14199 ( .A(n11503), .Z(n12736) );
  XNOR U14200 ( .A(n11913), .B(n13207), .Z(n11503) );
  XOR U14201 ( .A(n13208), .B(n13209), .Z(n11913) );
  XNOR U14202 ( .A(n13210), .B(n10404), .Z(n13209) );
  XOR U14203 ( .A(n13211), .B(n13212), .Z(n10404) );
  NOR U14204 ( .A(n13213), .B(n13214), .Z(n13211) );
  XNOR U14205 ( .A(n12405), .B(n13215), .Z(n13208) );
  XNOR U14206 ( .A(n11759), .B(n10299), .Z(n13215) );
  XNOR U14207 ( .A(n13216), .B(n13217), .Z(n10299) );
  ANDN U14208 ( .B(n13218), .A(n13219), .Z(n13216) );
  XNOR U14209 ( .A(n13220), .B(n13221), .Z(n11759) );
  ANDN U14210 ( .B(n13222), .A(n13223), .Z(n13220) );
  XOR U14211 ( .A(n13224), .B(n13225), .Z(n12405) );
  ANDN U14212 ( .B(n13226), .A(n13227), .Z(n13224) );
  XOR U14213 ( .A(n13228), .B(n9413), .Z(n12888) );
  AND U14214 ( .A(n5697), .B(n5699), .Z(n13045) );
  XOR U14215 ( .A(n11396), .B(n2092), .Z(n5699) );
  XNOR U14216 ( .A(n8236), .B(n9604), .Z(n2092) );
  XNOR U14217 ( .A(n13229), .B(n13230), .Z(n9604) );
  XOR U14218 ( .A(n5497), .B(n3633), .Z(n13230) );
  XNOR U14219 ( .A(n13231), .B(n13232), .Z(n3633) );
  ANDN U14220 ( .B(n8362), .A(n8363), .Z(n13231) );
  XOR U14221 ( .A(n10779), .B(n13233), .Z(n8363) );
  IV U14222 ( .A(n11356), .Z(n10779) );
  XOR U14223 ( .A(n13234), .B(n11531), .Z(n5497) );
  ANDN U14224 ( .B(n8358), .A(n8359), .Z(n13234) );
  XNOR U14225 ( .A(n13210), .B(n10300), .Z(n8359) );
  XOR U14226 ( .A(n13235), .B(n13236), .Z(n10300) );
  XNOR U14227 ( .A(n13237), .B(n13238), .Z(n13210) );
  ANDN U14228 ( .B(n13239), .A(n13240), .Z(n13237) );
  XNOR U14229 ( .A(n13241), .B(n11937), .Z(n8358) );
  XOR U14230 ( .A(n6304), .B(n13242), .Z(n13229) );
  XNOR U14231 ( .A(n2377), .B(n5604), .Z(n13242) );
  XNOR U14232 ( .A(n13243), .B(n11542), .Z(n5604) );
  ANDN U14233 ( .B(n9608), .A(n9606), .Z(n13243) );
  XOR U14234 ( .A(n13244), .B(n9793), .Z(n9606) );
  XNOR U14235 ( .A(n13245), .B(n12878), .Z(n9793) );
  XOR U14236 ( .A(n13246), .B(n13247), .Z(n12878) );
  XOR U14237 ( .A(n12113), .B(n11685), .Z(n13247) );
  XNOR U14238 ( .A(n13248), .B(n13249), .Z(n11685) );
  ANDN U14239 ( .B(n13250), .A(n13251), .Z(n13248) );
  XNOR U14240 ( .A(n13252), .B(n13253), .Z(n12113) );
  ANDN U14241 ( .B(n13254), .A(n13255), .Z(n13252) );
  XNOR U14242 ( .A(n11787), .B(n13256), .Z(n13246) );
  XOR U14243 ( .A(n12135), .B(n11728), .Z(n13256) );
  XNOR U14244 ( .A(n13257), .B(n13258), .Z(n11728) );
  ANDN U14245 ( .B(n13259), .A(n13260), .Z(n13257) );
  XNOR U14246 ( .A(n13261), .B(n13262), .Z(n12135) );
  ANDN U14247 ( .B(n13263), .A(n13264), .Z(n13261) );
  XNOR U14248 ( .A(n13265), .B(n13266), .Z(n11787) );
  ANDN U14249 ( .B(n13267), .A(n13268), .Z(n13265) );
  XNOR U14250 ( .A(n13269), .B(n11114), .Z(n9608) );
  XNOR U14251 ( .A(n13270), .B(n11534), .Z(n2377) );
  AND U14252 ( .A(n8348), .B(n8350), .Z(n13270) );
  XOR U14253 ( .A(n9101), .B(n13271), .Z(n8350) );
  XOR U14254 ( .A(n13175), .B(n11224), .Z(n8348) );
  XOR U14255 ( .A(n13272), .B(n13273), .Z(n13175) );
  NOR U14256 ( .A(n13274), .B(n12944), .Z(n13272) );
  XNOR U14257 ( .A(n13275), .B(n11539), .Z(n6304) );
  ANDN U14258 ( .B(n8354), .A(n8352), .Z(n13275) );
  XNOR U14259 ( .A(n13276), .B(n13277), .Z(n8352) );
  XNOR U14260 ( .A(n13278), .B(n11482), .Z(n8354) );
  XNOR U14261 ( .A(n13279), .B(n13280), .Z(n11482) );
  XOR U14262 ( .A(n13281), .B(n13282), .Z(n8236) );
  XOR U14263 ( .A(n3845), .B(n5158), .Z(n13282) );
  XOR U14264 ( .A(n13283), .B(n9501), .Z(n5158) );
  XNOR U14265 ( .A(n13284), .B(n9552), .Z(n9501) );
  ANDN U14266 ( .B(n11403), .A(n11404), .Z(n13283) );
  IV U14267 ( .A(n12907), .Z(n11404) );
  XOR U14268 ( .A(n10934), .B(n13285), .Z(n12907) );
  XNOR U14269 ( .A(n13286), .B(n13287), .Z(n10934) );
  XNOR U14270 ( .A(n13171), .B(n11224), .Z(n11403) );
  IV U14271 ( .A(n11929), .Z(n11224) );
  XOR U14272 ( .A(n13288), .B(n13289), .Z(n11929) );
  XNOR U14273 ( .A(n13290), .B(n13291), .Z(n13171) );
  NOR U14274 ( .A(n13166), .B(n13168), .Z(n13290) );
  IV U14275 ( .A(n13292), .Z(n13166) );
  XNOR U14276 ( .A(n13293), .B(n8296), .Z(n3845) );
  XOR U14277 ( .A(n13294), .B(n12299), .Z(n8296) );
  ANDN U14278 ( .B(n11393), .A(n11394), .Z(n13293) );
  IV U14279 ( .A(n12913), .Z(n11394) );
  XNOR U14280 ( .A(n13082), .B(n9866), .Z(n12913) );
  XNOR U14281 ( .A(n13297), .B(n13060), .Z(n13082) );
  ANDN U14282 ( .B(n13298), .A(n13299), .Z(n13297) );
  XOR U14283 ( .A(n13300), .B(n13301), .Z(n11393) );
  XNOR U14284 ( .A(n4786), .B(n13302), .Z(n13281) );
  XOR U14285 ( .A(n1740), .B(n11516), .Z(n13302) );
  XOR U14286 ( .A(n13303), .B(n8305), .Z(n11516) );
  XOR U14287 ( .A(n13304), .B(n10868), .Z(n8305) );
  ANDN U14288 ( .B(n11390), .A(n11389), .Z(n13303) );
  XNOR U14289 ( .A(n12687), .B(n13307), .Z(n11389) );
  XNOR U14290 ( .A(n12606), .B(n13308), .Z(n12687) );
  XOR U14291 ( .A(n13309), .B(n13310), .Z(n12606) );
  XNOR U14292 ( .A(n13311), .B(n13312), .Z(n13310) );
  XNOR U14293 ( .A(n12438), .B(n13313), .Z(n13309) );
  XOR U14294 ( .A(n9154), .B(n12514), .Z(n13313) );
  XNOR U14295 ( .A(n13314), .B(n13315), .Z(n12514) );
  ANDN U14296 ( .B(n13316), .A(n13317), .Z(n13314) );
  XNOR U14297 ( .A(n13318), .B(n13319), .Z(n9154) );
  ANDN U14298 ( .B(n13320), .A(n13321), .Z(n13318) );
  XOR U14299 ( .A(n13322), .B(n13323), .Z(n12438) );
  XNOR U14300 ( .A(n13326), .B(n10234), .Z(n11390) );
  XNOR U14301 ( .A(n13327), .B(n13328), .Z(n10234) );
  XNOR U14302 ( .A(n13329), .B(n8299), .Z(n1740) );
  XOR U14303 ( .A(n13330), .B(n11511), .Z(n8299) );
  IV U14304 ( .A(n11062), .Z(n11511) );
  NOR U14305 ( .A(n11399), .B(n11400), .Z(n13329) );
  XNOR U14306 ( .A(n13331), .B(n9927), .Z(n11400) );
  XNOR U14307 ( .A(n13332), .B(n9413), .Z(n11399) );
  XOR U14308 ( .A(n13333), .B(n12365), .Z(n9413) );
  XOR U14309 ( .A(n13334), .B(n13335), .Z(n12365) );
  XNOR U14310 ( .A(n13336), .B(n12780), .Z(n13335) );
  XOR U14311 ( .A(n13337), .B(n13338), .Z(n12780) );
  NOR U14312 ( .A(n13339), .B(n13340), .Z(n13337) );
  XOR U14313 ( .A(n13341), .B(n13342), .Z(n13334) );
  XNOR U14314 ( .A(n12312), .B(n11434), .Z(n13342) );
  XNOR U14315 ( .A(n13343), .B(n13344), .Z(n11434) );
  NOR U14316 ( .A(n13345), .B(n13346), .Z(n13343) );
  XNOR U14317 ( .A(n13347), .B(n13348), .Z(n12312) );
  ANDN U14318 ( .B(n13349), .A(n13350), .Z(n13347) );
  XNOR U14319 ( .A(n13351), .B(n8310), .Z(n4786) );
  XOR U14320 ( .A(n13352), .B(n11937), .Z(n8310) );
  ANDN U14321 ( .B(n11524), .A(n12900), .Z(n13351) );
  XOR U14322 ( .A(n13353), .B(n11524), .Z(n11396) );
  XNOR U14323 ( .A(n12796), .B(n9764), .Z(n11524) );
  XOR U14324 ( .A(n13130), .B(n13354), .Z(n9764) );
  XOR U14325 ( .A(n13355), .B(n13356), .Z(n13130) );
  XOR U14326 ( .A(n10825), .B(n12194), .Z(n13356) );
  XOR U14327 ( .A(n13357), .B(n13358), .Z(n12194) );
  AND U14328 ( .A(n13359), .B(n13360), .Z(n13357) );
  XNOR U14329 ( .A(n13361), .B(n13362), .Z(n10825) );
  ANDN U14330 ( .B(n12800), .A(n12798), .Z(n13361) );
  XNOR U14331 ( .A(n9619), .B(n13363), .Z(n13355) );
  XNOR U14332 ( .A(n9510), .B(n12372), .Z(n13363) );
  XOR U14333 ( .A(n13364), .B(n13365), .Z(n12372) );
  ANDN U14334 ( .B(n12955), .A(n12953), .Z(n13364) );
  XNOR U14335 ( .A(n13366), .B(n13367), .Z(n9510) );
  XNOR U14336 ( .A(n13368), .B(n13369), .Z(n9619) );
  ANDN U14337 ( .B(n12810), .A(n12808), .Z(n13368) );
  XOR U14338 ( .A(n13370), .B(n13360), .Z(n12796) );
  ANDN U14339 ( .B(n13371), .A(n13359), .Z(n13370) );
  XNOR U14340 ( .A(n13372), .B(n9136), .Z(n8308) );
  IV U14341 ( .A(n10060), .Z(n9136) );
  XNOR U14342 ( .A(n13373), .B(n13374), .Z(n10060) );
  XOR U14343 ( .A(n13375), .B(n12232), .Z(n12900) );
  XOR U14344 ( .A(n8805), .B(n5179), .Z(n5697) );
  XNOR U14345 ( .A(n13376), .B(n13377), .Z(n6477) );
  XOR U14346 ( .A(n5122), .B(n2521), .Z(n13377) );
  XOR U14347 ( .A(n13378), .B(n6527), .Z(n2521) );
  XOR U14348 ( .A(n13379), .B(n11648), .Z(n6527) );
  ANDN U14349 ( .B(n8812), .A(n8811), .Z(n13378) );
  IV U14350 ( .A(n8861), .Z(n8811) );
  XOR U14351 ( .A(n13380), .B(n10964), .Z(n8861) );
  XNOR U14352 ( .A(n13381), .B(n12706), .Z(n8812) );
  XNOR U14353 ( .A(n13382), .B(n6518), .Z(n5122) );
  XOR U14354 ( .A(n13383), .B(n10067), .Z(n6518) );
  IV U14355 ( .A(n11874), .Z(n10067) );
  XOR U14356 ( .A(n13384), .B(n13385), .Z(n11874) );
  NOR U14357 ( .A(n13386), .B(n13004), .Z(n13382) );
  XNOR U14358 ( .A(n3509), .B(n13387), .Z(n13376) );
  XOR U14359 ( .A(n8849), .B(n4886), .Z(n13387) );
  XOR U14360 ( .A(n13388), .B(n6512), .Z(n4886) );
  XOR U14361 ( .A(n12560), .B(n9142), .Z(n6512) );
  XNOR U14362 ( .A(n13389), .B(n13390), .Z(n12560) );
  NOR U14363 ( .A(n13391), .B(n13392), .Z(n13389) );
  NOR U14364 ( .A(n8854), .B(n8808), .Z(n13388) );
  XNOR U14365 ( .A(n13393), .B(n10182), .Z(n8808) );
  XNOR U14366 ( .A(n13394), .B(n12919), .Z(n10182) );
  XOR U14367 ( .A(n13395), .B(n13396), .Z(n12919) );
  XNOR U14368 ( .A(n10829), .B(n9781), .Z(n13396) );
  XNOR U14369 ( .A(n13397), .B(n13398), .Z(n9781) );
  NOR U14370 ( .A(n13399), .B(n13400), .Z(n13397) );
  XNOR U14371 ( .A(n13401), .B(n13402), .Z(n10829) );
  ANDN U14372 ( .B(n13403), .A(n13404), .Z(n13401) );
  XOR U14373 ( .A(n12948), .B(n13405), .Z(n13395) );
  XOR U14374 ( .A(n13406), .B(n12571), .Z(n13405) );
  XNOR U14375 ( .A(n13407), .B(n13408), .Z(n12571) );
  ANDN U14376 ( .B(n13409), .A(n13410), .Z(n13407) );
  XNOR U14377 ( .A(n13411), .B(n13412), .Z(n12948) );
  ANDN U14378 ( .B(n13413), .A(n13414), .Z(n13411) );
  XOR U14379 ( .A(n13415), .B(n11869), .Z(n8854) );
  XNOR U14380 ( .A(n13416), .B(n6509), .Z(n8849) );
  XNOR U14381 ( .A(n13417), .B(n9886), .Z(n6509) );
  XNOR U14382 ( .A(n13418), .B(n13419), .Z(n9886) );
  ANDN U14383 ( .B(n8802), .A(n8803), .Z(n13416) );
  XNOR U14384 ( .A(n13420), .B(n11099), .Z(n8803) );
  XNOR U14385 ( .A(n9242), .B(n13421), .Z(n8802) );
  XOR U14386 ( .A(n13423), .B(n13424), .Z(n11571) );
  XNOR U14387 ( .A(n13425), .B(n13124), .Z(n13424) );
  XNOR U14388 ( .A(n13426), .B(n13427), .Z(n13124) );
  ANDN U14389 ( .B(n13428), .A(n13429), .Z(n13426) );
  XOR U14390 ( .A(n13430), .B(n13431), .Z(n13423) );
  XNOR U14391 ( .A(n11738), .B(n11638), .Z(n13431) );
  XNOR U14392 ( .A(n13432), .B(n13433), .Z(n11638) );
  ANDN U14393 ( .B(n13434), .A(n13435), .Z(n13432) );
  XNOR U14394 ( .A(n13436), .B(n13437), .Z(n11738) );
  NOR U14395 ( .A(n13438), .B(n13439), .Z(n13436) );
  XNOR U14396 ( .A(n13440), .B(n6523), .Z(n3509) );
  XOR U14397 ( .A(n13441), .B(n9547), .Z(n6523) );
  XNOR U14398 ( .A(n13442), .B(n12765), .Z(n9547) );
  XNOR U14399 ( .A(n13443), .B(n13444), .Z(n12765) );
  XNOR U14400 ( .A(n12811), .B(n9965), .Z(n13444) );
  XNOR U14401 ( .A(n13445), .B(n13446), .Z(n9965) );
  ANDN U14402 ( .B(n13447), .A(n13448), .Z(n13445) );
  XNOR U14403 ( .A(n13449), .B(n13450), .Z(n12811) );
  ANDN U14404 ( .B(n13451), .A(n13452), .Z(n13449) );
  XOR U14405 ( .A(n13453), .B(n13454), .Z(n13443) );
  XNOR U14406 ( .A(n9228), .B(n12276), .Z(n13454) );
  XNOR U14407 ( .A(n13455), .B(n13456), .Z(n12276) );
  ANDN U14408 ( .B(n13457), .A(n13458), .Z(n13455) );
  XNOR U14409 ( .A(n13459), .B(n13460), .Z(n9228) );
  AND U14410 ( .A(n13461), .B(n13462), .Z(n13459) );
  NOR U14411 ( .A(n8859), .B(n8800), .Z(n13440) );
  XNOR U14412 ( .A(n13463), .B(n11960), .Z(n8800) );
  XNOR U14413 ( .A(n13464), .B(n9636), .Z(n8859) );
  XOR U14414 ( .A(n13465), .B(n13466), .Z(n6343) );
  XOR U14415 ( .A(n5469), .B(n3717), .Z(n13466) );
  XOR U14416 ( .A(n13467), .B(n13468), .Z(n3717) );
  ANDN U14417 ( .B(n6543), .A(n6544), .Z(n13467) );
  XNOR U14418 ( .A(n13469), .B(n10964), .Z(n6544) );
  XNOR U14419 ( .A(n13470), .B(n8869), .Z(n5469) );
  ANDN U14420 ( .B(n6534), .A(n6535), .Z(n13470) );
  XNOR U14421 ( .A(n13471), .B(n11960), .Z(n6535) );
  XNOR U14422 ( .A(n13472), .B(n13277), .Z(n6534) );
  XNOR U14423 ( .A(n4334), .B(n13473), .Z(n13465) );
  XOR U14424 ( .A(n5920), .B(n2125), .Z(n13473) );
  XOR U14425 ( .A(n13474), .B(n8866), .Z(n2125) );
  ANDN U14426 ( .B(n6548), .A(n6547), .Z(n13474) );
  XOR U14427 ( .A(n9506), .B(n13475), .Z(n6547) );
  IV U14428 ( .A(n12329), .Z(n9506) );
  XNOR U14429 ( .A(n13476), .B(n10637), .Z(n6548) );
  IV U14430 ( .A(n13477), .Z(n10637) );
  XNOR U14431 ( .A(n13478), .B(n8879), .Z(n5920) );
  IV U14432 ( .A(n13479), .Z(n8879) );
  ANDN U14433 ( .B(n6551), .A(n8925), .Z(n13478) );
  XNOR U14434 ( .A(n13480), .B(n11902), .Z(n8925) );
  IV U14435 ( .A(n8878), .Z(n6551) );
  XOR U14436 ( .A(n9138), .B(n13481), .Z(n8878) );
  XOR U14437 ( .A(n13482), .B(n8874), .Z(n4334) );
  NOR U14438 ( .A(n8875), .B(n6539), .Z(n13482) );
  XOR U14439 ( .A(n13483), .B(n9552), .Z(n6539) );
  XNOR U14440 ( .A(n13484), .B(n13485), .Z(n9552) );
  XOR U14441 ( .A(n13486), .B(n11099), .Z(n8875) );
  XOR U14442 ( .A(n13487), .B(n11898), .Z(n11099) );
  XOR U14443 ( .A(n13488), .B(n13489), .Z(n11898) );
  XOR U14444 ( .A(n13490), .B(n12308), .Z(n13489) );
  XOR U14445 ( .A(n13491), .B(n13492), .Z(n12308) );
  ANDN U14446 ( .B(n13493), .A(n13494), .Z(n13491) );
  XOR U14447 ( .A(n12339), .B(n13495), .Z(n13488) );
  XNOR U14448 ( .A(n9108), .B(n11353), .Z(n13495) );
  XNOR U14449 ( .A(n13496), .B(n13497), .Z(n11353) );
  ANDN U14450 ( .B(n13498), .A(n13499), .Z(n13496) );
  XNOR U14451 ( .A(n13500), .B(n13501), .Z(n9108) );
  ANDN U14452 ( .B(n13502), .A(n13503), .Z(n13500) );
  ANDN U14453 ( .B(n13506), .A(n13507), .Z(n13504) );
  XNOR U14454 ( .A(n13508), .B(n8857), .Z(n8805) );
  IV U14455 ( .A(n13386), .Z(n8857) );
  XNOR U14456 ( .A(n13509), .B(n12117), .Z(n13386) );
  XOR U14457 ( .A(n12096), .B(n13510), .Z(n6515) );
  IV U14458 ( .A(n11244), .Z(n12096) );
  XNOR U14459 ( .A(n13511), .B(n13512), .Z(n11244) );
  XNOR U14460 ( .A(n13513), .B(n10269), .Z(n13004) );
  XOR U14461 ( .A(n13514), .B(n6225), .Z(out[1002]) );
  XOR U14462 ( .A(n9057), .B(n2299), .Z(n6225) );
  XNOR U14463 ( .A(n6108), .B(n6189), .Z(n2299) );
  XNOR U14464 ( .A(n13515), .B(n13516), .Z(n6189) );
  XNOR U14465 ( .A(n2337), .B(n5486), .Z(n13516) );
  XNOR U14466 ( .A(n13517), .B(n7896), .Z(n5486) );
  XNOR U14467 ( .A(n13518), .B(n10231), .Z(n7896) );
  XOR U14468 ( .A(n13354), .B(n12773), .Z(n10231) );
  XOR U14469 ( .A(n13519), .B(n13520), .Z(n12773) );
  XNOR U14470 ( .A(n12961), .B(n10758), .Z(n13520) );
  XOR U14471 ( .A(n13521), .B(n13522), .Z(n10758) );
  AND U14472 ( .A(n13523), .B(n13524), .Z(n13521) );
  XNOR U14473 ( .A(n13525), .B(n13526), .Z(n12961) );
  NOR U14474 ( .A(n13527), .B(n13528), .Z(n13525) );
  XOR U14475 ( .A(n12168), .B(n13529), .Z(n13519) );
  XOR U14476 ( .A(n13530), .B(n13531), .Z(n13529) );
  XNOR U14477 ( .A(n13532), .B(n13533), .Z(n12168) );
  ANDN U14478 ( .B(n13534), .A(n13535), .Z(n13532) );
  XOR U14479 ( .A(n13536), .B(n13537), .Z(n13354) );
  XNOR U14480 ( .A(n12236), .B(n13073), .Z(n13537) );
  XNOR U14481 ( .A(n13538), .B(n13086), .Z(n13073) );
  ANDN U14482 ( .B(n13085), .A(n13539), .Z(n13538) );
  NOR U14483 ( .A(n13541), .B(n13065), .Z(n13540) );
  XOR U14484 ( .A(n11468), .B(n13542), .Z(n13536) );
  XOR U14485 ( .A(n12697), .B(n12704), .Z(n13542) );
  XNOR U14486 ( .A(n13543), .B(n13089), .Z(n12704) );
  ANDN U14487 ( .B(n13088), .A(n13054), .Z(n13543) );
  XNOR U14488 ( .A(n13544), .B(n13545), .Z(n12697) );
  NOR U14489 ( .A(n13546), .B(n13547), .Z(n13544) );
  XOR U14490 ( .A(n13548), .B(n13298), .Z(n11468) );
  ANDN U14491 ( .B(n13058), .A(n13549), .Z(n13548) );
  ANDN U14492 ( .B(n7895), .A(n9066), .Z(n13517) );
  XOR U14493 ( .A(n13550), .B(n9244), .Z(n9066) );
  XNOR U14494 ( .A(n13551), .B(n13477), .Z(n7895) );
  XNOR U14495 ( .A(n13552), .B(n8988), .Z(n2337) );
  XNOR U14496 ( .A(n13553), .B(n9149), .Z(n8988) );
  XOR U14497 ( .A(n13554), .B(n13555), .Z(n9149) );
  ANDN U14498 ( .B(n7900), .A(n9062), .Z(n13552) );
  XOR U14499 ( .A(n13556), .B(n13008), .Z(n9062) );
  XNOR U14500 ( .A(n12516), .B(n13328), .Z(n13008) );
  XNOR U14501 ( .A(n13557), .B(n13558), .Z(n13328) );
  XNOR U14502 ( .A(n11585), .B(n12118), .Z(n13558) );
  XNOR U14503 ( .A(n13559), .B(n13560), .Z(n12118) );
  XOR U14504 ( .A(n13563), .B(n13564), .Z(n11585) );
  ANDN U14505 ( .B(n13565), .A(n13566), .Z(n13563) );
  XOR U14506 ( .A(n13567), .B(n13568), .Z(n13557) );
  XNOR U14507 ( .A(n11794), .B(n13569), .Z(n13568) );
  XOR U14508 ( .A(n13570), .B(n13571), .Z(n11794) );
  ANDN U14509 ( .B(n13572), .A(n13573), .Z(n13570) );
  XOR U14510 ( .A(n13574), .B(n13575), .Z(n12516) );
  XNOR U14511 ( .A(n9931), .B(n13576), .Z(n13575) );
  XOR U14512 ( .A(n13577), .B(n13535), .Z(n9931) );
  ANDN U14513 ( .B(n13578), .A(n13579), .Z(n13577) );
  XOR U14514 ( .A(n11562), .B(n13580), .Z(n13574) );
  XOR U14515 ( .A(n10596), .B(n13581), .Z(n13580) );
  XOR U14516 ( .A(n13582), .B(n13583), .Z(n10596) );
  XNOR U14517 ( .A(n13586), .B(n13524), .Z(n11562) );
  ANDN U14518 ( .B(n13587), .A(n13588), .Z(n13586) );
  XNOR U14519 ( .A(n13589), .B(n10219), .Z(n7900) );
  IV U14520 ( .A(n10113), .Z(n10219) );
  XNOR U14521 ( .A(n3172), .B(n13590), .Z(n13515) );
  XOR U14522 ( .A(n6277), .B(n7889), .Z(n13590) );
  XNOR U14523 ( .A(n13591), .B(n7904), .Z(n7889) );
  XNOR U14524 ( .A(n13592), .B(n9274), .Z(n7904) );
  ANDN U14525 ( .B(n9064), .A(n7905), .Z(n13591) );
  XOR U14526 ( .A(n10950), .B(n13593), .Z(n7905) );
  IV U14527 ( .A(n11814), .Z(n10950) );
  XNOR U14528 ( .A(n13594), .B(n13595), .Z(n11814) );
  XOR U14529 ( .A(n13596), .B(n12381), .Z(n9064) );
  XNOR U14530 ( .A(n13597), .B(n7909), .Z(n6277) );
  XOR U14531 ( .A(n12558), .B(n9142), .Z(n7909) );
  XOR U14532 ( .A(n13598), .B(n13599), .Z(n12468) );
  XOR U14533 ( .A(n12049), .B(n13600), .Z(n13599) );
  XNOR U14534 ( .A(n13601), .B(n13602), .Z(n12049) );
  ANDN U14535 ( .B(n12553), .A(n12554), .Z(n13601) );
  IV U14536 ( .A(n13603), .Z(n12554) );
  XNOR U14537 ( .A(n9321), .B(n13604), .Z(n13598) );
  XOR U14538 ( .A(n9902), .B(n12710), .Z(n13604) );
  XNOR U14539 ( .A(n13605), .B(n13606), .Z(n12710) );
  ANDN U14540 ( .B(n12538), .A(n13607), .Z(n13605) );
  XNOR U14541 ( .A(n13608), .B(n13609), .Z(n9902) );
  NOR U14542 ( .A(n12549), .B(n12550), .Z(n13608) );
  XOR U14543 ( .A(n13610), .B(n13611), .Z(n9321) );
  AND U14544 ( .A(n12542), .B(n12540), .Z(n13610) );
  XOR U14545 ( .A(n13612), .B(n13613), .Z(n11122) );
  XNOR U14546 ( .A(n11895), .B(n11961), .Z(n13613) );
  XNOR U14547 ( .A(n13614), .B(n13615), .Z(n11961) );
  ANDN U14548 ( .B(n12872), .A(n13616), .Z(n13614) );
  XOR U14549 ( .A(n13617), .B(n13618), .Z(n11895) );
  NOR U14550 ( .A(n13619), .B(n13390), .Z(n13617) );
  XOR U14551 ( .A(n10747), .B(n13620), .Z(n13612) );
  XOR U14552 ( .A(n9770), .B(n11643), .Z(n13620) );
  XOR U14553 ( .A(n13621), .B(n13622), .Z(n11643) );
  ANDN U14554 ( .B(n12569), .A(n12567), .Z(n13621) );
  XOR U14555 ( .A(n13623), .B(n13624), .Z(n9770) );
  NOR U14556 ( .A(n12565), .B(n12563), .Z(n13623) );
  XNOR U14557 ( .A(n13625), .B(n13626), .Z(n10747) );
  NOR U14558 ( .A(n13627), .B(n13628), .Z(n13625) );
  XNOR U14559 ( .A(n13629), .B(n13627), .Z(n12558) );
  AND U14560 ( .A(n13630), .B(n13628), .Z(n13629) );
  ANDN U14561 ( .B(n13201), .A(n7908), .Z(n13597) );
  XOR U14562 ( .A(n13631), .B(n7912), .Z(n3172) );
  XOR U14563 ( .A(n11501), .B(n13632), .Z(n7912) );
  XNOR U14564 ( .A(n13633), .B(n13634), .Z(n11501) );
  ANDN U14565 ( .B(n7913), .A(n9059), .Z(n13631) );
  XOR U14566 ( .A(n11111), .B(n13635), .Z(n9059) );
  XOR U14567 ( .A(n12424), .B(n13636), .Z(n7913) );
  XOR U14568 ( .A(n13637), .B(n13638), .Z(n6108) );
  XNOR U14569 ( .A(n5292), .B(n1947), .Z(n13638) );
  XOR U14570 ( .A(n13639), .B(n9160), .Z(n1947) );
  NOR U14571 ( .A(n8019), .B(n9046), .Z(n13639) );
  XOR U14572 ( .A(n13640), .B(n9978), .Z(n9046) );
  XNOR U14573 ( .A(n13641), .B(n11614), .Z(n8019) );
  XOR U14574 ( .A(n13642), .B(n9165), .Z(n5292) );
  ANDN U14575 ( .B(n8011), .A(n9166), .Z(n13642) );
  XNOR U14576 ( .A(n13643), .B(n12713), .Z(n9166) );
  XOR U14577 ( .A(n13644), .B(n10836), .Z(n8011) );
  XNOR U14578 ( .A(n13645), .B(n13646), .Z(n10836) );
  XOR U14579 ( .A(n3742), .B(n13647), .Z(n13637) );
  XNOR U14580 ( .A(n9155), .B(n4207), .Z(n13647) );
  XNOR U14581 ( .A(n13648), .B(n9168), .Z(n4207) );
  ANDN U14582 ( .B(n8002), .A(n9054), .Z(n13648) );
  XNOR U14583 ( .A(n13649), .B(n13203), .Z(n9054) );
  XNOR U14584 ( .A(n13650), .B(n13651), .Z(n13203) );
  XOR U14585 ( .A(n9527), .B(n13652), .Z(n8002) );
  XNOR U14586 ( .A(n13653), .B(n9163), .Z(n9155) );
  AND U14587 ( .A(n9049), .B(n8006), .Z(n13653) );
  XOR U14588 ( .A(n13654), .B(n10343), .Z(n8006) );
  XNOR U14589 ( .A(n13655), .B(n11825), .Z(n9049) );
  IV U14590 ( .A(n9813), .Z(n11825) );
  XOR U14591 ( .A(n11726), .B(n13118), .Z(n9813) );
  XNOR U14592 ( .A(n13656), .B(n13657), .Z(n13118) );
  XNOR U14593 ( .A(n13658), .B(n12093), .Z(n13657) );
  XNOR U14594 ( .A(n13659), .B(n13660), .Z(n12093) );
  ANDN U14595 ( .B(n13661), .A(n13193), .Z(n13659) );
  XOR U14596 ( .A(n13662), .B(n13663), .Z(n13656) );
  XOR U14597 ( .A(n10874), .B(n11347), .Z(n13663) );
  XNOR U14598 ( .A(n13664), .B(n13665), .Z(n11347) );
  ANDN U14599 ( .B(n13666), .A(n13197), .Z(n13664) );
  XNOR U14600 ( .A(n13667), .B(n13668), .Z(n10874) );
  AND U14601 ( .A(n13184), .B(n13669), .Z(n13667) );
  XOR U14602 ( .A(n13670), .B(n13671), .Z(n11726) );
  XNOR U14603 ( .A(n12069), .B(n10086), .Z(n13671) );
  XOR U14604 ( .A(n13672), .B(n13673), .Z(n10086) );
  NOR U14605 ( .A(n13674), .B(n13675), .Z(n13672) );
  XOR U14606 ( .A(n13676), .B(n13677), .Z(n12069) );
  XOR U14607 ( .A(n11279), .B(n13680), .Z(n13670) );
  XOR U14608 ( .A(n9670), .B(n12644), .Z(n13680) );
  XNOR U14609 ( .A(n13681), .B(n13682), .Z(n12644) );
  ANDN U14610 ( .B(n13683), .A(n13684), .Z(n13681) );
  XOR U14611 ( .A(n13685), .B(n13686), .Z(n9670) );
  ANDN U14612 ( .B(n13687), .A(n13688), .Z(n13685) );
  XOR U14613 ( .A(n13689), .B(n13690), .Z(n11279) );
  ANDN U14614 ( .B(n13691), .A(n13692), .Z(n13689) );
  XNOR U14615 ( .A(n13693), .B(n13694), .Z(n3742) );
  ANDN U14616 ( .B(n8015), .A(n9052), .Z(n13693) );
  IV U14617 ( .A(n13695), .Z(n9052) );
  XOR U14618 ( .A(n12447), .B(n11942), .Z(n8015) );
  XOR U14619 ( .A(n13696), .B(n13697), .Z(n12447) );
  ANDN U14620 ( .B(n13698), .A(n13699), .Z(n13696) );
  XOR U14621 ( .A(n13700), .B(n7908), .Z(n9057) );
  XNOR U14622 ( .A(n11301), .B(n13701), .Z(n7908) );
  NOR U14623 ( .A(n13201), .B(n8990), .Z(n13700) );
  XOR U14624 ( .A(n13702), .B(n11614), .Z(n8990) );
  XNOR U14625 ( .A(n13703), .B(n11176), .Z(n11614) );
  XNOR U14626 ( .A(n13704), .B(n13705), .Z(n11176) );
  XOR U14627 ( .A(n13706), .B(n10607), .Z(n13705) );
  XNOR U14628 ( .A(n13707), .B(n13708), .Z(n10607) );
  NOR U14629 ( .A(n13709), .B(n13710), .Z(n13707) );
  XNOR U14630 ( .A(n10400), .B(n13711), .Z(n13704) );
  XNOR U14631 ( .A(n11107), .B(n12637), .Z(n13711) );
  XNOR U14632 ( .A(n13712), .B(n13713), .Z(n12637) );
  ANDN U14633 ( .B(n13714), .A(n13715), .Z(n13712) );
  XNOR U14634 ( .A(n13716), .B(n13717), .Z(n11107) );
  ANDN U14635 ( .B(n13718), .A(n13719), .Z(n13716) );
  XOR U14636 ( .A(n13720), .B(n13721), .Z(n10400) );
  ANDN U14637 ( .B(n13722), .A(n13723), .Z(n13720) );
  XNOR U14638 ( .A(n9509), .B(n13724), .Z(n13201) );
  IV U14639 ( .A(n9804), .Z(n9509) );
  ANDN U14640 ( .B(n5701), .A(n5703), .Z(n13514) );
  XOR U14641 ( .A(n11535), .B(n2095), .Z(n5703) );
  XNOR U14642 ( .A(n8290), .B(n9712), .Z(n2095) );
  XNOR U14643 ( .A(n13725), .B(n13726), .Z(n9712) );
  XNOR U14644 ( .A(n5501), .B(n3638), .Z(n13726) );
  XOR U14645 ( .A(n13727), .B(n13728), .Z(n3638) );
  ANDN U14646 ( .B(n8417), .A(n8419), .Z(n13727) );
  XOR U14647 ( .A(n12527), .B(n13729), .Z(n8419) );
  XNOR U14648 ( .A(n13730), .B(n13731), .Z(n12527) );
  XNOR U14649 ( .A(n13732), .B(n11664), .Z(n5501) );
  ANDN U14650 ( .B(n8414), .A(n8413), .Z(n13732) );
  IV U14651 ( .A(n11665), .Z(n8413) );
  XNOR U14652 ( .A(n13733), .B(n12099), .Z(n11665) );
  XOR U14653 ( .A(n10399), .B(n13706), .Z(n8414) );
  XNOR U14654 ( .A(n13734), .B(n13735), .Z(n13706) );
  NOR U14655 ( .A(n13736), .B(n13737), .Z(n13734) );
  XNOR U14656 ( .A(n13738), .B(n12992), .Z(n10399) );
  XOR U14657 ( .A(n13739), .B(n13740), .Z(n12992) );
  XOR U14658 ( .A(n13741), .B(n9663), .Z(n13740) );
  XNOR U14659 ( .A(n13742), .B(n13743), .Z(n9663) );
  ANDN U14660 ( .B(n13744), .A(n13745), .Z(n13742) );
  XOR U14661 ( .A(n11892), .B(n13746), .Z(n13739) );
  XOR U14662 ( .A(n10508), .B(n11292), .Z(n13746) );
  XOR U14663 ( .A(n13747), .B(n13748), .Z(n11292) );
  ANDN U14664 ( .B(n13749), .A(n13750), .Z(n13747) );
  XOR U14665 ( .A(n13751), .B(n13752), .Z(n10508) );
  ANDN U14666 ( .B(n13753), .A(n13754), .Z(n13751) );
  XNOR U14667 ( .A(n13755), .B(n13756), .Z(n11892) );
  ANDN U14668 ( .B(n13757), .A(n13758), .Z(n13755) );
  XOR U14669 ( .A(n6308), .B(n13759), .Z(n13725) );
  XOR U14670 ( .A(n2388), .B(n5648), .Z(n13759) );
  XNOR U14671 ( .A(n13760), .B(n11677), .Z(n5648) );
  ANDN U14672 ( .B(n9716), .A(n11678), .Z(n13760) );
  XNOR U14673 ( .A(n13761), .B(n9893), .Z(n11678) );
  XNOR U14674 ( .A(n13762), .B(n13161), .Z(n9893) );
  XNOR U14675 ( .A(n13763), .B(n13764), .Z(n13161) );
  XNOR U14676 ( .A(n12241), .B(n12018), .Z(n13764) );
  XNOR U14677 ( .A(n13765), .B(n13766), .Z(n12018) );
  ANDN U14678 ( .B(n13767), .A(n13768), .Z(n13765) );
  XNOR U14679 ( .A(n13769), .B(n13770), .Z(n12241) );
  ANDN U14680 ( .B(n13771), .A(n13772), .Z(n13769) );
  XOR U14681 ( .A(n12076), .B(n13773), .Z(n13763) );
  XOR U14682 ( .A(n11757), .B(n12264), .Z(n13773) );
  XNOR U14683 ( .A(n13774), .B(n13775), .Z(n12264) );
  ANDN U14684 ( .B(n13776), .A(n13777), .Z(n13774) );
  XOR U14685 ( .A(n13778), .B(n13779), .Z(n11757) );
  ANDN U14686 ( .B(n13780), .A(n13781), .Z(n13778) );
  XNOR U14687 ( .A(n13782), .B(n13783), .Z(n12076) );
  ANDN U14688 ( .B(n13784), .A(n13785), .Z(n13782) );
  XOR U14689 ( .A(n13786), .B(n11239), .Z(n9716) );
  XNOR U14690 ( .A(n13787), .B(n11669), .Z(n2388) );
  ANDN U14691 ( .B(n8404), .A(n8403), .Z(n13787) );
  IV U14692 ( .A(n11668), .Z(n8403) );
  XOR U14693 ( .A(n12092), .B(n13662), .Z(n11668) );
  XNOR U14694 ( .A(n13788), .B(n13789), .Z(n13662) );
  AND U14695 ( .A(n13790), .B(n13791), .Z(n13788) );
  XNOR U14696 ( .A(n13792), .B(n9260), .Z(n8404) );
  XNOR U14697 ( .A(n13793), .B(n11674), .Z(n6308) );
  ANDN U14698 ( .B(n8409), .A(n8407), .Z(n13793) );
  XOR U14699 ( .A(n13794), .B(n11704), .Z(n8407) );
  XOR U14700 ( .A(n13795), .B(n11630), .Z(n8409) );
  XNOR U14701 ( .A(n13796), .B(n13797), .Z(n11630) );
  XOR U14702 ( .A(n13798), .B(n13799), .Z(n8290) );
  XNOR U14703 ( .A(n3849), .B(n5160), .Z(n13799) );
  XOR U14704 ( .A(n13800), .B(n9607), .Z(n5160) );
  XNOR U14705 ( .A(n13801), .B(n9808), .Z(n9607) );
  XOR U14706 ( .A(n12092), .B(n13658), .Z(n11541) );
  XOR U14707 ( .A(n13802), .B(n13803), .Z(n13658) );
  ANDN U14708 ( .B(n13189), .A(n13804), .Z(n13802) );
  IV U14709 ( .A(n10873), .Z(n12092) );
  XOR U14710 ( .A(n12646), .B(n13805), .Z(n10873) );
  XOR U14711 ( .A(n13806), .B(n13807), .Z(n12646) );
  XOR U14712 ( .A(n13808), .B(n11086), .Z(n13807) );
  XNOR U14713 ( .A(n13809), .B(n13810), .Z(n11086) );
  NOR U14714 ( .A(n13679), .B(n13677), .Z(n13809) );
  XNOR U14715 ( .A(n12388), .B(n13811), .Z(n13806) );
  XOR U14716 ( .A(n11797), .B(n9909), .Z(n13811) );
  XOR U14717 ( .A(n13812), .B(n13813), .Z(n9909) );
  ANDN U14718 ( .B(n13690), .A(n13691), .Z(n13812) );
  XOR U14719 ( .A(n13814), .B(n13815), .Z(n11797) );
  NOR U14720 ( .A(n13687), .B(n13686), .Z(n13814) );
  XNOR U14721 ( .A(n13816), .B(n13817), .Z(n12388) );
  ANDN U14722 ( .B(n13674), .A(n13818), .Z(n13816) );
  XNOR U14723 ( .A(n13819), .B(n9949), .Z(n11542) );
  XOR U14724 ( .A(n13820), .B(n8349), .Z(n3849) );
  XOR U14725 ( .A(n10209), .B(n13821), .Z(n8349) );
  XNOR U14726 ( .A(n10722), .B(n13822), .Z(n10209) );
  XNOR U14727 ( .A(n13823), .B(n13824), .Z(n10722) );
  XNOR U14728 ( .A(n13825), .B(n11620), .Z(n13824) );
  XNOR U14729 ( .A(n13826), .B(n13827), .Z(n11620) );
  NOR U14730 ( .A(n13828), .B(n13829), .Z(n13826) );
  XOR U14731 ( .A(n10074), .B(n13830), .Z(n13823) );
  XOR U14732 ( .A(n11772), .B(n13831), .Z(n13830) );
  XOR U14733 ( .A(n13832), .B(n13833), .Z(n11772) );
  NOR U14734 ( .A(n13834), .B(n13835), .Z(n13832) );
  XNOR U14735 ( .A(n13836), .B(n13837), .Z(n10074) );
  ANDN U14736 ( .B(n13838), .A(n13839), .Z(n13836) );
  ANDN U14737 ( .B(n11534), .A(n11533), .Z(n13820) );
  XOR U14738 ( .A(n13840), .B(n10185), .Z(n11533) );
  XOR U14739 ( .A(n13581), .B(n9932), .Z(n11534) );
  XOR U14740 ( .A(n13841), .B(n13528), .Z(n13581) );
  ANDN U14741 ( .B(n13842), .A(n13843), .Z(n13841) );
  XOR U14742 ( .A(n5123), .B(n13844), .Z(n13798) );
  XNOR U14743 ( .A(n1744), .B(n11649), .Z(n13844) );
  XNOR U14744 ( .A(n13845), .B(n8360), .Z(n11649) );
  XNOR U14745 ( .A(n13846), .B(n10985), .Z(n8360) );
  XNOR U14746 ( .A(n12596), .B(n13847), .Z(n10985) );
  XOR U14747 ( .A(n13848), .B(n13849), .Z(n12596) );
  XOR U14748 ( .A(n13850), .B(n9430), .Z(n13849) );
  XNOR U14749 ( .A(n13851), .B(n13852), .Z(n9430) );
  ANDN U14750 ( .B(n13853), .A(n13854), .Z(n13851) );
  XNOR U14751 ( .A(n13855), .B(n13856), .Z(n13848) );
  XNOR U14752 ( .A(n10479), .B(n12340), .Z(n13856) );
  XNOR U14753 ( .A(n13857), .B(n13858), .Z(n12340) );
  XOR U14754 ( .A(n13861), .B(n13862), .Z(n10479) );
  NOR U14755 ( .A(n13863), .B(n13864), .Z(n13861) );
  XOR U14756 ( .A(n10386), .B(n13865), .Z(n11531) );
  XNOR U14757 ( .A(n13866), .B(n13867), .Z(n10386) );
  XOR U14758 ( .A(n13868), .B(n11039), .Z(n11530) );
  XOR U14759 ( .A(n13040), .B(n13869), .Z(n11039) );
  XOR U14760 ( .A(n13870), .B(n13871), .Z(n13040) );
  XOR U14761 ( .A(n10102), .B(n12066), .Z(n13871) );
  XOR U14762 ( .A(n13872), .B(n13873), .Z(n12066) );
  ANDN U14763 ( .B(n13874), .A(n13323), .Z(n13872) );
  XNOR U14764 ( .A(n13875), .B(n13876), .Z(n10102) );
  ANDN U14765 ( .B(n13877), .A(n13878), .Z(n13875) );
  XNOR U14766 ( .A(n10333), .B(n13879), .Z(n13870) );
  XNOR U14767 ( .A(n11884), .B(n10972), .Z(n13879) );
  XNOR U14768 ( .A(n13880), .B(n13881), .Z(n10972) );
  AND U14769 ( .A(n13882), .B(n13883), .Z(n13880) );
  XOR U14770 ( .A(n13884), .B(n13885), .Z(n11884) );
  AND U14771 ( .A(n13319), .B(n13886), .Z(n13884) );
  XOR U14772 ( .A(n13887), .B(n13888), .Z(n10333) );
  ANDN U14773 ( .B(n13889), .A(n13890), .Z(n13887) );
  XOR U14774 ( .A(n13891), .B(n8353), .Z(n1744) );
  XOR U14775 ( .A(n13892), .B(n10296), .Z(n8353) );
  IV U14776 ( .A(n11855), .Z(n10296) );
  XOR U14777 ( .A(n13487), .B(n13893), .Z(n11855) );
  XOR U14778 ( .A(n13894), .B(n13895), .Z(n13487) );
  XOR U14779 ( .A(n12980), .B(n11589), .Z(n13895) );
  XOR U14780 ( .A(n13896), .B(n13897), .Z(n11589) );
  ANDN U14781 ( .B(n13031), .A(n13898), .Z(n13896) );
  XNOR U14782 ( .A(n13899), .B(n13900), .Z(n12980) );
  ANDN U14783 ( .B(n13027), .A(n13901), .Z(n13899) );
  XOR U14784 ( .A(n12398), .B(n13902), .Z(n13894) );
  XOR U14785 ( .A(n11514), .B(n13903), .Z(n13902) );
  XNOR U14786 ( .A(n13904), .B(n13905), .Z(n11514) );
  ANDN U14787 ( .B(n13035), .A(n13906), .Z(n13904) );
  XNOR U14788 ( .A(n13907), .B(n13908), .Z(n12398) );
  ANDN U14789 ( .B(n13909), .A(n13910), .Z(n13907) );
  NOR U14790 ( .A(n11539), .B(n11538), .Z(n13891) );
  XOR U14791 ( .A(n9804), .B(n13911), .Z(n11538) );
  XNOR U14792 ( .A(n13912), .B(n13913), .Z(n9804) );
  XOR U14793 ( .A(n13914), .B(n10080), .Z(n11539) );
  XNOR U14794 ( .A(n13915), .B(n8364), .Z(n5123) );
  IV U14795 ( .A(n11657), .Z(n8364) );
  XOR U14796 ( .A(n13916), .B(n12099), .Z(n11657) );
  NOR U14797 ( .A(n13232), .B(n11656), .Z(n13915) );
  IV U14798 ( .A(n13917), .Z(n13232) );
  XNOR U14799 ( .A(n13918), .B(n11656), .Z(n11535) );
  XOR U14800 ( .A(n13077), .B(n9866), .Z(n11656) );
  XNOR U14801 ( .A(n13919), .B(n13920), .Z(n9866) );
  XNOR U14802 ( .A(n13921), .B(n13922), .Z(n13077) );
  ANDN U14803 ( .B(n13545), .A(n13923), .Z(n13921) );
  NOR U14804 ( .A(n13917), .B(n8362), .Z(n13918) );
  XNOR U14805 ( .A(n10163), .B(n13924), .Z(n8362) );
  XOR U14806 ( .A(n13555), .B(n13925), .Z(n10163) );
  XOR U14807 ( .A(n13926), .B(n13927), .Z(n13555) );
  XNOR U14808 ( .A(n13928), .B(n10694), .Z(n13927) );
  XNOR U14809 ( .A(n13929), .B(n13930), .Z(n10694) );
  ANDN U14810 ( .B(n13931), .A(n13932), .Z(n13929) );
  XNOR U14811 ( .A(n9857), .B(n13933), .Z(n13926) );
  XOR U14812 ( .A(n12272), .B(n13934), .Z(n13933) );
  XOR U14813 ( .A(n13935), .B(n13936), .Z(n12272) );
  ANDN U14814 ( .B(n13937), .A(n13938), .Z(n13935) );
  XOR U14815 ( .A(n13939), .B(n13940), .Z(n9857) );
  ANDN U14816 ( .B(n13941), .A(n13942), .Z(n13939) );
  XNOR U14817 ( .A(n13943), .B(n12117), .Z(n13917) );
  XOR U14818 ( .A(n8871), .B(n5187), .Z(n5701) );
  XNOR U14819 ( .A(n13944), .B(n13945), .Z(n6503) );
  XOR U14820 ( .A(n5509), .B(n2528), .Z(n13945) );
  XNOR U14821 ( .A(n13946), .B(n6552), .Z(n2528) );
  XNOR U14822 ( .A(n11972), .B(n13947), .Z(n6552) );
  ANDN U14823 ( .B(n8877), .A(n13479), .Z(n13946) );
  XOR U14824 ( .A(n10754), .B(n13948), .Z(n13479) );
  XOR U14825 ( .A(n13730), .B(n13949), .Z(n10754) );
  XOR U14826 ( .A(n13950), .B(n13951), .Z(n13730) );
  XNOR U14827 ( .A(n12177), .B(n12284), .Z(n13951) );
  NOR U14828 ( .A(n13953), .B(n13141), .Z(n13952) );
  XOR U14829 ( .A(n13954), .B(n13955), .Z(n12177) );
  NOR U14830 ( .A(n13956), .B(n13957), .Z(n13954) );
  XOR U14831 ( .A(n10625), .B(n13958), .Z(n13950) );
  XNOR U14832 ( .A(n10502), .B(n12305), .Z(n13958) );
  XNOR U14833 ( .A(n13959), .B(n13150), .Z(n12305) );
  ANDN U14834 ( .B(n13151), .A(n13960), .Z(n13959) );
  XNOR U14835 ( .A(n13961), .B(n13147), .Z(n10502) );
  ANDN U14836 ( .B(n13962), .A(n13146), .Z(n13961) );
  XOR U14837 ( .A(n13963), .B(n13154), .Z(n10625) );
  ANDN U14838 ( .B(n13155), .A(n13964), .Z(n13963) );
  XOR U14839 ( .A(n13965), .B(n11045), .Z(n8877) );
  XNOR U14840 ( .A(n13966), .B(n6545), .Z(n5509) );
  XOR U14841 ( .A(n10167), .B(n13098), .Z(n6545) );
  XOR U14842 ( .A(n13967), .B(n13968), .Z(n13098) );
  ANDN U14843 ( .B(n13969), .A(n13970), .Z(n13967) );
  IV U14844 ( .A(n11303), .Z(n10167) );
  XNOR U14845 ( .A(n13971), .B(n13972), .Z(n11303) );
  ANDN U14846 ( .B(n8922), .A(n13468), .Z(n13966) );
  XOR U14847 ( .A(n3512), .B(n13973), .Z(n13944) );
  XNOR U14848 ( .A(n8915), .B(n4890), .Z(n13973) );
  XNOR U14849 ( .A(n13974), .B(n6540), .Z(n4890) );
  XOR U14850 ( .A(n9238), .B(n13975), .Z(n6540) );
  ANDN U14851 ( .B(n8873), .A(n8874), .Z(n13974) );
  XNOR U14852 ( .A(n13976), .B(n10316), .Z(n8874) );
  XNOR U14853 ( .A(n11837), .B(n13280), .Z(n10316) );
  XNOR U14854 ( .A(n13977), .B(n13978), .Z(n13280) );
  XNOR U14855 ( .A(n10933), .B(n9881), .Z(n13978) );
  XOR U14856 ( .A(n13979), .B(n13980), .Z(n9881) );
  NOR U14857 ( .A(n13981), .B(n13982), .Z(n13979) );
  XOR U14858 ( .A(n13983), .B(n13984), .Z(n10933) );
  ANDN U14859 ( .B(n13985), .A(n13986), .Z(n13983) );
  XOR U14860 ( .A(n13285), .B(n13987), .Z(n13977) );
  XOR U14861 ( .A(n9115), .B(n12714), .Z(n13987) );
  XNOR U14862 ( .A(n13988), .B(n13989), .Z(n12714) );
  ANDN U14863 ( .B(n13990), .A(n13991), .Z(n13988) );
  XNOR U14864 ( .A(n13992), .B(n13993), .Z(n9115) );
  NOR U14865 ( .A(n13994), .B(n13995), .Z(n13992) );
  XOR U14866 ( .A(n13996), .B(n13997), .Z(n13285) );
  ANDN U14867 ( .B(n13998), .A(n13999), .Z(n13996) );
  XOR U14868 ( .A(n14000), .B(n14001), .Z(n11837) );
  XOR U14869 ( .A(n10635), .B(n10486), .Z(n14001) );
  XOR U14870 ( .A(n14002), .B(n14003), .Z(n10486) );
  NOR U14871 ( .A(n14004), .B(n14005), .Z(n14002) );
  XNOR U14872 ( .A(n14006), .B(n14007), .Z(n10635) );
  ANDN U14873 ( .B(n14008), .A(n14009), .Z(n14006) );
  XNOR U14874 ( .A(n9772), .B(n14010), .Z(n14000) );
  XNOR U14875 ( .A(n14011), .B(n10391), .Z(n14010) );
  XOR U14876 ( .A(n14012), .B(n14013), .Z(n10391) );
  ANDN U14877 ( .B(n14014), .A(n14015), .Z(n14012) );
  XNOR U14878 ( .A(n14016), .B(n14017), .Z(n9772) );
  ANDN U14879 ( .B(n14018), .A(n14019), .Z(n14016) );
  XOR U14880 ( .A(n11301), .B(n14020), .Z(n8873) );
  XNOR U14881 ( .A(n14021), .B(n6536), .Z(n8915) );
  XOR U14882 ( .A(n14022), .B(n11479), .Z(n6536) );
  XOR U14883 ( .A(n12633), .B(n14023), .Z(n11479) );
  XOR U14884 ( .A(n14024), .B(n14025), .Z(n12633) );
  XOR U14885 ( .A(n11076), .B(n10709), .Z(n14025) );
  XNOR U14886 ( .A(n14026), .B(n14027), .Z(n10709) );
  NOR U14887 ( .A(n14028), .B(n14029), .Z(n14026) );
  XNOR U14888 ( .A(n14030), .B(n13434), .Z(n11076) );
  ANDN U14889 ( .B(n13435), .A(n14031), .Z(n14030) );
  XNOR U14890 ( .A(n13421), .B(n14032), .Z(n14024) );
  XNOR U14891 ( .A(n9241), .B(n10152), .Z(n14032) );
  XNOR U14892 ( .A(n14033), .B(n14034), .Z(n10152) );
  XNOR U14893 ( .A(n14037), .B(n13439), .Z(n9241) );
  NOR U14894 ( .A(n14038), .B(n14039), .Z(n14037) );
  XNOR U14895 ( .A(n14040), .B(n13428), .Z(n13421) );
  ANDN U14896 ( .B(n14041), .A(n14042), .Z(n14040) );
  ANDN U14897 ( .B(n8868), .A(n8869), .Z(n14021) );
  XOR U14898 ( .A(n14043), .B(n11114), .Z(n8869) );
  XOR U14899 ( .A(n14044), .B(n9329), .Z(n8868) );
  XNOR U14900 ( .A(n13384), .B(n11707), .Z(n9329) );
  XNOR U14901 ( .A(n14045), .B(n14046), .Z(n11707) );
  XOR U14902 ( .A(n13635), .B(n10101), .Z(n14046) );
  XNOR U14903 ( .A(n14047), .B(n14048), .Z(n10101) );
  ANDN U14904 ( .B(n14049), .A(n14050), .Z(n14047) );
  XNOR U14905 ( .A(n14051), .B(n14052), .Z(n13635) );
  ANDN U14906 ( .B(n14053), .A(n14054), .Z(n14051) );
  XOR U14907 ( .A(n14055), .B(n14056), .Z(n14045) );
  XNOR U14908 ( .A(n11112), .B(n11965), .Z(n14056) );
  XOR U14909 ( .A(n14057), .B(n14058), .Z(n11965) );
  ANDN U14910 ( .B(n14059), .A(n14060), .Z(n14057) );
  XNOR U14911 ( .A(n14061), .B(n14062), .Z(n11112) );
  ANDN U14912 ( .B(n14063), .A(n14064), .Z(n14061) );
  XOR U14913 ( .A(n14065), .B(n14066), .Z(n13384) );
  XOR U14914 ( .A(n13094), .B(n10726), .Z(n14066) );
  XNOR U14915 ( .A(n14067), .B(n14068), .Z(n10726) );
  ANDN U14916 ( .B(n14069), .A(n14070), .Z(n14067) );
  XNOR U14917 ( .A(n14071), .B(n14072), .Z(n13094) );
  ANDN U14918 ( .B(n14073), .A(n14074), .Z(n14071) );
  XOR U14919 ( .A(n12702), .B(n14075), .Z(n14065) );
  XNOR U14920 ( .A(n12676), .B(n11799), .Z(n14075) );
  XNOR U14921 ( .A(n14076), .B(n14077), .Z(n11799) );
  ANDN U14922 ( .B(n14078), .A(n14079), .Z(n14076) );
  XNOR U14923 ( .A(n14080), .B(n14081), .Z(n12676) );
  AND U14924 ( .A(n14082), .B(n14083), .Z(n14080) );
  XNOR U14925 ( .A(n14084), .B(n14085), .Z(n12702) );
  ANDN U14926 ( .B(n14086), .A(n14087), .Z(n14084) );
  XNOR U14927 ( .A(n14088), .B(n6549), .Z(n3512) );
  XOR U14928 ( .A(n9652), .B(n14089), .Z(n6549) );
  XNOR U14929 ( .A(n14090), .B(n12959), .Z(n9652) );
  XOR U14930 ( .A(n14091), .B(n14092), .Z(n12959) );
  XNOR U14931 ( .A(n13090), .B(n14093), .Z(n14092) );
  XNOR U14932 ( .A(n14094), .B(n14095), .Z(n13090) );
  AND U14933 ( .A(n14096), .B(n14097), .Z(n14094) );
  XOR U14934 ( .A(n9335), .B(n14098), .Z(n14091) );
  XNOR U14935 ( .A(n12607), .B(n10119), .Z(n14098) );
  XNOR U14936 ( .A(n14099), .B(n14100), .Z(n10119) );
  ANDN U14937 ( .B(n14101), .A(n14102), .Z(n14099) );
  AND U14938 ( .A(n14105), .B(n14106), .Z(n14103) );
  XNOR U14939 ( .A(n14107), .B(n14108), .Z(n9335) );
  ANDN U14940 ( .B(n14109), .A(n14110), .Z(n14107) );
  ANDN U14941 ( .B(n8865), .A(n8866), .Z(n14088) );
  XOR U14942 ( .A(n14111), .B(n12122), .Z(n8866) );
  XOR U14943 ( .A(n9778), .B(n14112), .Z(n8865) );
  IV U14944 ( .A(n10050), .Z(n9778) );
  XOR U14945 ( .A(n14113), .B(n12597), .Z(n10050) );
  XOR U14946 ( .A(n14114), .B(n14115), .Z(n12597) );
  XOR U14947 ( .A(n14116), .B(n10107), .Z(n14115) );
  XNOR U14948 ( .A(n14117), .B(n14118), .Z(n10107) );
  AND U14949 ( .A(n14119), .B(n14120), .Z(n14117) );
  XNOR U14950 ( .A(n14121), .B(n14122), .Z(n14114) );
  XOR U14951 ( .A(n14123), .B(n14124), .Z(n14122) );
  XOR U14952 ( .A(n14125), .B(n14126), .Z(n6347) );
  XNOR U14953 ( .A(n5474), .B(n3722), .Z(n14126) );
  XOR U14954 ( .A(n14127), .B(n14128), .Z(n3722) );
  ANDN U14955 ( .B(n6569), .A(n6570), .Z(n14127) );
  XNOR U14956 ( .A(n14129), .B(n11877), .Z(n6570) );
  XNOR U14957 ( .A(n14130), .B(n8934), .Z(n5474) );
  ANDN U14958 ( .B(n6562), .A(n6560), .Z(n14130) );
  XOR U14959 ( .A(n14131), .B(n11704), .Z(n6560) );
  XOR U14960 ( .A(n14132), .B(n12122), .Z(n6562) );
  IV U14961 ( .A(n12843), .Z(n12122) );
  XOR U14962 ( .A(n4337), .B(n14133), .Z(n14125) );
  XNOR U14963 ( .A(n5925), .B(n2129), .Z(n14133) );
  XNOR U14964 ( .A(n14134), .B(n8930), .Z(n2129) );
  ANDN U14965 ( .B(n6575), .A(n8931), .Z(n14134) );
  XOR U14966 ( .A(n14135), .B(n9613), .Z(n8931) );
  XNOR U14967 ( .A(n14136), .B(n12137), .Z(n9613) );
  XNOR U14968 ( .A(n14137), .B(n14138), .Z(n12137) );
  XNOR U14969 ( .A(n13761), .B(n12257), .Z(n14138) );
  XOR U14970 ( .A(n14139), .B(n14140), .Z(n12257) );
  ANDN U14971 ( .B(n13253), .A(n13254), .Z(n14139) );
  XNOR U14972 ( .A(n14141), .B(n14142), .Z(n13761) );
  ANDN U14973 ( .B(n13251), .A(n13249), .Z(n14141) );
  XOR U14974 ( .A(n11923), .B(n14143), .Z(n14137) );
  XOR U14975 ( .A(n9892), .B(n12504), .Z(n14143) );
  XNOR U14976 ( .A(n14144), .B(n14145), .Z(n12504) );
  XNOR U14977 ( .A(n14146), .B(n14147), .Z(n9892) );
  ANDN U14978 ( .B(n13264), .A(n13262), .Z(n14146) );
  XNOR U14979 ( .A(n14148), .B(n14149), .Z(n11923) );
  XNOR U14980 ( .A(n10280), .B(n14150), .Z(n6575) );
  IV U14981 ( .A(n14151), .Z(n10280) );
  XNOR U14982 ( .A(n14152), .B(n8943), .Z(n5925) );
  NOR U14983 ( .A(n6578), .B(n6577), .Z(n14152) );
  XOR U14984 ( .A(n9623), .B(n14153), .Z(n6577) );
  XOR U14985 ( .A(n14155), .B(n14156), .Z(n11976) );
  XOR U14986 ( .A(n12016), .B(n12877), .Z(n14156) );
  XOR U14987 ( .A(n14157), .B(n13264), .Z(n12877) );
  XOR U14988 ( .A(n14158), .B(n14159), .Z(n13264) );
  NOR U14989 ( .A(n14160), .B(n13263), .Z(n14157) );
  XOR U14990 ( .A(n14161), .B(n13268), .Z(n12016) );
  XOR U14991 ( .A(n14162), .B(n14163), .Z(n13268) );
  NOR U14992 ( .A(n14164), .B(n13267), .Z(n14161) );
  XOR U14993 ( .A(n11346), .B(n14165), .Z(n14155) );
  XNOR U14994 ( .A(n10192), .B(n12665), .Z(n14165) );
  XNOR U14995 ( .A(n14166), .B(n13254), .Z(n12665) );
  XOR U14996 ( .A(n14167), .B(n14168), .Z(n13254) );
  XOR U14997 ( .A(n14170), .B(n13260), .Z(n10192) );
  XOR U14998 ( .A(n14171), .B(n14172), .Z(n13260) );
  NOR U14999 ( .A(n14173), .B(n13259), .Z(n14170) );
  XOR U15000 ( .A(n14175), .B(n14176), .Z(n13251) );
  NOR U15001 ( .A(n14177), .B(n13250), .Z(n14174) );
  XNOR U15002 ( .A(n14178), .B(n14179), .Z(n6578) );
  XNOR U15003 ( .A(n14180), .B(n8939), .Z(n4337) );
  ANDN U15004 ( .B(n6565), .A(n8940), .Z(n14180) );
  XNOR U15005 ( .A(n14181), .B(n11114), .Z(n8940) );
  XNOR U15006 ( .A(n14182), .B(n14183), .Z(n11114) );
  XNOR U15007 ( .A(n14184), .B(n9808), .Z(n6565) );
  XOR U15008 ( .A(n14185), .B(n14186), .Z(n9808) );
  XOR U15009 ( .A(n14187), .B(n8922), .Z(n8871) );
  XNOR U15010 ( .A(n12247), .B(n14188), .Z(n8922) );
  ANDN U15011 ( .B(n13468), .A(n6543), .Z(n14187) );
  XNOR U15012 ( .A(n14189), .B(n11369), .Z(n6543) );
  XNOR U15013 ( .A(n14190), .B(n14191), .Z(n11369) );
  XNOR U15014 ( .A(n13855), .B(n9431), .Z(n13468) );
  IV U15015 ( .A(n14192), .Z(n9431) );
  XOR U15016 ( .A(n14193), .B(n14194), .Z(n13855) );
  NOR U15017 ( .A(n14195), .B(n14196), .Z(n14193) );
  XOR U15018 ( .A(n14197), .B(n6235), .Z(out[1001]) );
  XOR U15019 ( .A(n9158), .B(n2306), .Z(n6235) );
  XNOR U15020 ( .A(n10042), .B(n6194), .Z(n2306) );
  XNOR U15021 ( .A(n14198), .B(n14199), .Z(n6194) );
  XNOR U15022 ( .A(n2344), .B(n5489), .Z(n14199) );
  XOR U15023 ( .A(n14200), .B(n8003), .Z(n5489) );
  XNOR U15024 ( .A(n14201), .B(n10357), .Z(n8003) );
  XOR U15025 ( .A(n12969), .B(n13919), .Z(n10357) );
  XOR U15026 ( .A(n14202), .B(n14203), .Z(n13919) );
  XNOR U15027 ( .A(n12998), .B(n13556), .Z(n14203) );
  ANDN U15028 ( .B(n14205), .A(n13585), .Z(n14204) );
  XOR U15029 ( .A(n14206), .B(n14207), .Z(n12998) );
  ANDN U15030 ( .B(n14208), .A(n14209), .Z(n14206) );
  XNOR U15031 ( .A(n13007), .B(n14210), .Z(n14202) );
  XNOR U15032 ( .A(n12406), .B(n11633), .Z(n14210) );
  XOR U15033 ( .A(n14211), .B(n13842), .Z(n11633) );
  AND U15034 ( .A(n13526), .B(n13843), .Z(n14211) );
  XOR U15035 ( .A(n14212), .B(n13578), .Z(n12406) );
  ANDN U15036 ( .B(n13579), .A(n14213), .Z(n14212) );
  XNOR U15037 ( .A(n14214), .B(n13588), .Z(n13007) );
  ANDN U15038 ( .B(n13522), .A(n13587), .Z(n14214) );
  XOR U15039 ( .A(n14215), .B(n14216), .Z(n12969) );
  XNOR U15040 ( .A(n13326), .B(n11786), .Z(n14216) );
  XOR U15041 ( .A(n14217), .B(n14218), .Z(n11786) );
  NOR U15042 ( .A(n14219), .B(n14220), .Z(n14217) );
  XOR U15043 ( .A(n14221), .B(n13561), .Z(n13326) );
  NOR U15044 ( .A(n13562), .B(n14222), .Z(n14221) );
  XOR U15045 ( .A(n12317), .B(n14223), .Z(n14215) );
  XOR U15046 ( .A(n10288), .B(n10233), .Z(n14223) );
  XOR U15047 ( .A(n14224), .B(n13565), .Z(n10233) );
  ANDN U15048 ( .B(n13566), .A(n14225), .Z(n14224) );
  XNOR U15049 ( .A(n14226), .B(n14227), .Z(n10288) );
  ANDN U15050 ( .B(n14228), .A(n13572), .Z(n14226) );
  XOR U15051 ( .A(n14229), .B(n14230), .Z(n12317) );
  ANDN U15052 ( .B(n14231), .A(n14232), .Z(n14229) );
  ANDN U15053 ( .B(n9168), .A(n8004), .Z(n14200) );
  XOR U15054 ( .A(n14151), .B(n14233), .Z(n8004) );
  XNOR U15055 ( .A(n11175), .B(n14234), .Z(n14151) );
  XOR U15056 ( .A(n14235), .B(n14236), .Z(n11175) );
  XOR U15057 ( .A(n9787), .B(n10616), .Z(n14236) );
  XNOR U15058 ( .A(n14237), .B(n13750), .Z(n10616) );
  IV U15059 ( .A(n14238), .Z(n13750) );
  NOR U15060 ( .A(n14239), .B(n13749), .Z(n14237) );
  XOR U15061 ( .A(n14240), .B(n14241), .Z(n9787) );
  ANDN U15062 ( .B(n14242), .A(n13744), .Z(n14240) );
  IV U15063 ( .A(n14243), .Z(n13744) );
  XOR U15064 ( .A(n12991), .B(n14244), .Z(n14235) );
  XOR U15065 ( .A(n12407), .B(n11208), .Z(n14244) );
  XNOR U15066 ( .A(n14245), .B(n13758), .Z(n11208) );
  IV U15067 ( .A(n14246), .Z(n13758) );
  NOR U15068 ( .A(n13757), .B(n14247), .Z(n14245) );
  NOR U15069 ( .A(n14249), .B(n14250), .Z(n14248) );
  XNOR U15070 ( .A(n14251), .B(n14252), .Z(n12991) );
  NOR U15071 ( .A(n14253), .B(n14254), .Z(n14251) );
  XNOR U15072 ( .A(n14124), .B(n10108), .Z(n9168) );
  XNOR U15073 ( .A(n14255), .B(n14256), .Z(n14124) );
  ANDN U15074 ( .B(n14257), .A(n14258), .Z(n14255) );
  XOR U15075 ( .A(n14259), .B(n9050), .Z(n2344) );
  XNOR U15076 ( .A(n14260), .B(n9244), .Z(n9050) );
  ANDN U15077 ( .B(n9163), .A(n8008), .Z(n14259) );
  XOR U15078 ( .A(n13000), .B(n14261), .Z(n8008) );
  XNOR U15079 ( .A(n14262), .B(n14263), .Z(n13000) );
  XOR U15080 ( .A(n14264), .B(n11960), .Z(n9163) );
  XNOR U15081 ( .A(n13867), .B(n12774), .Z(n11960) );
  XNOR U15082 ( .A(n14265), .B(n14266), .Z(n12774) );
  XNOR U15083 ( .A(n14267), .B(n14268), .Z(n14266) );
  XOR U15084 ( .A(n14269), .B(n14270), .Z(n14265) );
  XNOR U15085 ( .A(n11840), .B(n11699), .Z(n14270) );
  XNOR U15086 ( .A(n14271), .B(n14220), .Z(n11699) );
  ANDN U15087 ( .B(n14272), .A(n14273), .Z(n14271) );
  XNOR U15088 ( .A(n14274), .B(n14225), .Z(n11840) );
  NOR U15089 ( .A(n13564), .B(n14275), .Z(n14274) );
  XOR U15090 ( .A(n14276), .B(n14277), .Z(n13867) );
  XOR U15091 ( .A(n10943), .B(n12246), .Z(n14277) );
  XOR U15092 ( .A(n14278), .B(n14279), .Z(n12246) );
  AND U15093 ( .A(n14280), .B(n14281), .Z(n14278) );
  XNOR U15094 ( .A(n14282), .B(n14283), .Z(n10943) );
  XOR U15095 ( .A(n10171), .B(n14286), .Z(n14276) );
  XOR U15096 ( .A(n11721), .B(n14287), .Z(n14286) );
  XNOR U15097 ( .A(n14288), .B(n14289), .Z(n11721) );
  NOR U15098 ( .A(n14290), .B(n14291), .Z(n14288) );
  XNOR U15099 ( .A(n14292), .B(n14293), .Z(n10171) );
  ANDN U15100 ( .B(n14294), .A(n14295), .Z(n14292) );
  XNOR U15101 ( .A(n3176), .B(n14296), .Z(n14198) );
  XOR U15102 ( .A(n6322), .B(n7997), .Z(n14296) );
  XNOR U15103 ( .A(n14297), .B(n8013), .Z(n7997) );
  XOR U15104 ( .A(n9153), .B(n13312), .Z(n8013) );
  XNOR U15105 ( .A(n14298), .B(n13889), .Z(n13312) );
  NOR U15106 ( .A(n14299), .B(n14300), .Z(n14298) );
  NOR U15107 ( .A(n9165), .B(n8012), .Z(n14297) );
  XOR U15108 ( .A(n14301), .B(n10964), .Z(n8012) );
  XOR U15109 ( .A(n14302), .B(n12755), .Z(n10964) );
  XOR U15110 ( .A(n14303), .B(n14304), .Z(n12755) );
  XOR U15111 ( .A(n14305), .B(n11730), .Z(n14304) );
  XNOR U15112 ( .A(n14306), .B(n14307), .Z(n11730) );
  AND U15113 ( .A(n14308), .B(n14309), .Z(n14306) );
  XOR U15114 ( .A(n10481), .B(n14310), .Z(n14303) );
  XOR U15115 ( .A(n12630), .B(n11574), .Z(n14310) );
  XNOR U15116 ( .A(n14311), .B(n14312), .Z(n11574) );
  ANDN U15117 ( .B(n14313), .A(n14314), .Z(n14311) );
  XNOR U15118 ( .A(n14315), .B(n14316), .Z(n12630) );
  AND U15119 ( .A(n14317), .B(n14318), .Z(n14315) );
  XNOR U15120 ( .A(n14319), .B(n14320), .Z(n10481) );
  ANDN U15121 ( .B(n14321), .A(n14322), .Z(n14319) );
  XOR U15122 ( .A(n14323), .B(n9420), .Z(n9165) );
  XNOR U15123 ( .A(n14324), .B(n14325), .Z(n9420) );
  XNOR U15124 ( .A(n14326), .B(n8016), .Z(n6322) );
  XOR U15125 ( .A(n9238), .B(n14327), .Z(n8016) );
  XNOR U15126 ( .A(n14328), .B(n14329), .Z(n11865) );
  XNOR U15127 ( .A(n11284), .B(n12123), .Z(n14329) );
  XOR U15128 ( .A(n14330), .B(n12551), .Z(n12123) );
  NOR U15129 ( .A(n13609), .B(n14331), .Z(n14330) );
  IV U15130 ( .A(n14332), .Z(n13609) );
  XOR U15131 ( .A(n14333), .B(n14334), .Z(n11284) );
  NOR U15132 ( .A(n13602), .B(n14335), .Z(n14333) );
  XNOR U15133 ( .A(n11769), .B(n14336), .Z(n14328) );
  XOR U15134 ( .A(n9871), .B(n11969), .Z(n14336) );
  XNOR U15135 ( .A(n14337), .B(n14338), .Z(n11969) );
  XNOR U15136 ( .A(n14340), .B(n12546), .Z(n9871) );
  NOR U15137 ( .A(n14341), .B(n14342), .Z(n14340) );
  XOR U15138 ( .A(n14343), .B(n14344), .Z(n11769) );
  ANDN U15139 ( .B(n14345), .A(n14346), .Z(n14343) );
  XOR U15140 ( .A(n14347), .B(n14348), .Z(n12741) );
  XOR U15141 ( .A(n12179), .B(n10748), .Z(n14348) );
  XNOR U15142 ( .A(n14349), .B(n14350), .Z(n10748) );
  ANDN U15143 ( .B(n12482), .A(n14351), .Z(n14349) );
  XOR U15144 ( .A(n14352), .B(n14353), .Z(n12179) );
  NOR U15145 ( .A(n14354), .B(n14355), .Z(n14352) );
  XOR U15146 ( .A(n13014), .B(n14356), .Z(n14347) );
  XNOR U15147 ( .A(n14357), .B(n14358), .Z(n14356) );
  XNOR U15148 ( .A(n14359), .B(n14360), .Z(n13014) );
  ANDN U15149 ( .B(n12476), .A(n14361), .Z(n14359) );
  AND U15150 ( .A(n8017), .B(n13694), .Z(n14326) );
  XNOR U15151 ( .A(n14362), .B(n8020), .Z(n3176) );
  XNOR U15152 ( .A(n10965), .B(n14363), .Z(n8020) );
  XOR U15153 ( .A(n14364), .B(n14365), .Z(n10965) );
  ANDN U15154 ( .B(n8021), .A(n9160), .Z(n14362) );
  XOR U15155 ( .A(n12128), .B(n14366), .Z(n9160) );
  XNOR U15156 ( .A(n13594), .B(n14367), .Z(n12128) );
  XOR U15157 ( .A(n14368), .B(n14369), .Z(n13594) );
  XNOR U15158 ( .A(n11475), .B(n11050), .Z(n14369) );
  XOR U15159 ( .A(n14370), .B(n14371), .Z(n11050) );
  ANDN U15160 ( .B(n14372), .A(n13109), .Z(n14370) );
  XOR U15161 ( .A(n14373), .B(n14374), .Z(n11475) );
  XOR U15162 ( .A(n14376), .B(n14377), .Z(n14368) );
  XNOR U15163 ( .A(n9531), .B(n11845), .Z(n14377) );
  XOR U15164 ( .A(n14378), .B(n14379), .Z(n11845) );
  ANDN U15165 ( .B(n14380), .A(n13968), .Z(n14378) );
  XOR U15166 ( .A(n14381), .B(n14382), .Z(n9531) );
  ANDN U15167 ( .B(n14383), .A(n13113), .Z(n14381) );
  XOR U15168 ( .A(n12862), .B(n9224), .Z(n8021) );
  XNOR U15169 ( .A(n14384), .B(n14385), .Z(n12862) );
  ANDN U15170 ( .B(n14386), .A(n14387), .Z(n14384) );
  XOR U15171 ( .A(n14388), .B(n14389), .Z(n10042) );
  XOR U15172 ( .A(n5294), .B(n1952), .Z(n14389) );
  XNOR U15173 ( .A(n14390), .B(n9194), .Z(n1952) );
  NOR U15174 ( .A(n8070), .B(n9181), .Z(n14390) );
  XOR U15175 ( .A(n13062), .B(n10630), .Z(n9181) );
  IV U15176 ( .A(n12013), .Z(n10630) );
  XNOR U15177 ( .A(n14391), .B(n13547), .Z(n13062) );
  ANDN U15178 ( .B(n14392), .A(n13922), .Z(n14391) );
  XOR U15179 ( .A(n14393), .B(n11937), .Z(n8070) );
  XOR U15180 ( .A(n14394), .B(n9200), .Z(n5294) );
  NOR U15181 ( .A(n9179), .B(n8062), .Z(n14394) );
  XNOR U15182 ( .A(n14395), .B(n10971), .Z(n8062) );
  XNOR U15183 ( .A(n12720), .B(n13949), .Z(n10971) );
  XNOR U15184 ( .A(n14396), .B(n14397), .Z(n13949) );
  XNOR U15185 ( .A(n13652), .B(n14398), .Z(n14397) );
  XNOR U15186 ( .A(n14399), .B(n14400), .Z(n13652) );
  ANDN U15187 ( .B(n14401), .A(n14402), .Z(n14399) );
  XOR U15188 ( .A(n10169), .B(n14403), .Z(n14396) );
  XNOR U15189 ( .A(n9526), .B(n11793), .Z(n14403) );
  XNOR U15190 ( .A(n14404), .B(n14405), .Z(n11793) );
  ANDN U15191 ( .B(n14406), .A(n14407), .Z(n14404) );
  XOR U15192 ( .A(n14408), .B(n14409), .Z(n9526) );
  ANDN U15193 ( .B(n14410), .A(n14411), .Z(n14408) );
  XNOR U15194 ( .A(n14412), .B(n14413), .Z(n10169) );
  NOR U15195 ( .A(n14414), .B(n14415), .Z(n14412) );
  XOR U15196 ( .A(n14416), .B(n14417), .Z(n12720) );
  XOR U15197 ( .A(n11245), .B(n11887), .Z(n14417) );
  XNOR U15198 ( .A(n14418), .B(n14419), .Z(n11887) );
  ANDN U15199 ( .B(n14420), .A(n14421), .Z(n14418) );
  XNOR U15200 ( .A(n14422), .B(n14423), .Z(n11245) );
  XOR U15201 ( .A(n13510), .B(n14426), .Z(n14416) );
  XOR U15202 ( .A(n12610), .B(n12097), .Z(n14426) );
  XOR U15203 ( .A(n14427), .B(n14428), .Z(n12097) );
  ANDN U15204 ( .B(n14429), .A(n14430), .Z(n14427) );
  XNOR U15205 ( .A(n14431), .B(n14432), .Z(n12610) );
  XOR U15206 ( .A(n14435), .B(n14436), .Z(n13510) );
  XNOR U15207 ( .A(n4549), .B(n14437), .Z(n14436) );
  NANDN U15208 ( .A(n14438), .B(n14439), .Z(n14437) );
  XOR U15209 ( .A(n14440), .B(n10062), .Z(n9179) );
  XOR U15210 ( .A(n3746), .B(n14441), .Z(n14388) );
  XOR U15211 ( .A(n9189), .B(n4209), .Z(n14441) );
  XNOR U15212 ( .A(n14442), .B(n9203), .Z(n4209) );
  ANDN U15213 ( .B(n8053), .A(n9202), .Z(n14442) );
  XOR U15214 ( .A(n12444), .B(n14443), .Z(n9202) );
  XNOR U15215 ( .A(n14444), .B(n14445), .Z(n12444) );
  ANDN U15216 ( .B(n14446), .A(n14447), .Z(n14444) );
  XNOR U15217 ( .A(n9439), .B(n14448), .Z(n8053) );
  IV U15218 ( .A(n9632), .Z(n9439) );
  XOR U15219 ( .A(n14449), .B(n14191), .Z(n9632) );
  XNOR U15220 ( .A(n14450), .B(n14451), .Z(n14191) );
  XOR U15221 ( .A(n12198), .B(n10295), .Z(n14451) );
  XNOR U15222 ( .A(n14452), .B(n14453), .Z(n10295) );
  NOR U15223 ( .A(n14454), .B(n14455), .Z(n14452) );
  XNOR U15224 ( .A(n14456), .B(n14457), .Z(n12198) );
  XOR U15225 ( .A(n11854), .B(n14460), .Z(n14450) );
  XOR U15226 ( .A(n13892), .B(n11645), .Z(n14460) );
  XNOR U15227 ( .A(n14461), .B(n14462), .Z(n11645) );
  ANDN U15228 ( .B(n14463), .A(n14464), .Z(n14461) );
  XNOR U15229 ( .A(n14465), .B(n14466), .Z(n13892) );
  ANDN U15230 ( .B(n14467), .A(n14468), .Z(n14465) );
  XNOR U15231 ( .A(n14469), .B(n14470), .Z(n11854) );
  ANDN U15232 ( .B(n14471), .A(n14472), .Z(n14469) );
  NOR U15233 ( .A(n9173), .B(n8057), .Z(n14473) );
  XOR U15234 ( .A(n14474), .B(n13013), .Z(n8057) );
  XNOR U15235 ( .A(n13808), .B(n9910), .Z(n9173) );
  XOR U15236 ( .A(n14475), .B(n14476), .Z(n9910) );
  XOR U15237 ( .A(n14477), .B(n14478), .Z(n13808) );
  XNOR U15238 ( .A(n14479), .B(n14480), .Z(n3746) );
  NOR U15239 ( .A(n8066), .B(n9177), .Z(n14479) );
  XOR U15240 ( .A(n14481), .B(n12734), .Z(n8066) );
  XNOR U15241 ( .A(n14482), .B(n8017), .Z(n9158) );
  XOR U15242 ( .A(n11433), .B(n13336), .Z(n8017) );
  XNOR U15243 ( .A(n14483), .B(n14484), .Z(n13336) );
  ANDN U15244 ( .B(n14485), .A(n14486), .Z(n14483) );
  NOR U15245 ( .A(n13695), .B(n13694), .Z(n14482) );
  XOR U15246 ( .A(n9617), .B(n14487), .Z(n13694) );
  XNOR U15247 ( .A(n12588), .B(n14489), .Z(n11937) );
  XOR U15248 ( .A(n14490), .B(n14491), .Z(n12588) );
  XOR U15249 ( .A(n14492), .B(n13476), .Z(n14491) );
  XNOR U15250 ( .A(n14493), .B(n14494), .Z(n13476) );
  XOR U15251 ( .A(n13551), .B(n14496), .Z(n14490) );
  XOR U15252 ( .A(n10636), .B(n12285), .Z(n14496) );
  XNOR U15253 ( .A(n14497), .B(n14498), .Z(n12285) );
  NOR U15254 ( .A(n13717), .B(n14499), .Z(n14497) );
  XNOR U15255 ( .A(n14500), .B(n14501), .Z(n10636) );
  NOR U15256 ( .A(n13708), .B(n14502), .Z(n14500) );
  XNOR U15257 ( .A(n14503), .B(n14504), .Z(n13551) );
  ANDN U15258 ( .B(n5705), .A(n5707), .Z(n14197) );
  XOR U15259 ( .A(n11670), .B(n2098), .Z(n5707) );
  XNOR U15260 ( .A(n8344), .B(n9820), .Z(n2098) );
  XNOR U15261 ( .A(n14506), .B(n14507), .Z(n9820) );
  XOR U15262 ( .A(n5505), .B(n3644), .Z(n14507) );
  XOR U15263 ( .A(n14508), .B(n14509), .Z(n3644) );
  ANDN U15264 ( .B(n8504), .A(n8502), .Z(n14508) );
  IV U15265 ( .A(n14510), .Z(n8502) );
  XNOR U15266 ( .A(n11054), .B(n13138), .Z(n8504) );
  XNOR U15267 ( .A(n14511), .B(n14512), .Z(n13138) );
  NOR U15268 ( .A(n14513), .B(n13955), .Z(n14511) );
  XOR U15269 ( .A(n14514), .B(n14515), .Z(n11054) );
  XOR U15270 ( .A(n14516), .B(n11993), .Z(n5505) );
  NOR U15271 ( .A(n8498), .B(n8499), .Z(n14516) );
  XNOR U15272 ( .A(n10602), .B(n14517), .Z(n8499) );
  XOR U15273 ( .A(n14518), .B(n13419), .Z(n10602) );
  XNOR U15274 ( .A(n14519), .B(n14520), .Z(n13419) );
  XNOR U15275 ( .A(n10096), .B(n9810), .Z(n14520) );
  XNOR U15276 ( .A(n14521), .B(n14522), .Z(n9810) );
  AND U15277 ( .A(n14523), .B(n14524), .Z(n14521) );
  XNOR U15278 ( .A(n14525), .B(n14526), .Z(n10096) );
  ANDN U15279 ( .B(n14527), .A(n14528), .Z(n14525) );
  XOR U15280 ( .A(n11424), .B(n14529), .Z(n14519) );
  XNOR U15281 ( .A(n11432), .B(n14530), .Z(n14529) );
  XOR U15282 ( .A(n14531), .B(n14532), .Z(n11432) );
  ANDN U15283 ( .B(n14533), .A(n14534), .Z(n14531) );
  XNOR U15284 ( .A(n14535), .B(n14536), .Z(n11424) );
  ANDN U15285 ( .B(n14537), .A(n14538), .Z(n14535) );
  XOR U15286 ( .A(n14539), .B(n10287), .Z(n8498) );
  XOR U15287 ( .A(n6312), .B(n14540), .Z(n14506) );
  XOR U15288 ( .A(n2395), .B(n5692), .Z(n14540) );
  XNOR U15289 ( .A(n14541), .B(n12005), .Z(n5692) );
  ANDN U15290 ( .B(n9824), .A(n9822), .Z(n14541) );
  IV U15291 ( .A(n12006), .Z(n9822) );
  XNOR U15292 ( .A(n14542), .B(n9959), .Z(n12006) );
  XNOR U15293 ( .A(n14154), .B(n13651), .Z(n9959) );
  XNOR U15294 ( .A(n14543), .B(n14544), .Z(n13651) );
  XOR U15295 ( .A(n12412), .B(n12171), .Z(n14544) );
  XNOR U15296 ( .A(n14545), .B(n14546), .Z(n12171) );
  ANDN U15297 ( .B(n14547), .A(n14548), .Z(n14545) );
  XNOR U15298 ( .A(n14549), .B(n14550), .Z(n12412) );
  ANDN U15299 ( .B(n14551), .A(n14552), .Z(n14549) );
  XOR U15300 ( .A(n12207), .B(n14553), .Z(n14543) );
  XNOR U15301 ( .A(n11108), .B(n12439), .Z(n14553) );
  XOR U15302 ( .A(n14554), .B(n14555), .Z(n12439) );
  ANDN U15303 ( .B(n14556), .A(n14557), .Z(n14554) );
  XOR U15304 ( .A(n14558), .B(n14559), .Z(n11108) );
  ANDN U15305 ( .B(n14560), .A(n14561), .Z(n14558) );
  XOR U15306 ( .A(n14562), .B(n14563), .Z(n12207) );
  ANDN U15307 ( .B(n14564), .A(n14565), .Z(n14562) );
  XOR U15308 ( .A(n14566), .B(n14567), .Z(n14154) );
  XNOR U15309 ( .A(n12915), .B(n11222), .Z(n14567) );
  XNOR U15310 ( .A(n14568), .B(n14569), .Z(n11222) );
  ANDN U15311 ( .B(n13783), .A(n14570), .Z(n14568) );
  XNOR U15312 ( .A(n14571), .B(n14572), .Z(n12915) );
  XOR U15313 ( .A(n9855), .B(n14574), .Z(n14566) );
  XOR U15314 ( .A(n10352), .B(n14575), .Z(n14574) );
  XOR U15315 ( .A(n14576), .B(n14577), .Z(n10352) );
  XOR U15316 ( .A(n14579), .B(n14580), .Z(n9855) );
  NOR U15317 ( .A(n14581), .B(n13766), .Z(n14579) );
  XNOR U15318 ( .A(n14582), .B(n11364), .Z(n9824) );
  XNOR U15319 ( .A(n14583), .B(n11996), .Z(n2395) );
  ANDN U15320 ( .B(n8490), .A(n11997), .Z(n14583) );
  XNOR U15321 ( .A(n14584), .B(n10990), .Z(n11997) );
  XOR U15322 ( .A(n13825), .B(n10075), .Z(n8490) );
  XNOR U15323 ( .A(n14585), .B(n14586), .Z(n13825) );
  ANDN U15324 ( .B(n14587), .A(n14588), .Z(n14585) );
  XNOR U15325 ( .A(n14589), .B(n12002), .Z(n6312) );
  AND U15326 ( .A(n8493), .B(n8492), .Z(n14589) );
  XOR U15327 ( .A(n14590), .B(n11103), .Z(n8492) );
  XOR U15328 ( .A(n14591), .B(n12232), .Z(n8493) );
  XOR U15329 ( .A(n10537), .B(n14592), .Z(n12232) );
  XOR U15330 ( .A(n14593), .B(n14594), .Z(n10537) );
  XOR U15331 ( .A(n11835), .B(n11070), .Z(n14594) );
  XOR U15332 ( .A(n14595), .B(n14596), .Z(n11070) );
  ANDN U15333 ( .B(n14597), .A(n14598), .Z(n14595) );
  XNOR U15334 ( .A(n14599), .B(n14018), .Z(n11835) );
  ANDN U15335 ( .B(n14600), .A(n14601), .Z(n14599) );
  XOR U15336 ( .A(n10093), .B(n14602), .Z(n14593) );
  XNOR U15337 ( .A(n9245), .B(n10998), .Z(n14602) );
  XNOR U15338 ( .A(n14603), .B(n14009), .Z(n10998) );
  ANDN U15339 ( .B(n14604), .A(n14008), .Z(n14603) );
  XOR U15340 ( .A(n14605), .B(n14606), .Z(n9245) );
  ANDN U15341 ( .B(n14607), .A(n14608), .Z(n14605) );
  XNOR U15342 ( .A(n14609), .B(n14610), .Z(n10093) );
  ANDN U15343 ( .B(n14005), .A(n14611), .Z(n14609) );
  XOR U15344 ( .A(n14612), .B(n14613), .Z(n8344) );
  XNOR U15345 ( .A(n3853), .B(n5163), .Z(n14613) );
  XOR U15346 ( .A(n14614), .B(n9715), .Z(n5163) );
  XNOR U15347 ( .A(n14615), .B(n9907), .Z(n9715) );
  NOR U15348 ( .A(n11677), .B(n11676), .Z(n14614) );
  XNOR U15349 ( .A(n14616), .B(n10990), .Z(n11676) );
  XNOR U15350 ( .A(n11588), .B(n12850), .Z(n10990) );
  XNOR U15351 ( .A(n14617), .B(n14618), .Z(n12850) );
  XNOR U15352 ( .A(n14619), .B(n11214), .Z(n14618) );
  XOR U15353 ( .A(n14620), .B(n14621), .Z(n11214) );
  NOR U15354 ( .A(n14622), .B(n14623), .Z(n14620) );
  XOR U15355 ( .A(n9976), .B(n14624), .Z(n14617) );
  XNOR U15356 ( .A(n10948), .B(n12618), .Z(n14624) );
  XNOR U15357 ( .A(n14625), .B(n14626), .Z(n12618) );
  NOR U15358 ( .A(n14627), .B(n14628), .Z(n14625) );
  XNOR U15359 ( .A(n14629), .B(n14630), .Z(n10948) );
  NOR U15360 ( .A(n14631), .B(n14632), .Z(n14629) );
  XNOR U15361 ( .A(n14633), .B(n14634), .Z(n9976) );
  ANDN U15362 ( .B(n14635), .A(n14636), .Z(n14633) );
  XOR U15363 ( .A(n14637), .B(n14638), .Z(n11588) );
  XOR U15364 ( .A(n9419), .B(n12522), .Z(n14638) );
  XOR U15365 ( .A(n14639), .B(n13683), .Z(n12522) );
  AND U15366 ( .A(n14640), .B(n14478), .Z(n14639) );
  XOR U15367 ( .A(n14641), .B(n14642), .Z(n9419) );
  ANDN U15368 ( .B(n13813), .A(n14643), .Z(n14641) );
  XOR U15369 ( .A(n10938), .B(n14644), .Z(n14637) );
  XNOR U15370 ( .A(n14323), .B(n12359), .Z(n14644) );
  XOR U15371 ( .A(n14645), .B(n13678), .Z(n12359) );
  ANDN U15372 ( .B(n14646), .A(n13810), .Z(n14645) );
  XOR U15373 ( .A(n14647), .B(n13688), .Z(n14323) );
  AND U15374 ( .A(n13815), .B(n14648), .Z(n14647) );
  XOR U15375 ( .A(n14649), .B(n13675), .Z(n10938) );
  ANDN U15376 ( .B(n14650), .A(n13817), .Z(n14649) );
  XNOR U15377 ( .A(n14651), .B(n11902), .Z(n11677) );
  XNOR U15378 ( .A(n14652), .B(n8405), .Z(n3853) );
  XOR U15379 ( .A(n14653), .B(n10343), .Z(n8405) );
  XNOR U15380 ( .A(n14654), .B(n13236), .Z(n10343) );
  XNOR U15381 ( .A(n14655), .B(n14656), .Z(n13236) );
  XOR U15382 ( .A(n13641), .B(n12903), .Z(n14656) );
  XOR U15383 ( .A(n14657), .B(n14658), .Z(n12903) );
  ANDN U15384 ( .B(n13227), .A(n13225), .Z(n14657) );
  XOR U15385 ( .A(n14659), .B(n14660), .Z(n13641) );
  ANDN U15386 ( .B(n13219), .A(n13217), .Z(n14659) );
  XNOR U15387 ( .A(n11613), .B(n14661), .Z(n14655) );
  XOR U15388 ( .A(n13702), .B(n12972), .Z(n14661) );
  XNOR U15389 ( .A(n14662), .B(n14663), .Z(n12972) );
  AND U15390 ( .A(n13223), .B(n13221), .Z(n14662) );
  XNOR U15391 ( .A(n14664), .B(n14665), .Z(n13702) );
  NOR U15392 ( .A(n14666), .B(n13212), .Z(n14664) );
  XOR U15393 ( .A(n14667), .B(n14668), .Z(n11613) );
  ANDN U15394 ( .B(n13238), .A(n14669), .Z(n14667) );
  AND U15395 ( .A(n11667), .B(n11669), .Z(n14652) );
  XOR U15396 ( .A(n11698), .B(n14269), .Z(n11669) );
  XNOR U15397 ( .A(n14670), .B(n14222), .Z(n14269) );
  ANDN U15398 ( .B(n13560), .A(n14671), .Z(n14670) );
  XOR U15399 ( .A(n14672), .B(n10180), .Z(n11667) );
  XNOR U15400 ( .A(n5510), .B(n14673), .Z(n14612) );
  XNOR U15401 ( .A(n1748), .B(n11977), .Z(n14673) );
  XNOR U15402 ( .A(n14674), .B(n8415), .Z(n11977) );
  XOR U15403 ( .A(n14675), .B(n11085), .Z(n8415) );
  XNOR U15404 ( .A(n13554), .B(n14676), .Z(n11085) );
  XOR U15405 ( .A(n14677), .B(n14678), .Z(n13554) );
  XOR U15406 ( .A(n14679), .B(n14680), .Z(n14678) );
  XOR U15407 ( .A(n9635), .B(n14681), .Z(n14677) );
  XNOR U15408 ( .A(n13464), .B(n14682), .Z(n14681) );
  XOR U15409 ( .A(n14683), .B(n14684), .Z(n13464) );
  NOR U15410 ( .A(n14685), .B(n13852), .Z(n14683) );
  XNOR U15411 ( .A(n14686), .B(n14687), .Z(n9635) );
  NOR U15412 ( .A(n14688), .B(n14689), .Z(n14686) );
  ANDN U15413 ( .B(n11663), .A(n11664), .Z(n14674) );
  XOR U15414 ( .A(n11106), .B(n14690), .Z(n11664) );
  XNOR U15415 ( .A(n14691), .B(n11869), .Z(n11663) );
  XNOR U15416 ( .A(n14692), .B(n13485), .Z(n11869) );
  XNOR U15417 ( .A(n14693), .B(n14694), .Z(n13485) );
  XOR U15418 ( .A(n10215), .B(n12197), .Z(n14694) );
  XNOR U15419 ( .A(n14695), .B(n14696), .Z(n12197) );
  ANDN U15420 ( .B(n14697), .A(n14698), .Z(n14695) );
  XOR U15421 ( .A(n14699), .B(n14700), .Z(n10215) );
  ANDN U15422 ( .B(n14701), .A(n14702), .Z(n14699) );
  XOR U15423 ( .A(n14703), .B(n14704), .Z(n14693) );
  XNOR U15424 ( .A(n11295), .B(n11063), .Z(n14704) );
  XNOR U15425 ( .A(n14705), .B(n14706), .Z(n11063) );
  ANDN U15426 ( .B(n14707), .A(n14708), .Z(n14705) );
  XOR U15427 ( .A(n14709), .B(n14710), .Z(n11295) );
  ANDN U15428 ( .B(n14711), .A(n14712), .Z(n14709) );
  XNOR U15429 ( .A(n14713), .B(n8408), .Z(n1748) );
  IV U15430 ( .A(n11982), .Z(n8408) );
  XOR U15431 ( .A(n14714), .B(n12369), .Z(n11982) );
  IV U15432 ( .A(n10396), .Z(n12369) );
  XNOR U15433 ( .A(n14715), .B(n14716), .Z(n14183) );
  XNOR U15434 ( .A(n14717), .B(n12629), .Z(n14716) );
  XNOR U15435 ( .A(n14718), .B(n14719), .Z(n12629) );
  NOR U15436 ( .A(n14720), .B(n13492), .Z(n14718) );
  XOR U15437 ( .A(n13379), .B(n14721), .Z(n14715) );
  XNOR U15438 ( .A(n11723), .B(n11647), .Z(n14721) );
  XOR U15439 ( .A(n14722), .B(n14723), .Z(n11647) );
  NOR U15440 ( .A(n13505), .B(n14724), .Z(n14722) );
  XNOR U15441 ( .A(n14725), .B(n14726), .Z(n11723) );
  NOR U15442 ( .A(n14727), .B(n14728), .Z(n14725) );
  XNOR U15443 ( .A(n14729), .B(n14730), .Z(n13379) );
  AND U15444 ( .A(n14731), .B(n13497), .Z(n14729) );
  NOR U15445 ( .A(n11981), .B(n11674), .Z(n14713) );
  XNOR U15446 ( .A(n14733), .B(n10185), .Z(n11674) );
  IV U15447 ( .A(n11673), .Z(n11981) );
  XOR U15448 ( .A(n9617), .B(n14734), .Z(n11673) );
  XNOR U15449 ( .A(n14735), .B(n12764), .Z(n9617) );
  XOR U15450 ( .A(n14736), .B(n14737), .Z(n12764) );
  XNOR U15451 ( .A(n13372), .B(n12725), .Z(n14737) );
  XOR U15452 ( .A(n14738), .B(n14102), .Z(n12725) );
  ANDN U15453 ( .B(n14739), .A(n14740), .Z(n14738) );
  XOR U15454 ( .A(n14741), .B(n14110), .Z(n13372) );
  ANDN U15455 ( .B(n14742), .A(n14743), .Z(n14741) );
  XOR U15456 ( .A(n11708), .B(n14744), .Z(n14736) );
  XOR U15457 ( .A(n10059), .B(n9135), .Z(n14744) );
  XNOR U15458 ( .A(n14745), .B(n14105), .Z(n9135) );
  ANDN U15459 ( .B(n14746), .A(n14747), .Z(n14745) );
  XNOR U15460 ( .A(n14748), .B(n14096), .Z(n10059) );
  ANDN U15461 ( .B(n14749), .A(n14750), .Z(n14748) );
  XNOR U15462 ( .A(n14751), .B(n14752), .Z(n11708) );
  ANDN U15463 ( .B(n14753), .A(n14754), .Z(n14751) );
  XNOR U15464 ( .A(n14755), .B(n8418), .Z(n5510) );
  XNOR U15465 ( .A(n14756), .B(n10287), .Z(n8418) );
  XOR U15466 ( .A(n14757), .B(n11986), .Z(n11670) );
  XNOR U15467 ( .A(n13576), .B(n9932), .Z(n11986) );
  XNOR U15468 ( .A(n14758), .B(n14759), .Z(n9932) );
  XOR U15469 ( .A(n14760), .B(n14761), .Z(n13576) );
  ANDN U15470 ( .B(n14207), .A(n14762), .Z(n14760) );
  ANDN U15471 ( .B(n13728), .A(n8417), .Z(n14757) );
  XNOR U15472 ( .A(n14763), .B(n10269), .Z(n8417) );
  XNOR U15473 ( .A(n12247), .B(n14764), .Z(n13728) );
  XOR U15474 ( .A(n12022), .B(n11832), .Z(n12247) );
  XOR U15475 ( .A(n14765), .B(n14766), .Z(n11832) );
  XNOR U15476 ( .A(n10821), .B(n11321), .Z(n14766) );
  XOR U15477 ( .A(n14767), .B(n14768), .Z(n11321) );
  ANDN U15478 ( .B(n14769), .A(n14770), .Z(n14767) );
  XNOR U15479 ( .A(n14771), .B(n14772), .Z(n10821) );
  ANDN U15480 ( .B(n14773), .A(n14774), .Z(n14771) );
  XNOR U15481 ( .A(n10335), .B(n14775), .Z(n14765) );
  XOR U15482 ( .A(n9423), .B(n11200), .Z(n14775) );
  XOR U15483 ( .A(n14776), .B(n14777), .Z(n11200) );
  ANDN U15484 ( .B(n14778), .A(n14779), .Z(n14776) );
  XNOR U15485 ( .A(n14780), .B(n14781), .Z(n9423) );
  XNOR U15486 ( .A(n14784), .B(n14785), .Z(n10335) );
  ANDN U15487 ( .B(n14786), .A(n14787), .Z(n14784) );
  XNOR U15488 ( .A(n14788), .B(n14789), .Z(n12022) );
  XNOR U15489 ( .A(n11423), .B(n10203), .Z(n14789) );
  XNOR U15490 ( .A(n14790), .B(n14791), .Z(n10203) );
  ANDN U15491 ( .B(n14792), .A(n14793), .Z(n14790) );
  XNOR U15492 ( .A(n14794), .B(n14795), .Z(n11423) );
  ANDN U15493 ( .B(n14796), .A(n14797), .Z(n14794) );
  XOR U15494 ( .A(n14798), .B(n14799), .Z(n14788) );
  XOR U15495 ( .A(n9555), .B(n14800), .Z(n14799) );
  XOR U15496 ( .A(n14801), .B(n14802), .Z(n9555) );
  NOR U15497 ( .A(n14803), .B(n14804), .Z(n14801) );
  XNOR U15498 ( .A(n8936), .B(n4293), .Z(n5705) );
  XNOR U15499 ( .A(n14805), .B(n14806), .Z(n6530) );
  XNOR U15500 ( .A(n5868), .B(n2541), .Z(n14806) );
  XNOR U15501 ( .A(n14807), .B(n6579), .Z(n2541) );
  XNOR U15502 ( .A(n9113), .B(n14808), .Z(n6579) );
  XNOR U15503 ( .A(n13039), .B(n14809), .Z(n9113) );
  XOR U15504 ( .A(n14810), .B(n14811), .Z(n13039) );
  XNOR U15505 ( .A(n9117), .B(n11607), .Z(n14811) );
  XOR U15506 ( .A(n14812), .B(n14813), .Z(n11607) );
  NOR U15507 ( .A(n14814), .B(n14815), .Z(n14812) );
  XOR U15508 ( .A(n14816), .B(n14817), .Z(n9117) );
  ANDN U15509 ( .B(n14818), .A(n14819), .Z(n14816) );
  XNOR U15510 ( .A(n14820), .B(n14821), .Z(n14810) );
  XNOR U15511 ( .A(n14822), .B(n11507), .Z(n14821) );
  XNOR U15512 ( .A(n14823), .B(n14824), .Z(n11507) );
  ANDN U15513 ( .B(n14825), .A(n14826), .Z(n14823) );
  ANDN U15514 ( .B(n8943), .A(n9016), .Z(n14807) );
  XOR U15515 ( .A(n12830), .B(n10057), .Z(n9016) );
  XOR U15516 ( .A(n14827), .B(n14828), .Z(n12830) );
  NOR U15517 ( .A(n14829), .B(n14830), .Z(n14827) );
  XOR U15518 ( .A(n14831), .B(n13277), .Z(n8943) );
  IV U15519 ( .A(n10855), .Z(n13277) );
  XOR U15520 ( .A(n14515), .B(n14832), .Z(n10855) );
  XOR U15521 ( .A(n14833), .B(n14834), .Z(n14515) );
  XOR U15522 ( .A(n14835), .B(n10753), .Z(n14834) );
  XOR U15523 ( .A(n14836), .B(n14837), .Z(n10753) );
  ANDN U15524 ( .B(n14838), .A(n14409), .Z(n14836) );
  XNOR U15525 ( .A(n12327), .B(n14839), .Z(n14833) );
  XNOR U15526 ( .A(n12590), .B(n12579), .Z(n14839) );
  XNOR U15527 ( .A(n14840), .B(n14841), .Z(n12579) );
  AND U15528 ( .A(n14842), .B(n14400), .Z(n14840) );
  XOR U15529 ( .A(n14843), .B(n14844), .Z(n12590) );
  ANDN U15530 ( .B(n14845), .A(n14846), .Z(n14843) );
  XNOR U15531 ( .A(n14847), .B(n14848), .Z(n12327) );
  ANDN U15532 ( .B(n14413), .A(n14849), .Z(n14847) );
  XNOR U15533 ( .A(n14850), .B(n6571), .Z(n5868) );
  XOR U15534 ( .A(n14851), .B(n11440), .Z(n6571) );
  XOR U15535 ( .A(n14852), .B(n12662), .Z(n11440) );
  XNOR U15536 ( .A(n14853), .B(n14854), .Z(n12662) );
  XNOR U15537 ( .A(n12754), .B(n11496), .Z(n14854) );
  XOR U15538 ( .A(n14855), .B(n14318), .Z(n11496) );
  ANDN U15539 ( .B(n14856), .A(n14317), .Z(n14855) );
  XNOR U15540 ( .A(n14857), .B(n14308), .Z(n12754) );
  ANDN U15541 ( .B(n14858), .A(n14309), .Z(n14857) );
  XOR U15542 ( .A(n12744), .B(n14859), .Z(n14853) );
  XOR U15543 ( .A(n11748), .B(n10525), .Z(n14859) );
  XNOR U15544 ( .A(n14860), .B(n14313), .Z(n10525) );
  NOR U15545 ( .A(n14861), .B(n14862), .Z(n14860) );
  XNOR U15546 ( .A(n14863), .B(n14864), .Z(n11748) );
  ANDN U15547 ( .B(n14865), .A(n14866), .Z(n14863) );
  XNOR U15548 ( .A(n14867), .B(n14322), .Z(n12744) );
  ANDN U15549 ( .B(n14868), .A(n14321), .Z(n14867) );
  ANDN U15550 ( .B(n9013), .A(n14128), .Z(n14850) );
  XNOR U15551 ( .A(n3515), .B(n14869), .Z(n14805) );
  XOR U15552 ( .A(n9006), .B(n4893), .Z(n14869) );
  XNOR U15553 ( .A(n14870), .B(n6566), .Z(n4893) );
  XOR U15554 ( .A(n14871), .B(n12713), .Z(n6566) );
  ANDN U15555 ( .B(n8939), .A(n8938), .Z(n14870) );
  XOR U15556 ( .A(n12311), .B(n13341), .Z(n8938) );
  XNOR U15557 ( .A(n14872), .B(n14873), .Z(n13341) );
  ANDN U15558 ( .B(n14874), .A(n14875), .Z(n14872) );
  IV U15559 ( .A(n11433), .Z(n12311) );
  XOR U15560 ( .A(n14090), .B(n14876), .Z(n11433) );
  XOR U15561 ( .A(n14877), .B(n14878), .Z(n14090) );
  XOR U15562 ( .A(n9805), .B(n10264), .Z(n14878) );
  XNOR U15563 ( .A(n14879), .B(n14880), .Z(n10264) );
  ANDN U15564 ( .B(n14881), .A(n13460), .Z(n14879) );
  XNOR U15565 ( .A(n14882), .B(n14883), .Z(n9805) );
  ANDN U15566 ( .B(n14884), .A(n13446), .Z(n14882) );
  XOR U15567 ( .A(n13724), .B(n14885), .Z(n14877) );
  XNOR U15568 ( .A(n9508), .B(n13911), .Z(n14885) );
  XNOR U15569 ( .A(n14886), .B(n14887), .Z(n13911) );
  NOR U15570 ( .A(n14888), .B(n14889), .Z(n14886) );
  XNOR U15571 ( .A(n14890), .B(n14891), .Z(n9508) );
  ANDN U15572 ( .B(n13450), .A(n14892), .Z(n14890) );
  XNOR U15573 ( .A(n14893), .B(n14894), .Z(n13724) );
  ANDN U15574 ( .B(n14895), .A(n13456), .Z(n14893) );
  XNOR U15575 ( .A(n14896), .B(n10962), .Z(n8939) );
  XNOR U15576 ( .A(n14897), .B(n6561), .Z(n9006) );
  XOR U15577 ( .A(n11637), .B(n13430), .Z(n6561) );
  XNOR U15578 ( .A(n14898), .B(n14899), .Z(n13430) );
  ANDN U15579 ( .B(n14034), .A(n14035), .Z(n14898) );
  ANDN U15580 ( .B(n8934), .A(n8933), .Z(n14897) );
  XOR U15581 ( .A(n14900), .B(n10496), .Z(n8933) );
  XNOR U15582 ( .A(n14901), .B(n11352), .Z(n8934) );
  IV U15583 ( .A(n11239), .Z(n11352) );
  XNOR U15584 ( .A(n14902), .B(n6574), .Z(n3515) );
  XOR U15585 ( .A(n14903), .B(n9795), .Z(n6574) );
  IV U15586 ( .A(n9815), .Z(n9795) );
  XOR U15587 ( .A(n14904), .B(n13306), .Z(n9815) );
  XOR U15588 ( .A(n14905), .B(n14906), .Z(n13306) );
  XOR U15589 ( .A(n13589), .B(n10112), .Z(n14906) );
  XNOR U15590 ( .A(n14907), .B(n14908), .Z(n10112) );
  NOR U15591 ( .A(n14909), .B(n14910), .Z(n14907) );
  XNOR U15592 ( .A(n14911), .B(n14912), .Z(n13589) );
  ANDN U15593 ( .B(n14913), .A(n14914), .Z(n14911) );
  XOR U15594 ( .A(n10218), .B(n14915), .Z(n14905) );
  XNOR U15595 ( .A(n12696), .B(n14916), .Z(n14915) );
  XOR U15596 ( .A(n14917), .B(n14918), .Z(n12696) );
  ANDN U15597 ( .B(n14919), .A(n14920), .Z(n14917) );
  XNOR U15598 ( .A(n14921), .B(n14922), .Z(n10218) );
  ANDN U15599 ( .B(n14923), .A(n14924), .Z(n14921) );
  ANDN U15600 ( .B(n8930), .A(n8929), .Z(n14902) );
  XOR U15601 ( .A(n14925), .B(n9879), .Z(n8929) );
  XNOR U15602 ( .A(n14926), .B(n14927), .Z(n9879) );
  XOR U15603 ( .A(n14928), .B(n14929), .Z(n8930) );
  XOR U15604 ( .A(n14930), .B(n14931), .Z(n6352) );
  XOR U15605 ( .A(n5479), .B(n3729), .Z(n14931) );
  XOR U15606 ( .A(n14932), .B(n14933), .Z(n3729) );
  ANDN U15607 ( .B(n6590), .A(n6591), .Z(n14932) );
  XNOR U15608 ( .A(n12831), .B(n10057), .Z(n6591) );
  XOR U15609 ( .A(n14934), .B(n14935), .Z(n12661) );
  XOR U15610 ( .A(n11447), .B(n9869), .Z(n14935) );
  XOR U15611 ( .A(n14936), .B(n14937), .Z(n9869) );
  XNOR U15612 ( .A(n14940), .B(n14941), .Z(n11447) );
  XOR U15613 ( .A(n10922), .B(n14942), .Z(n14934) );
  XNOR U15614 ( .A(n12112), .B(n14943), .Z(n14942) );
  NOR U15615 ( .A(n12824), .B(n12822), .Z(n14944) );
  XNOR U15616 ( .A(n14946), .B(n14947), .Z(n10922) );
  ANDN U15617 ( .B(n12827), .A(n12826), .Z(n14946) );
  XOR U15618 ( .A(n14948), .B(n14949), .Z(n13289) );
  XOR U15619 ( .A(n9237), .B(n12210), .Z(n14949) );
  XNOR U15620 ( .A(n14950), .B(n14951), .Z(n12210) );
  NOR U15621 ( .A(n13292), .B(n13291), .Z(n14950) );
  XOR U15622 ( .A(n14952), .B(n14953), .Z(n13292) );
  XNOR U15623 ( .A(n14954), .B(n14955), .Z(n9237) );
  NOR U15624 ( .A(n14956), .B(n12940), .Z(n14954) );
  XOR U15625 ( .A(n14957), .B(n14958), .Z(n12940) );
  XOR U15626 ( .A(n12062), .B(n14959), .Z(n14948) );
  XNOR U15627 ( .A(n10702), .B(n13116), .Z(n14959) );
  XNOR U15628 ( .A(n14960), .B(n14961), .Z(n13116) );
  ANDN U15629 ( .B(n12936), .A(n13173), .Z(n14960) );
  XOR U15630 ( .A(n14962), .B(n14963), .Z(n12936) );
  XNOR U15631 ( .A(n14964), .B(n14965), .Z(n10702) );
  ANDN U15632 ( .B(n12944), .A(n13273), .Z(n14964) );
  XOR U15633 ( .A(n14966), .B(n14967), .Z(n12944) );
  XNOR U15634 ( .A(n14968), .B(n14969), .Z(n12062) );
  ANDN U15635 ( .B(n13179), .A(n12931), .Z(n14968) );
  XOR U15636 ( .A(n14970), .B(n14971), .Z(n12931) );
  XNOR U15637 ( .A(n14972), .B(n14938), .Z(n12831) );
  ANDN U15638 ( .B(n14973), .A(n14939), .Z(n14972) );
  XNOR U15639 ( .A(n14974), .B(n9024), .Z(n5479) );
  ANDN U15640 ( .B(n6599), .A(n6600), .Z(n14974) );
  XOR U15641 ( .A(n14975), .B(n14929), .Z(n6600) );
  XNOR U15642 ( .A(n14976), .B(n14977), .Z(n6599) );
  XOR U15643 ( .A(n4342), .B(n14978), .Z(n14930) );
  XOR U15644 ( .A(n5931), .B(n2132), .Z(n14978) );
  XOR U15645 ( .A(n14979), .B(n9021), .Z(n2132) );
  ANDN U15646 ( .B(n6595), .A(n6597), .Z(n14979) );
  XOR U15647 ( .A(n10380), .B(n14980), .Z(n6597) );
  XOR U15648 ( .A(n14981), .B(n9755), .Z(n6595) );
  XNOR U15649 ( .A(n14982), .B(n12265), .Z(n9755) );
  XOR U15650 ( .A(n14983), .B(n14984), .Z(n12265) );
  XNOR U15651 ( .A(n14542), .B(n12432), .Z(n14984) );
  XOR U15652 ( .A(n14985), .B(n14986), .Z(n12432) );
  NOR U15653 ( .A(n13771), .B(n13770), .Z(n14985) );
  XNOR U15654 ( .A(n14987), .B(n14581), .Z(n14542) );
  ANDN U15655 ( .B(n13766), .A(n13767), .Z(n14987) );
  XOR U15656 ( .A(n14988), .B(n14989), .Z(n13766) );
  XNOR U15657 ( .A(n12087), .B(n14990), .Z(n14983) );
  XOR U15658 ( .A(n9958), .B(n12758), .Z(n14990) );
  XNOR U15659 ( .A(n14991), .B(n14570), .Z(n12758) );
  XNOR U15660 ( .A(n14992), .B(n14993), .Z(n13783) );
  XNOR U15661 ( .A(n14994), .B(n14578), .Z(n9958) );
  ANDN U15662 ( .B(n13777), .A(n13775), .Z(n14994) );
  XOR U15663 ( .A(n14995), .B(n14996), .Z(n13775) );
  XOR U15664 ( .A(n14997), .B(n14573), .Z(n12087) );
  ANDN U15665 ( .B(n13779), .A(n13780), .Z(n14997) );
  XNOR U15666 ( .A(n14998), .B(n14999), .Z(n13779) );
  XOR U15667 ( .A(n15000), .B(n9032), .Z(n5931) );
  ANDN U15668 ( .B(n6588), .A(n6586), .Z(n15000) );
  XOR U15669 ( .A(n9765), .B(n15001), .Z(n6586) );
  XOR U15670 ( .A(n10202), .B(n14800), .Z(n6588) );
  XOR U15671 ( .A(n15002), .B(n15003), .Z(n14800) );
  ANDN U15672 ( .B(n15004), .A(n15005), .Z(n15002) );
  XNOR U15673 ( .A(n15006), .B(n9029), .Z(n4342) );
  ANDN U15674 ( .B(n6605), .A(n6603), .Z(n15006) );
  XOR U15675 ( .A(n15007), .B(n11239), .Z(n6603) );
  XOR U15676 ( .A(n15008), .B(n11580), .Z(n11239) );
  XNOR U15677 ( .A(n15009), .B(n15010), .Z(n11580) );
  XNOR U15678 ( .A(n12752), .B(n11609), .Z(n15010) );
  XNOR U15679 ( .A(n15011), .B(n15012), .Z(n11609) );
  ANDN U15680 ( .B(n15013), .A(n15014), .Z(n15011) );
  XNOR U15681 ( .A(n15015), .B(n15016), .Z(n12752) );
  ANDN U15682 ( .B(n15017), .A(n15018), .Z(n15015) );
  XNOR U15683 ( .A(n9460), .B(n15019), .Z(n15009) );
  XOR U15684 ( .A(n15020), .B(n12718), .Z(n15019) );
  XNOR U15685 ( .A(n15021), .B(n15022), .Z(n12718) );
  ANDN U15686 ( .B(n15023), .A(n15024), .Z(n15021) );
  XOR U15687 ( .A(n15025), .B(n15026), .Z(n9460) );
  AND U15688 ( .A(n15027), .B(n15028), .Z(n15025) );
  XNOR U15689 ( .A(n15029), .B(n9907), .Z(n6605) );
  IV U15690 ( .A(n9800), .Z(n9907) );
  XNOR U15691 ( .A(n15030), .B(n14876), .Z(n9800) );
  XNOR U15692 ( .A(n15031), .B(n15032), .Z(n14876) );
  XNOR U15693 ( .A(n11561), .B(n12509), .Z(n15032) );
  XNOR U15694 ( .A(n15033), .B(n15034), .Z(n12509) );
  XNOR U15695 ( .A(n15035), .B(n15036), .Z(n11561) );
  XOR U15696 ( .A(n10744), .B(n15037), .Z(n15031) );
  XNOR U15697 ( .A(n11315), .B(n15038), .Z(n15037) );
  XOR U15698 ( .A(n15039), .B(n15040), .Z(n11315) );
  AND U15699 ( .A(n13346), .B(n13344), .Z(n15039) );
  XNOR U15700 ( .A(n15041), .B(n15042), .Z(n10744) );
  AND U15701 ( .A(n13338), .B(n13340), .Z(n15041) );
  XNOR U15702 ( .A(n15043), .B(n9013), .Z(n8936) );
  XNOR U15703 ( .A(n15044), .B(n12419), .Z(n9013) );
  IV U15704 ( .A(n12685), .Z(n12419) );
  XOR U15705 ( .A(n13903), .B(n11515), .Z(n6569) );
  XOR U15706 ( .A(n15045), .B(n15046), .Z(n11515) );
  XNOR U15707 ( .A(n15047), .B(n15048), .Z(n13903) );
  NOR U15708 ( .A(n15049), .B(n15050), .Z(n15047) );
  XNOR U15709 ( .A(n15051), .B(n9524), .Z(n14128) );
  XOR U15710 ( .A(n15052), .B(n6240), .Z(out[1000]) );
  XOR U15711 ( .A(n9192), .B(n2317), .Z(n6240) );
  XNOR U15712 ( .A(n10145), .B(n6199), .Z(n2317) );
  XNOR U15713 ( .A(n15053), .B(n15054), .Z(n6199) );
  XOR U15714 ( .A(n2351), .B(n5493), .Z(n15054) );
  XNOR U15715 ( .A(n15055), .B(n10069), .Z(n5493) );
  IV U15716 ( .A(n8054), .Z(n10069) );
  XOR U15717 ( .A(n15056), .B(n13569), .Z(n8054) );
  XNOR U15718 ( .A(n15057), .B(n14272), .Z(n13569) );
  ANDN U15719 ( .B(n14219), .A(n14218), .Z(n15057) );
  AND U15720 ( .A(n9203), .B(n8055), .Z(n15055) );
  XNOR U15721 ( .A(n12692), .B(n15058), .Z(n8055) );
  IV U15722 ( .A(n10380), .Z(n12692) );
  XNOR U15723 ( .A(n13633), .B(n15059), .Z(n10380) );
  XOR U15724 ( .A(n15060), .B(n15061), .Z(n13633) );
  XNOR U15725 ( .A(n12400), .B(n10301), .Z(n15061) );
  XNOR U15726 ( .A(n15062), .B(n15063), .Z(n10301) );
  XOR U15727 ( .A(n15066), .B(n15067), .Z(n12400) );
  ANDN U15728 ( .B(n15068), .A(n15069), .Z(n15066) );
  XNOR U15729 ( .A(n10387), .B(n15070), .Z(n15060) );
  XOR U15730 ( .A(n15071), .B(n15072), .Z(n15070) );
  XOR U15731 ( .A(n15073), .B(n15074), .Z(n10387) );
  NOR U15732 ( .A(n15075), .B(n15076), .Z(n15073) );
  XOR U15733 ( .A(n15077), .B(n9426), .Z(n9203) );
  XOR U15734 ( .A(n13279), .B(n15078), .Z(n9426) );
  XOR U15735 ( .A(n15079), .B(n15080), .Z(n13279) );
  XNOR U15736 ( .A(n10260), .B(n10875), .Z(n15080) );
  XNOR U15737 ( .A(n15081), .B(n15082), .Z(n10875) );
  ANDN U15738 ( .B(n15083), .A(n15084), .Z(n15081) );
  XNOR U15739 ( .A(n15085), .B(n15086), .Z(n10260) );
  ANDN U15740 ( .B(n15087), .A(n13402), .Z(n15085) );
  XOR U15741 ( .A(n9945), .B(n15088), .Z(n15079) );
  XOR U15742 ( .A(n15089), .B(n11777), .Z(n15088) );
  ANDN U15743 ( .B(n15092), .A(n13412), .Z(n15090) );
  XNOR U15744 ( .A(n15093), .B(n15094), .Z(n9945) );
  ANDN U15745 ( .B(n15095), .A(n13408), .Z(n15093) );
  XNOR U15746 ( .A(n15096), .B(n9174), .Z(n2351) );
  XNOR U15747 ( .A(n14116), .B(n10108), .Z(n9174) );
  XNOR U15748 ( .A(n15097), .B(n15098), .Z(n14116) );
  AND U15749 ( .A(n15099), .B(n15100), .Z(n15097) );
  ANDN U15750 ( .B(n9198), .A(n9197), .Z(n15096) );
  XNOR U15751 ( .A(n14679), .B(n9636), .Z(n9197) );
  XOR U15752 ( .A(n15101), .B(n15102), .Z(n14679) );
  ANDN U15753 ( .B(n13862), .A(n15103), .Z(n15101) );
  XOR U15754 ( .A(n15104), .B(n12843), .Z(n9198) );
  XOR U15755 ( .A(n15105), .B(n12970), .Z(n12843) );
  XOR U15756 ( .A(n15106), .B(n15107), .Z(n12970) );
  XNOR U15757 ( .A(n10083), .B(n12279), .Z(n15107) );
  XOR U15758 ( .A(n15108), .B(n15109), .Z(n12279) );
  ANDN U15759 ( .B(n15110), .A(n14283), .Z(n15108) );
  XNOR U15760 ( .A(n15111), .B(n15112), .Z(n10083) );
  ANDN U15761 ( .B(n15113), .A(n15114), .Z(n15111) );
  XOR U15762 ( .A(n12053), .B(n15115), .Z(n15106) );
  XOR U15763 ( .A(n11807), .B(n15116), .Z(n15115) );
  XNOR U15764 ( .A(n15117), .B(n15118), .Z(n11807) );
  ANDN U15765 ( .B(n15119), .A(n15120), .Z(n15117) );
  XOR U15766 ( .A(n15121), .B(n15122), .Z(n12053) );
  ANDN U15767 ( .B(n15123), .A(n14293), .Z(n15121) );
  XOR U15768 ( .A(n3179), .B(n15124), .Z(n15053) );
  XOR U15769 ( .A(n6374), .B(n8048), .Z(n15124) );
  XNOR U15770 ( .A(n15125), .B(n8063), .Z(n8048) );
  XOR U15771 ( .A(n9252), .B(n15126), .Z(n8063) );
  XNOR U15772 ( .A(n15030), .B(n12067), .Z(n9252) );
  XOR U15773 ( .A(n15127), .B(n15128), .Z(n12067) );
  XOR U15774 ( .A(n12382), .B(n13205), .Z(n15128) );
  XOR U15775 ( .A(n15129), .B(n14712), .Z(n13205) );
  NOR U15776 ( .A(n14711), .B(n15130), .Z(n15129) );
  XNOR U15777 ( .A(n15131), .B(n15132), .Z(n12382) );
  NOR U15778 ( .A(n15133), .B(n15134), .Z(n15131) );
  XNOR U15779 ( .A(n11868), .B(n15135), .Z(n15127) );
  XNOR U15780 ( .A(n14691), .B(n13415), .Z(n15135) );
  XNOR U15781 ( .A(n15136), .B(n14697), .Z(n13415) );
  XOR U15782 ( .A(n15138), .B(n14702), .Z(n14691) );
  NOR U15783 ( .A(n15139), .B(n14701), .Z(n15138) );
  XOR U15784 ( .A(n15140), .B(n14708), .Z(n11868) );
  NOR U15785 ( .A(n15141), .B(n14707), .Z(n15140) );
  XOR U15786 ( .A(n15142), .B(n15143), .Z(n15030) );
  XNOR U15787 ( .A(n9449), .B(n12222), .Z(n15143) );
  XNOR U15788 ( .A(n15144), .B(n15145), .Z(n12222) );
  NOR U15789 ( .A(n15146), .B(n15147), .Z(n15144) );
  XOR U15790 ( .A(n15148), .B(n15149), .Z(n9449) );
  NOR U15791 ( .A(n15150), .B(n15151), .Z(n15148) );
  XOR U15792 ( .A(n12997), .B(n15152), .Z(n15142) );
  XNOR U15793 ( .A(n15153), .B(n12086), .Z(n15152) );
  XOR U15794 ( .A(n15154), .B(n15155), .Z(n12086) );
  NOR U15795 ( .A(n15156), .B(n15157), .Z(n15154) );
  XNOR U15796 ( .A(n15158), .B(n15159), .Z(n12997) );
  ANDN U15797 ( .B(n8064), .A(n9200), .Z(n15125) );
  XOR U15798 ( .A(n9515), .B(n15162), .Z(n9200) );
  XNOR U15799 ( .A(n12645), .B(n15163), .Z(n9515) );
  XOR U15800 ( .A(n15164), .B(n15165), .Z(n12645) );
  XOR U15801 ( .A(n11841), .B(n11713), .Z(n15165) );
  XOR U15802 ( .A(n15166), .B(n15167), .Z(n11713) );
  XOR U15803 ( .A(n15170), .B(n14636), .Z(n11841) );
  IV U15804 ( .A(n15171), .Z(n14636) );
  ANDN U15805 ( .B(n15172), .A(n15173), .Z(n15170) );
  XOR U15806 ( .A(n12073), .B(n15174), .Z(n15164) );
  XOR U15807 ( .A(n15175), .B(n15176), .Z(n15174) );
  XNOR U15808 ( .A(n15177), .B(n14622), .Z(n12073) );
  ANDN U15809 ( .B(n15178), .A(n15179), .Z(n15177) );
  XNOR U15810 ( .A(n15180), .B(n11877), .Z(n8064) );
  IV U15811 ( .A(n11045), .Z(n11877) );
  XNOR U15812 ( .A(n12926), .B(n15181), .Z(n11045) );
  XOR U15813 ( .A(n15182), .B(n15183), .Z(n12926) );
  XNOR U15814 ( .A(n12818), .B(n12078), .Z(n15183) );
  XNOR U15815 ( .A(n15184), .B(n12824), .Z(n12078) );
  XOR U15816 ( .A(n15185), .B(n15186), .Z(n12824) );
  NOR U15817 ( .A(n15187), .B(n12823), .Z(n15184) );
  XNOR U15818 ( .A(n15188), .B(n14829), .Z(n12818) );
  ANDN U15819 ( .B(n14830), .A(n15189), .Z(n15188) );
  XNOR U15820 ( .A(n11712), .B(n15190), .Z(n15182) );
  XOR U15821 ( .A(n9144), .B(n11823), .Z(n15190) );
  XNOR U15822 ( .A(n15191), .B(n14939), .Z(n11823) );
  XOR U15823 ( .A(n15192), .B(n15193), .Z(n14939) );
  NOR U15824 ( .A(n14973), .B(n15194), .Z(n15191) );
  XOR U15825 ( .A(n15195), .B(n12827), .Z(n9144) );
  XOR U15826 ( .A(n15196), .B(n15197), .Z(n12827) );
  ANDN U15827 ( .B(n12828), .A(n15198), .Z(n15195) );
  XNOR U15828 ( .A(n15199), .B(n12835), .Z(n11712) );
  XNOR U15829 ( .A(n15200), .B(n15201), .Z(n12835) );
  ANDN U15830 ( .B(n15202), .A(n12834), .Z(n15199) );
  XNOR U15831 ( .A(n15203), .B(n8068), .Z(n6374) );
  XNOR U15832 ( .A(n15204), .B(n12713), .Z(n8068) );
  ANDN U15833 ( .B(n14480), .A(n15205), .Z(n15203) );
  XNOR U15834 ( .A(n15206), .B(n8071), .Z(n3179) );
  XNOR U15835 ( .A(n15207), .B(n11043), .Z(n8071) );
  XNOR U15836 ( .A(n14367), .B(n13422), .Z(n11043) );
  XNOR U15837 ( .A(n15208), .B(n15209), .Z(n13422) );
  XOR U15838 ( .A(n12815), .B(n10605), .Z(n15209) );
  XNOR U15839 ( .A(n15210), .B(n14059), .Z(n10605) );
  AND U15840 ( .A(n15211), .B(n15212), .Z(n15210) );
  XOR U15841 ( .A(n15213), .B(n15214), .Z(n12815) );
  ANDN U15842 ( .B(n15215), .A(n15216), .Z(n15213) );
  XNOR U15843 ( .A(n10712), .B(n15217), .Z(n15208) );
  XOR U15844 ( .A(n12612), .B(n12583), .Z(n15217) );
  XOR U15845 ( .A(n15218), .B(n14064), .Z(n12583) );
  AND U15846 ( .A(n15219), .B(n15220), .Z(n15218) );
  XNOR U15847 ( .A(n15221), .B(n15222), .Z(n12612) );
  NOR U15848 ( .A(n15223), .B(n15224), .Z(n15221) );
  XOR U15849 ( .A(n15225), .B(n14050), .Z(n10712) );
  ANDN U15850 ( .B(n15226), .A(n15227), .Z(n15225) );
  XOR U15851 ( .A(n15228), .B(n15229), .Z(n14367) );
  XNOR U15852 ( .A(n15230), .B(n10121), .Z(n15229) );
  XOR U15853 ( .A(n15231), .B(n14078), .Z(n10121) );
  ANDN U15854 ( .B(n15232), .A(n15233), .Z(n15231) );
  XOR U15855 ( .A(n12190), .B(n15234), .Z(n15228) );
  XOR U15856 ( .A(n11100), .B(n12180), .Z(n15234) );
  XNOR U15857 ( .A(n15235), .B(n14086), .Z(n12180) );
  AND U15858 ( .A(n15236), .B(n15237), .Z(n15235) );
  XNOR U15859 ( .A(n15238), .B(n14082), .Z(n11100) );
  ANDN U15860 ( .B(n15239), .A(n15240), .Z(n15238) );
  XNOR U15861 ( .A(n15241), .B(n15242), .Z(n12190) );
  AND U15862 ( .A(n15243), .B(n15244), .Z(n15241) );
  ANDN U15863 ( .B(n9194), .A(n8072), .Z(n15206) );
  XOR U15864 ( .A(n9102), .B(n15245), .Z(n8072) );
  IV U15865 ( .A(n12880), .Z(n9102) );
  XNOR U15866 ( .A(n15246), .B(n14514), .Z(n12880) );
  XNOR U15867 ( .A(n15247), .B(n15248), .Z(n14514) );
  XOR U15868 ( .A(n10835), .B(n12771), .Z(n15248) );
  XNOR U15869 ( .A(n15249), .B(n15250), .Z(n12771) );
  NOR U15870 ( .A(n13147), .B(n13145), .Z(n15249) );
  XOR U15871 ( .A(n15251), .B(n15252), .Z(n13147) );
  XNOR U15872 ( .A(n15253), .B(n15254), .Z(n10835) );
  ANDN U15873 ( .B(n13154), .A(n13153), .Z(n15253) );
  XOR U15874 ( .A(n15255), .B(n15256), .Z(n13154) );
  XOR U15875 ( .A(n13644), .B(n15257), .Z(n15247) );
  XNOR U15876 ( .A(n11242), .B(n11582), .Z(n15257) );
  XOR U15877 ( .A(n15258), .B(n15259), .Z(n11582) );
  ANDN U15878 ( .B(n13142), .A(n13140), .Z(n15258) );
  XOR U15879 ( .A(n15260), .B(n15261), .Z(n13142) );
  XNOR U15880 ( .A(n15262), .B(n15263), .Z(n11242) );
  ANDN U15881 ( .B(n13955), .A(n14512), .Z(n15262) );
  XOR U15882 ( .A(n15264), .B(n15265), .Z(n13955) );
  XNOR U15883 ( .A(n15266), .B(n15267), .Z(n13644) );
  ANDN U15884 ( .B(n13149), .A(n13150), .Z(n15266) );
  XOR U15885 ( .A(n15268), .B(n15269), .Z(n13150) );
  XNOR U15886 ( .A(n15270), .B(n9277), .Z(n9194) );
  XOR U15887 ( .A(n15271), .B(n15272), .Z(n10145) );
  XNOR U15888 ( .A(n5104), .B(n1956), .Z(n15272) );
  XOR U15889 ( .A(n15273), .B(n7985), .Z(n1956) );
  XOR U15890 ( .A(n12351), .B(n10521), .Z(n7985) );
  XOR U15891 ( .A(n15274), .B(n15275), .Z(n12351) );
  ANDN U15892 ( .B(n15276), .A(n15277), .Z(n15274) );
  NOR U15893 ( .A(n9219), .B(n9218), .Z(n15273) );
  XOR U15894 ( .A(n13530), .B(n10759), .Z(n9218) );
  XNOR U15895 ( .A(n15278), .B(n14208), .Z(n13530) );
  NOR U15896 ( .A(n14761), .B(n15279), .Z(n15278) );
  XNOR U15897 ( .A(n15280), .B(n12099), .Z(n9219) );
  XNOR U15898 ( .A(n15281), .B(n8120), .Z(n5104) );
  XOR U15899 ( .A(n9620), .B(n15282), .Z(n8120) );
  XOR U15900 ( .A(n12849), .B(n13050), .Z(n9620) );
  XNOR U15901 ( .A(n15283), .B(n15284), .Z(n13050) );
  XNOR U15902 ( .A(n12608), .B(n12792), .Z(n15284) );
  XNOR U15903 ( .A(n15285), .B(n12806), .Z(n12792) );
  XOR U15904 ( .A(n15286), .B(n15265), .Z(n12806) );
  NOR U15905 ( .A(n15287), .B(n12805), .Z(n15285) );
  XNOR U15906 ( .A(n15288), .B(n13359), .Z(n12608) );
  XOR U15907 ( .A(n15289), .B(n15290), .Z(n13359) );
  ANDN U15908 ( .B(n15291), .A(n13371), .Z(n15288) );
  IV U15909 ( .A(n15292), .Z(n13371) );
  XOR U15910 ( .A(n12577), .B(n15293), .Z(n15283) );
  XOR U15911 ( .A(n12106), .B(n11324), .Z(n15293) );
  XNOR U15912 ( .A(n15294), .B(n12955), .Z(n11324) );
  XOR U15913 ( .A(n15295), .B(n15296), .Z(n12955) );
  ANDN U15914 ( .B(n12954), .A(n15297), .Z(n15294) );
  XNOR U15915 ( .A(n15298), .B(n12800), .Z(n12106) );
  XOR U15916 ( .A(n15299), .B(n15300), .Z(n12800) );
  XNOR U15917 ( .A(n15302), .B(n12810), .Z(n12577) );
  XOR U15918 ( .A(n15303), .B(n15304), .Z(n12810) );
  AND U15919 ( .A(n15305), .B(n12809), .Z(n15302) );
  XOR U15920 ( .A(n15306), .B(n15307), .Z(n12849) );
  XNOR U15921 ( .A(n10696), .B(n12063), .Z(n15307) );
  XNOR U15922 ( .A(n15308), .B(n15309), .Z(n12063) );
  XNOR U15923 ( .A(n15312), .B(n15313), .Z(n10696) );
  ANDN U15924 ( .B(n15314), .A(n15315), .Z(n15312) );
  XOR U15925 ( .A(n12203), .B(n15316), .Z(n15306) );
  XNOR U15926 ( .A(n9513), .B(n9415), .Z(n15316) );
  XNOR U15927 ( .A(n15317), .B(n15318), .Z(n9415) );
  NOR U15928 ( .A(n15319), .B(n15320), .Z(n15317) );
  XNOR U15929 ( .A(n15321), .B(n15322), .Z(n9513) );
  ANDN U15930 ( .B(n15323), .A(n15324), .Z(n15321) );
  XNOR U15931 ( .A(n15325), .B(n15326), .Z(n12203) );
  ANDN U15932 ( .B(n15327), .A(n15328), .Z(n15325) );
  AND U15933 ( .A(n9216), .B(n9215), .Z(n15281) );
  XNOR U15934 ( .A(n9138), .B(n15329), .Z(n9215) );
  XNOR U15935 ( .A(n15330), .B(n13762), .Z(n9138) );
  XOR U15936 ( .A(n15331), .B(n15332), .Z(n13762) );
  XNOR U15937 ( .A(n12745), .B(n11095), .Z(n15332) );
  XNOR U15938 ( .A(n15333), .B(n14173), .Z(n11095) );
  IV U15939 ( .A(n15334), .Z(n14173) );
  ANDN U15940 ( .B(n14145), .A(n13258), .Z(n15333) );
  XOR U15941 ( .A(n15335), .B(n15336), .Z(n13258) );
  XNOR U15942 ( .A(n15337), .B(n14164), .Z(n12745) );
  ANDN U15943 ( .B(n14149), .A(n13266), .Z(n15337) );
  XOR U15944 ( .A(n15338), .B(n15339), .Z(n13266) );
  XOR U15945 ( .A(n9754), .B(n15340), .Z(n15331) );
  XNOR U15946 ( .A(n10223), .B(n14981), .Z(n15340) );
  XOR U15947 ( .A(n15341), .B(n14169), .Z(n14981) );
  NOR U15948 ( .A(n14140), .B(n13253), .Z(n15341) );
  XOR U15949 ( .A(n15342), .B(n15343), .Z(n13253) );
  XNOR U15950 ( .A(n15344), .B(n14160), .Z(n10223) );
  IV U15951 ( .A(n15345), .Z(n14160) );
  ANDN U15952 ( .B(n13262), .A(n14147), .Z(n15344) );
  XNOR U15953 ( .A(n15346), .B(n15347), .Z(n13262) );
  XNOR U15954 ( .A(n15348), .B(n15349), .Z(n9754) );
  ANDN U15955 ( .B(n13249), .A(n14142), .Z(n15348) );
  XOR U15956 ( .A(n15350), .B(n15351), .Z(n13249) );
  XOR U15957 ( .A(n15352), .B(n11062), .Z(n9216) );
  XNOR U15958 ( .A(n13020), .B(n14832), .Z(n11062) );
  XNOR U15959 ( .A(n15353), .B(n15354), .Z(n14832) );
  XNOR U15960 ( .A(n9633), .B(n14448), .Z(n15354) );
  XNOR U15961 ( .A(n15355), .B(n15356), .Z(n14448) );
  ANDN U15962 ( .B(n14435), .A(n15357), .Z(n15355) );
  XNOR U15963 ( .A(n15358), .B(n15359), .Z(n9633) );
  ANDN U15964 ( .B(n15360), .A(n14428), .Z(n15358) );
  XNOR U15965 ( .A(n9440), .B(n15361), .Z(n15353) );
  XOR U15966 ( .A(n10942), .B(n10272), .Z(n15361) );
  XOR U15967 ( .A(n15362), .B(n15363), .Z(n10272) );
  ANDN U15968 ( .B(n15364), .A(n14432), .Z(n15362) );
  AND U15969 ( .A(n15367), .B(n14423), .Z(n15365) );
  XNOR U15970 ( .A(n15368), .B(n15369), .Z(n9440) );
  ANDN U15971 ( .B(n14419), .A(n15370), .Z(n15368) );
  XOR U15972 ( .A(n15371), .B(n15372), .Z(n13020) );
  XOR U15973 ( .A(n12675), .B(n11451), .Z(n15372) );
  XOR U15974 ( .A(n15373), .B(n14458), .Z(n11451) );
  ANDN U15975 ( .B(n15374), .A(n14459), .Z(n15373) );
  XNOR U15976 ( .A(n15375), .B(n14464), .Z(n12675) );
  ANDN U15977 ( .B(n15376), .A(n14463), .Z(n15375) );
  XOR U15978 ( .A(n12227), .B(n15377), .Z(n15371) );
  XOR U15979 ( .A(n11368), .B(n14189), .Z(n15377) );
  XNOR U15980 ( .A(n15378), .B(n14455), .Z(n14189) );
  ANDN U15981 ( .B(n14454), .A(n15379), .Z(n15378) );
  XNOR U15982 ( .A(n15380), .B(n14468), .Z(n11368) );
  ANDN U15983 ( .B(n15381), .A(n14467), .Z(n15380) );
  XOR U15984 ( .A(n15382), .B(n14471), .Z(n12227) );
  NOR U15985 ( .A(n15383), .B(n15384), .Z(n15382) );
  XOR U15986 ( .A(n3750), .B(n15385), .Z(n15271) );
  XNOR U15987 ( .A(n9288), .B(n4211), .Z(n15385) );
  XNOR U15988 ( .A(n15386), .B(n7995), .Z(n4211) );
  XOR U15989 ( .A(n10359), .B(n15387), .Z(n7995) );
  NOR U15990 ( .A(n10046), .B(n9295), .Z(n15386) );
  XOR U15991 ( .A(n15388), .B(n12734), .Z(n9295) );
  XOR U15992 ( .A(n15389), .B(n13296), .Z(n12734) );
  XOR U15993 ( .A(n15390), .B(n15391), .Z(n13296) );
  XNOR U15994 ( .A(n12847), .B(n12463), .Z(n15391) );
  XOR U15995 ( .A(n15392), .B(n13839), .Z(n12463) );
  ANDN U15996 ( .B(n15393), .A(n15394), .Z(n15392) );
  XNOR U15997 ( .A(n15395), .B(n15396), .Z(n12847) );
  ANDN U15998 ( .B(n15397), .A(n15398), .Z(n15395) );
  XNOR U15999 ( .A(n11359), .B(n15399), .Z(n15390) );
  XNOR U16000 ( .A(n12894), .B(n12519), .Z(n15399) );
  XNOR U16001 ( .A(n15400), .B(n13829), .Z(n12519) );
  ANDN U16002 ( .B(n15401), .A(n15402), .Z(n15400) );
  XOR U16003 ( .A(n15403), .B(n15404), .Z(n12894) );
  ANDN U16004 ( .B(n15405), .A(n15406), .Z(n15403) );
  XOR U16005 ( .A(n15407), .B(n14587), .Z(n11359) );
  NOR U16006 ( .A(n15408), .B(n15409), .Z(n15407) );
  XNOR U16007 ( .A(n9539), .B(n15410), .Z(n10046) );
  XNOR U16008 ( .A(n15045), .B(n12721), .Z(n9539) );
  XOR U16009 ( .A(n15411), .B(n15412), .Z(n12721) );
  XNOR U16010 ( .A(n14976), .B(n14590), .Z(n15412) );
  XOR U16011 ( .A(n15413), .B(n15384), .Z(n14590) );
  ANDN U16012 ( .B(n15414), .A(n14470), .Z(n15413) );
  XOR U16013 ( .A(n15415), .B(n15379), .Z(n14976) );
  ANDN U16014 ( .B(n15416), .A(n14453), .Z(n15415) );
  XOR U16015 ( .A(n11102), .B(n15417), .Z(n15411) );
  XOR U16016 ( .A(n15418), .B(n12057), .Z(n15417) );
  XNOR U16017 ( .A(n15419), .B(n15381), .Z(n12057) );
  ANDN U16018 ( .B(n15420), .A(n14466), .Z(n15419) );
  IV U16019 ( .A(n15421), .Z(n14466) );
  XNOR U16020 ( .A(n15422), .B(n15376), .Z(n11102) );
  NOR U16021 ( .A(n14462), .B(n15423), .Z(n15422) );
  IV U16022 ( .A(n15424), .Z(n14462) );
  XOR U16023 ( .A(n15425), .B(n15426), .Z(n15045) );
  XOR U16024 ( .A(n12368), .B(n10395), .Z(n15426) );
  XNOR U16025 ( .A(n15427), .B(n15428), .Z(n10395) );
  ANDN U16026 ( .B(n15048), .A(n15429), .Z(n15427) );
  XNOR U16027 ( .A(n15430), .B(n13033), .Z(n12368) );
  NOR U16028 ( .A(n15431), .B(n13897), .Z(n15430) );
  XNOR U16029 ( .A(n11316), .B(n15432), .Z(n15425) );
  XNOR U16030 ( .A(n14714), .B(n11971), .Z(n15432) );
  XOR U16031 ( .A(n15433), .B(n13029), .Z(n11971) );
  XOR U16032 ( .A(n15434), .B(n13037), .Z(n14714) );
  AND U16033 ( .A(n13906), .B(n13905), .Z(n15434) );
  XNOR U16034 ( .A(n15435), .B(n15436), .Z(n11316) );
  ANDN U16035 ( .B(n15437), .A(n15438), .Z(n15435) );
  XOR U16036 ( .A(n15439), .B(n7990), .Z(n9288) );
  XNOR U16037 ( .A(n15440), .B(n12255), .Z(n7990) );
  IV U16038 ( .A(n14929), .Z(n12255) );
  XOR U16039 ( .A(n15441), .B(n15442), .Z(n14929) );
  ANDN U16040 ( .B(n9208), .A(n9209), .Z(n15439) );
  XNOR U16041 ( .A(n14492), .B(n13477), .Z(n9209) );
  XNOR U16042 ( .A(n11914), .B(n14518), .Z(n13477) );
  XOR U16043 ( .A(n15443), .B(n15444), .Z(n14518) );
  XNOR U16044 ( .A(n12098), .B(n15445), .Z(n15444) );
  XNOR U16045 ( .A(n15446), .B(n14254), .Z(n12098) );
  XNOR U16046 ( .A(n13733), .B(n15449), .Z(n15443) );
  XOR U16047 ( .A(n13916), .B(n15280), .Z(n15449) );
  NOR U16048 ( .A(n15451), .B(n13743), .Z(n15450) );
  XNOR U16049 ( .A(n15452), .B(n14250), .Z(n13916) );
  NOR U16050 ( .A(n15453), .B(n13752), .Z(n15452) );
  XNOR U16051 ( .A(n15454), .B(n14239), .Z(n13733) );
  ANDN U16052 ( .B(n13748), .A(n15455), .Z(n15454) );
  XOR U16053 ( .A(n15456), .B(n15457), .Z(n11914) );
  XOR U16054 ( .A(n15458), .B(n9646), .Z(n15457) );
  XOR U16055 ( .A(n15459), .B(n13722), .Z(n9646) );
  ANDN U16056 ( .B(n15460), .A(n15461), .Z(n15459) );
  XNOR U16057 ( .A(n12690), .B(n15462), .Z(n15456) );
  XNOR U16058 ( .A(n12237), .B(n11080), .Z(n15462) );
  XNOR U16059 ( .A(n15463), .B(n13710), .Z(n11080) );
  ANDN U16060 ( .B(n14502), .A(n14501), .Z(n15463) );
  IV U16061 ( .A(n15464), .Z(n14501) );
  XOR U16062 ( .A(n15465), .B(n13718), .Z(n12237) );
  ANDN U16063 ( .B(n14499), .A(n14498), .Z(n15465) );
  IV U16064 ( .A(n15466), .Z(n14498) );
  XNOR U16065 ( .A(n15467), .B(n13737), .Z(n12690) );
  ANDN U16066 ( .B(n14505), .A(n14504), .Z(n15467) );
  XNOR U16067 ( .A(n15468), .B(n15461), .Z(n14492) );
  ANDN U16068 ( .B(n13721), .A(n15460), .Z(n15468) );
  XOR U16069 ( .A(n10947), .B(n14619), .Z(n9208) );
  XNOR U16070 ( .A(n15469), .B(n15470), .Z(n14619) );
  NOR U16071 ( .A(n15471), .B(n15167), .Z(n15469) );
  XOR U16072 ( .A(n12204), .B(n14325), .Z(n10947) );
  XNOR U16073 ( .A(n15472), .B(n15473), .Z(n14325) );
  XNOR U16074 ( .A(n15474), .B(n12394), .Z(n15473) );
  XOR U16075 ( .A(n15475), .B(n15476), .Z(n12394) );
  XOR U16076 ( .A(n11068), .B(n15477), .Z(n15472) );
  XOR U16077 ( .A(n11621), .B(n15478), .Z(n15477) );
  XNOR U16078 ( .A(n15479), .B(n15173), .Z(n11621) );
  NOR U16079 ( .A(n14634), .B(n14635), .Z(n15479) );
  XOR U16080 ( .A(n15480), .B(n15179), .Z(n11068) );
  AND U16081 ( .A(n14621), .B(n14623), .Z(n15480) );
  XOR U16082 ( .A(n15481), .B(n15482), .Z(n12204) );
  XOR U16083 ( .A(n12367), .B(n10327), .Z(n15482) );
  XOR U16084 ( .A(n15483), .B(n15484), .Z(n10327) );
  ANDN U16085 ( .B(n15324), .A(n15322), .Z(n15483) );
  IV U16086 ( .A(n15485), .Z(n15322) );
  XOR U16087 ( .A(n15486), .B(n15487), .Z(n12367) );
  ANDN U16088 ( .B(n15328), .A(n15326), .Z(n15486) );
  XOR U16089 ( .A(n11547), .B(n15488), .Z(n15481) );
  XNOR U16090 ( .A(n13129), .B(n9911), .Z(n15488) );
  XOR U16091 ( .A(n15489), .B(n15490), .Z(n9911) );
  ANDN U16092 ( .B(n15320), .A(n15318), .Z(n15489) );
  XOR U16093 ( .A(n15491), .B(n15492), .Z(n13129) );
  NOR U16094 ( .A(n15310), .B(n15309), .Z(n15491) );
  XNOR U16095 ( .A(n15493), .B(n15494), .Z(n11547) );
  NOR U16096 ( .A(n15314), .B(n15313), .Z(n15493) );
  XNOR U16097 ( .A(n15495), .B(n7981), .Z(n3750) );
  XOR U16098 ( .A(n13934), .B(n10695), .Z(n7981) );
  XNOR U16099 ( .A(n15496), .B(n15497), .Z(n13934) );
  ANDN U16100 ( .B(n15498), .A(n15499), .Z(n15496) );
  ANDN U16101 ( .B(n9212), .A(n9213), .Z(n15495) );
  XOR U16102 ( .A(n15500), .B(n10305), .Z(n9213) );
  IV U16103 ( .A(n10860), .Z(n10305) );
  XOR U16104 ( .A(n12589), .B(n13822), .Z(n10860) );
  XNOR U16105 ( .A(n15501), .B(n15502), .Z(n13822) );
  XOR U16106 ( .A(n13132), .B(n12735), .Z(n15502) );
  XOR U16107 ( .A(n15503), .B(n15504), .Z(n12735) );
  AND U16108 ( .A(n15505), .B(n15506), .Z(n15503) );
  XNOR U16109 ( .A(n15507), .B(n15508), .Z(n13132) );
  NOR U16110 ( .A(n15509), .B(n15510), .Z(n15507) );
  XNOR U16111 ( .A(n11502), .B(n15511), .Z(n15501) );
  XNOR U16112 ( .A(n13206), .B(n12777), .Z(n15511) );
  XNOR U16113 ( .A(n15512), .B(n15513), .Z(n12777) );
  XOR U16114 ( .A(n15516), .B(n15517), .Z(n13206) );
  NOR U16115 ( .A(n15518), .B(n15519), .Z(n15516) );
  XOR U16116 ( .A(n15520), .B(n15521), .Z(n11502) );
  NOR U16117 ( .A(n15522), .B(n15523), .Z(n15520) );
  XOR U16118 ( .A(n15524), .B(n15525), .Z(n12589) );
  XOR U16119 ( .A(n10188), .B(n9880), .Z(n15525) );
  XOR U16120 ( .A(n15526), .B(n14669), .Z(n9880) );
  IV U16121 ( .A(n13240), .Z(n14669) );
  XOR U16122 ( .A(n15527), .B(n15528), .Z(n13240) );
  NOR U16123 ( .A(n13239), .B(n15529), .Z(n15526) );
  XNOR U16124 ( .A(n15530), .B(n13223), .Z(n10188) );
  XOR U16125 ( .A(n15531), .B(n15532), .Z(n13223) );
  NOR U16126 ( .A(n13222), .B(n15533), .Z(n15530) );
  XOR U16127 ( .A(n11037), .B(n15534), .Z(n15524) );
  XOR U16128 ( .A(n9457), .B(n11912), .Z(n15534) );
  XNOR U16129 ( .A(n15535), .B(n13227), .Z(n11912) );
  XOR U16130 ( .A(n15536), .B(n15537), .Z(n13227) );
  NOR U16131 ( .A(n13226), .B(n15538), .Z(n15535) );
  XNOR U16132 ( .A(n15539), .B(n13219), .Z(n9457) );
  XNOR U16133 ( .A(n15540), .B(n15541), .Z(n13219) );
  ANDN U16134 ( .B(n15542), .A(n13218), .Z(n15539) );
  XNOR U16135 ( .A(n15543), .B(n13213), .Z(n11037) );
  IV U16136 ( .A(n14666), .Z(n13213) );
  XOR U16137 ( .A(n15544), .B(n15545), .Z(n14666) );
  ANDN U16138 ( .B(n13214), .A(n15546), .Z(n15543) );
  XNOR U16139 ( .A(n15547), .B(n10287), .Z(n9212) );
  XOR U16140 ( .A(n11570), .B(n12993), .Z(n10287) );
  XNOR U16141 ( .A(n15548), .B(n15549), .Z(n12993) );
  XOR U16142 ( .A(n10381), .B(n14980), .Z(n15549) );
  XNOR U16143 ( .A(n15550), .B(n14537), .Z(n14980) );
  NOR U16144 ( .A(n15551), .B(n15552), .Z(n15550) );
  XNOR U16145 ( .A(n15553), .B(n14523), .Z(n10381) );
  ANDN U16146 ( .B(n15554), .A(n15555), .Z(n15553) );
  XNOR U16147 ( .A(n12693), .B(n15556), .Z(n15548) );
  XNOR U16148 ( .A(n10865), .B(n15058), .Z(n15556) );
  XNOR U16149 ( .A(n15557), .B(n14527), .Z(n15058) );
  ANDN U16150 ( .B(n15558), .A(n15559), .Z(n15557) );
  XNOR U16151 ( .A(n15560), .B(n14534), .Z(n10865) );
  IV U16152 ( .A(n15561), .Z(n14534) );
  ANDN U16153 ( .B(n15562), .A(n15563), .Z(n15560) );
  XNOR U16154 ( .A(n15564), .B(n15565), .Z(n12693) );
  ANDN U16155 ( .B(n15566), .A(n15567), .Z(n15564) );
  XOR U16156 ( .A(n15568), .B(n15569), .Z(n11570) );
  XNOR U16157 ( .A(n13632), .B(n11500), .Z(n15569) );
  XNOR U16158 ( .A(n15570), .B(n15571), .Z(n11500) );
  XNOR U16159 ( .A(n15574), .B(n15575), .Z(n13632) );
  XOR U16160 ( .A(n11813), .B(n15578), .Z(n15568) );
  XOR U16161 ( .A(n12600), .B(n10969), .Z(n15578) );
  XOR U16162 ( .A(n15579), .B(n15064), .Z(n10969) );
  ANDN U16163 ( .B(n15580), .A(n15065), .Z(n15579) );
  XNOR U16164 ( .A(n15581), .B(n15069), .Z(n12600) );
  NOR U16165 ( .A(n15582), .B(n15068), .Z(n15581) );
  XNOR U16166 ( .A(n15583), .B(n15076), .Z(n11813) );
  AND U16167 ( .A(n15584), .B(n15075), .Z(n15583) );
  XNOR U16168 ( .A(n15585), .B(n15205), .Z(n9192) );
  IV U16169 ( .A(n8067), .Z(n15205) );
  XOR U16170 ( .A(n15586), .B(n11568), .Z(n8067) );
  ANDN U16171 ( .B(n9177), .A(n14480), .Z(n15585) );
  XNOR U16172 ( .A(n15587), .B(n9757), .Z(n14480) );
  XNOR U16173 ( .A(n15445), .B(n12099), .Z(n9177) );
  XNOR U16174 ( .A(n15588), .B(n15589), .Z(n12099) );
  XOR U16175 ( .A(n15590), .B(n14247), .Z(n15445) );
  NOR U16176 ( .A(n15591), .B(n13756), .Z(n15590) );
  NOR U16177 ( .A(n5711), .B(n5709), .Z(n15052) );
  XOR U16178 ( .A(n9026), .B(n5192), .Z(n5709) );
  XOR U16179 ( .A(n6356), .B(n6556), .Z(n5192) );
  XNOR U16180 ( .A(n15592), .B(n15593), .Z(n6556) );
  XOR U16181 ( .A(n6369), .B(n2546), .Z(n15593) );
  XOR U16182 ( .A(n15594), .B(n6587), .Z(n2546) );
  XOR U16183 ( .A(n15595), .B(n9274), .Z(n6587) );
  XOR U16184 ( .A(n13484), .B(n11579), .Z(n9274) );
  XOR U16185 ( .A(n15596), .B(n15597), .Z(n11579) );
  XOR U16186 ( .A(n13307), .B(n12667), .Z(n15597) );
  XNOR U16187 ( .A(n15598), .B(n15599), .Z(n12667) );
  NOR U16188 ( .A(n15600), .B(n15601), .Z(n15598) );
  XNOR U16189 ( .A(n15602), .B(n15603), .Z(n13307) );
  NOR U16190 ( .A(n15604), .B(n15605), .Z(n15602) );
  XNOR U16191 ( .A(n12686), .B(n15606), .Z(n15596) );
  XOR U16192 ( .A(n10957), .B(n12080), .Z(n15606) );
  XOR U16193 ( .A(n15607), .B(n15608), .Z(n12080) );
  ANDN U16194 ( .B(n14813), .A(n15609), .Z(n15607) );
  XNOR U16195 ( .A(n15610), .B(n15611), .Z(n10957) );
  ANDN U16196 ( .B(n15612), .A(n14817), .Z(n15610) );
  XNOR U16197 ( .A(n15613), .B(n15614), .Z(n12686) );
  ANDN U16198 ( .B(n14824), .A(n15615), .Z(n15613) );
  XOR U16199 ( .A(n15616), .B(n15617), .Z(n13484) );
  XNOR U16200 ( .A(n9270), .B(n11927), .Z(n15617) );
  XNOR U16201 ( .A(n15618), .B(n14300), .Z(n11927) );
  ANDN U16202 ( .B(n14299), .A(n13888), .Z(n15618) );
  XOR U16203 ( .A(n15619), .B(n15620), .Z(n9270) );
  ANDN U16204 ( .B(n13881), .A(n15621), .Z(n15619) );
  XOR U16205 ( .A(n11605), .B(n15622), .Z(n15616) );
  XOR U16206 ( .A(n9278), .B(n12604), .Z(n15622) );
  XNOR U16207 ( .A(n15623), .B(n13321), .Z(n12604) );
  NOR U16208 ( .A(n15624), .B(n13320), .Z(n15623) );
  XOR U16209 ( .A(n15625), .B(n13316), .Z(n9278) );
  AND U16210 ( .A(n13317), .B(n13876), .Z(n15625) );
  XNOR U16211 ( .A(n15626), .B(n13324), .Z(n11605) );
  ANDN U16212 ( .B(n13873), .A(n13325), .Z(n15626) );
  NOR U16213 ( .A(n9032), .B(n9031), .Z(n15594) );
  XNOR U16214 ( .A(n11904), .B(n15627), .Z(n9031) );
  XNOR U16215 ( .A(n15628), .B(n11704), .Z(n9032) );
  XNOR U16216 ( .A(n15629), .B(n13893), .Z(n11704) );
  XNOR U16217 ( .A(n15630), .B(n15631), .Z(n13893) );
  XNOR U16218 ( .A(n10483), .B(n11048), .Z(n15631) );
  XNOR U16219 ( .A(n15632), .B(n15420), .Z(n11048) );
  ANDN U16220 ( .B(n14468), .A(n15421), .Z(n15632) );
  XOR U16221 ( .A(n15633), .B(n15541), .Z(n15421) );
  XOR U16222 ( .A(n15634), .B(n15635), .Z(n14468) );
  XNOR U16223 ( .A(n15636), .B(n15423), .Z(n10483) );
  ANDN U16224 ( .B(n14464), .A(n15424), .Z(n15636) );
  XOR U16225 ( .A(n15637), .B(n15638), .Z(n15424) );
  XNOR U16226 ( .A(n15639), .B(n15640), .Z(n14464) );
  XNOR U16227 ( .A(n15410), .B(n15641), .Z(n15630) );
  XNOR U16228 ( .A(n9540), .B(n9775), .Z(n15641) );
  XNOR U16229 ( .A(n15642), .B(n15414), .Z(n9775) );
  ANDN U16230 ( .B(n14470), .A(n14471), .Z(n15642) );
  XNOR U16231 ( .A(n15643), .B(n15644), .Z(n14471) );
  XOR U16232 ( .A(n15645), .B(n15646), .Z(n14470) );
  XOR U16233 ( .A(n15647), .B(n15648), .Z(n9540) );
  ANDN U16234 ( .B(n14457), .A(n14458), .Z(n15647) );
  XNOR U16235 ( .A(n15649), .B(n15650), .Z(n14458) );
  XNOR U16236 ( .A(n15651), .B(n15416), .Z(n15410) );
  AND U16237 ( .A(n14453), .B(n14455), .Z(n15651) );
  XNOR U16238 ( .A(n15652), .B(n15653), .Z(n14455) );
  XOR U16239 ( .A(n15654), .B(n15655), .Z(n14453) );
  XNOR U16240 ( .A(n15656), .B(n6592), .Z(n6369) );
  XNOR U16241 ( .A(n14305), .B(n10482), .Z(n6592) );
  XNOR U16242 ( .A(n12886), .B(n11859), .Z(n10482) );
  XNOR U16243 ( .A(n15657), .B(n15658), .Z(n11859) );
  XOR U16244 ( .A(n15180), .B(n11044), .Z(n15658) );
  XOR U16245 ( .A(n15659), .B(n15660), .Z(n11044) );
  ANDN U16246 ( .B(n15661), .A(n14308), .Z(n15659) );
  XOR U16247 ( .A(n15662), .B(n15663), .Z(n14308) );
  XNOR U16248 ( .A(n15664), .B(n15665), .Z(n15180) );
  XNOR U16249 ( .A(n14129), .B(n15667), .Z(n15657) );
  XOR U16250 ( .A(n13965), .B(n11876), .Z(n15667) );
  XNOR U16251 ( .A(n15668), .B(n15669), .Z(n11876) );
  NOR U16252 ( .A(n14313), .B(n14312), .Z(n15668) );
  XNOR U16253 ( .A(n15670), .B(n15671), .Z(n14313) );
  XNOR U16254 ( .A(n15672), .B(n15673), .Z(n13965) );
  NOR U16255 ( .A(n14316), .B(n14318), .Z(n15672) );
  XNOR U16256 ( .A(n15674), .B(n15675), .Z(n14318) );
  XOR U16257 ( .A(n15676), .B(n15677), .Z(n14129) );
  ANDN U16258 ( .B(n14322), .A(n14320), .Z(n15676) );
  XOR U16259 ( .A(n15678), .B(n15679), .Z(n14322) );
  XOR U16260 ( .A(n15680), .B(n15681), .Z(n12886) );
  XOR U16261 ( .A(n12925), .B(n11608), .Z(n15681) );
  XOR U16262 ( .A(n15682), .B(n14830), .Z(n11608) );
  XOR U16263 ( .A(n15645), .B(n15683), .Z(n14830) );
  NOR U16264 ( .A(n15684), .B(n15685), .Z(n15682) );
  XOR U16265 ( .A(n15686), .B(n12823), .Z(n12925) );
  XNOR U16266 ( .A(n15687), .B(n15688), .Z(n12823) );
  XOR U16267 ( .A(n12914), .B(n15689), .Z(n15680) );
  XOR U16268 ( .A(n11094), .B(n10645), .Z(n15689) );
  XOR U16269 ( .A(n15690), .B(n12834), .Z(n10645) );
  XOR U16270 ( .A(n15691), .B(n15692), .Z(n12834) );
  NOR U16271 ( .A(n14941), .B(n15202), .Z(n15690) );
  XNOR U16272 ( .A(n15693), .B(n12828), .Z(n11094) );
  XOR U16273 ( .A(n15694), .B(n15695), .Z(n12828) );
  ANDN U16274 ( .B(n15198), .A(n14947), .Z(n15693) );
  XOR U16275 ( .A(n15697), .B(n15698), .Z(n14973) );
  AND U16276 ( .A(n14937), .B(n15194), .Z(n15696) );
  XOR U16277 ( .A(n15699), .B(n15666), .Z(n14305) );
  NOR U16278 ( .A(n15700), .B(n14864), .Z(n15699) );
  XNOR U16279 ( .A(n15701), .B(n15702), .Z(n14864) );
  ANDN U16280 ( .B(n9075), .A(n14933), .Z(n15656) );
  XOR U16281 ( .A(n3518), .B(n15703), .Z(n15592) );
  XNOR U16282 ( .A(n9068), .B(n4896), .Z(n15703) );
  XNOR U16283 ( .A(n15704), .B(n6604), .Z(n4896) );
  XOR U16284 ( .A(n15705), .B(n10062), .Z(n6604) );
  IV U16285 ( .A(n9418), .Z(n10062) );
  XNOR U16286 ( .A(n15706), .B(n13245), .Z(n9418) );
  XOR U16287 ( .A(n15707), .B(n15708), .Z(n13245) );
  XOR U16288 ( .A(n12491), .B(n11749), .Z(n15708) );
  XNOR U16289 ( .A(n15709), .B(n15710), .Z(n11749) );
  XNOR U16290 ( .A(n15713), .B(n15714), .Z(n12491) );
  NOR U16291 ( .A(n15715), .B(n15716), .Z(n15713) );
  XOR U16292 ( .A(n9612), .B(n15717), .Z(n15707) );
  XOR U16293 ( .A(n10115), .B(n14135), .Z(n15717) );
  XNOR U16294 ( .A(n15718), .B(n15719), .Z(n14135) );
  ANDN U16295 ( .B(n15720), .A(n15721), .Z(n15718) );
  XNOR U16296 ( .A(n15722), .B(n15723), .Z(n10115) );
  ANDN U16297 ( .B(n15724), .A(n15725), .Z(n15722) );
  XNOR U16298 ( .A(n15726), .B(n15727), .Z(n9612) );
  ANDN U16299 ( .B(n15728), .A(n15729), .Z(n15726) );
  ANDN U16300 ( .B(n9029), .A(n9028), .Z(n15704) );
  XNOR U16301 ( .A(n15731), .B(n14904), .Z(n11568) );
  XOR U16302 ( .A(n15732), .B(n15733), .Z(n14904) );
  XNOR U16303 ( .A(n9901), .B(n10490), .Z(n15733) );
  XOR U16304 ( .A(n15734), .B(n14742), .Z(n10490) );
  ANDN U16305 ( .B(n14108), .A(n15735), .Z(n15734) );
  XNOR U16306 ( .A(n14754), .B(n15736), .Z(n9901) );
  XNOR U16307 ( .A(n4687), .B(n15737), .Z(n15736) );
  NANDN U16308 ( .A(n14753), .B(n15738), .Z(n15737) );
  XOR U16309 ( .A(n14487), .B(n15739), .Z(n15732) );
  XNOR U16310 ( .A(n9616), .B(n14734), .Z(n15739) );
  XNOR U16311 ( .A(n15740), .B(n14740), .Z(n14734) );
  NOR U16312 ( .A(n14100), .B(n14739), .Z(n15740) );
  XOR U16313 ( .A(n15741), .B(n14750), .Z(n9616) );
  NOR U16314 ( .A(n15742), .B(n14749), .Z(n15741) );
  XNOR U16315 ( .A(n15743), .B(n14746), .Z(n14487) );
  ANDN U16316 ( .B(n14104), .A(n15744), .Z(n15743) );
  XOR U16317 ( .A(n10878), .B(n15745), .Z(n9029) );
  XOR U16318 ( .A(n15746), .B(n6601), .Z(n9068) );
  XOR U16319 ( .A(n11111), .B(n14055), .Z(n6601) );
  XNOR U16320 ( .A(n15747), .B(n15748), .Z(n14055) );
  NOR U16321 ( .A(n15214), .B(n15749), .Z(n15747) );
  XOR U16322 ( .A(n13095), .B(n14365), .Z(n11111) );
  XNOR U16323 ( .A(n15750), .B(n15751), .Z(n14365) );
  XOR U16324 ( .A(n15752), .B(n15753), .Z(n15751) );
  XOR U16325 ( .A(n12058), .B(n15754), .Z(n15750) );
  XNOR U16326 ( .A(n11753), .B(n12050), .Z(n15754) );
  XOR U16327 ( .A(n15755), .B(n15219), .Z(n12050) );
  NOR U16328 ( .A(n14062), .B(n14063), .Z(n15755) );
  XNOR U16329 ( .A(n15756), .B(n15224), .Z(n11753) );
  ANDN U16330 ( .B(n15757), .A(n14052), .Z(n15756) );
  XOR U16331 ( .A(n15758), .B(n15211), .Z(n12058) );
  ANDN U16332 ( .B(n14058), .A(n15759), .Z(n15758) );
  XOR U16333 ( .A(n15760), .B(n15761), .Z(n13095) );
  XOR U16334 ( .A(n15762), .B(n10944), .Z(n15761) );
  XNOR U16335 ( .A(n15763), .B(n15233), .Z(n10944) );
  XOR U16336 ( .A(n10495), .B(n15764), .Z(n15760) );
  XOR U16337 ( .A(n11332), .B(n14900), .Z(n15764) );
  XNOR U16338 ( .A(n15765), .B(n15240), .Z(n14900) );
  NOR U16339 ( .A(n14083), .B(n14081), .Z(n15765) );
  XNOR U16340 ( .A(n15766), .B(n15243), .Z(n11332) );
  ANDN U16341 ( .B(n14068), .A(n14069), .Z(n15766) );
  XNOR U16342 ( .A(n15767), .B(n15768), .Z(n10495) );
  ANDN U16343 ( .B(n14072), .A(n14073), .Z(n15767) );
  ANDN U16344 ( .B(n9023), .A(n9024), .Z(n15746) );
  XOR U16345 ( .A(n15769), .B(n11364), .Z(n9024) );
  XOR U16346 ( .A(n9530), .B(n14376), .Z(n9023) );
  XNOR U16347 ( .A(n15770), .B(n15771), .Z(n14376) );
  ANDN U16348 ( .B(n13100), .A(n15772), .Z(n15770) );
  XNOR U16349 ( .A(n15773), .B(n14852), .Z(n9530) );
  XOR U16350 ( .A(n15774), .B(n15775), .Z(n14852) );
  XOR U16351 ( .A(n14301), .B(n10963), .Z(n15775) );
  XOR U16352 ( .A(n15776), .B(n12431), .Z(n10963) );
  ANDN U16353 ( .B(n15777), .A(n15778), .Z(n15776) );
  XOR U16354 ( .A(n15779), .B(n15780), .Z(n14301) );
  NOR U16355 ( .A(n15781), .B(n15782), .Z(n15779) );
  XOR U16356 ( .A(n13469), .B(n15783), .Z(n15774) );
  XNOR U16357 ( .A(n13380), .B(n11053), .Z(n15783) );
  XOR U16358 ( .A(n15784), .B(n12348), .Z(n11053) );
  ANDN U16359 ( .B(n15785), .A(n15786), .Z(n15784) );
  XNOR U16360 ( .A(n15787), .B(n15276), .Z(n13380) );
  ANDN U16361 ( .B(n15788), .A(n15789), .Z(n15787) );
  XNOR U16362 ( .A(n15790), .B(n12356), .Z(n13469) );
  IV U16363 ( .A(n15791), .Z(n12356) );
  ANDN U16364 ( .B(n15792), .A(n15793), .Z(n15790) );
  XNOR U16365 ( .A(n15794), .B(n6596), .Z(n3518) );
  XNOR U16366 ( .A(n15795), .B(n9891), .Z(n6596) );
  XNOR U16367 ( .A(n13374), .B(n13847), .Z(n9891) );
  XNOR U16368 ( .A(n15796), .B(n15797), .Z(n13847) );
  XNOR U16369 ( .A(n14261), .B(n10228), .Z(n15797) );
  XNOR U16370 ( .A(n15798), .B(n15799), .Z(n10228) );
  ANDN U16371 ( .B(n15800), .A(n15801), .Z(n15798) );
  XNOR U16372 ( .A(n15802), .B(n13941), .Z(n14261) );
  NOR U16373 ( .A(n15803), .B(n15804), .Z(n15802) );
  XOR U16374 ( .A(n10349), .B(n15805), .Z(n15796) );
  XOR U16375 ( .A(n9519), .B(n12999), .Z(n15805) );
  XOR U16376 ( .A(n15806), .B(n15499), .Z(n12999) );
  AND U16377 ( .A(n15807), .B(n15808), .Z(n15806) );
  XOR U16378 ( .A(n15809), .B(n15810), .Z(n9519) );
  XNOR U16379 ( .A(n15813), .B(n13937), .Z(n10349) );
  ANDN U16380 ( .B(n15814), .A(n15815), .Z(n15813) );
  XOR U16381 ( .A(n15816), .B(n15817), .Z(n13374) );
  XOR U16382 ( .A(n9969), .B(n11839), .Z(n15817) );
  XOR U16383 ( .A(n15818), .B(n15819), .Z(n11839) );
  NOR U16384 ( .A(n15820), .B(n15821), .Z(n15818) );
  XNOR U16385 ( .A(n15822), .B(n15823), .Z(n9969) );
  ANDN U16386 ( .B(n15824), .A(n14908), .Z(n15822) );
  XNOR U16387 ( .A(n9756), .B(n15825), .Z(n15816) );
  XOR U16388 ( .A(n15826), .B(n15587), .Z(n15825) );
  XOR U16389 ( .A(n15827), .B(n15828), .Z(n15587) );
  ANDN U16390 ( .B(n15829), .A(n15830), .Z(n15827) );
  XOR U16391 ( .A(n15831), .B(n15832), .Z(n9756) );
  NOR U16392 ( .A(n14912), .B(n15833), .Z(n15831) );
  NOR U16393 ( .A(n9021), .B(n9020), .Z(n15794) );
  XOR U16394 ( .A(n15089), .B(n11778), .Z(n9020) );
  IV U16395 ( .A(n9946), .Z(n11778) );
  XNOR U16396 ( .A(n13287), .B(n15834), .Z(n9946) );
  XOR U16397 ( .A(n15835), .B(n15836), .Z(n13287) );
  XOR U16398 ( .A(n13795), .B(n12975), .Z(n15836) );
  XNOR U16399 ( .A(n15837), .B(n15838), .Z(n12975) );
  AND U16400 ( .A(n13999), .B(n13997), .Z(n15837) );
  XNOR U16401 ( .A(n15839), .B(n15840), .Z(n13795) );
  ANDN U16402 ( .B(n13986), .A(n13984), .Z(n15839) );
  XNOR U16403 ( .A(n12102), .B(n15841), .Z(n15835) );
  XNOR U16404 ( .A(n12723), .B(n11629), .Z(n15841) );
  XNOR U16405 ( .A(n15842), .B(n15843), .Z(n11629) );
  ANDN U16406 ( .B(n13995), .A(n13993), .Z(n15842) );
  IV U16407 ( .A(n15844), .Z(n13993) );
  XNOR U16408 ( .A(n15845), .B(n15846), .Z(n12723) );
  ANDN U16409 ( .B(n13982), .A(n15847), .Z(n15845) );
  XNOR U16410 ( .A(n15848), .B(n15849), .Z(n12102) );
  NOR U16411 ( .A(n13990), .B(n13989), .Z(n15848) );
  XNOR U16412 ( .A(n15850), .B(n15851), .Z(n15089) );
  ANDN U16413 ( .B(n13398), .A(n15852), .Z(n15850) );
  XOR U16414 ( .A(n10278), .B(n15853), .Z(n9021) );
  XNOR U16415 ( .A(n15854), .B(n15855), .Z(n6356) );
  XNOR U16416 ( .A(n3735), .B(n5484), .Z(n15855) );
  XOR U16417 ( .A(n15856), .B(n9083), .Z(n5484) );
  XOR U16418 ( .A(n14822), .B(n11508), .Z(n9083) );
  IV U16419 ( .A(n9118), .Z(n11508) );
  XOR U16420 ( .A(n15857), .B(n15605), .Z(n14822) );
  ANDN U16421 ( .B(n15858), .A(n15859), .Z(n15857) );
  ANDN U16422 ( .B(n6625), .A(n9129), .Z(n15856) );
  IV U16423 ( .A(n6626), .Z(n9129) );
  XOR U16424 ( .A(n10278), .B(n15860), .Z(n6626) );
  IV U16425 ( .A(n12424), .Z(n10278) );
  XNOR U16426 ( .A(n15861), .B(n15862), .Z(n12424) );
  XOR U16427 ( .A(n11228), .B(n13023), .Z(n6625) );
  XNOR U16428 ( .A(n15863), .B(n15050), .Z(n13023) );
  ANDN U16429 ( .B(n15428), .A(n15864), .Z(n15863) );
  XNOR U16430 ( .A(n15865), .B(n7092), .Z(n3735) );
  XOR U16431 ( .A(n9780), .B(n13406), .Z(n7092) );
  XNOR U16432 ( .A(n15866), .B(n15084), .Z(n13406) );
  NOR U16433 ( .A(n15867), .B(n15868), .Z(n15866) );
  IV U16434 ( .A(n12947), .Z(n9780) );
  XNOR U16435 ( .A(n10536), .B(n14926), .Z(n12947) );
  XOR U16436 ( .A(n15869), .B(n15870), .Z(n14926) );
  XOR U16437 ( .A(n13278), .B(n12781), .Z(n15870) );
  XOR U16438 ( .A(n15871), .B(n15092), .Z(n12781) );
  ANDN U16439 ( .B(n13412), .A(n13413), .Z(n15871) );
  XNOR U16440 ( .A(n15872), .B(n15873), .Z(n13412) );
  XOR U16441 ( .A(n15874), .B(n15087), .Z(n13278) );
  AND U16442 ( .A(n13404), .B(n13402), .Z(n15874) );
  XNOR U16443 ( .A(n15875), .B(n15876), .Z(n13402) );
  XOR U16444 ( .A(n11939), .B(n15877), .Z(n15869) );
  XNOR U16445 ( .A(n12602), .B(n11481), .Z(n15877) );
  XOR U16446 ( .A(n15878), .B(n15083), .Z(n11481) );
  XOR U16447 ( .A(n15879), .B(n15880), .Z(n15084) );
  XOR U16448 ( .A(n15881), .B(n15852), .Z(n12602) );
  ANDN U16449 ( .B(n13400), .A(n13398), .Z(n15881) );
  XOR U16450 ( .A(n15882), .B(n15883), .Z(n13398) );
  XOR U16451 ( .A(n15884), .B(n15095), .Z(n11939) );
  ANDN U16452 ( .B(n13408), .A(n13409), .Z(n15884) );
  XNOR U16453 ( .A(n15885), .B(n15886), .Z(n13408) );
  XOR U16454 ( .A(n15887), .B(n15888), .Z(n10536) );
  XNOR U16455 ( .A(n10648), .B(n11289), .Z(n15888) );
  XOR U16456 ( .A(n15889), .B(n13990), .Z(n11289) );
  XOR U16457 ( .A(n15890), .B(n15891), .Z(n13990) );
  ANDN U16458 ( .B(n13991), .A(n15892), .Z(n15889) );
  XNOR U16459 ( .A(n15893), .B(n13999), .Z(n10648) );
  XOR U16460 ( .A(n15894), .B(n15638), .Z(n13999) );
  ANDN U16461 ( .B(n15895), .A(n13998), .Z(n15893) );
  XNOR U16462 ( .A(n10315), .B(n15896), .Z(n15887) );
  XOR U16463 ( .A(n13976), .B(n11812), .Z(n15896) );
  XNOR U16464 ( .A(n15897), .B(n13982), .Z(n11812) );
  XOR U16465 ( .A(n15898), .B(n15899), .Z(n13982) );
  ANDN U16466 ( .B(n15900), .A(n15901), .Z(n15897) );
  XNOR U16467 ( .A(n15902), .B(n13995), .Z(n13976) );
  XOR U16468 ( .A(n15903), .B(n15904), .Z(n13995) );
  ANDN U16469 ( .B(n13994), .A(n15905), .Z(n15902) );
  XNOR U16470 ( .A(n15906), .B(n13986), .Z(n10315) );
  XOR U16471 ( .A(n15879), .B(n15907), .Z(n13986) );
  NOR U16472 ( .A(n13985), .B(n15908), .Z(n15906) );
  ANDN U16473 ( .B(n6618), .A(n6616), .Z(n15865) );
  XOR U16474 ( .A(n15909), .B(n11972), .Z(n6616) );
  XNOR U16475 ( .A(n11897), .B(n15910), .Z(n11972) );
  XOR U16476 ( .A(n15911), .B(n15912), .Z(n11897) );
  XOR U16477 ( .A(n10723), .B(n12767), .Z(n15912) );
  XOR U16478 ( .A(n15913), .B(n15914), .Z(n12767) );
  ANDN U16479 ( .B(n15915), .A(n15916), .Z(n15913) );
  XNOR U16480 ( .A(n15917), .B(n15918), .Z(n10723) );
  ANDN U16481 ( .B(n15919), .A(n15920), .Z(n15917) );
  XOR U16482 ( .A(n11596), .B(n15921), .Z(n15911) );
  XNOR U16483 ( .A(n12271), .B(n12263), .Z(n15921) );
  XNOR U16484 ( .A(n15922), .B(n15923), .Z(n12263) );
  AND U16485 ( .A(n15924), .B(n15925), .Z(n15922) );
  XOR U16486 ( .A(n15926), .B(n15927), .Z(n12271) );
  ANDN U16487 ( .B(n15928), .A(n15929), .Z(n15926) );
  XNOR U16488 ( .A(n15930), .B(n15931), .Z(n11596) );
  ANDN U16489 ( .B(n15932), .A(n15933), .Z(n15930) );
  XOR U16490 ( .A(n11904), .B(n15934), .Z(n6618) );
  XNOR U16491 ( .A(n12885), .B(n13805), .Z(n11904) );
  XNOR U16492 ( .A(n15935), .B(n15936), .Z(n13805) );
  XNOR U16493 ( .A(n15937), .B(n12380), .Z(n15936) );
  XOR U16494 ( .A(n15938), .B(n13190), .Z(n12380) );
  ANDN U16495 ( .B(n13804), .A(n13803), .Z(n15938) );
  XNOR U16496 ( .A(n10832), .B(n15939), .Z(n15935) );
  XOR U16497 ( .A(n13596), .B(n12193), .Z(n15939) );
  NOR U16498 ( .A(n13668), .B(n13669), .Z(n15940) );
  XNOR U16499 ( .A(n15941), .B(n13194), .Z(n13596) );
  NOR U16500 ( .A(n13660), .B(n13661), .Z(n15941) );
  XNOR U16501 ( .A(n15942), .B(n15943), .Z(n10832) );
  NOR U16502 ( .A(n13789), .B(n13791), .Z(n15942) );
  XOR U16503 ( .A(n15944), .B(n15945), .Z(n12885) );
  XNOR U16504 ( .A(n11581), .B(n9936), .Z(n15945) );
  XNOR U16505 ( .A(n15946), .B(n13274), .Z(n9936) );
  IV U16506 ( .A(n12946), .Z(n13274) );
  XOR U16507 ( .A(n15947), .B(n15948), .Z(n12946) );
  NOR U16508 ( .A(n12945), .B(n14965), .Z(n15946) );
  XNOR U16509 ( .A(n12932), .B(n15949), .Z(n11581) );
  XNOR U16510 ( .A(n11417), .B(n15950), .Z(n15949) );
  NANDN U16511 ( .A(n14969), .B(n12933), .Z(n15950) );
  XOR U16512 ( .A(n15951), .B(n15952), .Z(n12932) );
  XNOR U16513 ( .A(n11853), .B(n15953), .Z(n15944) );
  XNOR U16514 ( .A(n12242), .B(n9465), .Z(n15953) );
  XOR U16515 ( .A(n15954), .B(n12938), .Z(n9465) );
  NOR U16516 ( .A(n12937), .B(n14961), .Z(n15954) );
  XNOR U16517 ( .A(n15957), .B(n13168), .Z(n12242) );
  XNOR U16518 ( .A(n15958), .B(n15959), .Z(n13168) );
  NOR U16519 ( .A(n13167), .B(n14951), .Z(n15957) );
  XOR U16520 ( .A(n15960), .B(n12942), .Z(n11853) );
  XNOR U16521 ( .A(n15961), .B(n15962), .Z(n12942) );
  NOR U16522 ( .A(n14955), .B(n12941), .Z(n15960) );
  XOR U16523 ( .A(n4344), .B(n15963), .Z(n15854) );
  XOR U16524 ( .A(n5936), .B(n2135), .Z(n15963) );
  XNOR U16525 ( .A(n15964), .B(n7084), .Z(n2135) );
  XNOR U16526 ( .A(n12856), .B(n9224), .Z(n7084) );
  XOR U16527 ( .A(n13731), .B(n15965), .Z(n9224) );
  XOR U16528 ( .A(n15966), .B(n15967), .Z(n13731) );
  XNOR U16529 ( .A(n12513), .B(n13134), .Z(n15967) );
  XOR U16530 ( .A(n15968), .B(n15969), .Z(n13134) );
  AND U16531 ( .A(n15970), .B(n15971), .Z(n15968) );
  XNOR U16532 ( .A(n15972), .B(n15973), .Z(n12513) );
  NOR U16533 ( .A(n15974), .B(n15975), .Z(n15972) );
  XNOR U16534 ( .A(n11446), .B(n15976), .Z(n15966) );
  XNOR U16535 ( .A(n11119), .B(n11844), .Z(n15976) );
  XNOR U16536 ( .A(n15977), .B(n15978), .Z(n11844) );
  XNOR U16537 ( .A(n15981), .B(n15982), .Z(n11119) );
  NOR U16538 ( .A(n15983), .B(n15984), .Z(n15981) );
  XOR U16539 ( .A(n15985), .B(n15986), .Z(n11446) );
  NOR U16540 ( .A(n15987), .B(n15988), .Z(n15985) );
  XNOR U16541 ( .A(n15989), .B(n15990), .Z(n12856) );
  ANDN U16542 ( .B(n15991), .A(n15992), .Z(n15989) );
  ANDN U16543 ( .B(n6623), .A(n6621), .Z(n15964) );
  XNOR U16544 ( .A(n14575), .B(n9856), .Z(n6621) );
  XNOR U16545 ( .A(n12440), .B(n12879), .Z(n9856) );
  XNOR U16546 ( .A(n15993), .B(n15994), .Z(n12879) );
  XNOR U16547 ( .A(n9766), .B(n15001), .Z(n15994) );
  XOR U16548 ( .A(n15995), .B(n13772), .Z(n15001) );
  ANDN U16549 ( .B(n14986), .A(n15996), .Z(n15995) );
  XOR U16550 ( .A(n15997), .B(n13784), .Z(n9766) );
  ANDN U16551 ( .B(n14570), .A(n15998), .Z(n15997) );
  XNOR U16552 ( .A(n15999), .B(n16000), .Z(n14570) );
  XNOR U16553 ( .A(n10478), .B(n16001), .Z(n15993) );
  XOR U16554 ( .A(n10394), .B(n16002), .Z(n16001) );
  XOR U16555 ( .A(n16003), .B(n13776), .Z(n10394) );
  ANDN U16556 ( .B(n14578), .A(n14577), .Z(n16003) );
  XOR U16557 ( .A(n16004), .B(n16005), .Z(n14578) );
  XOR U16558 ( .A(n16006), .B(n13768), .Z(n10478) );
  ANDN U16559 ( .B(n14581), .A(n14580), .Z(n16006) );
  XOR U16560 ( .A(n16007), .B(n16008), .Z(n14581) );
  XOR U16561 ( .A(n16009), .B(n16010), .Z(n12440) );
  XNOR U16562 ( .A(n16011), .B(n12659), .Z(n16010) );
  XNOR U16563 ( .A(n16012), .B(n16013), .Z(n12659) );
  XOR U16564 ( .A(n12219), .B(n16014), .Z(n16009) );
  XOR U16565 ( .A(n16015), .B(n12950), .Z(n16014) );
  XOR U16566 ( .A(n16016), .B(n16017), .Z(n12950) );
  ANDN U16567 ( .B(n14563), .A(n14564), .Z(n16016) );
  ANDN U16568 ( .B(n14561), .A(n14559), .Z(n16018) );
  XOR U16569 ( .A(n16020), .B(n15996), .Z(n14575) );
  IV U16570 ( .A(n16021), .Z(n15996) );
  ANDN U16571 ( .B(n13770), .A(n14986), .Z(n16020) );
  XNOR U16572 ( .A(n16022), .B(n16023), .Z(n14986) );
  XNOR U16573 ( .A(n16024), .B(n16025), .Z(n13770) );
  XNOR U16574 ( .A(n16026), .B(n10980), .Z(n6623) );
  XNOR U16575 ( .A(n16027), .B(n14364), .Z(n10980) );
  XOR U16576 ( .A(n16028), .B(n16029), .Z(n14364) );
  XNOR U16577 ( .A(n12631), .B(n10401), .Z(n16029) );
  ANDN U16578 ( .B(n16033), .A(n16034), .Z(n16030) );
  XOR U16579 ( .A(n16035), .B(n14035), .Z(n12631) );
  XNOR U16580 ( .A(n16036), .B(n16037), .Z(n14035) );
  ANDN U16581 ( .B(n16038), .A(n14036), .Z(n16035) );
  XOR U16582 ( .A(n12291), .B(n16039), .Z(n16028) );
  XOR U16583 ( .A(n12281), .B(n10591), .Z(n16039) );
  XNOR U16584 ( .A(n16040), .B(n16041), .Z(n10591) );
  AND U16585 ( .A(n14029), .B(n16042), .Z(n16040) );
  XNOR U16586 ( .A(n16043), .B(n13429), .Z(n12281) );
  IV U16587 ( .A(n14042), .Z(n13429) );
  XOR U16588 ( .A(n16044), .B(n15545), .Z(n14042) );
  IV U16589 ( .A(n16045), .Z(n15545) );
  NOR U16590 ( .A(n14041), .B(n16046), .Z(n16043) );
  XNOR U16591 ( .A(n16047), .B(n13438), .Z(n12291) );
  IV U16592 ( .A(n14038), .Z(n13438) );
  XOR U16593 ( .A(n16048), .B(n16049), .Z(n14038) );
  ANDN U16594 ( .B(n14039), .A(n16050), .Z(n16047) );
  XNOR U16595 ( .A(n16051), .B(n7089), .Z(n5936) );
  XNOR U16596 ( .A(n15418), .B(n11103), .Z(n7089) );
  IV U16597 ( .A(n14977), .Z(n11103) );
  XOR U16598 ( .A(n13512), .B(n14732), .Z(n14977) );
  XOR U16599 ( .A(n16052), .B(n16053), .Z(n14732) );
  XOR U16600 ( .A(n9644), .B(n11159), .Z(n16053) );
  XOR U16601 ( .A(n16054), .B(n13036), .Z(n11159) );
  XOR U16602 ( .A(n16055), .B(n16056), .Z(n13905) );
  XNOR U16603 ( .A(n16057), .B(n16058), .Z(n13037) );
  XNOR U16604 ( .A(n16059), .B(n13032), .Z(n9644) );
  AND U16605 ( .A(n13033), .B(n13897), .Z(n16059) );
  XOR U16606 ( .A(n16060), .B(n16061), .Z(n13897) );
  XOR U16607 ( .A(n16062), .B(n16063), .Z(n13033) );
  XNOR U16608 ( .A(n9876), .B(n16064), .Z(n16052) );
  XOR U16609 ( .A(n11826), .B(n10308), .Z(n16064) );
  XNOR U16610 ( .A(n16065), .B(n16066), .Z(n10308) );
  NOR U16611 ( .A(n15048), .B(n15428), .Z(n16065) );
  XNOR U16612 ( .A(n16067), .B(n16068), .Z(n15428) );
  XNOR U16613 ( .A(n16069), .B(n14958), .Z(n15048) );
  XNOR U16614 ( .A(n16070), .B(n13028), .Z(n11826) );
  NOR U16615 ( .A(n13900), .B(n13029), .Z(n16070) );
  XOR U16616 ( .A(n16071), .B(n16072), .Z(n13029) );
  XOR U16617 ( .A(n16073), .B(n16074), .Z(n13900) );
  XOR U16618 ( .A(n16075), .B(n16076), .Z(n9876) );
  NOR U16619 ( .A(n15437), .B(n15436), .Z(n16075) );
  IV U16620 ( .A(n13908), .Z(n15437) );
  XOR U16621 ( .A(n16077), .B(n16078), .Z(n13908) );
  XOR U16622 ( .A(n16079), .B(n16080), .Z(n13512) );
  XNOR U16623 ( .A(n12742), .B(n12995), .Z(n16080) );
  XNOR U16624 ( .A(n16081), .B(n14459), .Z(n12995) );
  XOR U16625 ( .A(n16082), .B(n16083), .Z(n14459) );
  NOR U16626 ( .A(n15648), .B(n15374), .Z(n16081) );
  XOR U16627 ( .A(n16084), .B(n14463), .Z(n12742) );
  XOR U16628 ( .A(n16085), .B(n16086), .Z(n14463) );
  ANDN U16629 ( .B(n15423), .A(n15376), .Z(n16084) );
  XOR U16630 ( .A(n16087), .B(n16088), .Z(n15376) );
  XNOR U16631 ( .A(n16089), .B(n16090), .Z(n15423) );
  XOR U16632 ( .A(n11751), .B(n16091), .Z(n16079) );
  XOR U16633 ( .A(n10841), .B(n13019), .Z(n16091) );
  XNOR U16634 ( .A(n16092), .B(n14454), .Z(n13019) );
  XOR U16635 ( .A(n16093), .B(n16094), .Z(n14454) );
  ANDN U16636 ( .B(n15379), .A(n15416), .Z(n16092) );
  XOR U16637 ( .A(n16095), .B(n16096), .Z(n15416) );
  XNOR U16638 ( .A(n16097), .B(n16098), .Z(n15379) );
  XOR U16639 ( .A(n16099), .B(n14467), .Z(n10841) );
  XOR U16640 ( .A(n16100), .B(n16101), .Z(n14467) );
  NOR U16641 ( .A(n15381), .B(n15420), .Z(n16099) );
  XOR U16642 ( .A(n16102), .B(n16103), .Z(n15420) );
  XNOR U16643 ( .A(n16104), .B(n16105), .Z(n15381) );
  XNOR U16644 ( .A(n16106), .B(n15383), .Z(n11751) );
  IV U16645 ( .A(n14472), .Z(n15383) );
  XOR U16646 ( .A(n16107), .B(n16108), .Z(n14472) );
  ANDN U16647 ( .B(n15384), .A(n15414), .Z(n16106) );
  XNOR U16648 ( .A(n16109), .B(n16110), .Z(n15414) );
  XNOR U16649 ( .A(n16111), .B(n16112), .Z(n15384) );
  XNOR U16650 ( .A(n16113), .B(n15374), .Z(n15418) );
  XNOR U16651 ( .A(n16114), .B(n16115), .Z(n15374) );
  ANDN U16652 ( .B(n15648), .A(n14457), .Z(n16113) );
  XNOR U16653 ( .A(n16116), .B(n16117), .Z(n14457) );
  XOR U16654 ( .A(n16118), .B(n16119), .Z(n15648) );
  AND U16655 ( .A(n6614), .B(n6612), .Z(n16051) );
  XNOR U16656 ( .A(n16120), .B(n9864), .Z(n6612) );
  XOR U16657 ( .A(n12266), .B(n13295), .Z(n9864) );
  XNOR U16658 ( .A(n16121), .B(n16122), .Z(n13295) );
  XOR U16659 ( .A(n13792), .B(n11492), .Z(n16122) );
  XNOR U16660 ( .A(n16123), .B(n16124), .Z(n11492) );
  ANDN U16661 ( .B(n16125), .A(n16126), .Z(n16123) );
  XNOR U16662 ( .A(n16127), .B(n12462), .Z(n13792) );
  ANDN U16663 ( .B(n16128), .A(n16129), .Z(n16127) );
  XOR U16664 ( .A(n9259), .B(n16130), .Z(n16121) );
  XNOR U16665 ( .A(n10649), .B(n16131), .Z(n16130) );
  XOR U16666 ( .A(n16132), .B(n16133), .Z(n10649) );
  XNOR U16667 ( .A(n16136), .B(n13699), .Z(n9259) );
  XOR U16668 ( .A(n16139), .B(n16140), .Z(n12266) );
  XOR U16669 ( .A(n12320), .B(n13649), .Z(n16140) );
  XNOR U16670 ( .A(n16141), .B(n14556), .Z(n13649) );
  XNOR U16671 ( .A(n16143), .B(n14561), .Z(n12320) );
  XNOR U16672 ( .A(n16144), .B(n15541), .Z(n14561) );
  XOR U16673 ( .A(n11619), .B(n16146), .Z(n16139) );
  XOR U16674 ( .A(n10511), .B(n13202), .Z(n16146) );
  XNOR U16675 ( .A(n16147), .B(n14551), .Z(n13202) );
  XNOR U16676 ( .A(n16148), .B(n16149), .Z(n14551) );
  NOR U16677 ( .A(n16150), .B(n16151), .Z(n16147) );
  XNOR U16678 ( .A(n16152), .B(n14564), .Z(n10511) );
  XOR U16679 ( .A(n16153), .B(n16154), .Z(n14564) );
  ANDN U16680 ( .B(n16155), .A(n16156), .Z(n16152) );
  XNOR U16681 ( .A(n16157), .B(n14547), .Z(n11619) );
  ANDN U16682 ( .B(n14548), .A(n16158), .Z(n16157) );
  XOR U16683 ( .A(n9659), .B(n16159), .Z(n6614) );
  IV U16684 ( .A(n11558), .Z(n9659) );
  XNOR U16685 ( .A(n16160), .B(n11864), .Z(n11558) );
  XOR U16686 ( .A(n16161), .B(n16162), .Z(n11864) );
  XOR U16687 ( .A(n11335), .B(n12324), .Z(n16162) );
  XOR U16688 ( .A(n16163), .B(n13630), .Z(n12324) );
  NOR U16689 ( .A(n13626), .B(n16164), .Z(n16163) );
  IV U16690 ( .A(n16165), .Z(n13626) );
  XNOR U16691 ( .A(n16166), .B(n12568), .Z(n11335) );
  ANDN U16692 ( .B(n13622), .A(n16167), .Z(n16166) );
  XNOR U16693 ( .A(n11115), .B(n16168), .Z(n16161) );
  XNOR U16694 ( .A(n16169), .B(n11573), .Z(n16168) );
  XOR U16695 ( .A(n16170), .B(n12564), .Z(n11573) );
  AND U16696 ( .A(n13624), .B(n16171), .Z(n16170) );
  XNOR U16697 ( .A(n16172), .B(n13392), .Z(n11115) );
  ANDN U16698 ( .B(n13618), .A(n16173), .Z(n16172) );
  XNOR U16699 ( .A(n16174), .B(n7079), .Z(n4344) );
  XOR U16700 ( .A(n16175), .B(n10741), .Z(n7079) );
  ANDN U16701 ( .B(n6631), .A(n9086), .Z(n16174) );
  XOR U16702 ( .A(n16178), .B(n11364), .Z(n9086) );
  XNOR U16703 ( .A(n12769), .B(n16179), .Z(n11364) );
  XOR U16704 ( .A(n16180), .B(n16181), .Z(n12769) );
  XNOR U16705 ( .A(n12202), .B(n13093), .Z(n16181) );
  XOR U16706 ( .A(n16182), .B(n16183), .Z(n13093) );
  NOR U16707 ( .A(n16184), .B(n16185), .Z(n16182) );
  XNOR U16708 ( .A(n16186), .B(n16187), .Z(n12202) );
  ANDN U16709 ( .B(n16188), .A(n15026), .Z(n16186) );
  XNOR U16710 ( .A(n12138), .B(n16189), .Z(n16180) );
  XOR U16711 ( .A(n9112), .B(n14808), .Z(n16189) );
  XNOR U16712 ( .A(n16190), .B(n16191), .Z(n14808) );
  NOR U16713 ( .A(n16192), .B(n15012), .Z(n16190) );
  XNOR U16714 ( .A(n16193), .B(n16194), .Z(n9112) );
  ANDN U16715 ( .B(n16195), .A(n16196), .Z(n16193) );
  XNOR U16716 ( .A(n16197), .B(n16198), .Z(n12138) );
  ANDN U16717 ( .B(n16199), .A(n16200), .Z(n16197) );
  XOR U16718 ( .A(n16201), .B(n16202), .Z(n6631) );
  XNOR U16719 ( .A(n16203), .B(n9075), .Z(n9026) );
  XOR U16720 ( .A(n16204), .B(n12652), .Z(n9075) );
  ANDN U16721 ( .B(n14933), .A(n6590), .Z(n16203) );
  XOR U16722 ( .A(n14717), .B(n11648), .Z(n6590) );
  XNOR U16723 ( .A(n16205), .B(n11828), .Z(n11648) );
  XNOR U16724 ( .A(n16206), .B(n16207), .Z(n11828) );
  XOR U16725 ( .A(n12511), .B(n10598), .Z(n16207) );
  XNOR U16726 ( .A(n16208), .B(n16209), .Z(n10598) );
  ANDN U16727 ( .B(n16210), .A(n16211), .Z(n16208) );
  XNOR U16728 ( .A(n16212), .B(n16213), .Z(n12511) );
  AND U16729 ( .A(n14726), .B(n14728), .Z(n16212) );
  XOR U16730 ( .A(n11459), .B(n16214), .Z(n16206) );
  XNOR U16731 ( .A(n16215), .B(n12134), .Z(n16214) );
  XNOR U16732 ( .A(n16216), .B(n13498), .Z(n12134) );
  NOR U16733 ( .A(n16217), .B(n14731), .Z(n16216) );
  XNOR U16734 ( .A(n16218), .B(n13493), .Z(n11459) );
  ANDN U16735 ( .B(n14719), .A(n16219), .Z(n16218) );
  XOR U16736 ( .A(n16220), .B(n16211), .Z(n14717) );
  NOR U16737 ( .A(n13501), .B(n16210), .Z(n16220) );
  XNOR U16738 ( .A(n9639), .B(n16221), .Z(n14933) );
  IV U16739 ( .A(n10698), .Z(n9639) );
  XNOR U16740 ( .A(n16222), .B(n14113), .Z(n10698) );
  XOR U16741 ( .A(n16223), .B(n16224), .Z(n14113) );
  XNOR U16742 ( .A(n12918), .B(n12524), .Z(n16224) );
  XOR U16743 ( .A(n16225), .B(n16226), .Z(n12524) );
  NOR U16744 ( .A(n16227), .B(n16228), .Z(n16225) );
  XOR U16745 ( .A(n16229), .B(n16230), .Z(n12918) );
  NOR U16746 ( .A(n16231), .B(n16232), .Z(n16229) );
  XNOR U16747 ( .A(n11617), .B(n16233), .Z(n16223) );
  XOR U16748 ( .A(n12310), .B(n11339), .Z(n16233) );
  XOR U16749 ( .A(n16234), .B(n16235), .Z(n11339) );
  ANDN U16750 ( .B(n16236), .A(n16237), .Z(n16234) );
  XOR U16751 ( .A(n16238), .B(n16239), .Z(n12310) );
  NOR U16752 ( .A(n16240), .B(n16241), .Z(n16238) );
  XOR U16753 ( .A(n16242), .B(n16243), .Z(n11617) );
  NOR U16754 ( .A(n16244), .B(n16245), .Z(n16242) );
  XOR U16755 ( .A(n11998), .B(n2101), .Z(n5711) );
  XNOR U16756 ( .A(n8399), .B(n9916), .Z(n2101) );
  XNOR U16757 ( .A(n16246), .B(n16247), .Z(n9916) );
  XNOR U16758 ( .A(n5519), .B(n3648), .Z(n16247) );
  XOR U16759 ( .A(n16248), .B(n8524), .Z(n3648) );
  XNOR U16760 ( .A(n16249), .B(n12652), .Z(n8524) );
  IV U16761 ( .A(n13121), .Z(n12652) );
  XNOR U16762 ( .A(n16250), .B(n16251), .Z(n13121) );
  ANDN U16763 ( .B(n8577), .A(n8578), .Z(n16248) );
  XOR U16764 ( .A(n16252), .B(n11124), .Z(n8578) );
  XNOR U16765 ( .A(n16253), .B(n15629), .Z(n11124) );
  XOR U16766 ( .A(n16254), .B(n16255), .Z(n15629) );
  XNOR U16767 ( .A(n10739), .B(n12466), .Z(n16255) );
  XNOR U16768 ( .A(n16256), .B(n14433), .Z(n12466) );
  NOR U16769 ( .A(n14434), .B(n15363), .Z(n16256) );
  XNOR U16770 ( .A(n16257), .B(n14425), .Z(n10739) );
  ANDN U16771 ( .B(n14424), .A(n15366), .Z(n16257) );
  XNOR U16772 ( .A(n12719), .B(n16258), .Z(n16254) );
  XNOR U16773 ( .A(n12691), .B(n11773), .Z(n16258) );
  XNOR U16774 ( .A(n16259), .B(n14430), .Z(n11773) );
  ANDN U16775 ( .B(n15359), .A(n14429), .Z(n16259) );
  XOR U16776 ( .A(n16260), .B(n14420), .Z(n12691) );
  XOR U16777 ( .A(n16261), .B(n14438), .Z(n12719) );
  ANDN U16778 ( .B(n15356), .A(n14439), .Z(n16261) );
  XNOR U16779 ( .A(n16262), .B(n9524), .Z(n8577) );
  XOR U16780 ( .A(n16264), .B(n16265), .Z(n15078) );
  XOR U16781 ( .A(n16266), .B(n11870), .Z(n16265) );
  XOR U16782 ( .A(n16267), .B(n16244), .Z(n11870) );
  AND U16783 ( .A(n16268), .B(n16269), .Z(n16267) );
  XOR U16784 ( .A(n10076), .B(n16270), .Z(n16264) );
  XNOR U16785 ( .A(n12988), .B(n10601), .Z(n16270) );
  XOR U16786 ( .A(n16271), .B(n16240), .Z(n10601) );
  ANDN U16787 ( .B(n16272), .A(n16273), .Z(n16271) );
  XOR U16788 ( .A(n16274), .B(n16236), .Z(n12988) );
  ANDN U16789 ( .B(n16275), .A(n16276), .Z(n16274) );
  XNOR U16790 ( .A(n16277), .B(n16231), .Z(n10076) );
  ANDN U16791 ( .B(n16278), .A(n16279), .Z(n16277) );
  XOR U16792 ( .A(n16280), .B(n12155), .Z(n5519) );
  XOR U16793 ( .A(n16281), .B(n11356), .Z(n12155) );
  XNOR U16794 ( .A(n15862), .B(n16282), .Z(n11356) );
  XOR U16795 ( .A(n16283), .B(n16284), .Z(n15862) );
  XOR U16796 ( .A(n11899), .B(n12852), .Z(n16284) );
  XNOR U16797 ( .A(n16285), .B(n12866), .Z(n12852) );
  NOR U16798 ( .A(n12865), .B(n16286), .Z(n16285) );
  XOR U16799 ( .A(n16287), .B(n15991), .Z(n11899) );
  XNOR U16800 ( .A(n10608), .B(n16289), .Z(n16283) );
  XNOR U16801 ( .A(n12371), .B(n11744), .Z(n16289) );
  XNOR U16802 ( .A(n16290), .B(n14387), .Z(n11744) );
  ANDN U16803 ( .B(n16291), .A(n14386), .Z(n16290) );
  XOR U16804 ( .A(n16292), .B(n12860), .Z(n12371) );
  ANDN U16805 ( .B(n16293), .A(n12859), .Z(n16292) );
  XOR U16806 ( .A(n16294), .B(n12869), .Z(n10608) );
  ANDN U16807 ( .B(n16295), .A(n12870), .Z(n16294) );
  ANDN U16808 ( .B(n8573), .A(n8575), .Z(n16280) );
  XOR U16809 ( .A(n16296), .B(n11805), .Z(n8575) );
  IV U16810 ( .A(n10729), .Z(n11805) );
  XOR U16811 ( .A(n14234), .B(n14023), .Z(n10729) );
  XNOR U16812 ( .A(n16297), .B(n16298), .Z(n14023) );
  XOR U16813 ( .A(n10204), .B(n9904), .Z(n16298) );
  XOR U16814 ( .A(n16299), .B(n15075), .Z(n9904) );
  XNOR U16815 ( .A(n16300), .B(n16301), .Z(n15075) );
  ANDN U16816 ( .B(n16302), .A(n15584), .Z(n16299) );
  XNOR U16817 ( .A(n16303), .B(n15068), .Z(n10204) );
  XOR U16818 ( .A(n16304), .B(n16305), .Z(n15068) );
  ANDN U16819 ( .B(n15582), .A(n16306), .Z(n16303) );
  XOR U16820 ( .A(n11569), .B(n16307), .Z(n16297) );
  XNOR U16821 ( .A(n10756), .B(n11557), .Z(n16307) );
  XNOR U16822 ( .A(n16308), .B(n15576), .Z(n11557) );
  NOR U16823 ( .A(n15577), .B(n16309), .Z(n16308) );
  XNOR U16824 ( .A(n16310), .B(n15572), .Z(n10756) );
  ANDN U16825 ( .B(n16311), .A(n15573), .Z(n16310) );
  XNOR U16826 ( .A(n16312), .B(n15065), .Z(n11569) );
  XOR U16827 ( .A(n16313), .B(n16314), .Z(n15065) );
  NOR U16828 ( .A(n16315), .B(n15580), .Z(n16312) );
  XOR U16829 ( .A(n16316), .B(n16317), .Z(n14234) );
  XOR U16830 ( .A(n12228), .B(n15547), .Z(n16317) );
  XOR U16831 ( .A(n16318), .B(n15563), .Z(n15547) );
  ANDN U16832 ( .B(n14532), .A(n15562), .Z(n16318) );
  XNOR U16833 ( .A(n16319), .B(n16320), .Z(n12228) );
  NOR U16834 ( .A(n15558), .B(n14526), .Z(n16319) );
  XOR U16835 ( .A(n14539), .B(n16321), .Z(n16316) );
  XOR U16836 ( .A(n14756), .B(n10286), .Z(n16321) );
  ANDN U16837 ( .B(n14522), .A(n15554), .Z(n16322) );
  XNOR U16838 ( .A(n16323), .B(n16324), .Z(n14756) );
  ANDN U16839 ( .B(n16325), .A(n15566), .Z(n16323) );
  IV U16840 ( .A(n16326), .Z(n15566) );
  XOR U16841 ( .A(n16327), .B(n15552), .Z(n14539) );
  AND U16842 ( .A(n15551), .B(n14536), .Z(n16327) );
  XNOR U16843 ( .A(n15072), .B(n10388), .Z(n8573) );
  XNOR U16844 ( .A(n16328), .B(n16329), .Z(n15072) );
  NOR U16845 ( .A(n15576), .B(n15575), .Z(n16328) );
  XOR U16846 ( .A(n16330), .B(n16331), .Z(n15576) );
  XOR U16847 ( .A(n6316), .B(n16332), .Z(n16246) );
  XOR U16848 ( .A(n2402), .B(n5727), .Z(n16332) );
  XNOR U16849 ( .A(n16333), .B(n8509), .Z(n5727) );
  XOR U16850 ( .A(n10202), .B(n14798), .Z(n8509) );
  XNOR U16851 ( .A(n16334), .B(n16335), .Z(n14798) );
  ANDN U16852 ( .B(n16336), .A(n16337), .Z(n16334) );
  XNOR U16853 ( .A(n11322), .B(n11121), .Z(n10202) );
  XOR U16854 ( .A(n16338), .B(n16339), .Z(n11121) );
  XNOR U16855 ( .A(n11209), .B(n12176), .Z(n16339) );
  XNOR U16856 ( .A(n16340), .B(n16341), .Z(n12176) );
  ANDN U16857 ( .B(n12044), .A(n16342), .Z(n16340) );
  XOR U16858 ( .A(n16343), .B(n16344), .Z(n11209) );
  NOR U16859 ( .A(n16345), .B(n12035), .Z(n16343) );
  XNOR U16860 ( .A(n11740), .B(n16346), .Z(n16338) );
  XNOR U16861 ( .A(n16347), .B(n11436), .Z(n16346) );
  XNOR U16862 ( .A(n16348), .B(n16349), .Z(n11436) );
  XOR U16863 ( .A(n16350), .B(n16351), .Z(n11740) );
  NOR U16864 ( .A(n12031), .B(n12030), .Z(n16350) );
  XOR U16865 ( .A(n16352), .B(n16353), .Z(n11322) );
  XNOR U16866 ( .A(n12418), .B(n12838), .Z(n16353) );
  XNOR U16867 ( .A(n16354), .B(n16355), .Z(n12838) );
  XNOR U16868 ( .A(n16356), .B(n16357), .Z(n12418) );
  ANDN U16869 ( .B(n14803), .A(n14802), .Z(n16356) );
  IV U16870 ( .A(n16358), .Z(n14803) );
  XOR U16871 ( .A(n12684), .B(n16359), .Z(n16352) );
  XNOR U16872 ( .A(n16360), .B(n15044), .Z(n16359) );
  XNOR U16873 ( .A(n16361), .B(n16362), .Z(n15044) );
  ANDN U16874 ( .B(n14791), .A(n14792), .Z(n16361) );
  XOR U16875 ( .A(n16363), .B(n16364), .Z(n12684) );
  NOR U16876 ( .A(n14795), .B(n14796), .Z(n16363) );
  ANDN U16877 ( .B(n9919), .A(n12161), .Z(n16333) );
  XNOR U16878 ( .A(n16011), .B(n12220), .Z(n12161) );
  XNOR U16879 ( .A(n16365), .B(n16366), .Z(n16011) );
  NOR U16880 ( .A(n14547), .B(n14546), .Z(n16365) );
  XOR U16881 ( .A(n16367), .B(n16368), .Z(n14547) );
  IV U16882 ( .A(n12274), .Z(n9919) );
  XOR U16883 ( .A(n14820), .B(n9118), .Z(n12274) );
  XNOR U16884 ( .A(n16369), .B(n16370), .Z(n12963) );
  XOR U16885 ( .A(n9273), .B(n13592), .Z(n16370) );
  XNOR U16886 ( .A(n16371), .B(n15609), .Z(n13592) );
  IV U16887 ( .A(n16372), .Z(n15609) );
  NOR U16888 ( .A(n16373), .B(n14813), .Z(n16371) );
  XOR U16889 ( .A(n16374), .B(n16375), .Z(n14813) );
  XOR U16890 ( .A(n16376), .B(n15612), .Z(n9273) );
  ANDN U16891 ( .B(n14817), .A(n14818), .Z(n16376) );
  XOR U16892 ( .A(n14952), .B(n16377), .Z(n14817) );
  XOR U16893 ( .A(n15595), .B(n16378), .Z(n16369) );
  XOR U16894 ( .A(n12375), .B(n12267), .Z(n16378) );
  XOR U16895 ( .A(n16379), .B(n15615), .Z(n12267) );
  NOR U16896 ( .A(n14825), .B(n14824), .Z(n16379) );
  XNOR U16897 ( .A(n16380), .B(n16119), .Z(n14824) );
  XNOR U16898 ( .A(n16381), .B(n15604), .Z(n12375) );
  IV U16899 ( .A(n16382), .Z(n15604) );
  ANDN U16900 ( .B(n15605), .A(n15858), .Z(n16381) );
  XNOR U16901 ( .A(n16383), .B(n16301), .Z(n15605) );
  XNOR U16902 ( .A(n16384), .B(n16385), .Z(n15595) );
  ANDN U16903 ( .B(n15601), .A(n16386), .Z(n16384) );
  XOR U16904 ( .A(n16387), .B(n16388), .Z(n12068) );
  XOR U16905 ( .A(n12091), .B(n9551), .Z(n16388) );
  XOR U16906 ( .A(n16389), .B(n15621), .Z(n9551) );
  NOR U16907 ( .A(n13881), .B(n13883), .Z(n16389) );
  XNOR U16908 ( .A(n16390), .B(n16391), .Z(n13881) );
  XNOR U16909 ( .A(n16392), .B(n13320), .Z(n12091) );
  XOR U16910 ( .A(n16393), .B(n16032), .Z(n13320) );
  NOR U16911 ( .A(n13885), .B(n13886), .Z(n16392) );
  IV U16912 ( .A(n15624), .Z(n13885) );
  XOR U16913 ( .A(n15654), .B(n16394), .Z(n15624) );
  XNOR U16914 ( .A(n13483), .B(n16395), .Z(n16387) );
  XNOR U16915 ( .A(n13284), .B(n9665), .Z(n16395) );
  XNOR U16916 ( .A(n16396), .B(n13317), .Z(n9665) );
  XOR U16917 ( .A(n16397), .B(n16398), .Z(n13317) );
  NOR U16918 ( .A(n13876), .B(n13877), .Z(n16396) );
  XNOR U16919 ( .A(n16399), .B(n16400), .Z(n13876) );
  XOR U16920 ( .A(n16401), .B(n13325), .Z(n13284) );
  XOR U16921 ( .A(n16402), .B(n15537), .Z(n13325) );
  NOR U16922 ( .A(n13873), .B(n13874), .Z(n16401) );
  XOR U16923 ( .A(n16403), .B(n16404), .Z(n13873) );
  XNOR U16924 ( .A(n16405), .B(n14299), .Z(n13483) );
  XOR U16925 ( .A(n16406), .B(n16407), .Z(n14299) );
  AND U16926 ( .A(n13888), .B(n13890), .Z(n16405) );
  XOR U16927 ( .A(n16408), .B(n16409), .Z(n13888) );
  XOR U16928 ( .A(n16410), .B(n15601), .Z(n14820) );
  XOR U16929 ( .A(n16411), .B(n16412), .Z(n15601) );
  ANDN U16930 ( .B(n16413), .A(n16414), .Z(n16410) );
  XNOR U16931 ( .A(n16415), .B(n8514), .Z(n2402) );
  IV U16932 ( .A(n12157), .Z(n8514) );
  XOR U16933 ( .A(n10186), .B(n16416), .Z(n12157) );
  IV U16934 ( .A(n12182), .Z(n10186) );
  XNOR U16935 ( .A(n13866), .B(n12649), .Z(n12182) );
  XOR U16936 ( .A(n16417), .B(n16418), .Z(n12649) );
  XOR U16937 ( .A(n15853), .B(n10279), .Z(n16418) );
  XNOR U16938 ( .A(n16419), .B(n16420), .Z(n10279) );
  XOR U16939 ( .A(n16423), .B(n16424), .Z(n15853) );
  ANDN U16940 ( .B(n16425), .A(n16426), .Z(n16423) );
  XOR U16941 ( .A(n12425), .B(n16427), .Z(n16417) );
  XOR U16942 ( .A(n15860), .B(n13636), .Z(n16427) );
  XOR U16943 ( .A(n16428), .B(n16429), .Z(n13636) );
  NOR U16944 ( .A(n16430), .B(n16431), .Z(n16428) );
  XNOR U16945 ( .A(n16432), .B(n16433), .Z(n15860) );
  XNOR U16946 ( .A(n16436), .B(n16437), .Z(n12425) );
  ANDN U16947 ( .B(n16438), .A(n16439), .Z(n16436) );
  XOR U16948 ( .A(n16440), .B(n16441), .Z(n13866) );
  XOR U16949 ( .A(n11421), .B(n13300), .Z(n16441) );
  XOR U16950 ( .A(n16442), .B(n16443), .Z(n13300) );
  ANDN U16951 ( .B(n16444), .A(n16445), .Z(n16442) );
  XNOR U16952 ( .A(n16446), .B(n16447), .Z(n11421) );
  NOR U16953 ( .A(n16448), .B(n16449), .Z(n16446) );
  XOR U16954 ( .A(n10079), .B(n16450), .Z(n16440) );
  XOR U16955 ( .A(n16451), .B(n13914), .Z(n16450) );
  XOR U16956 ( .A(n16452), .B(n16453), .Z(n13914) );
  NOR U16957 ( .A(n16454), .B(n16455), .Z(n16452) );
  XOR U16958 ( .A(n16456), .B(n16457), .Z(n10079) );
  ANDN U16959 ( .B(n16458), .A(n16459), .Z(n16456) );
  ANDN U16960 ( .B(n8564), .A(n8565), .Z(n16415) );
  XNOR U16961 ( .A(n9438), .B(n16460), .Z(n8565) );
  XNOR U16962 ( .A(n15389), .B(n13703), .Z(n9438) );
  XOR U16963 ( .A(n16461), .B(n16462), .Z(n13703) );
  XOR U16964 ( .A(n14474), .B(n13012), .Z(n16462) );
  XOR U16965 ( .A(n16463), .B(n15538), .Z(n13012) );
  XOR U16966 ( .A(n16464), .B(n16465), .Z(n13225) );
  ANDN U16967 ( .B(n13217), .A(n14660), .Z(n16466) );
  XOR U16968 ( .A(n15885), .B(n16467), .Z(n13217) );
  XOR U16969 ( .A(n13068), .B(n16468), .Z(n16461) );
  XNOR U16970 ( .A(n16469), .B(n16470), .Z(n16468) );
  XNOR U16971 ( .A(n16471), .B(n15529), .Z(n13068) );
  NOR U16972 ( .A(n16472), .B(n13238), .Z(n16471) );
  XNOR U16973 ( .A(n16473), .B(n16301), .Z(n13238) );
  XOR U16974 ( .A(n16474), .B(n16475), .Z(n15389) );
  XNOR U16975 ( .A(n9782), .B(n16476), .Z(n16475) );
  XNOR U16976 ( .A(n16477), .B(n15522), .Z(n9782) );
  ANDN U16977 ( .B(n16478), .A(n16479), .Z(n16477) );
  XNOR U16978 ( .A(n10935), .B(n16480), .Z(n16474) );
  XOR U16979 ( .A(n16481), .B(n10959), .Z(n16480) );
  XNOR U16980 ( .A(n16482), .B(n15518), .Z(n10959) );
  IV U16981 ( .A(n16483), .Z(n15518) );
  AND U16982 ( .A(n16484), .B(n16485), .Z(n16482) );
  XOR U16983 ( .A(n16486), .B(n15506), .Z(n10935) );
  ANDN U16984 ( .B(n16487), .A(n16488), .Z(n16486) );
  XOR U16985 ( .A(n15478), .B(n12395), .Z(n8564) );
  XNOR U16986 ( .A(n16489), .B(n16490), .Z(n15478) );
  XNOR U16987 ( .A(n16491), .B(n8519), .Z(n6316) );
  XOR U16988 ( .A(n16492), .B(n16493), .Z(n8519) );
  ANDN U16989 ( .B(n8568), .A(n8567), .Z(n16491) );
  XOR U16990 ( .A(n11228), .B(n13024), .Z(n8567) );
  XNOR U16991 ( .A(n16494), .B(n13909), .Z(n13024) );
  ANDN U16992 ( .B(n15436), .A(n16076), .Z(n16494) );
  XOR U16993 ( .A(n16495), .B(n15650), .Z(n15436) );
  XNOR U16994 ( .A(n14190), .B(n16496), .Z(n11228) );
  XOR U16995 ( .A(n16497), .B(n16498), .Z(n14190) );
  XOR U16996 ( .A(n12911), .B(n13420), .Z(n16498) );
  XNOR U16997 ( .A(n16499), .B(n15431), .Z(n13420) );
  IV U16998 ( .A(n13898), .Z(n15431) );
  XOR U16999 ( .A(n16500), .B(n15541), .Z(n13898) );
  NOR U17000 ( .A(n13031), .B(n13032), .Z(n16499) );
  XOR U17001 ( .A(n16501), .B(n16502), .Z(n13032) );
  XNOR U17002 ( .A(n16503), .B(n16504), .Z(n13031) );
  XOR U17003 ( .A(n16505), .B(n13901), .Z(n12911) );
  XOR U17004 ( .A(n16506), .B(n16507), .Z(n13901) );
  NOR U17005 ( .A(n13028), .B(n13027), .Z(n16505) );
  XNOR U17006 ( .A(n16508), .B(n16509), .Z(n13027) );
  XOR U17007 ( .A(n16510), .B(n16511), .Z(n13028) );
  XOR U17008 ( .A(n11098), .B(n16512), .Z(n16497) );
  XOR U17009 ( .A(n11739), .B(n13486), .Z(n16512) );
  XNOR U17010 ( .A(n16513), .B(n15429), .Z(n13486) );
  IV U17011 ( .A(n15049), .Z(n15429) );
  XOR U17012 ( .A(n16514), .B(n16110), .Z(n15049) );
  ANDN U17013 ( .B(n15050), .A(n16066), .Z(n16513) );
  IV U17014 ( .A(n15864), .Z(n16066) );
  XOR U17015 ( .A(n16515), .B(n16516), .Z(n15864) );
  XNOR U17016 ( .A(n16517), .B(n14967), .Z(n15050) );
  XOR U17017 ( .A(n16518), .B(n13906), .Z(n11739) );
  XNOR U17018 ( .A(n16519), .B(n16520), .Z(n13906) );
  NOR U17019 ( .A(n13035), .B(n13036), .Z(n16518) );
  XOR U17020 ( .A(n16521), .B(n16522), .Z(n13036) );
  XOR U17021 ( .A(n16523), .B(n16524), .Z(n13035) );
  XNOR U17022 ( .A(n16525), .B(n13910), .Z(n11098) );
  IV U17023 ( .A(n15438), .Z(n13910) );
  XOR U17024 ( .A(n16526), .B(n15186), .Z(n15438) );
  IV U17025 ( .A(n16527), .Z(n15186) );
  ANDN U17026 ( .B(n16076), .A(n13909), .Z(n16525) );
  XNOR U17027 ( .A(n16528), .B(n16529), .Z(n13909) );
  XOR U17028 ( .A(n16530), .B(n16531), .Z(n16076) );
  XNOR U17029 ( .A(n16532), .B(n12117), .Z(n8568) );
  XNOR U17030 ( .A(n16176), .B(n16533), .Z(n12117) );
  XOR U17031 ( .A(n16534), .B(n16535), .Z(n16176) );
  XNOR U17032 ( .A(n9453), .B(n16536), .Z(n16535) );
  XNOR U17033 ( .A(n16537), .B(n14770), .Z(n9453) );
  ANDN U17034 ( .B(n16538), .A(n16539), .Z(n16537) );
  XNOR U17035 ( .A(n16540), .B(n16541), .Z(n16534) );
  XOR U17036 ( .A(n11291), .B(n14179), .Z(n16541) );
  XNOR U17037 ( .A(n16542), .B(n14787), .Z(n14179) );
  IV U17038 ( .A(n16543), .Z(n14787) );
  ANDN U17039 ( .B(n16544), .A(n16545), .Z(n16542) );
  XNOR U17040 ( .A(n16546), .B(n16547), .Z(n11291) );
  ANDN U17041 ( .B(n16548), .A(n16549), .Z(n16546) );
  XOR U17042 ( .A(n16550), .B(n16551), .Z(n8399) );
  XNOR U17043 ( .A(n3857), .B(n5165), .Z(n16551) );
  XNOR U17044 ( .A(n16552), .B(n9823), .Z(n5165) );
  IV U17045 ( .A(n12144), .Z(n9823) );
  XOR U17046 ( .A(n16553), .B(n16202), .Z(n12144) );
  IV U17047 ( .A(n9899), .Z(n16202) );
  XNOR U17048 ( .A(n16554), .B(n15731), .Z(n9899) );
  XNOR U17049 ( .A(n16555), .B(n16556), .Z(n15731) );
  XOR U17050 ( .A(n11697), .B(n12763), .Z(n16556) );
  XNOR U17051 ( .A(n16557), .B(n13457), .Z(n12763) );
  NOR U17052 ( .A(n16558), .B(n14894), .Z(n16557) );
  XNOR U17053 ( .A(n16559), .B(n13452), .Z(n11697) );
  NOR U17054 ( .A(n13451), .B(n14891), .Z(n16559) );
  XOR U17055 ( .A(n11779), .B(n16560), .Z(n16555) );
  XNOR U17056 ( .A(n10639), .B(n11457), .Z(n16560) );
  XNOR U17057 ( .A(n16561), .B(n16562), .Z(n11457) );
  ANDN U17058 ( .B(n14883), .A(n13447), .Z(n16561) );
  XNOR U17059 ( .A(n16563), .B(n16564), .Z(n10639) );
  ANDN U17060 ( .B(n16565), .A(n14887), .Z(n16563) );
  XNOR U17061 ( .A(n16566), .B(n13461), .Z(n11779) );
  NOR U17062 ( .A(n13462), .B(n14880), .Z(n16566) );
  ANDN U17063 ( .B(n12004), .A(n12005), .Z(n16552) );
  XOR U17064 ( .A(n9452), .B(n16540), .Z(n12005) );
  XNOR U17065 ( .A(n16567), .B(n14779), .Z(n16540) );
  ANDN U17066 ( .B(n16568), .A(n16569), .Z(n16567) );
  XOR U17067 ( .A(n15474), .B(n11069), .Z(n12004) );
  IV U17068 ( .A(n12395), .Z(n11069) );
  XNOR U17069 ( .A(n11725), .B(n13131), .Z(n12395) );
  XNOR U17070 ( .A(n16570), .B(n16571), .Z(n13131) );
  XNOR U17071 ( .A(n12786), .B(n11338), .Z(n16571) );
  XNOR U17072 ( .A(n16572), .B(n16573), .Z(n11338) );
  AND U17073 ( .A(n15326), .B(n15487), .Z(n16572) );
  XOR U17074 ( .A(n16574), .B(n16575), .Z(n15326) );
  XNOR U17075 ( .A(n16576), .B(n16577), .Z(n12786) );
  ANDN U17076 ( .B(n15484), .A(n15485), .Z(n16576) );
  XNOR U17077 ( .A(n16578), .B(n16579), .Z(n15485) );
  XOR U17078 ( .A(n16580), .B(n16581), .Z(n16570) );
  XNOR U17079 ( .A(n10283), .B(n11052), .Z(n16581) );
  XOR U17080 ( .A(n16582), .B(n16583), .Z(n11052) );
  ANDN U17081 ( .B(n15318), .A(n15490), .Z(n16582) );
  XOR U17082 ( .A(n16584), .B(n16585), .Z(n15318) );
  XNOR U17083 ( .A(n16586), .B(n16587), .Z(n10283) );
  AND U17084 ( .A(n15492), .B(n15309), .Z(n16586) );
  XNOR U17085 ( .A(n16588), .B(n16589), .Z(n15309) );
  XOR U17086 ( .A(n16590), .B(n16591), .Z(n11725) );
  XNOR U17087 ( .A(n15162), .B(n12779), .Z(n16591) );
  XNOR U17088 ( .A(n16592), .B(n15169), .Z(n12779) );
  ANDN U17089 ( .B(n15470), .A(n15168), .Z(n16592) );
  XNOR U17090 ( .A(n16593), .B(n16594), .Z(n15162) );
  ANDN U17091 ( .B(n15476), .A(n14630), .Z(n16593) );
  XOR U17092 ( .A(n16595), .B(n16596), .Z(n14630) );
  XNOR U17093 ( .A(n12505), .B(n16597), .Z(n16590) );
  XOR U17094 ( .A(n9516), .B(n11879), .Z(n16597) );
  XNOR U17095 ( .A(n16598), .B(n16599), .Z(n11879) );
  ANDN U17096 ( .B(n16490), .A(n14626), .Z(n16598) );
  XOR U17097 ( .A(n16600), .B(n16601), .Z(n14626) );
  XOR U17098 ( .A(n16602), .B(n15172), .Z(n9516) );
  AND U17099 ( .A(n14634), .B(n15173), .Z(n16602) );
  XNOR U17100 ( .A(n16603), .B(n16604), .Z(n15173) );
  XNOR U17101 ( .A(n16605), .B(n16529), .Z(n14634) );
  XOR U17102 ( .A(n16606), .B(n15178), .Z(n12505) );
  ANDN U17103 ( .B(n15179), .A(n14621), .Z(n16606) );
  XOR U17104 ( .A(n16607), .B(n16608), .Z(n14621) );
  XOR U17105 ( .A(n16609), .B(n16610), .Z(n15179) );
  XNOR U17106 ( .A(n16611), .B(n15168), .Z(n15474) );
  XNOR U17107 ( .A(n16612), .B(n16613), .Z(n15168) );
  NOR U17108 ( .A(n16614), .B(n15470), .Z(n16611) );
  XNOR U17109 ( .A(n16615), .B(n16616), .Z(n15470) );
  XNOR U17110 ( .A(n16617), .B(n8489), .Z(n3857) );
  XOR U17111 ( .A(n16470), .B(n13013), .Z(n8489) );
  IV U17112 ( .A(n13069), .Z(n13013) );
  XNOR U17113 ( .A(n16618), .B(n15533), .Z(n16470) );
  ANDN U17114 ( .B(n14663), .A(n13221), .Z(n16618) );
  XOR U17115 ( .A(n16619), .B(n16620), .Z(n13221) );
  XOR U17116 ( .A(n10317), .B(n16621), .Z(n11995) );
  IV U17117 ( .A(n16493), .Z(n10317) );
  XOR U17118 ( .A(n12280), .B(n15116), .Z(n11996) );
  XNOR U17119 ( .A(n16622), .B(n16623), .Z(n15116) );
  ANDN U17120 ( .B(n16624), .A(n14279), .Z(n16622) );
  XNOR U17121 ( .A(n13327), .B(n12416), .Z(n12280) );
  XOR U17122 ( .A(n16625), .B(n16626), .Z(n12416) );
  XNOR U17123 ( .A(n14928), .B(n15440), .Z(n16626) );
  XOR U17124 ( .A(n16627), .B(n16628), .Z(n15440) );
  ANDN U17125 ( .B(n16629), .A(n16630), .Z(n16627) );
  XNOR U17126 ( .A(n16631), .B(n16445), .Z(n14928) );
  NOR U17127 ( .A(n16632), .B(n16633), .Z(n16631) );
  XOR U17128 ( .A(n14975), .B(n16634), .Z(n16625) );
  XOR U17129 ( .A(n13125), .B(n12254), .Z(n16634) );
  XNOR U17130 ( .A(n16635), .B(n16455), .Z(n12254) );
  ANDN U17131 ( .B(n16636), .A(n16637), .Z(n16635) );
  XNOR U17132 ( .A(n16638), .B(n16449), .Z(n13125) );
  NOR U17133 ( .A(n16639), .B(n16640), .Z(n16638) );
  XNOR U17134 ( .A(n16641), .B(n16458), .Z(n14975) );
  AND U17135 ( .A(n16642), .B(n16643), .Z(n16641) );
  XOR U17136 ( .A(n16644), .B(n16645), .Z(n13327) );
  XNOR U17137 ( .A(n9926), .B(n12951), .Z(n16645) );
  XNOR U17138 ( .A(n16646), .B(n14285), .Z(n12951) );
  XOR U17139 ( .A(n16647), .B(n14291), .Z(n9926) );
  ANDN U17140 ( .B(n15118), .A(n16648), .Z(n16647) );
  XNOR U17141 ( .A(n16649), .B(n16650), .Z(n16644) );
  XOR U17142 ( .A(n13331), .B(n11287), .Z(n16650) );
  XOR U17143 ( .A(n16651), .B(n16652), .Z(n11287) );
  ANDN U17144 ( .B(n15114), .A(n15112), .Z(n16651) );
  XNOR U17145 ( .A(n16653), .B(n14281), .Z(n13331) );
  ANDN U17146 ( .B(n16623), .A(n16624), .Z(n16653) );
  XOR U17147 ( .A(n5867), .B(n16654), .Z(n16550) );
  XNOR U17148 ( .A(n1753), .B(n12139), .Z(n16654) );
  XNOR U17149 ( .A(n16655), .B(n8500), .Z(n12139) );
  XOR U17150 ( .A(n16656), .B(n11213), .Z(n8500) );
  XNOR U17151 ( .A(n16657), .B(n16658), .Z(n11213) );
  ANDN U17152 ( .B(n11993), .A(n11992), .Z(n16655) );
  IV U17153 ( .A(n12150), .Z(n11992) );
  XOR U17154 ( .A(n11301), .B(n16659), .Z(n12150) );
  XOR U17155 ( .A(n16660), .B(n16661), .Z(n13442) );
  XNOR U17156 ( .A(n9661), .B(n10158), .Z(n16661) );
  XOR U17157 ( .A(n16662), .B(n13340), .Z(n10158) );
  XOR U17158 ( .A(n16663), .B(n16664), .Z(n13340) );
  AND U17159 ( .A(n16665), .B(n13339), .Z(n16662) );
  XOR U17160 ( .A(n16666), .B(n13346), .Z(n9661) );
  XNOR U17161 ( .A(n16667), .B(n16407), .Z(n13346) );
  IV U17162 ( .A(n16668), .Z(n16407) );
  ANDN U17163 ( .B(n16669), .A(n16670), .Z(n16666) );
  XOR U17164 ( .A(n9412), .B(n16671), .Z(n16660) );
  XOR U17165 ( .A(n13332), .B(n13228), .Z(n16671) );
  XNOR U17166 ( .A(n16672), .B(n14874), .Z(n13228) );
  XNOR U17167 ( .A(n16673), .B(n16674), .Z(n14874) );
  XNOR U17168 ( .A(n16676), .B(n13349), .Z(n13332) );
  ANDN U17169 ( .B(n16677), .A(n16678), .Z(n16676) );
  XOR U17170 ( .A(n16679), .B(n14485), .Z(n9412) );
  XOR U17171 ( .A(n16680), .B(n16105), .Z(n14485) );
  ANDN U17172 ( .B(n16681), .A(n16682), .Z(n16679) );
  XOR U17173 ( .A(n16683), .B(n16684), .Z(n14186) );
  XNOR U17174 ( .A(n11427), .B(n12364), .Z(n16684) );
  XOR U17175 ( .A(n16685), .B(n15157), .Z(n12364) );
  XOR U17176 ( .A(n16688), .B(n15161), .Z(n11427) );
  NOR U17177 ( .A(n16689), .B(n16690), .Z(n16688) );
  XOR U17178 ( .A(n10618), .B(n16691), .Z(n16683) );
  XNOR U17179 ( .A(n10345), .B(n11852), .Z(n16691) );
  XNOR U17180 ( .A(n16692), .B(n15150), .Z(n11852) );
  XNOR U17181 ( .A(n16695), .B(n16696), .Z(n10345) );
  ANDN U17182 ( .B(n16697), .A(n16698), .Z(n16695) );
  XNOR U17183 ( .A(n16699), .B(n15147), .Z(n10618) );
  ANDN U17184 ( .B(n16700), .A(n16701), .Z(n16699) );
  XOR U17185 ( .A(n16702), .B(n16703), .Z(n11993) );
  XNOR U17186 ( .A(n16704), .B(n8494), .Z(n1753) );
  XNOR U17187 ( .A(n16215), .B(n11460), .Z(n8494) );
  XNOR U17188 ( .A(n16496), .B(n15008), .Z(n11460) );
  XOR U17189 ( .A(n16705), .B(n16706), .Z(n15008) );
  XOR U17190 ( .A(n12074), .B(n12814), .Z(n16706) );
  XOR U17191 ( .A(n16707), .B(n15932), .Z(n12814) );
  ANDN U17192 ( .B(n16708), .A(n16709), .Z(n16707) );
  XNOR U17193 ( .A(n16710), .B(n15915), .Z(n12074) );
  ANDN U17194 ( .B(n16711), .A(n16712), .Z(n16710) );
  XNOR U17195 ( .A(n11973), .B(n16713), .Z(n16705) );
  XNOR U17196 ( .A(n15909), .B(n13947), .Z(n16713) );
  XNOR U17197 ( .A(n16714), .B(n15925), .Z(n13947) );
  ANDN U17198 ( .B(n16715), .A(n15924), .Z(n16714) );
  XOR U17199 ( .A(n16716), .B(n15919), .Z(n15909) );
  AND U17200 ( .A(n16717), .B(n15920), .Z(n16716) );
  XOR U17201 ( .A(n16718), .B(n15928), .Z(n11973) );
  ANDN U17202 ( .B(n16719), .A(n16720), .Z(n16718) );
  XOR U17203 ( .A(n16721), .B(n16722), .Z(n16496) );
  XOR U17204 ( .A(n9789), .B(n11896), .Z(n16722) );
  XNOR U17205 ( .A(n16723), .B(n16724), .Z(n11896) );
  XNOR U17206 ( .A(n16725), .B(n16726), .Z(n9789) );
  ANDN U17207 ( .B(n16213), .A(n14726), .Z(n16725) );
  XOR U17208 ( .A(n16727), .B(n16728), .Z(n14726) );
  XOR U17209 ( .A(n9943), .B(n16729), .Z(n16721) );
  XOR U17210 ( .A(n10704), .B(n10407), .Z(n16729) );
  XNOR U17211 ( .A(n16730), .B(n13502), .Z(n10407) );
  ANDN U17212 ( .B(n16211), .A(n16209), .Z(n16730) );
  IV U17213 ( .A(n13503), .Z(n16209) );
  XOR U17214 ( .A(n16731), .B(n16732), .Z(n13503) );
  XOR U17215 ( .A(n16733), .B(n16734), .Z(n16211) );
  XOR U17216 ( .A(n16735), .B(n13499), .Z(n10704) );
  ANDN U17217 ( .B(n16217), .A(n13498), .Z(n16735) );
  XOR U17218 ( .A(n16736), .B(n16737), .Z(n13498) );
  IV U17219 ( .A(n14730), .Z(n16217) );
  XOR U17220 ( .A(n16738), .B(n16063), .Z(n14730) );
  IV U17221 ( .A(n16739), .Z(n16063) );
  XNOR U17222 ( .A(n16740), .B(n13494), .Z(n9943) );
  IV U17223 ( .A(n16741), .Z(n13494) );
  NOR U17224 ( .A(n14719), .B(n13493), .Z(n16740) );
  XOR U17225 ( .A(n16742), .B(n16061), .Z(n13493) );
  XNOR U17226 ( .A(n16743), .B(n16744), .Z(n14719) );
  XNOR U17227 ( .A(n16745), .B(n13506), .Z(n16215) );
  XNOR U17228 ( .A(n16746), .B(n16008), .Z(n13506) );
  ANDN U17229 ( .B(n14724), .A(n14723), .Z(n16745) );
  XOR U17230 ( .A(n16747), .B(n16748), .Z(n14723) );
  AND U17231 ( .A(n12001), .B(n12002), .Z(n16704) );
  XNOR U17232 ( .A(n16749), .B(n10180), .Z(n12002) );
  XNOR U17233 ( .A(n15246), .B(n12650), .Z(n10180) );
  XNOR U17234 ( .A(n16750), .B(n16751), .Z(n12650) );
  XNOR U17235 ( .A(n11798), .B(n11357), .Z(n16751) );
  XOR U17236 ( .A(n16752), .B(n12870), .Z(n11357) );
  XOR U17237 ( .A(n16753), .B(n16754), .Z(n12870) );
  ANDN U17238 ( .B(n16755), .A(n16295), .Z(n16752) );
  XNOR U17239 ( .A(n16756), .B(n15992), .Z(n11798) );
  XOR U17240 ( .A(n16757), .B(n16758), .Z(n15992) );
  ANDN U17241 ( .B(n16759), .A(n16288), .Z(n16756) );
  XOR U17242 ( .A(n10780), .B(n16760), .Z(n16750) );
  XNOR U17243 ( .A(n16281), .B(n13233), .Z(n16760) );
  XOR U17244 ( .A(n16761), .B(n14386), .Z(n13233) );
  XOR U17245 ( .A(n16762), .B(n16763), .Z(n14386) );
  ANDN U17246 ( .B(n16764), .A(n16291), .Z(n16761) );
  XOR U17247 ( .A(n16765), .B(n12865), .Z(n16281) );
  XNOR U17248 ( .A(n16766), .B(n16767), .Z(n12865) );
  ANDN U17249 ( .B(n16286), .A(n16768), .Z(n16765) );
  XNOR U17250 ( .A(n16769), .B(n12859), .Z(n10780) );
  XOR U17251 ( .A(n16770), .B(n16771), .Z(n12859) );
  ANDN U17252 ( .B(n16772), .A(n16293), .Z(n16769) );
  XOR U17253 ( .A(n16773), .B(n16774), .Z(n15246) );
  XNOR U17254 ( .A(n16775), .B(n13381), .Z(n16774) );
  NOR U17255 ( .A(n15986), .B(n16778), .Z(n16776) );
  XOR U17256 ( .A(n12748), .B(n16779), .Z(n16773) );
  XOR U17257 ( .A(n11890), .B(n12705), .Z(n16779) );
  XNOR U17258 ( .A(n16780), .B(n16781), .Z(n12705) );
  ANDN U17259 ( .B(n16782), .A(n15969), .Z(n16780) );
  XNOR U17260 ( .A(n16783), .B(n16784), .Z(n11890) );
  NOR U17261 ( .A(n16785), .B(n15973), .Z(n16783) );
  XOR U17262 ( .A(n16786), .B(n16787), .Z(n12748) );
  AND U17263 ( .A(n15978), .B(n16788), .Z(n16786) );
  XOR U17264 ( .A(n15826), .B(n9757), .Z(n12001) );
  XNOR U17265 ( .A(n14263), .B(n12960), .Z(n9757) );
  XNOR U17266 ( .A(n16789), .B(n16790), .Z(n12960) );
  XNOR U17267 ( .A(n10164), .B(n13924), .Z(n16790) );
  XNOR U17268 ( .A(n16791), .B(n16792), .Z(n13924) );
  ANDN U17269 ( .B(n15821), .A(n15819), .Z(n16791) );
  XNOR U17270 ( .A(n16793), .B(n14913), .Z(n10164) );
  ANDN U17271 ( .B(n15833), .A(n15832), .Z(n16793) );
  IV U17272 ( .A(n16794), .Z(n15832) );
  XOR U17273 ( .A(n13044), .B(n16795), .Z(n16789) );
  XNOR U17274 ( .A(n9232), .B(n12059), .Z(n16795) );
  XNOR U17275 ( .A(n16796), .B(n14910), .Z(n12059) );
  ANDN U17276 ( .B(n15823), .A(n15824), .Z(n16796) );
  XOR U17277 ( .A(n16797), .B(n14919), .Z(n9232) );
  NOR U17278 ( .A(n15829), .B(n15828), .Z(n16797) );
  XNOR U17279 ( .A(n16798), .B(n14924), .Z(n13044) );
  ANDN U17280 ( .B(n16799), .A(n16800), .Z(n16798) );
  XOR U17281 ( .A(n16801), .B(n16802), .Z(n14263) );
  XOR U17282 ( .A(n9960), .B(n13553), .Z(n16802) );
  XOR U17283 ( .A(n16803), .B(n13931), .Z(n13553) );
  ANDN U17284 ( .B(n13932), .A(n15812), .Z(n16803) );
  IV U17285 ( .A(n15810), .Z(n13932) );
  XOR U17286 ( .A(n16313), .B(n16804), .Z(n15810) );
  XNOR U17287 ( .A(n16805), .B(n16806), .Z(n9960) );
  ANDN U17288 ( .B(n15799), .A(n15800), .Z(n16805) );
  XNOR U17289 ( .A(n9148), .B(n16807), .Z(n16801) );
  XNOR U17290 ( .A(n9979), .B(n13070), .Z(n16807) );
  XOR U17291 ( .A(n16808), .B(n15498), .Z(n13070) );
  ANDN U17292 ( .B(n15499), .A(n15807), .Z(n16808) );
  XOR U17293 ( .A(n16809), .B(n16810), .Z(n15499) );
  XNOR U17294 ( .A(n16811), .B(n13938), .Z(n9979) );
  NOR U17295 ( .A(n15814), .B(n13937), .Z(n16811) );
  XNOR U17296 ( .A(n16812), .B(n16813), .Z(n13937) );
  XNOR U17297 ( .A(n16814), .B(n13942), .Z(n9148) );
  ANDN U17298 ( .B(n15803), .A(n13941), .Z(n16814) );
  XOR U17299 ( .A(n16815), .B(n16816), .Z(n13941) );
  XNOR U17300 ( .A(n16817), .B(n16799), .Z(n15826) );
  ANDN U17301 ( .B(n16800), .A(n14922), .Z(n16817) );
  XNOR U17302 ( .A(n16818), .B(n8503), .Z(n5867) );
  XOR U17303 ( .A(n15071), .B(n10388), .Z(n8503) );
  XNOR U17304 ( .A(n11706), .B(n13418), .Z(n10388) );
  XOR U17305 ( .A(n16819), .B(n16820), .Z(n13418) );
  XNOR U17306 ( .A(n10981), .B(n10585), .Z(n16820) );
  XNOR U17307 ( .A(n16821), .B(n16302), .Z(n10585) );
  ANDN U17308 ( .B(n15076), .A(n15074), .Z(n16821) );
  XNOR U17309 ( .A(n16822), .B(n16823), .Z(n15076) );
  ANDN U17310 ( .B(n15064), .A(n15063), .Z(n16824) );
  XOR U17311 ( .A(n16825), .B(n16826), .Z(n15064) );
  XOR U17312 ( .A(n12994), .B(n16827), .Z(n16819) );
  XNOR U17313 ( .A(n16026), .B(n10048), .Z(n16827) );
  XNOR U17314 ( .A(n16828), .B(n16306), .Z(n10048) );
  AND U17315 ( .A(n15067), .B(n15069), .Z(n16828) );
  XNOR U17316 ( .A(n16829), .B(n16830), .Z(n15069) );
  XOR U17317 ( .A(n16831), .B(n16309), .Z(n16026) );
  XOR U17318 ( .A(n16832), .B(n16502), .Z(n15575) );
  XNOR U17319 ( .A(n16833), .B(n16311), .Z(n12994) );
  ANDN U17320 ( .B(n15571), .A(n16834), .Z(n16833) );
  XOR U17321 ( .A(n16835), .B(n16836), .Z(n11706) );
  XOR U17322 ( .A(n12681), .B(n11060), .Z(n16836) );
  XNOR U17323 ( .A(n16837), .B(n16034), .Z(n11060) );
  IV U17324 ( .A(n14031), .Z(n16034) );
  XOR U17325 ( .A(n16838), .B(n16068), .Z(n14031) );
  ANDN U17326 ( .B(n13433), .A(n16033), .Z(n16837) );
  XNOR U17327 ( .A(n16839), .B(n14036), .Z(n12681) );
  XOR U17328 ( .A(n16840), .B(n16841), .Z(n14036) );
  ANDN U17329 ( .B(n14899), .A(n16038), .Z(n16839) );
  XOR U17330 ( .A(n14363), .B(n16842), .Z(n16835) );
  XNOR U17331 ( .A(n10966), .B(n11615), .Z(n16842) );
  XNOR U17332 ( .A(n16843), .B(n14041), .Z(n11615) );
  XOR U17333 ( .A(n16844), .B(n16845), .Z(n14041) );
  AND U17334 ( .A(n13427), .B(n16046), .Z(n16843) );
  XOR U17335 ( .A(n16846), .B(n14029), .Z(n10966) );
  XOR U17336 ( .A(n16847), .B(n16848), .Z(n14029) );
  NOR U17337 ( .A(n16849), .B(n16042), .Z(n16846) );
  XNOR U17338 ( .A(n16850), .B(n14039), .Z(n14363) );
  XOR U17339 ( .A(n16851), .B(n16852), .Z(n14039) );
  ANDN U17340 ( .B(n16050), .A(n16853), .Z(n16850) );
  XNOR U17341 ( .A(n16854), .B(n16834), .Z(n15071) );
  NOR U17342 ( .A(n15572), .B(n15571), .Z(n16854) );
  XOR U17343 ( .A(n16855), .B(n16856), .Z(n15571) );
  XOR U17344 ( .A(n16857), .B(n16858), .Z(n15572) );
  AND U17345 ( .A(n14509), .B(n12147), .Z(n16818) );
  XOR U17346 ( .A(n16859), .B(n12147), .Z(n11998) );
  XOR U17347 ( .A(n11698), .B(n14268), .Z(n12147) );
  XNOR U17348 ( .A(n16860), .B(n14228), .Z(n14268) );
  ANDN U17349 ( .B(n13571), .A(n16861), .Z(n16860) );
  NOR U17350 ( .A(n14510), .B(n14509), .Z(n16859) );
  XOR U17351 ( .A(n16360), .B(n12685), .Z(n14509) );
  XOR U17352 ( .A(n11847), .B(n16862), .Z(n12685) );
  XOR U17353 ( .A(n16863), .B(n16864), .Z(n11847) );
  XNOR U17354 ( .A(n10924), .B(n11465), .Z(n16864) );
  XNOR U17355 ( .A(n16865), .B(n16866), .Z(n11465) );
  ANDN U17356 ( .B(n14802), .A(n16357), .Z(n16865) );
  XNOR U17357 ( .A(n16867), .B(n16868), .Z(n14802) );
  XNOR U17358 ( .A(n16869), .B(n16870), .Z(n10924) );
  AND U17359 ( .A(n16364), .B(n14795), .Z(n16869) );
  XOR U17360 ( .A(n16871), .B(n16872), .Z(n14795) );
  XNOR U17361 ( .A(n11328), .B(n16873), .Z(n16863) );
  XNOR U17362 ( .A(n9534), .B(n16874), .Z(n16873) );
  XNOR U17363 ( .A(n16875), .B(n16876), .Z(n9534) );
  ANDN U17364 ( .B(n16362), .A(n14791), .Z(n16875) );
  XOR U17365 ( .A(n16879), .B(n16880), .Z(n11328) );
  AND U17366 ( .A(n16881), .B(n16335), .Z(n16879) );
  XOR U17367 ( .A(n16882), .B(n16881), .Z(n16360) );
  NOR U17368 ( .A(n16335), .B(n16336), .Z(n16882) );
  XOR U17369 ( .A(n16883), .B(n16674), .Z(n16335) );
  XOR U17370 ( .A(n13850), .B(n14192), .Z(n14510) );
  XNOR U17371 ( .A(n14262), .B(n16884), .Z(n14192) );
  XOR U17372 ( .A(n16885), .B(n16886), .Z(n14262) );
  XNOR U17373 ( .A(n12495), .B(n14675), .Z(n16886) );
  XNOR U17374 ( .A(n16887), .B(n14685), .Z(n14675) );
  ANDN U17375 ( .B(n13852), .A(n13853), .Z(n16887) );
  XNOR U17376 ( .A(n16888), .B(n16889), .Z(n13852) );
  XNOR U17377 ( .A(n16890), .B(n15103), .Z(n12495) );
  ANDN U17378 ( .B(n13863), .A(n13862), .Z(n16890) );
  XOR U17379 ( .A(n16891), .B(n14176), .Z(n13862) );
  IV U17380 ( .A(n16892), .Z(n14176) );
  XOR U17381 ( .A(n11344), .B(n16893), .Z(n16885) );
  XNOR U17382 ( .A(n11084), .B(n12212), .Z(n16893) );
  XNOR U17383 ( .A(n16894), .B(n16895), .Z(n12212) );
  ANDN U17384 ( .B(n13858), .A(n13860), .Z(n16894) );
  XNOR U17385 ( .A(n16896), .B(n16897), .Z(n11084) );
  ANDN U17386 ( .B(n14195), .A(n14194), .Z(n16896) );
  XNOR U17387 ( .A(n16898), .B(n14688), .Z(n11344) );
  ANDN U17388 ( .B(n14689), .A(n16899), .Z(n16898) );
  XNOR U17389 ( .A(n16900), .B(n14689), .Z(n13850) );
  XOR U17390 ( .A(n16901), .B(n16412), .Z(n14689) );
  ANDN U17391 ( .B(n16899), .A(n16902), .Z(n16900) );
  XOR U17392 ( .A(n16903), .B(n2608), .Z(out[0]) );
  XOR U17393 ( .A(n3363), .B(n10500), .Z(n2608) );
  XNOR U17394 ( .A(n16904), .B(n8616), .Z(n10500) );
  IV U17395 ( .A(n16905), .Z(n8616) );
  AND U17396 ( .A(n10354), .B(n10534), .Z(n16904) );
  XOR U17397 ( .A(n10589), .B(n16906), .Z(n10354) );
  IV U17398 ( .A(n11106), .Z(n10589) );
  XNOR U17399 ( .A(n12678), .B(n15105), .Z(n11106) );
  XOR U17400 ( .A(n16907), .B(n16908), .Z(n15105) );
  XOR U17401 ( .A(n11049), .B(n12415), .Z(n16908) );
  XOR U17402 ( .A(n16909), .B(n16636), .Z(n12415) );
  AND U17403 ( .A(n16637), .B(n16453), .Z(n16909) );
  XNOR U17404 ( .A(n16910), .B(n16633), .Z(n11049) );
  ANDN U17405 ( .B(n16632), .A(n16443), .Z(n16910) );
  XNOR U17406 ( .A(n10306), .B(n16911), .Z(n16907) );
  XOR U17407 ( .A(n12072), .B(n10778), .Z(n16911) );
  XNOR U17408 ( .A(n16912), .B(n16639), .Z(n10778) );
  IV U17409 ( .A(n16913), .Z(n16639) );
  ANDN U17410 ( .B(n16640), .A(n16447), .Z(n16912) );
  IV U17411 ( .A(n16914), .Z(n16447) );
  XNOR U17412 ( .A(n16915), .B(n16629), .Z(n12072) );
  ANDN U17413 ( .B(n16630), .A(n16916), .Z(n16915) );
  XNOR U17414 ( .A(n16917), .B(n16642), .Z(n10306) );
  NOR U17415 ( .A(n16457), .B(n16643), .Z(n16917) );
  XOR U17416 ( .A(n16918), .B(n16919), .Z(n12678) );
  XOR U17417 ( .A(n11554), .B(n13840), .Z(n16919) );
  XOR U17418 ( .A(n16920), .B(n16921), .Z(n13840) );
  NOR U17419 ( .A(n16922), .B(n16424), .Z(n16920) );
  XNOR U17420 ( .A(n16923), .B(n16924), .Z(n11554) );
  ANDN U17421 ( .B(n16429), .A(n16925), .Z(n16923) );
  XOR U17422 ( .A(n10184), .B(n16926), .Z(n16918) );
  XOR U17423 ( .A(n16927), .B(n14733), .Z(n16926) );
  XNOR U17424 ( .A(n16928), .B(n16929), .Z(n14733) );
  ANDN U17425 ( .B(n16930), .A(n16931), .Z(n16928) );
  XOR U17426 ( .A(n16932), .B(n16933), .Z(n10184) );
  ANDN U17427 ( .B(n16934), .A(n16433), .Z(n16932) );
  IV U17428 ( .A(n2210), .Z(n3363) );
  XOR U17429 ( .A(n8045), .B(n6003), .Z(n2210) );
  XOR U17430 ( .A(n16935), .B(n16936), .Z(n6003) );
  XNOR U17431 ( .A(n5302), .B(n3751), .Z(n16936) );
  XOR U17432 ( .A(n16938), .B(n10850), .Z(n8619) );
  XNOR U17433 ( .A(n11950), .B(n13595), .Z(n10850) );
  XNOR U17434 ( .A(n16939), .B(n16940), .Z(n13595) );
  XOR U17435 ( .A(n14851), .B(n11593), .Z(n16940) );
  XOR U17436 ( .A(n16941), .B(n15777), .Z(n11593) );
  ANDN U17437 ( .B(n15778), .A(n12429), .Z(n16941) );
  XNOR U17438 ( .A(n16942), .B(n15781), .Z(n14851) );
  IV U17439 ( .A(n16943), .Z(n15781) );
  AND U17440 ( .A(n16944), .B(n15782), .Z(n16942) );
  XOR U17441 ( .A(n10273), .B(n16945), .Z(n16939) );
  XOR U17442 ( .A(n12401), .B(n11439), .Z(n16945) );
  XOR U17443 ( .A(n16946), .B(n15786), .Z(n11439) );
  ANDN U17444 ( .B(n12347), .A(n15785), .Z(n16946) );
  IV U17445 ( .A(n16947), .Z(n15785) );
  XNOR U17446 ( .A(n16948), .B(n15788), .Z(n12401) );
  ANDN U17447 ( .B(n15789), .A(n15275), .Z(n16948) );
  XNOR U17448 ( .A(n16949), .B(n15792), .Z(n10273) );
  XOR U17449 ( .A(n16950), .B(n16951), .Z(n11950) );
  XNOR U17450 ( .A(n12660), .B(n10641), .Z(n16951) );
  XNOR U17451 ( .A(n16952), .B(n14314), .Z(n10641) );
  IV U17452 ( .A(n14861), .Z(n14314) );
  XNOR U17453 ( .A(n16953), .B(n16954), .Z(n14861) );
  ANDN U17454 ( .B(n14862), .A(n15669), .Z(n16952) );
  IV U17455 ( .A(n16955), .Z(n15669) );
  XOR U17456 ( .A(n16956), .B(n14309), .Z(n12660) );
  XOR U17457 ( .A(n16957), .B(n16958), .Z(n14309) );
  NOR U17458 ( .A(n14858), .B(n15660), .Z(n16956) );
  XOR U17459 ( .A(n11601), .B(n16959), .Z(n16950) );
  XOR U17460 ( .A(n10285), .B(n9462), .Z(n16959) );
  XNOR U17461 ( .A(n16960), .B(n15700), .Z(n9462) );
  IV U17462 ( .A(n14866), .Z(n15700) );
  XOR U17463 ( .A(n16961), .B(n16962), .Z(n14866) );
  NOR U17464 ( .A(n14865), .B(n15665), .Z(n16960) );
  XOR U17465 ( .A(n16963), .B(n14317), .Z(n10285) );
  XOR U17466 ( .A(n16964), .B(n16664), .Z(n14317) );
  NOR U17467 ( .A(n15673), .B(n14856), .Z(n16963) );
  XOR U17468 ( .A(n16965), .B(n14321), .Z(n11601) );
  XOR U17469 ( .A(n16966), .B(n16967), .Z(n14321) );
  ANDN U17470 ( .B(n8620), .A(n7933), .Z(n16937) );
  XOR U17471 ( .A(n16968), .B(n10962), .Z(n7933) );
  XNOR U17472 ( .A(n16969), .B(n13797), .Z(n10962) );
  XNOR U17473 ( .A(n16970), .B(n16971), .Z(n13797) );
  XNOR U17474 ( .A(n11916), .B(n9948), .Z(n16971) );
  XNOR U17475 ( .A(n16972), .B(n14607), .Z(n9948) );
  NOR U17476 ( .A(n14013), .B(n16973), .Z(n16972) );
  XOR U17477 ( .A(n16974), .B(n16975), .Z(n11916) );
  ANDN U17478 ( .B(n14017), .A(n16976), .Z(n16974) );
  XOR U17479 ( .A(n13016), .B(n16977), .Z(n16970) );
  XNOR U17480 ( .A(n16978), .B(n13819), .Z(n16977) );
  XNOR U17481 ( .A(n16979), .B(n14604), .Z(n13819) );
  AND U17482 ( .A(n14007), .B(n16980), .Z(n16979) );
  XNOR U17483 ( .A(n16981), .B(n14611), .Z(n13016) );
  ANDN U17484 ( .B(n14003), .A(n16982), .Z(n16981) );
  XOR U17485 ( .A(n15458), .B(n11081), .Z(n8620) );
  XOR U17486 ( .A(n13235), .B(n15589), .Z(n11081) );
  XNOR U17487 ( .A(n16983), .B(n16984), .Z(n15589) );
  XNOR U17488 ( .A(n11766), .B(n14150), .Z(n16984) );
  XOR U17489 ( .A(n16985), .B(n13749), .Z(n14150) );
  XOR U17490 ( .A(n16986), .B(n16841), .Z(n13749) );
  AND U17491 ( .A(n14239), .B(n15455), .Z(n16985) );
  XOR U17492 ( .A(n15999), .B(n16987), .Z(n14239) );
  XNOR U17493 ( .A(n16988), .B(n13757), .Z(n11766) );
  XNOR U17494 ( .A(n16989), .B(n15339), .Z(n13757) );
  ANDN U17495 ( .B(n14247), .A(n16990), .Z(n16988) );
  XOR U17496 ( .A(n16991), .B(n16992), .Z(n14247) );
  XOR U17497 ( .A(n14233), .B(n16993), .Z(n16983) );
  XOR U17498 ( .A(n12591), .B(n10281), .Z(n16993) );
  XNOR U17499 ( .A(n16994), .B(n14243), .Z(n10281) );
  XOR U17500 ( .A(n16995), .B(n16996), .Z(n14243) );
  ANDN U17501 ( .B(n15451), .A(n14242), .Z(n16994) );
  XNOR U17502 ( .A(n16997), .B(n16998), .Z(n14242) );
  XNOR U17503 ( .A(n16999), .B(n13754), .Z(n12591) );
  IV U17504 ( .A(n14249), .Z(n13754) );
  XOR U17505 ( .A(n17000), .B(n17001), .Z(n14249) );
  AND U17506 ( .A(n14250), .B(n15453), .Z(n16999) );
  XNOR U17507 ( .A(n17002), .B(n16668), .Z(n14250) );
  XOR U17508 ( .A(n17003), .B(n14253), .Z(n14233) );
  AND U17509 ( .A(n14254), .B(n15447), .Z(n17003) );
  XOR U17510 ( .A(n16097), .B(n17004), .Z(n14254) );
  XOR U17511 ( .A(n17005), .B(n17006), .Z(n13235) );
  XNOR U17512 ( .A(n9947), .B(n9560), .Z(n17006) );
  XNOR U17513 ( .A(n17007), .B(n13723), .Z(n9560) );
  ANDN U17514 ( .B(n15461), .A(n13722), .Z(n17007) );
  XOR U17515 ( .A(n17008), .B(n17009), .Z(n13722) );
  XNOR U17516 ( .A(n17010), .B(n16101), .Z(n15461) );
  XNOR U17517 ( .A(n17011), .B(n13736), .Z(n9947) );
  AND U17518 ( .A(n14504), .B(n13737), .Z(n17011) );
  XOR U17519 ( .A(n17012), .B(n17013), .Z(n13737) );
  XNOR U17520 ( .A(n17014), .B(n17015), .Z(n14504) );
  XOR U17521 ( .A(n11168), .B(n17016), .Z(n17005) );
  XNOR U17522 ( .A(n11174), .B(n10322), .Z(n17016) );
  XNOR U17523 ( .A(n17017), .B(n13719), .Z(n10322) );
  NOR U17524 ( .A(n15466), .B(n13718), .Z(n17017) );
  XOR U17525 ( .A(n17018), .B(n15644), .Z(n13718) );
  XOR U17526 ( .A(n17019), .B(n17020), .Z(n15466) );
  XNOR U17527 ( .A(n17021), .B(n13714), .Z(n11174) );
  XOR U17528 ( .A(n17022), .B(n13709), .Z(n11168) );
  ANDN U17529 ( .B(n13710), .A(n15464), .Z(n17022) );
  XOR U17530 ( .A(n17023), .B(n17024), .Z(n15464) );
  XNOR U17531 ( .A(n17025), .B(n17026), .Z(n13710) );
  XOR U17532 ( .A(n17027), .B(n13715), .Z(n15458) );
  XOR U17533 ( .A(n17028), .B(n17029), .Z(n13715) );
  ANDN U17534 ( .B(n14495), .A(n14494), .Z(n17027) );
  XOR U17535 ( .A(n17030), .B(n17031), .Z(n14494) );
  XNOR U17536 ( .A(n17032), .B(n8612), .Z(n5302) );
  XNOR U17537 ( .A(n16266), .B(n10077), .Z(n8612) );
  XNOR U17538 ( .A(n15834), .B(n16658), .Z(n10077) );
  XNOR U17539 ( .A(n17033), .B(n17034), .Z(n16658) );
  XNOR U17540 ( .A(n12753), .B(n16221), .Z(n17034) );
  XNOR U17541 ( .A(n17035), .B(n16237), .Z(n16221) );
  NOR U17542 ( .A(n16236), .B(n16275), .Z(n17035) );
  XOR U17543 ( .A(n15885), .B(n17036), .Z(n16236) );
  XNOR U17544 ( .A(n17037), .B(n16228), .Z(n12753) );
  AND U17545 ( .A(n17038), .B(n16227), .Z(n17037) );
  XNOR U17546 ( .A(n12302), .B(n17039), .Z(n17033) );
  XOR U17547 ( .A(n9640), .B(n10699), .Z(n17039) );
  XOR U17548 ( .A(n17040), .B(n16232), .Z(n10699) );
  XNOR U17549 ( .A(n17041), .B(n16998), .Z(n16231) );
  XNOR U17550 ( .A(n17042), .B(n16241), .Z(n9640) );
  ANDN U17551 ( .B(n16240), .A(n17043), .Z(n17042) );
  XOR U17552 ( .A(n17044), .B(n17045), .Z(n16240) );
  XOR U17553 ( .A(n17046), .B(n16245), .Z(n12302) );
  ANDN U17554 ( .B(n16244), .A(n16268), .Z(n17046) );
  XNOR U17555 ( .A(n17047), .B(n17048), .Z(n16244) );
  XOR U17556 ( .A(n17049), .B(n17050), .Z(n15834) );
  XNOR U17557 ( .A(n17051), .B(n10154), .Z(n17050) );
  XOR U17558 ( .A(n17052), .B(n13410), .Z(n10154) );
  NOR U17559 ( .A(n17053), .B(n15095), .Z(n17052) );
  XNOR U17560 ( .A(n17054), .B(n17055), .Z(n15095) );
  XOR U17561 ( .A(n15387), .B(n17056), .Z(n17049) );
  XNOR U17562 ( .A(n9533), .B(n10358), .Z(n17056) );
  XNOR U17563 ( .A(n17057), .B(n15867), .Z(n10358) );
  ANDN U17564 ( .B(n15082), .A(n15083), .Z(n17057) );
  XOR U17565 ( .A(n17058), .B(n17059), .Z(n15083) );
  XNOR U17566 ( .A(n17060), .B(n13403), .Z(n9533) );
  NOR U17567 ( .A(n17061), .B(n15087), .Z(n17060) );
  XNOR U17568 ( .A(n17062), .B(n17063), .Z(n15087) );
  XNOR U17569 ( .A(n17064), .B(n17065), .Z(n15387) );
  AND U17570 ( .A(n15851), .B(n15852), .Z(n17064) );
  XOR U17571 ( .A(n17066), .B(n17067), .Z(n15852) );
  XNOR U17572 ( .A(n17068), .B(n16227), .Z(n16266) );
  XOR U17573 ( .A(n16313), .B(n17069), .Z(n16227) );
  NOR U17574 ( .A(n17038), .B(n17070), .Z(n17068) );
  AND U17575 ( .A(n8613), .B(n7925), .Z(n17032) );
  XNOR U17576 ( .A(n11166), .B(n17071), .Z(n7925) );
  IV U17577 ( .A(n12493), .Z(n11166) );
  XNOR U17578 ( .A(n17072), .B(n13135), .Z(n12493) );
  XOR U17579 ( .A(n17073), .B(n17074), .Z(n13135) );
  XNOR U17580 ( .A(n15245), .B(n10584), .Z(n17074) );
  XNOR U17581 ( .A(n17075), .B(n16785), .Z(n10584) );
  AND U17582 ( .A(n15975), .B(n15973), .Z(n17075) );
  XNOR U17583 ( .A(n17076), .B(n15261), .Z(n15973) );
  XNOR U17584 ( .A(n17077), .B(n17078), .Z(n15245) );
  ANDN U17585 ( .B(n15984), .A(n15982), .Z(n17077) );
  XOR U17586 ( .A(n12881), .B(n17079), .Z(n17073) );
  XNOR U17587 ( .A(n9103), .B(n9332), .Z(n17079) );
  XOR U17588 ( .A(n17080), .B(n16788), .Z(n9332) );
  NOR U17589 ( .A(n15978), .B(n15979), .Z(n17080) );
  XNOR U17590 ( .A(n16757), .B(n17081), .Z(n15978) );
  XNOR U17591 ( .A(n17082), .B(n16778), .Z(n9103) );
  AND U17592 ( .A(n15988), .B(n15986), .Z(n17082) );
  XNOR U17593 ( .A(n17083), .B(n17055), .Z(n15986) );
  XNOR U17594 ( .A(n17084), .B(n17085), .Z(n12881) );
  ANDN U17595 ( .B(n15969), .A(n15970), .Z(n17084) );
  XOR U17596 ( .A(n15956), .B(n17086), .Z(n15969) );
  XOR U17597 ( .A(n16493), .B(n17087), .Z(n8613) );
  XOR U17598 ( .A(n17088), .B(n12853), .Z(n16493) );
  XNOR U17599 ( .A(n17089), .B(n17090), .Z(n12853) );
  XNOR U17600 ( .A(n10886), .B(n13729), .Z(n17090) );
  XNOR U17601 ( .A(n17091), .B(n15984), .Z(n13729) );
  XOR U17602 ( .A(n17092), .B(n17093), .Z(n15984) );
  ANDN U17603 ( .B(n15983), .A(n17094), .Z(n17091) );
  IV U17604 ( .A(n17095), .Z(n15983) );
  XNOR U17605 ( .A(n17096), .B(n15975), .Z(n10886) );
  XNOR U17606 ( .A(n17097), .B(n17098), .Z(n15975) );
  ANDN U17607 ( .B(n15974), .A(n16784), .Z(n17096) );
  XOR U17608 ( .A(n11499), .B(n17099), .Z(n17089) );
  XOR U17609 ( .A(n10951), .B(n12526), .Z(n17099) );
  XNOR U17610 ( .A(n17100), .B(n15970), .Z(n12526) );
  XOR U17611 ( .A(n17101), .B(n17102), .Z(n15970) );
  NOR U17612 ( .A(n15971), .B(n16781), .Z(n17100) );
  XOR U17613 ( .A(n17103), .B(n15988), .Z(n10951) );
  XNOR U17614 ( .A(n17104), .B(n17105), .Z(n15988) );
  XNOR U17615 ( .A(n17106), .B(n15979), .Z(n11499) );
  XNOR U17616 ( .A(n17107), .B(n17108), .Z(n15979) );
  NOR U17617 ( .A(n15980), .B(n16787), .Z(n17106) );
  XOR U17618 ( .A(n6417), .B(n17109), .Z(n16935) );
  XNOR U17619 ( .A(n2557), .B(n8598), .Z(n17109) );
  XOR U17620 ( .A(n17110), .B(n8604), .Z(n8598) );
  XOR U17621 ( .A(n17111), .B(n9277), .Z(n8604) );
  XNOR U17622 ( .A(n14302), .B(n13385), .Z(n9277) );
  XNOR U17623 ( .A(n17112), .B(n17113), .Z(n13385) );
  XOR U17624 ( .A(n12341), .B(n11230), .Z(n17113) );
  XNOR U17625 ( .A(n17114), .B(n17115), .Z(n11230) );
  ANDN U17626 ( .B(n13102), .A(n15771), .Z(n17114) );
  IV U17627 ( .A(n17116), .Z(n15771) );
  XNOR U17628 ( .A(n17117), .B(n13107), .Z(n12341) );
  ANDN U17629 ( .B(n14374), .A(n13106), .Z(n17117) );
  XNOR U17630 ( .A(n12331), .B(n17118), .Z(n17112) );
  XNOR U17631 ( .A(n10750), .B(n10220), .Z(n17118) );
  XNOR U17632 ( .A(n17119), .B(n13110), .Z(n10220) );
  ANDN U17633 ( .B(n13111), .A(n14371), .Z(n17119) );
  XNOR U17634 ( .A(n17120), .B(n13969), .Z(n10750) );
  XOR U17635 ( .A(n17121), .B(n13114), .Z(n12331) );
  ANDN U17636 ( .B(n13115), .A(n14382), .Z(n17121) );
  XOR U17637 ( .A(n17122), .B(n17123), .Z(n14302) );
  XOR U17638 ( .A(n11857), .B(n9626), .Z(n17123) );
  XNOR U17639 ( .A(n17124), .B(n12355), .Z(n9626) );
  NOR U17640 ( .A(n15791), .B(n15792), .Z(n17124) );
  XOR U17641 ( .A(n16399), .B(n17125), .Z(n15792) );
  XOR U17642 ( .A(n17126), .B(n17001), .Z(n15791) );
  XNOR U17643 ( .A(n17127), .B(n12349), .Z(n11857) );
  IV U17644 ( .A(n17128), .Z(n12349) );
  ANDN U17645 ( .B(n15786), .A(n12348), .Z(n17127) );
  XOR U17646 ( .A(n17129), .B(n16868), .Z(n12348) );
  XOR U17647 ( .A(n17130), .B(n17131), .Z(n15786) );
  XNOR U17648 ( .A(n11625), .B(n17132), .Z(n17122) );
  XOR U17649 ( .A(n9130), .B(n10687), .Z(n17132) );
  XOR U17650 ( .A(n17133), .B(n17134), .Z(n10687) );
  NOR U17651 ( .A(n16943), .B(n15780), .Z(n17133) );
  XOR U17652 ( .A(n17135), .B(n17136), .Z(n16943) );
  XOR U17653 ( .A(n17137), .B(n17138), .Z(n9130) );
  XOR U17654 ( .A(n16313), .B(n17141), .Z(n15276) );
  XOR U17655 ( .A(n17142), .B(n12430), .Z(n11625) );
  ANDN U17656 ( .B(n12431), .A(n15777), .Z(n17142) );
  XNOR U17657 ( .A(n17143), .B(n17144), .Z(n15777) );
  XOR U17658 ( .A(n17145), .B(n17146), .Z(n12431) );
  NOR U17659 ( .A(n10510), .B(n7929), .Z(n17110) );
  XOR U17660 ( .A(n12479), .B(n11283), .Z(n7929) );
  XNOR U17661 ( .A(n15706), .B(n17147), .Z(n11283) );
  XOR U17662 ( .A(n17148), .B(n17149), .Z(n15706) );
  XNOR U17663 ( .A(n11550), .B(n12423), .Z(n17149) );
  XOR U17664 ( .A(n17150), .B(n17151), .Z(n12423) );
  ANDN U17665 ( .B(n17152), .A(n17153), .Z(n17150) );
  XOR U17666 ( .A(n17154), .B(n17155), .Z(n11550) );
  XNOR U17667 ( .A(n12261), .B(n17158), .Z(n17148) );
  XNOR U17668 ( .A(n11093), .B(n17159), .Z(n17158) );
  XNOR U17669 ( .A(n17160), .B(n17161), .Z(n11093) );
  ANDN U17670 ( .B(n17162), .A(n17163), .Z(n17160) );
  XNOR U17671 ( .A(n17164), .B(n17165), .Z(n12261) );
  NOR U17672 ( .A(n17166), .B(n17167), .Z(n17164) );
  XNOR U17673 ( .A(n17168), .B(n14354), .Z(n12479) );
  ANDN U17674 ( .B(n17169), .A(n17170), .Z(n17168) );
  XNOR U17675 ( .A(n17171), .B(n9978), .Z(n10510) );
  XNOR U17676 ( .A(n12624), .B(n13920), .Z(n9978) );
  XNOR U17677 ( .A(n17172), .B(n17173), .Z(n13920) );
  XNOR U17678 ( .A(n10930), .B(n12361), .Z(n17173) );
  XNOR U17679 ( .A(n17174), .B(n14392), .Z(n12361) );
  ANDN U17680 ( .B(n13922), .A(n13545), .Z(n17174) );
  XOR U17681 ( .A(n17175), .B(n16023), .Z(n13545) );
  XOR U17682 ( .A(n17176), .B(n17177), .Z(n13922) );
  XNOR U17683 ( .A(n17178), .B(n17179), .Z(n10930) );
  ANDN U17684 ( .B(n13067), .A(n13079), .Z(n17178) );
  XOR U17685 ( .A(n17180), .B(n17181), .Z(n13079) );
  XOR U17686 ( .A(n17182), .B(n16878), .Z(n13067) );
  XOR U17687 ( .A(n12515), .B(n17183), .Z(n17172) );
  XNOR U17688 ( .A(n9615), .B(n9762), .Z(n17183) );
  XNOR U17689 ( .A(n17184), .B(n13055), .Z(n9762) );
  AND U17690 ( .A(n13056), .B(n13089), .Z(n17184) );
  XNOR U17691 ( .A(n17185), .B(n17186), .Z(n13089) );
  XOR U17692 ( .A(n17187), .B(n17188), .Z(n13056) );
  XOR U17693 ( .A(n17189), .B(n17190), .Z(n9615) );
  ANDN U17694 ( .B(n13086), .A(n13084), .Z(n17189) );
  IV U17695 ( .A(n17191), .Z(n13084) );
  XNOR U17696 ( .A(n17192), .B(n17193), .Z(n13086) );
  XNOR U17697 ( .A(n17194), .B(n13059), .Z(n12515) );
  NOR U17698 ( .A(n13060), .B(n13298), .Z(n17194) );
  XOR U17699 ( .A(n17195), .B(n17196), .Z(n13298) );
  XOR U17700 ( .A(n17197), .B(n17198), .Z(n13060) );
  XOR U17701 ( .A(n17199), .B(n17200), .Z(n12624) );
  XOR U17702 ( .A(n10382), .B(n11483), .Z(n17200) );
  XOR U17703 ( .A(n17201), .B(n12954), .Z(n11483) );
  XNOR U17704 ( .A(n17202), .B(n17203), .Z(n12954) );
  XNOR U17705 ( .A(n17204), .B(n15292), .Z(n10382) );
  XOR U17706 ( .A(n17205), .B(n17140), .Z(n15292) );
  ANDN U17707 ( .B(n13358), .A(n15291), .Z(n17204) );
  XOR U17708 ( .A(n13049), .B(n17206), .Z(n17199) );
  XOR U17709 ( .A(n11163), .B(n10124), .Z(n17206) );
  XNOR U17710 ( .A(n17207), .B(n12799), .Z(n10124) );
  XNOR U17711 ( .A(n17208), .B(n17209), .Z(n12799) );
  NOR U17712 ( .A(n15301), .B(n13362), .Z(n17207) );
  XNOR U17713 ( .A(n17210), .B(n12805), .Z(n11163) );
  XOR U17714 ( .A(n17211), .B(n17048), .Z(n12805) );
  IV U17715 ( .A(n17212), .Z(n17048) );
  ANDN U17716 ( .B(n15287), .A(n13367), .Z(n17210) );
  XNOR U17717 ( .A(n17213), .B(n12809), .Z(n13049) );
  XNOR U17718 ( .A(n17214), .B(n17215), .Z(n12809) );
  NOR U17719 ( .A(n13369), .B(n15305), .Z(n17213) );
  XNOR U17720 ( .A(n17216), .B(n8617), .Z(n2557) );
  XNOR U17721 ( .A(n14680), .B(n9636), .Z(n8617) );
  XNOR U17722 ( .A(n17217), .B(n17218), .Z(n14680) );
  NOR U17723 ( .A(n13858), .B(n16895), .Z(n17217) );
  XOR U17724 ( .A(n17219), .B(n16056), .Z(n13858) );
  NOR U17725 ( .A(n16905), .B(n10534), .Z(n17216) );
  XOR U17726 ( .A(n11584), .B(n13567), .Z(n10534) );
  XNOR U17727 ( .A(n17220), .B(n17221), .Z(n13567) );
  NOR U17728 ( .A(n14231), .B(n14230), .Z(n17220) );
  IV U17729 ( .A(n15056), .Z(n11584) );
  XNOR U17730 ( .A(n17222), .B(n14758), .Z(n15056) );
  XOR U17731 ( .A(n17223), .B(n17224), .Z(n14758) );
  XNOR U17732 ( .A(n13463), .B(n14264), .Z(n17224) );
  XOR U17733 ( .A(n17225), .B(n14275), .Z(n14264) );
  ANDN U17734 ( .B(n13564), .A(n13565), .Z(n17225) );
  XOR U17735 ( .A(n17226), .B(n17227), .Z(n13565) );
  XOR U17736 ( .A(n17230), .B(n16861), .Z(n13463) );
  NOR U17737 ( .A(n14227), .B(n13571), .Z(n17230) );
  XOR U17738 ( .A(n17231), .B(n17232), .Z(n13571) );
  IV U17739 ( .A(n13573), .Z(n14227) );
  XOR U17740 ( .A(n17233), .B(n17234), .Z(n13573) );
  XOR U17741 ( .A(n13471), .B(n17235), .Z(n17223) );
  XNOR U17742 ( .A(n12639), .B(n11959), .Z(n17235) );
  XOR U17743 ( .A(n17236), .B(n14671), .Z(n11959) );
  ANDN U17744 ( .B(n13561), .A(n13560), .Z(n17236) );
  XNOR U17745 ( .A(n17237), .B(n17238), .Z(n13560) );
  XOR U17746 ( .A(n17239), .B(n17240), .Z(n13561) );
  XOR U17747 ( .A(n17241), .B(n17242), .Z(n12639) );
  ANDN U17748 ( .B(n14230), .A(n17221), .Z(n17241) );
  XOR U17749 ( .A(n17243), .B(n17244), .Z(n14230) );
  XOR U17750 ( .A(n17245), .B(n14273), .Z(n13471) );
  ANDN U17751 ( .B(n14218), .A(n14272), .Z(n17245) );
  XNOR U17752 ( .A(n17246), .B(n17247), .Z(n14272) );
  XNOR U17753 ( .A(n17248), .B(n17249), .Z(n14218) );
  XOR U17754 ( .A(n10214), .B(n14703), .Z(n16905) );
  XOR U17755 ( .A(n17250), .B(n17251), .Z(n14703) );
  AND U17756 ( .A(n15132), .B(n15134), .Z(n17250) );
  IV U17757 ( .A(n11294), .Z(n10214) );
  XOR U17758 ( .A(n12605), .B(n17252), .Z(n11294) );
  XOR U17759 ( .A(n17253), .B(n17254), .Z(n12605) );
  XNOR U17760 ( .A(n12224), .B(n9656), .Z(n17254) );
  XOR U17761 ( .A(n17255), .B(n17256), .Z(n9656) );
  XOR U17762 ( .A(n17257), .B(n16527), .Z(n14708) );
  XOR U17763 ( .A(n17258), .B(n17259), .Z(n12224) );
  AND U17764 ( .A(n14712), .B(n14710), .Z(n17258) );
  XNOR U17765 ( .A(n17260), .B(n17261), .Z(n14712) );
  XNOR U17766 ( .A(n14184), .B(n17262), .Z(n17253) );
  XOR U17767 ( .A(n13801), .B(n9807), .Z(n17262) );
  XOR U17768 ( .A(n17263), .B(n17264), .Z(n9807) );
  XNOR U17769 ( .A(n17265), .B(n15342), .Z(n14702) );
  XOR U17770 ( .A(n17266), .B(n17267), .Z(n13801) );
  NOR U17771 ( .A(n14696), .B(n14697), .Z(n17266) );
  XOR U17772 ( .A(n17268), .B(n17269), .Z(n14697) );
  XNOR U17773 ( .A(n17270), .B(n17271), .Z(n14184) );
  ANDN U17774 ( .B(n17251), .A(n15132), .Z(n17270) );
  XOR U17775 ( .A(n17272), .B(n17273), .Z(n15132) );
  XNOR U17776 ( .A(n17274), .B(n8608), .Z(n6417) );
  XOR U17777 ( .A(n10359), .B(n17051), .Z(n8608) );
  XNOR U17778 ( .A(n17275), .B(n13414), .Z(n17051) );
  NOR U17779 ( .A(n15091), .B(n15092), .Z(n17275) );
  XNOR U17780 ( .A(n17276), .B(n17277), .Z(n15092) );
  XNOR U17781 ( .A(n13796), .B(n16222), .Z(n10359) );
  XOR U17782 ( .A(n17278), .B(n17279), .Z(n16222) );
  XNOR U17783 ( .A(n10529), .B(n11186), .Z(n17279) );
  XOR U17784 ( .A(n17280), .B(n13409), .Z(n11186) );
  XOR U17785 ( .A(n17281), .B(n17282), .Z(n13409) );
  ANDN U17786 ( .B(n13410), .A(n15094), .Z(n17280) );
  IV U17787 ( .A(n17053), .Z(n15094) );
  XOR U17788 ( .A(n17283), .B(n16737), .Z(n17053) );
  XOR U17789 ( .A(n17284), .B(n17285), .Z(n13410) );
  XNOR U17790 ( .A(n17286), .B(n13413), .Z(n10529) );
  XOR U17791 ( .A(n17287), .B(n17288), .Z(n13413) );
  XOR U17792 ( .A(n17289), .B(n17093), .Z(n13414) );
  XOR U17793 ( .A(n15674), .B(n17290), .Z(n15091) );
  XNOR U17794 ( .A(n10181), .B(n17291), .Z(n17278) );
  XNOR U17795 ( .A(n13393), .B(n11820), .Z(n17291) );
  XOR U17796 ( .A(n17292), .B(n13400), .Z(n11820) );
  XOR U17797 ( .A(n17293), .B(n17294), .Z(n13400) );
  ANDN U17798 ( .B(n13399), .A(n15851), .Z(n17292) );
  XOR U17799 ( .A(n17295), .B(n15698), .Z(n15851) );
  IV U17800 ( .A(n17065), .Z(n13399) );
  XOR U17801 ( .A(n17296), .B(n17297), .Z(n17065) );
  XNOR U17802 ( .A(n17298), .B(n15868), .Z(n13393) );
  XNOR U17803 ( .A(n17299), .B(n16103), .Z(n15868) );
  ANDN U17804 ( .B(n15867), .A(n15082), .Z(n17298) );
  XOR U17805 ( .A(n17300), .B(n17301), .Z(n15082) );
  XOR U17806 ( .A(n17302), .B(n17303), .Z(n15867) );
  XOR U17807 ( .A(n17304), .B(n13404), .Z(n10181) );
  XOR U17808 ( .A(n17305), .B(n17306), .Z(n13404) );
  NOR U17809 ( .A(n15086), .B(n13403), .Z(n17304) );
  XOR U17810 ( .A(n17307), .B(n17131), .Z(n13403) );
  IV U17811 ( .A(n17061), .Z(n15086) );
  XOR U17812 ( .A(n17308), .B(n16589), .Z(n17061) );
  XOR U17813 ( .A(n17309), .B(n17310), .Z(n13796) );
  XOR U17814 ( .A(n10487), .B(n10988), .Z(n17310) );
  XOR U17815 ( .A(n17311), .B(n15905), .Z(n10988) );
  ANDN U17816 ( .B(n15843), .A(n15844), .Z(n17311) );
  XOR U17817 ( .A(n17312), .B(n16331), .Z(n15844) );
  XNOR U17818 ( .A(n17313), .B(n15908), .Z(n10487) );
  ANDN U17819 ( .B(n13984), .A(n17314), .Z(n17313) );
  XNOR U17820 ( .A(n17315), .B(n16101), .Z(n13984) );
  XOR U17821 ( .A(n10882), .B(n17316), .Z(n17309) );
  XOR U17822 ( .A(n9146), .B(n17317), .Z(n17316) );
  XOR U17823 ( .A(n17318), .B(n15900), .Z(n9146) );
  NOR U17824 ( .A(n13980), .B(n15846), .Z(n17318) );
  IV U17825 ( .A(n15847), .Z(n13980) );
  XNOR U17826 ( .A(n17195), .B(n17319), .Z(n15847) );
  XNOR U17827 ( .A(n17320), .B(n15895), .Z(n10882) );
  ANDN U17828 ( .B(n15838), .A(n13997), .Z(n17320) );
  XNOR U17829 ( .A(n17321), .B(n17322), .Z(n13997) );
  ANDN U17830 ( .B(n7920), .A(n8609), .Z(n17274) );
  XOR U17831 ( .A(n16874), .B(n9535), .Z(n8609) );
  IV U17832 ( .A(n11466), .Z(n9535) );
  XOR U17833 ( .A(n16160), .B(n16177), .Z(n11466) );
  XOR U17834 ( .A(n17323), .B(n17324), .Z(n16177) );
  XNOR U17835 ( .A(n10820), .B(n17325), .Z(n17324) );
  XNOR U17836 ( .A(n17326), .B(n15004), .Z(n10820) );
  ANDN U17837 ( .B(n17327), .A(n16355), .Z(n17326) );
  IV U17838 ( .A(n17328), .Z(n16355) );
  XNOR U17839 ( .A(n10979), .B(n17329), .Z(n17323) );
  XOR U17840 ( .A(n11000), .B(n11802), .Z(n17329) );
  XNOR U17841 ( .A(n17330), .B(n14793), .Z(n11802) );
  NOR U17842 ( .A(n17331), .B(n16362), .Z(n17330) );
  XNOR U17843 ( .A(n17332), .B(n17333), .Z(n16362) );
  XOR U17844 ( .A(n17334), .B(n14804), .Z(n11000) );
  AND U17845 ( .A(n16866), .B(n16357), .Z(n17334) );
  XOR U17846 ( .A(n17335), .B(n17336), .Z(n16357) );
  XOR U17847 ( .A(n17337), .B(n16337), .Z(n10979) );
  NOR U17848 ( .A(n16880), .B(n16881), .Z(n17337) );
  XNOR U17849 ( .A(n17338), .B(n17339), .Z(n16881) );
  XOR U17850 ( .A(n17340), .B(n17341), .Z(n16160) );
  XOR U17851 ( .A(n12651), .B(n13120), .Z(n17341) );
  XNOR U17852 ( .A(n17342), .B(n12045), .Z(n13120) );
  ANDN U17853 ( .B(n17343), .A(n16341), .Z(n17342) );
  XNOR U17854 ( .A(n17344), .B(n12028), .Z(n12651) );
  NOR U17855 ( .A(n17345), .B(n17346), .Z(n17344) );
  XNOR U17856 ( .A(n12987), .B(n17347), .Z(n17340) );
  XNOR U17857 ( .A(n16249), .B(n16204), .Z(n17347) );
  XNOR U17858 ( .A(n17348), .B(n12041), .Z(n16204) );
  NOR U17859 ( .A(n16349), .B(n17349), .Z(n17348) );
  XNOR U17860 ( .A(n17350), .B(n12037), .Z(n16249) );
  ANDN U17861 ( .B(n16344), .A(n17351), .Z(n17350) );
  XNOR U17862 ( .A(n17352), .B(n12032), .Z(n12987) );
  XNOR U17863 ( .A(n17354), .B(n17327), .Z(n16874) );
  NOR U17864 ( .A(n17328), .B(n15003), .Z(n17354) );
  XNOR U17865 ( .A(n17355), .B(n16848), .Z(n15003) );
  XOR U17866 ( .A(n17356), .B(n16739), .Z(n17328) );
  XOR U17867 ( .A(n15752), .B(n11754), .Z(n7920) );
  XNOR U17868 ( .A(n17357), .B(n15215), .Z(n15752) );
  ANDN U17869 ( .B(n15749), .A(n15748), .Z(n17357) );
  XOR U17870 ( .A(n17358), .B(n17359), .Z(n8045) );
  XNOR U17871 ( .A(n4955), .B(n10612), .Z(n17359) );
  XOR U17872 ( .A(n17360), .B(n6981), .Z(n10612) );
  XOR U17873 ( .A(n14287), .B(n10172), .Z(n6981) );
  IV U17874 ( .A(n11722), .Z(n10172) );
  XNOR U17875 ( .A(n17363), .B(n15113), .Z(n14287) );
  NOR U17876 ( .A(n16652), .B(n17364), .Z(n17363) );
  AND U17877 ( .A(n10531), .B(n9364), .Z(n17360) );
  XNOR U17878 ( .A(n14011), .B(n9773), .Z(n9364) );
  XOR U17879 ( .A(n13286), .B(n16533), .Z(n9773) );
  XNOR U17880 ( .A(n17365), .B(n17366), .Z(n16533) );
  XOR U17881 ( .A(n17367), .B(n11197), .Z(n17366) );
  XNOR U17882 ( .A(n17368), .B(n17369), .Z(n11197) );
  NOR U17883 ( .A(n17370), .B(n17371), .Z(n17368) );
  XOR U17884 ( .A(n11073), .B(n17372), .Z(n17365) );
  XNOR U17885 ( .A(n10691), .B(n10201), .Z(n17372) );
  XNOR U17886 ( .A(n17373), .B(n17374), .Z(n10201) );
  ANDN U17887 ( .B(n17375), .A(n17376), .Z(n17373) );
  XOR U17888 ( .A(n17377), .B(n17378), .Z(n10691) );
  AND U17889 ( .A(n17379), .B(n17380), .Z(n17377) );
  XNOR U17890 ( .A(n17381), .B(n17382), .Z(n11073) );
  ANDN U17891 ( .B(n17383), .A(n17384), .Z(n17381) );
  XOR U17892 ( .A(n17385), .B(n17386), .Z(n13286) );
  XOR U17893 ( .A(n11774), .B(n11420), .Z(n17386) );
  XNOR U17894 ( .A(n17387), .B(n17388), .Z(n11420) );
  NOR U17895 ( .A(n14610), .B(n14003), .Z(n17387) );
  XNOR U17896 ( .A(n17389), .B(n17390), .Z(n14003) );
  IV U17897 ( .A(n14004), .Z(n14610) );
  XOR U17898 ( .A(n17391), .B(n17392), .Z(n14004) );
  XNOR U17899 ( .A(n17393), .B(n16980), .Z(n11774) );
  ANDN U17900 ( .B(n14009), .A(n14007), .Z(n17393) );
  XNOR U17901 ( .A(n17396), .B(n15650), .Z(n14009) );
  XOR U17902 ( .A(n16968), .B(n17397), .Z(n17385) );
  XNOR U17903 ( .A(n14896), .B(n10961), .Z(n17397) );
  XOR U17904 ( .A(n17398), .B(n16973), .Z(n10961) );
  ANDN U17905 ( .B(n14013), .A(n14014), .Z(n17398) );
  IV U17906 ( .A(n14606), .Z(n14014) );
  XOR U17907 ( .A(n17399), .B(n17400), .Z(n14606) );
  XOR U17908 ( .A(n17401), .B(n17402), .Z(n14013) );
  XOR U17909 ( .A(n17403), .B(n17404), .Z(n14896) );
  ANDN U17910 ( .B(n14596), .A(n17405), .Z(n17403) );
  XOR U17911 ( .A(n17406), .B(n16976), .Z(n16968) );
  NOR U17912 ( .A(n14018), .B(n14017), .Z(n17406) );
  XOR U17913 ( .A(n17407), .B(n15201), .Z(n14017) );
  XOR U17914 ( .A(n17408), .B(n17212), .Z(n14018) );
  XNOR U17915 ( .A(n17409), .B(n17405), .Z(n14011) );
  NOR U17916 ( .A(n14597), .B(n14596), .Z(n17409) );
  XOR U17917 ( .A(n16603), .B(n17410), .Z(n14596) );
  XOR U17918 ( .A(n17411), .B(n10714), .Z(n10531) );
  IV U17919 ( .A(n16703), .Z(n10714) );
  XNOR U17920 ( .A(n17072), .B(n15442), .Z(n16703) );
  XNOR U17921 ( .A(n17412), .B(n17413), .Z(n15442) );
  XOR U17922 ( .A(n11160), .B(n12648), .Z(n17413) );
  XOR U17923 ( .A(n17414), .B(n16438), .Z(n12648) );
  ANDN U17924 ( .B(n16439), .A(n16929), .Z(n17414) );
  XNOR U17925 ( .A(n17415), .B(n16425), .Z(n11160) );
  ANDN U17926 ( .B(n16921), .A(n17416), .Z(n17415) );
  XOR U17927 ( .A(n10405), .B(n17417), .Z(n17412) );
  XNOR U17928 ( .A(n12201), .B(n10884), .Z(n17417) );
  XNOR U17929 ( .A(n17418), .B(n16431), .Z(n10884) );
  ANDN U17930 ( .B(n16430), .A(n16924), .Z(n17418) );
  IV U17931 ( .A(n17419), .Z(n16924) );
  IV U17932 ( .A(n17420), .Z(n16430) );
  XOR U17933 ( .A(n17421), .B(n16421), .Z(n12201) );
  ANDN U17934 ( .B(n16422), .A(n17422), .Z(n17421) );
  XNOR U17935 ( .A(n17423), .B(n16435), .Z(n10405) );
  NOR U17936 ( .A(n17424), .B(n16933), .Z(n17423) );
  XOR U17937 ( .A(n17425), .B(n17426), .Z(n17072) );
  XOR U17938 ( .A(n11691), .B(n14672), .Z(n17426) );
  XOR U17939 ( .A(n17427), .B(n16288), .Z(n14672) );
  XNOR U17940 ( .A(n17428), .B(n17429), .Z(n16288) );
  NOR U17941 ( .A(n15990), .B(n16759), .Z(n17427) );
  XNOR U17942 ( .A(n17430), .B(n16291), .Z(n11691) );
  XNOR U17943 ( .A(n17431), .B(n17432), .Z(n16291) );
  NOR U17944 ( .A(n16764), .B(n14385), .Z(n17430) );
  XNOR U17945 ( .A(n10320), .B(n17433), .Z(n17425) );
  XOR U17946 ( .A(n10179), .B(n16749), .Z(n17433) );
  XNOR U17947 ( .A(n17434), .B(n16286), .Z(n16749) );
  XOR U17948 ( .A(n17435), .B(n17436), .Z(n16286) );
  XNOR U17949 ( .A(n17438), .B(n16293), .Z(n10179) );
  XNOR U17950 ( .A(n17439), .B(n17440), .Z(n16293) );
  NOR U17951 ( .A(n16772), .B(n12858), .Z(n17438) );
  XOR U17952 ( .A(n17441), .B(n16295), .Z(n10320) );
  XNOR U17953 ( .A(n17442), .B(n16068), .Z(n16295) );
  NOR U17954 ( .A(n12868), .B(n16755), .Z(n17441) );
  XNOR U17955 ( .A(n17443), .B(n6985), .Z(n4955) );
  IV U17956 ( .A(n10623), .Z(n6985) );
  XOR U17957 ( .A(n15230), .B(n11101), .Z(n10623) );
  IV U17958 ( .A(n10122), .Z(n11101) );
  XNOR U17959 ( .A(n15773), .B(n12816), .Z(n10122) );
  XNOR U17960 ( .A(n17444), .B(n17445), .Z(n12816) );
  XNOR U17961 ( .A(n13383), .B(n11909), .Z(n17445) );
  XNOR U17962 ( .A(n17447), .B(n15256), .Z(n14069) );
  NOR U17963 ( .A(n15242), .B(n15244), .Z(n17446) );
  IV U17964 ( .A(n14070), .Z(n15242) );
  XNOR U17965 ( .A(n16071), .B(n17448), .Z(n14070) );
  XOR U17966 ( .A(n17449), .B(n14073), .Z(n13383) );
  XNOR U17967 ( .A(n17450), .B(n17451), .Z(n14073) );
  XOR U17968 ( .A(n10066), .B(n17453), .Z(n17444) );
  XOR U17969 ( .A(n12100), .B(n11873), .Z(n17453) );
  XNOR U17970 ( .A(n17454), .B(n14079), .Z(n11873) );
  XOR U17971 ( .A(n17455), .B(n16404), .Z(n14079) );
  NOR U17972 ( .A(n14078), .B(n15232), .Z(n17454) );
  XOR U17973 ( .A(n17456), .B(n17457), .Z(n14078) );
  XNOR U17974 ( .A(n17458), .B(n14083), .Z(n12100) );
  XNOR U17975 ( .A(n17459), .B(n16616), .Z(n14083) );
  NOR U17976 ( .A(n14082), .B(n15239), .Z(n17458) );
  XOR U17977 ( .A(n16757), .B(n17460), .Z(n14082) );
  XNOR U17978 ( .A(n17461), .B(n14087), .Z(n10066) );
  NOR U17979 ( .A(n14086), .B(n15237), .Z(n17461) );
  XOR U17980 ( .A(n17462), .B(n17463), .Z(n14086) );
  XOR U17981 ( .A(n17464), .B(n17465), .Z(n15773) );
  XOR U17982 ( .A(n15270), .B(n17111), .Z(n17465) );
  XOR U17983 ( .A(n17466), .B(n13111), .Z(n17111) );
  XOR U17984 ( .A(n17467), .B(n17468), .Z(n13111) );
  ANDN U17985 ( .B(n14371), .A(n14372), .Z(n17466) );
  XOR U17986 ( .A(n17469), .B(n17470), .Z(n14371) );
  XOR U17987 ( .A(n17471), .B(n13102), .Z(n15270) );
  XNOR U17988 ( .A(n17472), .B(n17473), .Z(n13102) );
  ANDN U17989 ( .B(n15772), .A(n17116), .Z(n17471) );
  XOR U17990 ( .A(n17474), .B(n17475), .Z(n17116) );
  XOR U17991 ( .A(n11362), .B(n17476), .Z(n17464) );
  XNOR U17992 ( .A(n12258), .B(n9276), .Z(n17476) );
  XOR U17993 ( .A(n17477), .B(n13970), .Z(n9276) );
  XOR U17994 ( .A(n17478), .B(n17479), .Z(n13970) );
  ANDN U17995 ( .B(n14379), .A(n14380), .Z(n17477) );
  XOR U17996 ( .A(n17480), .B(n16094), .Z(n14379) );
  XOR U17997 ( .A(n17481), .B(n13106), .Z(n12258) );
  XNOR U17998 ( .A(n17482), .B(n16620), .Z(n13106) );
  NOR U17999 ( .A(n14375), .B(n14374), .Z(n17481) );
  XNOR U18000 ( .A(n17483), .B(n17484), .Z(n14374) );
  XOR U18001 ( .A(n17485), .B(n13115), .Z(n11362) );
  XOR U18002 ( .A(n17486), .B(n17487), .Z(n13115) );
  ANDN U18003 ( .B(n14382), .A(n14383), .Z(n17485) );
  IV U18004 ( .A(n17488), .Z(n14383) );
  XNOR U18005 ( .A(n17489), .B(n15196), .Z(n14382) );
  XOR U18006 ( .A(n17490), .B(n14074), .Z(n15230) );
  XOR U18007 ( .A(n17491), .B(n14989), .Z(n14074) );
  IV U18008 ( .A(n17009), .Z(n14989) );
  ANDN U18009 ( .B(n15768), .A(n17452), .Z(n17490) );
  ANDN U18010 ( .B(n10516), .A(n9358), .Z(n17443) );
  XNOR U18011 ( .A(n16469), .B(n13069), .Z(n9358) );
  XOR U18012 ( .A(n13738), .B(n17492), .Z(n13069) );
  XOR U18013 ( .A(n17493), .B(n17494), .Z(n13738) );
  XNOR U18014 ( .A(n11936), .B(n14488), .Z(n17494) );
  XOR U18015 ( .A(n17495), .B(n14502), .Z(n14488) );
  XNOR U18016 ( .A(n16390), .B(n17496), .Z(n14502) );
  AND U18017 ( .A(n13709), .B(n13708), .Z(n17495) );
  XOR U18018 ( .A(n17497), .B(n17498), .Z(n13708) );
  XOR U18019 ( .A(n17499), .B(n17500), .Z(n13709) );
  XOR U18020 ( .A(n17501), .B(n14505), .Z(n11936) );
  XOR U18021 ( .A(n17502), .B(n17503), .Z(n14505) );
  AND U18022 ( .A(n13735), .B(n13736), .Z(n17501) );
  XOR U18023 ( .A(n17504), .B(n17294), .Z(n13736) );
  XOR U18024 ( .A(n17505), .B(n17506), .Z(n13735) );
  XNOR U18025 ( .A(n13241), .B(n17507), .Z(n17493) );
  XNOR U18026 ( .A(n13352), .B(n14393), .Z(n17507) );
  XNOR U18027 ( .A(n17508), .B(n15460), .Z(n14393) );
  XOR U18028 ( .A(n17509), .B(n15537), .Z(n15460) );
  ANDN U18029 ( .B(n13723), .A(n13721), .Z(n17508) );
  XNOR U18030 ( .A(n17510), .B(n16103), .Z(n13721) );
  XOR U18031 ( .A(n17511), .B(n16058), .Z(n13723) );
  XNOR U18032 ( .A(n17512), .B(n14499), .Z(n13352) );
  XNOR U18033 ( .A(n17513), .B(n17514), .Z(n14499) );
  AND U18034 ( .A(n13717), .B(n13719), .Z(n17512) );
  XOR U18035 ( .A(n17515), .B(n17516), .Z(n13719) );
  XOR U18036 ( .A(n17517), .B(n16531), .Z(n13717) );
  XOR U18037 ( .A(n17518), .B(n14495), .Z(n13241) );
  XOR U18038 ( .A(n17519), .B(n17520), .Z(n14495) );
  ANDN U18039 ( .B(n13713), .A(n13714), .Z(n17518) );
  XOR U18040 ( .A(n17521), .B(n16998), .Z(n13714) );
  XOR U18041 ( .A(n17522), .B(n17523), .Z(n13713) );
  XNOR U18042 ( .A(n17524), .B(n15546), .Z(n16469) );
  ANDN U18043 ( .B(n13212), .A(n14665), .Z(n17524) );
  XNOR U18044 ( .A(n15956), .B(n17525), .Z(n13212) );
  XOR U18045 ( .A(n13600), .B(n9322), .Z(n10516) );
  XNOR U18046 ( .A(n11962), .B(n17147), .Z(n9322) );
  XNOR U18047 ( .A(n17526), .B(n17527), .Z(n17147) );
  XNOR U18048 ( .A(n11639), .B(n12739), .Z(n17527) );
  XNOR U18049 ( .A(n17528), .B(n17529), .Z(n12739) );
  NOR U18050 ( .A(n17530), .B(n12473), .Z(n17528) );
  XNOR U18051 ( .A(n17531), .B(n14361), .Z(n11639) );
  ANDN U18052 ( .B(n12478), .A(n12476), .Z(n17531) );
  XNOR U18053 ( .A(n17532), .B(n17533), .Z(n12476) );
  XOR U18054 ( .A(n12061), .B(n17534), .Z(n17526) );
  XNOR U18055 ( .A(n9545), .B(n11365), .Z(n17534) );
  XNOR U18056 ( .A(n17535), .B(n14355), .Z(n11365) );
  ANDN U18057 ( .B(n14354), .A(n17169), .Z(n17535) );
  XOR U18058 ( .A(n17197), .B(n17536), .Z(n14354) );
  XOR U18059 ( .A(n17537), .B(n17538), .Z(n9545) );
  NOR U18060 ( .A(n12487), .B(n12486), .Z(n17537) );
  XNOR U18061 ( .A(n17539), .B(n14351), .Z(n12061) );
  NOR U18062 ( .A(n12483), .B(n12482), .Z(n17539) );
  XNOR U18063 ( .A(n17540), .B(n17541), .Z(n12482) );
  XOR U18064 ( .A(n17542), .B(n17543), .Z(n11962) );
  XNOR U18065 ( .A(n13156), .B(n14327), .Z(n17543) );
  XOR U18066 ( .A(n17544), .B(n14345), .Z(n14327) );
  NOR U18067 ( .A(n13611), .B(n12540), .Z(n17544) );
  XOR U18068 ( .A(n17545), .B(n17546), .Z(n12540) );
  IV U18069 ( .A(n14346), .Z(n13611) );
  XOR U18070 ( .A(n17547), .B(n17548), .Z(n14346) );
  XNOR U18071 ( .A(n17549), .B(n14331), .Z(n13156) );
  ANDN U18072 ( .B(n12549), .A(n14332), .Z(n17549) );
  XOR U18073 ( .A(n17550), .B(n15698), .Z(n14332) );
  XNOR U18074 ( .A(n17551), .B(n17552), .Z(n12549) );
  XOR U18075 ( .A(n13975), .B(n17553), .Z(n17542) );
  XOR U18076 ( .A(n9239), .B(n12572), .Z(n17553) );
  XOR U18077 ( .A(n17554), .B(n14339), .Z(n12572) );
  ANDN U18078 ( .B(n13607), .A(n13606), .Z(n17554) );
  XOR U18079 ( .A(n17555), .B(n17390), .Z(n13606) );
  IV U18080 ( .A(n12536), .Z(n13607) );
  XOR U18081 ( .A(n17556), .B(n17261), .Z(n12536) );
  XOR U18082 ( .A(n17557), .B(n14342), .Z(n9239) );
  NOR U18083 ( .A(n17558), .B(n12545), .Z(n17557) );
  XNOR U18084 ( .A(n17559), .B(n14335), .Z(n13975) );
  ANDN U18085 ( .B(n13602), .A(n12553), .Z(n17559) );
  XNOR U18086 ( .A(n17560), .B(n15679), .Z(n12553) );
  XOR U18087 ( .A(n17561), .B(n17470), .Z(n13602) );
  XNOR U18088 ( .A(n17562), .B(n14341), .Z(n13600) );
  IV U18089 ( .A(n17558), .Z(n14341) );
  XNOR U18090 ( .A(n17563), .B(n17564), .Z(n17558) );
  AND U18091 ( .A(n12547), .B(n12545), .Z(n17562) );
  XOR U18092 ( .A(n17565), .B(n16813), .Z(n12545) );
  XNOR U18093 ( .A(n2654), .B(n17566), .Z(n17358) );
  XNOR U18094 ( .A(n3569), .B(n5757), .Z(n17566) );
  XOR U18095 ( .A(n17567), .B(n10627), .Z(n5757) );
  IV U18096 ( .A(n6976), .Z(n10627) );
  XOR U18097 ( .A(n16775), .B(n12706), .Z(n6976) );
  IV U18098 ( .A(n11891), .Z(n12706) );
  XOR U18099 ( .A(n13646), .B(n16282), .Z(n11891) );
  XNOR U18100 ( .A(n17568), .B(n17569), .Z(n16282) );
  XNOR U18101 ( .A(n12046), .B(n16621), .Z(n17569) );
  XOR U18102 ( .A(n17570), .B(n15987), .Z(n16621) );
  XOR U18103 ( .A(n17571), .B(n17572), .Z(n15987) );
  ANDN U18104 ( .B(n16778), .A(n16777), .Z(n17570) );
  XOR U18105 ( .A(n17573), .B(n17574), .Z(n16777) );
  XNOR U18106 ( .A(n17575), .B(n16996), .Z(n16778) );
  XNOR U18107 ( .A(n17576), .B(n17095), .Z(n12046) );
  XNOR U18108 ( .A(n17577), .B(n17578), .Z(n17095) );
  AND U18109 ( .A(n17094), .B(n17078), .Z(n17576) );
  XOR U18110 ( .A(n17087), .B(n17579), .Z(n17568) );
  XNOR U18111 ( .A(n16492), .B(n10318), .Z(n17579) );
  XOR U18112 ( .A(n17580), .B(n15974), .Z(n10318) );
  XOR U18113 ( .A(n17581), .B(n16892), .Z(n15974) );
  AND U18114 ( .A(n16785), .B(n16784), .Z(n17580) );
  XNOR U18115 ( .A(n17582), .B(n17533), .Z(n16784) );
  XOR U18116 ( .A(n17583), .B(n16412), .Z(n16785) );
  XNOR U18117 ( .A(n17584), .B(n15971), .Z(n16492) );
  XNOR U18118 ( .A(n17585), .B(n17586), .Z(n15971) );
  ANDN U18119 ( .B(n16781), .A(n16782), .Z(n17584) );
  IV U18120 ( .A(n17085), .Z(n16782) );
  XNOR U18121 ( .A(n17587), .B(n17564), .Z(n17085) );
  XOR U18122 ( .A(n17588), .B(n17589), .Z(n16781) );
  XNOR U18123 ( .A(n17590), .B(n15980), .Z(n17087) );
  XOR U18124 ( .A(n17591), .B(n17592), .Z(n15980) );
  ANDN U18125 ( .B(n16787), .A(n16788), .Z(n17590) );
  XOR U18126 ( .A(n17593), .B(n15269), .Z(n16788) );
  XNOR U18127 ( .A(n16961), .B(n17594), .Z(n16787) );
  XOR U18128 ( .A(n17595), .B(n17596), .Z(n13646) );
  XNOR U18129 ( .A(n17597), .B(n11834), .Z(n17596) );
  XOR U18130 ( .A(n17598), .B(n13962), .Z(n11834) );
  ANDN U18131 ( .B(n13145), .A(n17599), .Z(n17598) );
  XNOR U18132 ( .A(n17600), .B(n17601), .Z(n13145) );
  XOR U18133 ( .A(n13162), .B(n17602), .Z(n17595) );
  XNOR U18134 ( .A(n10064), .B(n17603), .Z(n17602) );
  XNOR U18135 ( .A(n17604), .B(n13957), .Z(n10064) );
  ANDN U18136 ( .B(n14512), .A(n15263), .Z(n17604) );
  XOR U18137 ( .A(n17605), .B(n17606), .Z(n14512) );
  XNOR U18138 ( .A(n17607), .B(n13960), .Z(n13162) );
  ANDN U18139 ( .B(n15267), .A(n13149), .Z(n17607) );
  XOR U18140 ( .A(n17608), .B(n17479), .Z(n13149) );
  XNOR U18141 ( .A(n17609), .B(n17094), .Z(n16775) );
  XOR U18142 ( .A(n17610), .B(n14996), .Z(n17094) );
  XOR U18143 ( .A(n14158), .B(n17611), .Z(n17078) );
  XOR U18144 ( .A(n17612), .B(n17613), .Z(n15982) );
  ANDN U18145 ( .B(n9361), .A(n10528), .Z(n17567) );
  XOR U18146 ( .A(n10095), .B(n14530), .Z(n10528) );
  XNOR U18147 ( .A(n17614), .B(n16325), .Z(n14530) );
  AND U18148 ( .A(n17615), .B(n15565), .Z(n17614) );
  XNOR U18149 ( .A(n16027), .B(n15588), .Z(n10095) );
  XOR U18150 ( .A(n17616), .B(n17617), .Z(n15588) );
  XNOR U18151 ( .A(n16296), .B(n11804), .Z(n17617) );
  XOR U18152 ( .A(n17618), .B(n15562), .Z(n11804) );
  XNOR U18153 ( .A(n17619), .B(n17620), .Z(n15562) );
  NOR U18154 ( .A(n14533), .B(n14532), .Z(n17618) );
  XOR U18155 ( .A(n17621), .B(n17622), .Z(n14532) );
  XNOR U18156 ( .A(n17623), .B(n15558), .Z(n16296) );
  XNOR U18157 ( .A(n17456), .B(n17624), .Z(n15558) );
  AND U18158 ( .A(n14528), .B(n14526), .Z(n17623) );
  XNOR U18159 ( .A(n17625), .B(n17626), .Z(n14526) );
  XOR U18160 ( .A(n13123), .B(n17627), .Z(n17616) );
  XNOR U18161 ( .A(n11358), .B(n10728), .Z(n17627) );
  XNOR U18162 ( .A(n17628), .B(n15554), .Z(n10728) );
  XNOR U18163 ( .A(n17629), .B(n17630), .Z(n15554) );
  NOR U18164 ( .A(n14524), .B(n14522), .Z(n17628) );
  XNOR U18165 ( .A(n17631), .B(n17632), .Z(n14522) );
  XOR U18166 ( .A(n17633), .B(n16326), .Z(n11358) );
  XNOR U18167 ( .A(n15962), .B(n17634), .Z(n16326) );
  NOR U18168 ( .A(n17615), .B(n16325), .Z(n17633) );
  XNOR U18169 ( .A(n17635), .B(n17636), .Z(n16325) );
  XOR U18170 ( .A(n17637), .B(n15551), .Z(n13123) );
  XOR U18171 ( .A(n17638), .B(n16119), .Z(n15551) );
  NOR U18172 ( .A(n17639), .B(n14536), .Z(n17637) );
  XOR U18173 ( .A(n17640), .B(n17641), .Z(n14536) );
  XOR U18174 ( .A(n17642), .B(n17643), .Z(n16027) );
  XOR U18175 ( .A(n12841), .B(n9955), .Z(n17643) );
  XOR U18176 ( .A(n17644), .B(n15584), .Z(n9955) );
  XOR U18177 ( .A(n17645), .B(n17646), .Z(n15584) );
  ANDN U18178 ( .B(n15074), .A(n16302), .Z(n17644) );
  XOR U18179 ( .A(n17647), .B(n17648), .Z(n16302) );
  XNOR U18180 ( .A(n15879), .B(n17649), .Z(n15074) );
  XOR U18181 ( .A(n17650), .B(n15573), .Z(n12841) );
  XOR U18182 ( .A(n17651), .B(n16032), .Z(n15573) );
  ANDN U18183 ( .B(n16834), .A(n16311), .Z(n17650) );
  XNOR U18184 ( .A(n17652), .B(n17203), .Z(n16311) );
  XNOR U18185 ( .A(n17653), .B(n17654), .Z(n16834) );
  XOR U18186 ( .A(n11782), .B(n17655), .Z(n17642) );
  XNOR U18187 ( .A(n11478), .B(n14022), .Z(n17655) );
  XNOR U18188 ( .A(n17656), .B(n15582), .Z(n14022) );
  XOR U18189 ( .A(n17657), .B(n17658), .Z(n15582) );
  ANDN U18190 ( .B(n16306), .A(n15067), .Z(n17656) );
  XOR U18191 ( .A(n17659), .B(n17660), .Z(n15067) );
  XNOR U18192 ( .A(n17661), .B(n17586), .Z(n16306) );
  XOR U18193 ( .A(n17662), .B(n15580), .Z(n11478) );
  XOR U18194 ( .A(n17663), .B(n16154), .Z(n15580) );
  XNOR U18195 ( .A(n17664), .B(n16744), .Z(n15063) );
  XOR U18196 ( .A(n17665), .B(n17333), .Z(n16315) );
  XNOR U18197 ( .A(n17666), .B(n15577), .Z(n11782) );
  XOR U18198 ( .A(n17667), .B(n14999), .Z(n15577) );
  ANDN U18199 ( .B(n16309), .A(n16329), .Z(n17666) );
  XNOR U18200 ( .A(n17668), .B(n16954), .Z(n16329) );
  XOR U18201 ( .A(n17669), .B(n15692), .Z(n16309) );
  IV U18202 ( .A(n17451), .Z(n15692) );
  XOR U18203 ( .A(n9101), .B(n17670), .Z(n9361) );
  XNOR U18204 ( .A(n13160), .B(n12671), .Z(n9101) );
  XNOR U18205 ( .A(n17671), .B(n17672), .Z(n12671) );
  XOR U18206 ( .A(n12883), .B(n12298), .Z(n17672) );
  XOR U18207 ( .A(n17673), .B(n17674), .Z(n12298) );
  XNOR U18208 ( .A(n17676), .B(n16137), .Z(n12883) );
  ANDN U18209 ( .B(n13697), .A(n16138), .Z(n17676) );
  XOR U18210 ( .A(n12389), .B(n17677), .Z(n17671) );
  XOR U18211 ( .A(n10105), .B(n13294), .Z(n17677) );
  XNOR U18212 ( .A(n17678), .B(n16126), .Z(n13294) );
  IV U18213 ( .A(n17679), .Z(n16126) );
  NOR U18214 ( .A(n16125), .B(n17680), .Z(n17678) );
  XNOR U18215 ( .A(n17681), .B(n16134), .Z(n10105) );
  IV U18216 ( .A(n17682), .Z(n16134) );
  ANDN U18217 ( .B(n16135), .A(n17683), .Z(n17681) );
  XOR U18218 ( .A(n17684), .B(n16128), .Z(n12389) );
  ANDN U18219 ( .B(n16129), .A(n12460), .Z(n17684) );
  XOR U18220 ( .A(n17685), .B(n17686), .Z(n13160) );
  XNOR U18221 ( .A(n9432), .B(n16120), .Z(n17686) );
  XNOR U18222 ( .A(n17687), .B(n14552), .Z(n16120) );
  IV U18223 ( .A(n16150), .Z(n14552) );
  XOR U18224 ( .A(n17688), .B(n15261), .Z(n16150) );
  ANDN U18225 ( .B(n16151), .A(n16013), .Z(n17687) );
  XOR U18226 ( .A(n17689), .B(n14560), .Z(n9432) );
  XOR U18227 ( .A(n17690), .B(n16115), .Z(n14560) );
  ANDN U18228 ( .B(n16019), .A(n16145), .Z(n17689) );
  XOR U18229 ( .A(n11819), .B(n17691), .Z(n17685) );
  XNOR U18230 ( .A(n9863), .B(n10597), .Z(n17691) );
  XOR U18231 ( .A(n17692), .B(n14557), .Z(n10597) );
  XOR U18232 ( .A(n17693), .B(n17514), .Z(n14557) );
  XNOR U18233 ( .A(n17695), .B(n14565), .Z(n9863) );
  IV U18234 ( .A(n16156), .Z(n14565) );
  XOR U18235 ( .A(n16036), .B(n17696), .Z(n16156) );
  XNOR U18236 ( .A(n17698), .B(n17699), .Z(n14548) );
  ANDN U18237 ( .B(n16158), .A(n16366), .Z(n17697) );
  XNOR U18238 ( .A(n17700), .B(n9370), .Z(n3569) );
  IV U18239 ( .A(n10631), .Z(n9370) );
  XOR U18240 ( .A(n17701), .B(n11414), .Z(n10631) );
  XNOR U18241 ( .A(n15330), .B(n17702), .Z(n11414) );
  XOR U18242 ( .A(n17703), .B(n17704), .Z(n15330) );
  XOR U18243 ( .A(n11687), .B(n12655), .Z(n17704) );
  XNOR U18244 ( .A(n17705), .B(n17706), .Z(n12655) );
  AND U18245 ( .A(n17707), .B(n15723), .Z(n17705) );
  XOR U18246 ( .A(n17708), .B(n17709), .Z(n11687) );
  NOR U18247 ( .A(n17710), .B(n17711), .Z(n17708) );
  XOR U18248 ( .A(n11220), .B(n17712), .Z(n17703) );
  XOR U18249 ( .A(n17713), .B(n12435), .Z(n17712) );
  XNOR U18250 ( .A(n17714), .B(n17715), .Z(n12435) );
  ANDN U18251 ( .B(n17716), .A(n15719), .Z(n17714) );
  XNOR U18252 ( .A(n17717), .B(n17718), .Z(n11220) );
  ANDN U18253 ( .B(n15727), .A(n17719), .Z(n17717) );
  NOR U18254 ( .A(n9354), .B(n10519), .Z(n17700) );
  XOR U18255 ( .A(n12446), .B(n11942), .Z(n10519) );
  IV U18256 ( .A(n14443), .Z(n11942) );
  XNOR U18257 ( .A(n17720), .B(n17721), .Z(n14443) );
  XNOR U18258 ( .A(n17722), .B(n17680), .Z(n12446) );
  NOR U18259 ( .A(n16124), .B(n17723), .Z(n17722) );
  XOR U18260 ( .A(n10743), .B(n15038), .Z(n9354) );
  XNOR U18261 ( .A(n17724), .B(n17725), .Z(n15038) );
  NOR U18262 ( .A(n13348), .B(n13349), .Z(n17724) );
  XNOR U18263 ( .A(n17726), .B(n16507), .Z(n13349) );
  XNOR U18264 ( .A(n13913), .B(n17727), .Z(n10743) );
  XOR U18265 ( .A(n17728), .B(n17729), .Z(n13913) );
  XOR U18266 ( .A(n12976), .B(n12601), .Z(n17729) );
  XOR U18267 ( .A(n17730), .B(n16565), .Z(n12601) );
  AND U18268 ( .A(n14888), .B(n14887), .Z(n17730) );
  XOR U18269 ( .A(n17731), .B(n17732), .Z(n14887) );
  XNOR U18270 ( .A(n17733), .B(n13462), .Z(n12976) );
  XNOR U18271 ( .A(n17734), .B(n17735), .Z(n13462) );
  ANDN U18272 ( .B(n14880), .A(n14881), .Z(n17733) );
  XNOR U18273 ( .A(n16815), .B(n17736), .Z(n14880) );
  XNOR U18274 ( .A(n11567), .B(n17737), .Z(n17728) );
  XOR U18275 ( .A(n15586), .B(n15730), .Z(n17737) );
  XNOR U18276 ( .A(n17738), .B(n16558), .Z(n15730) );
  IV U18277 ( .A(n13458), .Z(n16558) );
  XOR U18278 ( .A(n17739), .B(n17740), .Z(n13458) );
  ANDN U18279 ( .B(n14894), .A(n14895), .Z(n17738) );
  XOR U18280 ( .A(n17284), .B(n17741), .Z(n14894) );
  XNOR U18281 ( .A(n17742), .B(n13451), .Z(n15586) );
  XOR U18282 ( .A(n17743), .B(n17744), .Z(n13451) );
  AND U18283 ( .A(n14891), .B(n14892), .Z(n17742) );
  XOR U18284 ( .A(n17745), .B(n17746), .Z(n14891) );
  XNOR U18285 ( .A(n17747), .B(n13447), .Z(n11567) );
  XOR U18286 ( .A(n17748), .B(n17601), .Z(n13447) );
  NOR U18287 ( .A(n14883), .B(n14884), .Z(n17747) );
  XOR U18288 ( .A(n17749), .B(n17750), .Z(n14883) );
  XNOR U18289 ( .A(n17751), .B(n6972), .Z(n2654) );
  XNOR U18290 ( .A(n10878), .B(n17752), .Z(n6972) );
  XNOR U18291 ( .A(n17753), .B(n17754), .Z(n14592) );
  XNOR U18292 ( .A(n11901), .B(n17755), .Z(n17754) );
  XNOR U18293 ( .A(n17756), .B(n17379), .Z(n11901) );
  AND U18294 ( .A(n17757), .B(n17758), .Z(n17756) );
  XNOR U18295 ( .A(n13480), .B(n17759), .Z(n17753) );
  XOR U18296 ( .A(n17760), .B(n14651), .Z(n17759) );
  ANDN U18297 ( .B(n17762), .A(n17763), .Z(n17761) );
  XOR U18298 ( .A(n17764), .B(n17376), .Z(n13480) );
  ANDN U18299 ( .B(n17765), .A(n17766), .Z(n17764) );
  XOR U18300 ( .A(n17767), .B(n17768), .Z(n11323) );
  XNOR U18301 ( .A(n9938), .B(n11776), .Z(n17768) );
  XOR U18302 ( .A(n17769), .B(n16539), .Z(n11776) );
  ANDN U18303 ( .B(n14768), .A(n14769), .Z(n17769) );
  XNOR U18304 ( .A(n17770), .B(n16549), .Z(n9938) );
  ANDN U18305 ( .B(n14772), .A(n17771), .Z(n17770) );
  XNOR U18306 ( .A(n10689), .B(n17772), .Z(n17767) );
  XOR U18307 ( .A(n11846), .B(n10864), .Z(n17772) );
  XNOR U18308 ( .A(n17773), .B(n16568), .Z(n10864) );
  ANDN U18309 ( .B(n14777), .A(n14778), .Z(n17773) );
  XOR U18310 ( .A(n17774), .B(n17775), .Z(n11846) );
  ANDN U18311 ( .B(n14781), .A(n14782), .Z(n17774) );
  XOR U18312 ( .A(n17776), .B(n16544), .Z(n10689) );
  ANDN U18313 ( .B(n14785), .A(n14786), .Z(n17776) );
  ANDN U18314 ( .B(n9367), .A(n10524), .Z(n17751) );
  XOR U18315 ( .A(n10752), .B(n14835), .Z(n10524) );
  XOR U18316 ( .A(n17777), .B(n17778), .Z(n14835) );
  NOR U18317 ( .A(n17779), .B(n14405), .Z(n17777) );
  IV U18318 ( .A(n12326), .Z(n10752) );
  XNOR U18319 ( .A(n13645), .B(n14449), .Z(n12326) );
  XOR U18320 ( .A(n17780), .B(n17781), .Z(n14449) );
  XOR U18321 ( .A(n14131), .B(n13794), .Z(n17781) );
  XOR U18322 ( .A(n17782), .B(n14429), .Z(n13794) );
  XNOR U18323 ( .A(n14992), .B(n17783), .Z(n14429) );
  NOR U18324 ( .A(n15359), .B(n15360), .Z(n17782) );
  XOR U18325 ( .A(n17784), .B(n16094), .Z(n15359) );
  XOR U18326 ( .A(n17785), .B(n14439), .Z(n14131) );
  XOR U18327 ( .A(n17786), .B(n17503), .Z(n14439) );
  ANDN U18328 ( .B(n15357), .A(n15356), .Z(n17785) );
  XOR U18329 ( .A(n17787), .B(n17788), .Z(n15356) );
  XNOR U18330 ( .A(n11752), .B(n17789), .Z(n17780) );
  XOR U18331 ( .A(n15628), .B(n11703), .Z(n17789) );
  XOR U18332 ( .A(n17790), .B(n14424), .Z(n11703) );
  XOR U18333 ( .A(n15342), .B(n17791), .Z(n14424) );
  ANDN U18334 ( .B(n15366), .A(n15367), .Z(n17790) );
  XNOR U18335 ( .A(n15885), .B(n17792), .Z(n15366) );
  XNOR U18336 ( .A(n17793), .B(n14421), .Z(n15628) );
  XOR U18337 ( .A(n17794), .B(n17795), .Z(n14421) );
  ANDN U18338 ( .B(n15370), .A(n15369), .Z(n17793) );
  XOR U18339 ( .A(n17796), .B(n16872), .Z(n15369) );
  XOR U18340 ( .A(n17797), .B(n14434), .Z(n11752) );
  XOR U18341 ( .A(n17798), .B(n17108), .Z(n14434) );
  ANDN U18342 ( .B(n15363), .A(n15364), .Z(n17797) );
  XNOR U18343 ( .A(n17799), .B(n16579), .Z(n15363) );
  XOR U18344 ( .A(n17800), .B(n17801), .Z(n13645) );
  XOR U18345 ( .A(n16252), .B(n11164), .Z(n17801) );
  XOR U18346 ( .A(n17802), .B(n17803), .Z(n11164) );
  ANDN U18347 ( .B(n14844), .A(n14845), .Z(n17802) );
  XOR U18348 ( .A(n17804), .B(n14415), .Z(n16252) );
  ANDN U18349 ( .B(n14849), .A(n14848), .Z(n17804) );
  XOR U18350 ( .A(n11934), .B(n17805), .Z(n17800) );
  XOR U18351 ( .A(n11123), .B(n13043), .Z(n17805) );
  XNOR U18352 ( .A(n17806), .B(n14402), .Z(n13043) );
  IV U18353 ( .A(n17807), .Z(n14402) );
  NOR U18354 ( .A(n14841), .B(n14842), .Z(n17806) );
  XOR U18355 ( .A(n17808), .B(n14406), .Z(n11123) );
  XNOR U18356 ( .A(n17809), .B(n17810), .Z(n11934) );
  ANDN U18357 ( .B(n14837), .A(n14838), .Z(n17809) );
  XOR U18358 ( .A(n14682), .B(n9636), .Z(n9367) );
  XNOR U18359 ( .A(n17811), .B(n16263), .Z(n9636) );
  XNOR U18360 ( .A(n17812), .B(n17813), .Z(n16263) );
  XNOR U18361 ( .A(n12747), .B(n12383), .Z(n17813) );
  XOR U18362 ( .A(n17814), .B(n14120), .Z(n12383) );
  NOR U18363 ( .A(n17815), .B(n17816), .Z(n17814) );
  XOR U18364 ( .A(n17817), .B(n17818), .Z(n12747) );
  ANDN U18365 ( .B(n17819), .A(n17820), .Z(n17817) );
  XNOR U18366 ( .A(n11487), .B(n17821), .Z(n17812) );
  XOR U18367 ( .A(n16656), .B(n11212), .Z(n17821) );
  XOR U18368 ( .A(n17822), .B(n17823), .Z(n11212) );
  NOR U18369 ( .A(n17824), .B(n17825), .Z(n17822) );
  XOR U18370 ( .A(n17826), .B(n14257), .Z(n16656) );
  NOR U18371 ( .A(n17827), .B(n17828), .Z(n17826) );
  XOR U18372 ( .A(n17829), .B(n15100), .Z(n11487) );
  NOR U18373 ( .A(n17830), .B(n17831), .Z(n17829) );
  XNOR U18374 ( .A(n17832), .B(n17833), .Z(n14682) );
  ANDN U18375 ( .B(n14194), .A(n16897), .Z(n17832) );
  XOR U18376 ( .A(n17834), .B(n15537), .Z(n14194) );
  IV U18377 ( .A(n17835), .Z(n15537) );
  AND U18378 ( .A(n4105), .B(n2607), .Z(n16903) );
  XOR U18379 ( .A(n7669), .B(n2622), .Z(n2607) );
  XNOR U18380 ( .A(n5992), .B(n6413), .Z(n2622) );
  XNOR U18381 ( .A(n17836), .B(n17837), .Z(n6413) );
  XNOR U18382 ( .A(n2656), .B(n5381), .Z(n17837) );
  XNOR U18383 ( .A(n17838), .B(n6859), .Z(n5381) );
  XNOR U18384 ( .A(n16131), .B(n9260), .Z(n6859) );
  XNOR U18385 ( .A(n13650), .B(n12896), .Z(n9260) );
  XNOR U18386 ( .A(n17839), .B(n17840), .Z(n12896) );
  XNOR U18387 ( .A(n10210), .B(n13164), .Z(n17840) );
  XNOR U18388 ( .A(n17841), .B(n17842), .Z(n13164) );
  ANDN U18389 ( .B(n15396), .A(n15397), .Z(n17841) );
  XNOR U18390 ( .A(n17843), .B(n13835), .Z(n10210) );
  ANDN U18391 ( .B(n13834), .A(n15405), .Z(n17843) );
  IV U18392 ( .A(n15404), .Z(n13834) );
  XOR U18393 ( .A(n17844), .B(n17845), .Z(n15404) );
  XNOR U18394 ( .A(n13821), .B(n17846), .Z(n17839) );
  XOR U18395 ( .A(n12531), .B(n12620), .Z(n17846) );
  XNOR U18396 ( .A(n17847), .B(n14588), .Z(n12620) );
  ANDN U18397 ( .B(n15409), .A(n14587), .Z(n17847) );
  XNOR U18398 ( .A(n17848), .B(n17589), .Z(n14587) );
  XNOR U18399 ( .A(n17849), .B(n13838), .Z(n12531) );
  AND U18400 ( .A(n15394), .B(n13839), .Z(n17849) );
  XOR U18401 ( .A(n17850), .B(n15702), .Z(n13839) );
  XNOR U18402 ( .A(n17851), .B(n13828), .Z(n13821) );
  ANDN U18403 ( .B(n13829), .A(n15401), .Z(n17851) );
  XNOR U18404 ( .A(n17852), .B(n17853), .Z(n13829) );
  XOR U18405 ( .A(n17854), .B(n17855), .Z(n13650) );
  XOR U18406 ( .A(n10720), .B(n9933), .Z(n17855) );
  XNOR U18407 ( .A(n17856), .B(n17723), .Z(n9933) );
  ANDN U18408 ( .B(n16124), .A(n17679), .Z(n17856) );
  XOR U18409 ( .A(n17857), .B(n16954), .Z(n17679) );
  XOR U18410 ( .A(n17858), .B(n17845), .Z(n16124) );
  IV U18411 ( .A(n17108), .Z(n17845) );
  XOR U18412 ( .A(n17859), .B(n14446), .Z(n10720) );
  ANDN U18413 ( .B(n14447), .A(n17682), .Z(n17859) );
  XNOR U18414 ( .A(n17860), .B(n17861), .Z(n17682) );
  IV U18415 ( .A(n16133), .Z(n14447) );
  XOR U18416 ( .A(n17862), .B(n17186), .Z(n16133) );
  XNOR U18417 ( .A(n10700), .B(n17863), .Z(n17854) );
  XOR U18418 ( .A(n9521), .B(n9123), .Z(n17863) );
  XNOR U18419 ( .A(n17864), .B(n13698), .Z(n9123) );
  ANDN U18420 ( .B(n13699), .A(n16137), .Z(n17864) );
  XOR U18421 ( .A(n17865), .B(n16892), .Z(n16137) );
  XNOR U18422 ( .A(n17866), .B(n17626), .Z(n13699) );
  XOR U18423 ( .A(n17867), .B(n12461), .Z(n9521) );
  XNOR U18424 ( .A(n17868), .B(n15304), .Z(n16128) );
  XOR U18425 ( .A(n17869), .B(n17870), .Z(n12462) );
  XNOR U18426 ( .A(n17871), .B(n12451), .Z(n10700) );
  ANDN U18427 ( .B(n17674), .A(n12450), .Z(n17871) );
  XNOR U18428 ( .A(n17872), .B(n12450), .Z(n16131) );
  XOR U18429 ( .A(n17873), .B(n17874), .Z(n12450) );
  NOR U18430 ( .A(n17675), .B(n17674), .Z(n17872) );
  XNOR U18431 ( .A(n17875), .B(n16301), .Z(n17674) );
  ANDN U18432 ( .B(n7678), .A(n6860), .Z(n17838) );
  XOR U18433 ( .A(n10224), .B(n17876), .Z(n6860) );
  IV U18434 ( .A(n10928), .Z(n10224) );
  XOR U18435 ( .A(n14927), .B(n14676), .Z(n10928) );
  XNOR U18436 ( .A(n17877), .B(n17878), .Z(n14676) );
  XOR U18437 ( .A(n11821), .B(n9523), .Z(n17878) );
  XNOR U18438 ( .A(n17879), .B(n17828), .Z(n9523) );
  ANDN U18439 ( .B(n17827), .A(n17880), .Z(n17879) );
  XNOR U18440 ( .A(n17881), .B(n17820), .Z(n11821) );
  IV U18441 ( .A(n17882), .Z(n17820) );
  NOR U18442 ( .A(n17819), .B(n17883), .Z(n17881) );
  IV U18443 ( .A(n17884), .Z(n17819) );
  XNOR U18444 ( .A(n16262), .B(n17885), .Z(n17877) );
  XNOR U18445 ( .A(n15051), .B(n12501), .Z(n17885) );
  XNOR U18446 ( .A(n17886), .B(n17815), .Z(n12501) );
  IV U18447 ( .A(n17887), .Z(n17815) );
  ANDN U18448 ( .B(n17816), .A(n14118), .Z(n17886) );
  XNOR U18449 ( .A(n17888), .B(n17825), .Z(n15051) );
  ANDN U18450 ( .B(n17824), .A(n17889), .Z(n17888) );
  XNOR U18451 ( .A(n17890), .B(n17831), .Z(n16262) );
  ANDN U18452 ( .B(n17830), .A(n17891), .Z(n17890) );
  XNOR U18453 ( .A(n17892), .B(n17893), .Z(n14927) );
  XNOR U18454 ( .A(n10211), .B(n10052), .Z(n17893) );
  XNOR U18455 ( .A(n17894), .B(n16268), .Z(n10052) );
  XOR U18456 ( .A(n17895), .B(n16674), .Z(n16268) );
  ANDN U18457 ( .B(n16243), .A(n16269), .Z(n17894) );
  XNOR U18458 ( .A(n17896), .B(n17038), .Z(n10211) );
  XOR U18459 ( .A(n17897), .B(n17898), .Z(n17038) );
  AND U18460 ( .A(n17070), .B(n16226), .Z(n17896) );
  XNOR U18461 ( .A(n9425), .B(n17899), .Z(n17892) );
  XOR U18462 ( .A(n10232), .B(n15077), .Z(n17899) );
  XNOR U18463 ( .A(n17900), .B(n17043), .Z(n15077) );
  IV U18464 ( .A(n16273), .Z(n17043) );
  XOR U18465 ( .A(n17901), .B(n17902), .Z(n16273) );
  ANDN U18466 ( .B(n16239), .A(n16272), .Z(n17900) );
  XOR U18467 ( .A(n17903), .B(n16275), .Z(n10232) );
  XOR U18468 ( .A(n16609), .B(n17904), .Z(n16275) );
  IV U18469 ( .A(n15196), .Z(n16609) );
  AND U18470 ( .A(n16276), .B(n16235), .Z(n17903) );
  XNOR U18471 ( .A(n17905), .B(n16278), .Z(n9425) );
  XNOR U18472 ( .A(n17906), .B(n17907), .Z(n16278) );
  AND U18473 ( .A(n16279), .B(n16230), .Z(n17905) );
  XOR U18474 ( .A(n16451), .B(n10080), .Z(n7678) );
  IV U18475 ( .A(n13301), .Z(n10080) );
  XOR U18476 ( .A(n15861), .B(n17362), .Z(n13301) );
  XOR U18477 ( .A(n17908), .B(n17909), .Z(n17362) );
  XOR U18478 ( .A(n10590), .B(n14690), .Z(n17909) );
  XNOR U18479 ( .A(n17910), .B(n16637), .Z(n14690) );
  XOR U18480 ( .A(n17911), .B(n17658), .Z(n16637) );
  NOR U18481 ( .A(n17912), .B(n16453), .Z(n17910) );
  XOR U18482 ( .A(n17913), .B(n17015), .Z(n16453) );
  XNOR U18483 ( .A(n17914), .B(n16632), .Z(n10590) );
  XOR U18484 ( .A(n17915), .B(n17916), .Z(n16632) );
  ANDN U18485 ( .B(n16443), .A(n16444), .Z(n17914) );
  XNOR U18486 ( .A(n17917), .B(n17918), .Z(n16443) );
  XOR U18487 ( .A(n16906), .B(n17919), .Z(n17908) );
  XNOR U18488 ( .A(n11105), .B(n12731), .Z(n17919) );
  XNOR U18489 ( .A(n17920), .B(n16640), .Z(n12731) );
  XNOR U18490 ( .A(n17921), .B(n17922), .Z(n16640) );
  ANDN U18491 ( .B(n16448), .A(n16914), .Z(n17920) );
  XOR U18492 ( .A(n17923), .B(n16061), .Z(n16914) );
  XOR U18493 ( .A(n17924), .B(n16643), .Z(n11105) );
  XOR U18494 ( .A(n17925), .B(n16096), .Z(n16643) );
  AND U18495 ( .A(n16459), .B(n16457), .Z(n17924) );
  XOR U18496 ( .A(n17926), .B(n17927), .Z(n16457) );
  XNOR U18497 ( .A(n17928), .B(n16630), .Z(n16906) );
  XOR U18498 ( .A(n17929), .B(n16108), .Z(n16630) );
  AND U18499 ( .A(n16916), .B(n17930), .Z(n17928) );
  XOR U18500 ( .A(n17931), .B(n17932), .Z(n15861) );
  XOR U18501 ( .A(n10323), .B(n12677), .Z(n17932) );
  XNOR U18502 ( .A(n17933), .B(n16922), .Z(n12677) );
  ANDN U18503 ( .B(n16424), .A(n16425), .Z(n17933) );
  XOR U18504 ( .A(n17934), .B(n16763), .Z(n16425) );
  IV U18505 ( .A(n17898), .Z(n16763) );
  XOR U18506 ( .A(n15875), .B(n17935), .Z(n16424) );
  XNOR U18507 ( .A(n17936), .B(n16925), .Z(n10323) );
  ANDN U18508 ( .B(n16431), .A(n16429), .Z(n17936) );
  XOR U18509 ( .A(n17938), .B(n16045), .Z(n16431) );
  XNOR U18510 ( .A(n12335), .B(n17939), .Z(n17931) );
  XNOR U18511 ( .A(n11036), .B(n12293), .Z(n17939) );
  NOR U18512 ( .A(n16437), .B(n16438), .Z(n17940) );
  XNOR U18513 ( .A(n17941), .B(n17942), .Z(n16438) );
  IV U18514 ( .A(n16931), .Z(n16437) );
  XOR U18515 ( .A(n17943), .B(n17944), .Z(n16931) );
  XNOR U18516 ( .A(n17945), .B(n17946), .Z(n11036) );
  ANDN U18517 ( .B(n16420), .A(n16421), .Z(n17945) );
  XOR U18518 ( .A(n17947), .B(n17429), .Z(n16421) );
  XOR U18519 ( .A(n17948), .B(n16934), .Z(n12335) );
  XOR U18520 ( .A(n17949), .B(n17436), .Z(n16433) );
  XNOR U18521 ( .A(n17950), .B(n17916), .Z(n16435) );
  XOR U18522 ( .A(n17951), .B(n16916), .Z(n16451) );
  XNOR U18523 ( .A(n17952), .B(n15290), .Z(n16916) );
  NOR U18524 ( .A(n16628), .B(n17930), .Z(n17951) );
  XNOR U18525 ( .A(n17953), .B(n6864), .Z(n2656) );
  XNOR U18526 ( .A(n16649), .B(n9927), .Z(n6864) );
  XNOR U18527 ( .A(n17222), .B(n15441), .Z(n9927) );
  XOR U18528 ( .A(n17954), .B(n17955), .Z(n15441) );
  XNOR U18529 ( .A(n16416), .B(n10187), .Z(n17955) );
  XNOR U18530 ( .A(n17956), .B(n16448), .Z(n10187) );
  XNOR U18531 ( .A(n17957), .B(n17958), .Z(n16448) );
  ANDN U18532 ( .B(n16449), .A(n16913), .Z(n17956) );
  XNOR U18533 ( .A(n17959), .B(n17654), .Z(n16913) );
  XOR U18534 ( .A(n17960), .B(n17961), .Z(n16449) );
  XNOR U18535 ( .A(n17962), .B(n16454), .Z(n16416) );
  IV U18536 ( .A(n17912), .Z(n16454) );
  XOR U18537 ( .A(n17963), .B(n14999), .Z(n17912) );
  ANDN U18538 ( .B(n16455), .A(n16636), .Z(n17962) );
  XNOR U18539 ( .A(n17964), .B(n16579), .Z(n16636) );
  XNOR U18540 ( .A(n17965), .B(n16878), .Z(n16455) );
  XNOR U18541 ( .A(n12183), .B(n17966), .Z(n17954) );
  XNOR U18542 ( .A(n12613), .B(n10956), .Z(n17966) );
  XNOR U18543 ( .A(n17967), .B(n17930), .Z(n10956) );
  XOR U18544 ( .A(n17968), .B(n16739), .Z(n17930) );
  ANDN U18545 ( .B(n16628), .A(n16629), .Z(n17967) );
  XNOR U18546 ( .A(n17969), .B(n17970), .Z(n16629) );
  XOR U18547 ( .A(n17971), .B(n14168), .Z(n16628) );
  XOR U18548 ( .A(n17972), .B(n16444), .Z(n12613) );
  XNOR U18549 ( .A(n17321), .B(n17973), .Z(n16444) );
  AND U18550 ( .A(n16633), .B(n16445), .Z(n17972) );
  XNOR U18551 ( .A(n17974), .B(n17975), .Z(n16445) );
  XOR U18552 ( .A(n17976), .B(n17977), .Z(n16633) );
  XNOR U18553 ( .A(n17978), .B(n16459), .Z(n12183) );
  XOR U18554 ( .A(n17979), .B(n17980), .Z(n16459) );
  NOR U18555 ( .A(n16458), .B(n16642), .Z(n17978) );
  XOR U18556 ( .A(n17981), .B(n16858), .Z(n16642) );
  IV U18557 ( .A(n17982), .Z(n16858) );
  XOR U18558 ( .A(n17026), .B(n17983), .Z(n16458) );
  XOR U18559 ( .A(n17984), .B(n17985), .Z(n17222) );
  XNOR U18560 ( .A(n10385), .B(n13865), .Z(n17985) );
  XNOR U18561 ( .A(n17986), .B(n14280), .Z(n13865) );
  NOR U18562 ( .A(n16623), .B(n14281), .Z(n17986) );
  XOR U18563 ( .A(n17987), .B(n17988), .Z(n14281) );
  XNOR U18564 ( .A(n17989), .B(n15339), .Z(n16623) );
  XNOR U18565 ( .A(n17990), .B(n17991), .Z(n10385) );
  ANDN U18566 ( .B(n15109), .A(n14285), .Z(n17990) );
  XOR U18567 ( .A(n17992), .B(n17229), .Z(n14285) );
  XOR U18568 ( .A(n17993), .B(n15873), .Z(n15109) );
  IV U18569 ( .A(n17994), .Z(n15873) );
  XNOR U18570 ( .A(n10361), .B(n17995), .Z(n17984) );
  XNOR U18571 ( .A(n11756), .B(n12457), .Z(n17995) );
  XOR U18572 ( .A(n17996), .B(n17364), .Z(n12457) );
  XOR U18573 ( .A(n17997), .B(n15650), .Z(n16652) );
  XNOR U18574 ( .A(n17998), .B(n17564), .Z(n15112) );
  XNOR U18575 ( .A(n17999), .B(n14294), .Z(n11756) );
  XOR U18576 ( .A(n18000), .B(n14290), .Z(n10361) );
  ANDN U18577 ( .B(n14291), .A(n15118), .Z(n18000) );
  XOR U18578 ( .A(n18001), .B(n16074), .Z(n15118) );
  XNOR U18579 ( .A(n18002), .B(n17744), .Z(n14291) );
  XOR U18580 ( .A(n18003), .B(n14295), .Z(n16649) );
  XOR U18581 ( .A(n18004), .B(n18005), .Z(n14295) );
  ANDN U18582 ( .B(n15122), .A(n15123), .Z(n18003) );
  XOR U18583 ( .A(n18006), .B(n16767), .Z(n15122) );
  ANDN U18584 ( .B(n9968), .A(n6863), .Z(n17953) );
  XNOR U18585 ( .A(n3345), .B(n18007), .Z(n17836) );
  XOR U18586 ( .A(n5364), .B(n6853), .Z(n18007) );
  XNOR U18587 ( .A(n18008), .B(n7559), .Z(n6853) );
  IV U18588 ( .A(n6868), .Z(n7559) );
  XOR U18589 ( .A(n9565), .B(n13182), .Z(n6868) );
  XNOR U18590 ( .A(n18009), .B(n13790), .Z(n13182) );
  ANDN U18591 ( .B(n18010), .A(n15943), .Z(n18009) );
  IV U18592 ( .A(n11907), .Z(n9565) );
  XNOR U18593 ( .A(n14324), .B(n13288), .Z(n11907) );
  XOR U18594 ( .A(n18011), .B(n18012), .Z(n13288) );
  XNOR U18595 ( .A(n13655), .B(n10983), .Z(n18012) );
  XOR U18596 ( .A(n18013), .B(n13669), .Z(n10983) );
  XOR U18597 ( .A(n18014), .B(n18015), .Z(n13669) );
  ANDN U18598 ( .B(n13186), .A(n13184), .Z(n18013) );
  XOR U18599 ( .A(n18016), .B(n18017), .Z(n13184) );
  XOR U18600 ( .A(n18018), .B(n13804), .Z(n13655) );
  XOR U18601 ( .A(n18019), .B(n16844), .Z(n13804) );
  NOR U18602 ( .A(n18020), .B(n13189), .Z(n18018) );
  XOR U18603 ( .A(n18021), .B(n16036), .Z(n13189) );
  XOR U18604 ( .A(n12217), .B(n18022), .Z(n18011) );
  XNOR U18605 ( .A(n11824), .B(n9812), .Z(n18022) );
  XNOR U18606 ( .A(n18023), .B(n13666), .Z(n9812) );
  ANDN U18607 ( .B(n13197), .A(n18024), .Z(n18023) );
  XNOR U18608 ( .A(n18025), .B(n16855), .Z(n13197) );
  XNOR U18609 ( .A(n18026), .B(n13661), .Z(n11824) );
  XOR U18610 ( .A(n18027), .B(n18028), .Z(n13661) );
  AND U18611 ( .A(n13193), .B(n13195), .Z(n18026) );
  XOR U18612 ( .A(n18029), .B(n17498), .Z(n13193) );
  XNOR U18613 ( .A(n18030), .B(n13791), .Z(n12217) );
  XNOR U18614 ( .A(n15958), .B(n18031), .Z(n13791) );
  NOR U18615 ( .A(n13790), .B(n18010), .Z(n18030) );
  XOR U18616 ( .A(n18032), .B(n18033), .Z(n13790) );
  XOR U18617 ( .A(n18034), .B(n18035), .Z(n14324) );
  XOR U18618 ( .A(n10492), .B(n11575), .Z(n18035) );
  XNOR U18619 ( .A(n18036), .B(n13684), .Z(n11575) );
  NOR U18620 ( .A(n13683), .B(n14640), .Z(n18036) );
  XOR U18621 ( .A(n18039), .B(n13691), .Z(n10492) );
  XOR U18622 ( .A(n18040), .B(n17916), .Z(n13691) );
  ANDN U18623 ( .B(n14643), .A(n14642), .Z(n18039) );
  IV U18624 ( .A(n13692), .Z(n14642) );
  XOR U18625 ( .A(n18041), .B(n17195), .Z(n13692) );
  XOR U18626 ( .A(n9325), .B(n18042), .Z(n18034) );
  XOR U18627 ( .A(n9250), .B(n11724), .Z(n18042) );
  XOR U18628 ( .A(n18043), .B(n13679), .Z(n11724) );
  XOR U18629 ( .A(n17399), .B(n18044), .Z(n13679) );
  ANDN U18630 ( .B(n13678), .A(n14646), .Z(n18043) );
  XOR U18631 ( .A(n18045), .B(n18046), .Z(n13678) );
  XNOR U18632 ( .A(n18047), .B(n13687), .Z(n9250) );
  XOR U18633 ( .A(n18048), .B(n18049), .Z(n13687) );
  XOR U18634 ( .A(n18050), .B(n18051), .Z(n13688) );
  XNOR U18635 ( .A(n18052), .B(n13674), .Z(n9325) );
  XOR U18636 ( .A(n18053), .B(n18054), .Z(n13674) );
  ANDN U18637 ( .B(n13675), .A(n14650), .Z(n18052) );
  XOR U18638 ( .A(n17901), .B(n18055), .Z(n13675) );
  AND U18639 ( .A(n7676), .B(n6869), .Z(n18008) );
  XNOR U18640 ( .A(n10978), .B(n17325), .Z(n6869) );
  XNOR U18641 ( .A(n18056), .B(n14797), .Z(n17325) );
  ANDN U18642 ( .B(n16870), .A(n16364), .Z(n18056) );
  XNOR U18643 ( .A(n18057), .B(n18058), .Z(n16364) );
  XOR U18644 ( .A(n18059), .B(n16251), .Z(n10978) );
  XNOR U18645 ( .A(n18060), .B(n18061), .Z(n16251) );
  XNOR U18646 ( .A(n11860), .B(n11635), .Z(n18061) );
  XNOR U18647 ( .A(n18062), .B(n12027), .Z(n11635) );
  AND U18648 ( .A(n12028), .B(n17346), .Z(n18062) );
  XOR U18649 ( .A(n18063), .B(n18064), .Z(n12028) );
  XNOR U18650 ( .A(n18065), .B(n12031), .Z(n11860) );
  XNOR U18651 ( .A(n18066), .B(n17918), .Z(n12031) );
  ANDN U18652 ( .B(n12032), .A(n17353), .Z(n18065) );
  XNOR U18653 ( .A(n18067), .B(n17994), .Z(n12032) );
  XOR U18654 ( .A(n11471), .B(n18068), .Z(n18060) );
  XNOR U18655 ( .A(n9628), .B(n10622), .Z(n18068) );
  XNOR U18656 ( .A(n18069), .B(n12044), .Z(n10622) );
  XOR U18657 ( .A(n18070), .B(n18071), .Z(n12044) );
  ANDN U18658 ( .B(n12045), .A(n17343), .Z(n18069) );
  IV U18659 ( .A(n18072), .Z(n17343) );
  XNOR U18660 ( .A(n18073), .B(n18074), .Z(n12045) );
  XOR U18661 ( .A(n18075), .B(n12040), .Z(n9628) );
  XOR U18662 ( .A(n18076), .B(n15304), .Z(n12040) );
  AND U18663 ( .A(n12041), .B(n17349), .Z(n18075) );
  XOR U18664 ( .A(n18077), .B(n18078), .Z(n12041) );
  XNOR U18665 ( .A(n18079), .B(n12036), .Z(n11471) );
  IV U18666 ( .A(n16345), .Z(n12036) );
  XOR U18667 ( .A(n18080), .B(n17578), .Z(n16345) );
  AND U18668 ( .A(n17351), .B(n12037), .Z(n18079) );
  XOR U18669 ( .A(n18081), .B(n17212), .Z(n12037) );
  XOR U18670 ( .A(n11092), .B(n17159), .Z(n7676) );
  XNOR U18671 ( .A(n18082), .B(n18083), .Z(n17159) );
  ANDN U18672 ( .B(n18084), .A(n18085), .Z(n18082) );
  IV U18673 ( .A(n12422), .Z(n11092) );
  XNOR U18674 ( .A(n12740), .B(n14136), .Z(n12422) );
  XOR U18675 ( .A(n18086), .B(n18087), .Z(n14136) );
  XNOR U18676 ( .A(n9514), .B(n13481), .Z(n18087) );
  XOR U18677 ( .A(n18088), .B(n17716), .Z(n13481) );
  ANDN U18678 ( .B(n15719), .A(n18089), .Z(n18088) );
  XOR U18679 ( .A(n18090), .B(n18091), .Z(n15719) );
  XNOR U18680 ( .A(n18092), .B(n18093), .Z(n9514) );
  ANDN U18681 ( .B(n18094), .A(n15710), .Z(n18092) );
  XNOR U18682 ( .A(n15329), .B(n18095), .Z(n18086) );
  XOR U18683 ( .A(n9137), .B(n10162), .Z(n18095) );
  XNOR U18684 ( .A(n18096), .B(n17719), .Z(n10162) );
  NOR U18685 ( .A(n18097), .B(n15727), .Z(n18096) );
  XOR U18686 ( .A(n18098), .B(n15201), .Z(n15727) );
  XNOR U18687 ( .A(n18099), .B(n17711), .Z(n9137) );
  ANDN U18688 ( .B(n15716), .A(n15714), .Z(n18099) );
  IV U18689 ( .A(n17710), .Z(n15714) );
  XOR U18690 ( .A(n18100), .B(n18101), .Z(n17710) );
  XOR U18691 ( .A(n18102), .B(n17707), .Z(n15329) );
  NOR U18692 ( .A(n15724), .B(n15723), .Z(n18102) );
  XOR U18693 ( .A(n18103), .B(n18104), .Z(n15723) );
  XOR U18694 ( .A(n18105), .B(n18106), .Z(n12740) );
  XNOR U18695 ( .A(n11626), .B(n11413), .Z(n18106) );
  XOR U18696 ( .A(n18107), .B(n18108), .Z(n11413) );
  XNOR U18697 ( .A(n18109), .B(n18110), .Z(n11626) );
  ANDN U18698 ( .B(n17166), .A(n17165), .Z(n18109) );
  XOR U18699 ( .A(n17701), .B(n18111), .Z(n18105) );
  XOR U18700 ( .A(n11646), .B(n11454), .Z(n18111) );
  XNOR U18701 ( .A(n18112), .B(n18113), .Z(n11454) );
  NOR U18702 ( .A(n18083), .B(n18084), .Z(n18112) );
  XOR U18703 ( .A(n18114), .B(n18115), .Z(n11646) );
  NOR U18704 ( .A(n17151), .B(n17152), .Z(n18114) );
  XNOR U18705 ( .A(n18116), .B(n18117), .Z(n17701) );
  NOR U18706 ( .A(n17155), .B(n17156), .Z(n18116) );
  XNOR U18707 ( .A(n18118), .B(n7565), .Z(n5364) );
  IV U18708 ( .A(n6872), .Z(n7565) );
  XOR U18709 ( .A(n18119), .B(n11444), .Z(n6872) );
  IV U18710 ( .A(n9888), .Z(n11444) );
  XNOR U18711 ( .A(n14809), .B(n14182), .Z(n9888) );
  XOR U18712 ( .A(n18120), .B(n18121), .Z(n14182) );
  XOR U18713 ( .A(n11497), .B(n9264), .Z(n18121) );
  XNOR U18714 ( .A(n18122), .B(n16717), .Z(n9264) );
  ANDN U18715 ( .B(n15918), .A(n18123), .Z(n18122) );
  XNOR U18716 ( .A(n18124), .B(n16715), .Z(n11497) );
  AND U18717 ( .A(n18125), .B(n15923), .Z(n18124) );
  XOR U18718 ( .A(n18126), .B(n18127), .Z(n18120) );
  XOR U18719 ( .A(n12580), .B(n12500), .Z(n18127) );
  XNOR U18720 ( .A(n18128), .B(n16719), .Z(n12500) );
  ANDN U18721 ( .B(n18129), .A(n15927), .Z(n18128) );
  XOR U18722 ( .A(n18130), .B(n16708), .Z(n12580) );
  ANDN U18723 ( .B(n18131), .A(n15931), .Z(n18130) );
  XOR U18724 ( .A(n18132), .B(n18133), .Z(n14809) );
  XOR U18725 ( .A(n11732), .B(n12594), .Z(n18133) );
  XOR U18726 ( .A(n18134), .B(n15018), .Z(n12594) );
  NOR U18727 ( .A(n16198), .B(n16199), .Z(n18134) );
  IV U18728 ( .A(n18135), .Z(n16198) );
  XNOR U18729 ( .A(n18136), .B(n18137), .Z(n11732) );
  AND U18730 ( .A(n16183), .B(n16185), .Z(n18136) );
  XNOR U18731 ( .A(n12962), .B(n18138), .Z(n18132) );
  XOR U18732 ( .A(n12437), .B(n11810), .Z(n18138) );
  XNOR U18733 ( .A(n18139), .B(n18140), .Z(n11810) );
  ANDN U18734 ( .B(n16196), .A(n16194), .Z(n18139) );
  IV U18735 ( .A(n18141), .Z(n16196) );
  ANDN U18736 ( .B(n16191), .A(n18143), .Z(n18142) );
  IV U18737 ( .A(n16192), .Z(n18143) );
  XNOR U18738 ( .A(n18144), .B(n15028), .Z(n12962) );
  NOR U18739 ( .A(n16188), .B(n16187), .Z(n18144) );
  ANDN U18740 ( .B(n6873), .A(n9963), .Z(n18118) );
  XNOR U18741 ( .A(n13063), .B(n12013), .Z(n9963) );
  XOR U18742 ( .A(n12793), .B(n14759), .Z(n12013) );
  XNOR U18743 ( .A(n18145), .B(n18146), .Z(n14759) );
  XNOR U18744 ( .A(n11871), .B(n12506), .Z(n18146) );
  XOR U18745 ( .A(n18147), .B(n15279), .Z(n12506) );
  ANDN U18746 ( .B(n14761), .A(n14207), .Z(n18147) );
  XNOR U18747 ( .A(n18148), .B(n17440), .Z(n14207) );
  XOR U18748 ( .A(n18149), .B(n16748), .Z(n14761) );
  IV U18749 ( .A(n18150), .Z(n16748) );
  XNOR U18750 ( .A(n18151), .B(n13534), .Z(n11871) );
  ANDN U18751 ( .B(n13535), .A(n13578), .Z(n18151) );
  XOR U18752 ( .A(n18014), .B(n18152), .Z(n13578) );
  XOR U18753 ( .A(n18153), .B(n18154), .Z(n13535) );
  XNOR U18754 ( .A(n9862), .B(n18155), .Z(n18145) );
  XNOR U18755 ( .A(n9758), .B(n12772), .Z(n18155) );
  XOR U18756 ( .A(n18156), .B(n13527), .Z(n12772) );
  ANDN U18757 ( .B(n13528), .A(n13842), .Z(n18156) );
  XNOR U18758 ( .A(n18157), .B(n15948), .Z(n13842) );
  XOR U18759 ( .A(n17028), .B(n18158), .Z(n13528) );
  XNOR U18760 ( .A(n18159), .B(n18160), .Z(n9758) );
  ANDN U18761 ( .B(n13583), .A(n13584), .Z(n18159) );
  XOR U18762 ( .A(n18161), .B(n18162), .Z(n13584) );
  XNOR U18763 ( .A(n18163), .B(n13523), .Z(n9862) );
  ANDN U18764 ( .B(n13588), .A(n13524), .Z(n18163) );
  XOR U18765 ( .A(n18164), .B(n18165), .Z(n13524) );
  XOR U18766 ( .A(n18166), .B(n18167), .Z(n13588) );
  XOR U18767 ( .A(n18168), .B(n18169), .Z(n12793) );
  XNOR U18768 ( .A(n10586), .B(n11628), .Z(n18169) );
  XNOR U18769 ( .A(n18170), .B(n13299), .Z(n11628) );
  IV U18770 ( .A(n13549), .Z(n13299) );
  XNOR U18771 ( .A(n18171), .B(n18172), .Z(n13549) );
  ANDN U18772 ( .B(n13059), .A(n13058), .Z(n18170) );
  XOR U18773 ( .A(n18173), .B(n17297), .Z(n13058) );
  XNOR U18774 ( .A(n18174), .B(n15304), .Z(n13059) );
  XNOR U18775 ( .A(n18175), .B(n13546), .Z(n10586) );
  IV U18776 ( .A(n13923), .Z(n13546) );
  XOR U18777 ( .A(n18176), .B(n18177), .Z(n13923) );
  ANDN U18778 ( .B(n13547), .A(n14392), .Z(n18175) );
  XOR U18779 ( .A(n18178), .B(n17212), .Z(n14392) );
  XNOR U18780 ( .A(n18179), .B(n18180), .Z(n17212) );
  XOR U18781 ( .A(n18181), .B(n18182), .Z(n13547) );
  XOR U18782 ( .A(n13518), .B(n18183), .Z(n18168) );
  XOR U18783 ( .A(n11886), .B(n10230), .Z(n18183) );
  XNOR U18784 ( .A(n18184), .B(n13541), .Z(n10230) );
  IV U18785 ( .A(n13080), .Z(n13541) );
  XNOR U18786 ( .A(n18185), .B(n18186), .Z(n13080) );
  ANDN U18787 ( .B(n13065), .A(n17179), .Z(n18184) );
  IV U18788 ( .A(n13066), .Z(n17179) );
  XNOR U18789 ( .A(n18187), .B(n18188), .Z(n13066) );
  XNOR U18790 ( .A(n18189), .B(n17140), .Z(n13065) );
  XNOR U18791 ( .A(n18190), .B(n13085), .Z(n11886) );
  XNOR U18792 ( .A(n18191), .B(n18192), .Z(n13085) );
  ANDN U18793 ( .B(n13539), .A(n17190), .Z(n18190) );
  XNOR U18794 ( .A(n18193), .B(n13088), .Z(n13518) );
  XOR U18795 ( .A(n18194), .B(n18195), .Z(n13088) );
  ANDN U18796 ( .B(n13054), .A(n13055), .Z(n18193) );
  XNOR U18797 ( .A(n18196), .B(n18197), .Z(n13055) );
  XOR U18798 ( .A(n18198), .B(n17564), .Z(n13054) );
  XOR U18799 ( .A(n18199), .B(n13539), .Z(n13063) );
  XOR U18800 ( .A(n18200), .B(n16732), .Z(n13539) );
  ANDN U18801 ( .B(n17190), .A(n17191), .Z(n18199) );
  XOR U18802 ( .A(n17395), .B(n18201), .Z(n17191) );
  XOR U18803 ( .A(n18202), .B(n17261), .Z(n17190) );
  IV U18804 ( .A(n18203), .Z(n17261) );
  XOR U18805 ( .A(n12787), .B(n16580), .Z(n6873) );
  XOR U18806 ( .A(n18204), .B(n18205), .Z(n16580) );
  ANDN U18807 ( .B(n15313), .A(n15494), .Z(n18204) );
  XOR U18808 ( .A(n18206), .B(n18207), .Z(n15313) );
  XNOR U18809 ( .A(n15163), .B(n12374), .Z(n12787) );
  XNOR U18810 ( .A(n18208), .B(n18209), .Z(n12374) );
  XNOR U18811 ( .A(n12510), .B(n17171), .Z(n18209) );
  XOR U18812 ( .A(n18210), .B(n15305), .Z(n17171) );
  XNOR U18813 ( .A(n18211), .B(n18212), .Z(n15305) );
  AND U18814 ( .A(n13369), .B(n12808), .Z(n18210) );
  XOR U18815 ( .A(n18213), .B(n17240), .Z(n12808) );
  XOR U18816 ( .A(n18214), .B(n16090), .Z(n13369) );
  XOR U18817 ( .A(n18215), .B(n15297), .Z(n12510) );
  XOR U18818 ( .A(n18216), .B(n18217), .Z(n15297) );
  ANDN U18819 ( .B(n12953), .A(n13365), .Z(n18215) );
  XOR U18820 ( .A(n18218), .B(n18219), .Z(n13365) );
  XOR U18821 ( .A(n11683), .B(n18222), .Z(n18208) );
  XOR U18822 ( .A(n13640), .B(n9977), .Z(n18222) );
  XNOR U18823 ( .A(n18223), .B(n15287), .Z(n9977) );
  XOR U18824 ( .A(n18224), .B(n16068), .Z(n15287) );
  ANDN U18825 ( .B(n13367), .A(n12804), .Z(n18223) );
  XOR U18826 ( .A(n18225), .B(n17055), .Z(n12804) );
  XOR U18827 ( .A(n18226), .B(n18227), .Z(n13367) );
  XNOR U18828 ( .A(n18228), .B(n15291), .Z(n13640) );
  XNOR U18829 ( .A(n18229), .B(n18195), .Z(n15291) );
  NOR U18830 ( .A(n13358), .B(n13360), .Z(n18228) );
  XNOR U18831 ( .A(n18230), .B(n15635), .Z(n13360) );
  XOR U18832 ( .A(n17338), .B(n18231), .Z(n13358) );
  XNOR U18833 ( .A(n18232), .B(n15301), .Z(n11683) );
  XNOR U18834 ( .A(n18233), .B(n18234), .Z(n15301) );
  AND U18835 ( .A(n12798), .B(n13362), .Z(n18232) );
  XNOR U18836 ( .A(n18235), .B(n17105), .Z(n13362) );
  XOR U18837 ( .A(n18236), .B(n18237), .Z(n12798) );
  XOR U18838 ( .A(n18238), .B(n18239), .Z(n15163) );
  XOR U18839 ( .A(n12275), .B(n12623), .Z(n18239) );
  XNOR U18840 ( .A(n18240), .B(n15319), .Z(n12623) );
  IV U18841 ( .A(n18241), .Z(n15319) );
  ANDN U18842 ( .B(n15490), .A(n16583), .Z(n18240) );
  XOR U18843 ( .A(n18242), .B(n16825), .Z(n15490) );
  XOR U18844 ( .A(n18243), .B(n15311), .Z(n12275) );
  ANDN U18845 ( .B(n16587), .A(n15492), .Z(n18243) );
  XOR U18846 ( .A(n18244), .B(n17215), .Z(n15492) );
  XNOR U18847 ( .A(n12294), .B(n18245), .Z(n18238) );
  XOR U18848 ( .A(n11943), .B(n11195), .Z(n18245) );
  XOR U18849 ( .A(n18246), .B(n15327), .Z(n11195) );
  ANDN U18850 ( .B(n16573), .A(n15487), .Z(n18246) );
  XOR U18851 ( .A(n18247), .B(n18248), .Z(n15487) );
  XNOR U18852 ( .A(n18249), .B(n15315), .Z(n11943) );
  IV U18853 ( .A(n18250), .Z(n15315) );
  ANDN U18854 ( .B(n15494), .A(n18205), .Z(n18249) );
  XOR U18855 ( .A(n18251), .B(n16616), .Z(n15494) );
  XOR U18856 ( .A(n18252), .B(n15323), .Z(n12294) );
  ANDN U18857 ( .B(n16577), .A(n15484), .Z(n18252) );
  XNOR U18858 ( .A(n18253), .B(n18154), .Z(n15484) );
  XNOR U18859 ( .A(n18254), .B(n6877), .Z(n3345) );
  XOR U18860 ( .A(n17317), .B(n9147), .Z(n6877) );
  IV U18861 ( .A(n10488), .Z(n9147) );
  XNOR U18862 ( .A(n18255), .B(n13394), .Z(n10488) );
  XOR U18863 ( .A(n18256), .B(n18257), .Z(n13394) );
  XNOR U18864 ( .A(n10517), .B(n10261), .Z(n18257) );
  XNOR U18865 ( .A(n18258), .B(n13991), .Z(n10261) );
  XOR U18866 ( .A(n18259), .B(n18260), .Z(n13991) );
  ANDN U18867 ( .B(n15892), .A(n15849), .Z(n18258) );
  XNOR U18868 ( .A(n18261), .B(n13998), .Z(n10517) );
  XNOR U18869 ( .A(n18262), .B(n17606), .Z(n13998) );
  IV U18870 ( .A(n17055), .Z(n17606) );
  NOR U18871 ( .A(n15838), .B(n15895), .Z(n18261) );
  XNOR U18872 ( .A(n15645), .B(n18265), .Z(n15895) );
  XOR U18873 ( .A(n18266), .B(n18267), .Z(n15838) );
  XOR U18874 ( .A(n10291), .B(n18268), .Z(n18256) );
  XOR U18875 ( .A(n9629), .B(n10535), .Z(n18268) );
  XNOR U18876 ( .A(n18269), .B(n13994), .Z(n10535) );
  XOR U18877 ( .A(n18270), .B(n15883), .Z(n13994) );
  ANDN U18878 ( .B(n15905), .A(n15843), .Z(n18269) );
  XOR U18879 ( .A(n18271), .B(n16767), .Z(n15843) );
  XNOR U18880 ( .A(n17467), .B(n18272), .Z(n15905) );
  XNOR U18881 ( .A(n18273), .B(n13985), .Z(n9629) );
  XOR U18882 ( .A(n18274), .B(n18275), .Z(n13985) );
  ANDN U18883 ( .B(n15908), .A(n15840), .Z(n18273) );
  IV U18884 ( .A(n17314), .Z(n15840) );
  XOR U18885 ( .A(n17338), .B(n18278), .Z(n15908) );
  XNOR U18886 ( .A(n18279), .B(n15901), .Z(n10291) );
  IV U18887 ( .A(n13981), .Z(n15901) );
  XNOR U18888 ( .A(n18280), .B(n17013), .Z(n13981) );
  ANDN U18889 ( .B(n15846), .A(n15900), .Z(n18279) );
  XNOR U18890 ( .A(n18281), .B(n18282), .Z(n15900) );
  XOR U18891 ( .A(n18283), .B(n18284), .Z(n15846) );
  XNOR U18892 ( .A(n18285), .B(n15892), .Z(n17317) );
  XOR U18893 ( .A(n18286), .B(n18287), .Z(n15892) );
  AND U18894 ( .A(n15849), .B(n13989), .Z(n18285) );
  XNOR U18895 ( .A(n18288), .B(n18289), .Z(n13989) );
  XOR U18896 ( .A(n17395), .B(n18290), .Z(n15849) );
  ANDN U18897 ( .B(n7672), .A(n7671), .Z(n18254) );
  XOR U18898 ( .A(n13741), .B(n9664), .Z(n7671) );
  XNOR U18899 ( .A(n15059), .B(n14489), .Z(n9664) );
  XNOR U18900 ( .A(n18291), .B(n18292), .Z(n14489) );
  XNOR U18901 ( .A(n11233), .B(n14517), .Z(n18292) );
  XNOR U18902 ( .A(n18293), .B(n15447), .Z(n14517) );
  XOR U18903 ( .A(n18294), .B(n18295), .Z(n15447) );
  ANDN U18904 ( .B(n14252), .A(n15448), .Z(n18293) );
  XNOR U18905 ( .A(n18296), .B(n15453), .Z(n11233) );
  XNOR U18906 ( .A(n16957), .B(n18297), .Z(n15453) );
  ANDN U18907 ( .B(n13752), .A(n13753), .Z(n18296) );
  XNOR U18908 ( .A(n18298), .B(n16078), .Z(n13753) );
  XOR U18909 ( .A(n17246), .B(n18299), .Z(n13752) );
  XOR U18910 ( .A(n12840), .B(n18300), .Z(n18291) );
  XOR U18911 ( .A(n10603), .B(n10731), .Z(n18300) );
  XNOR U18912 ( .A(n18301), .B(n15591), .Z(n10731) );
  IV U18913 ( .A(n16990), .Z(n15591) );
  XOR U18914 ( .A(n18302), .B(n18303), .Z(n16990) );
  ANDN U18915 ( .B(n13756), .A(n14246), .Z(n18301) );
  XOR U18916 ( .A(n18304), .B(n17436), .Z(n14246) );
  IV U18917 ( .A(n14172), .Z(n17436) );
  XNOR U18918 ( .A(n18305), .B(n17613), .Z(n13756) );
  XOR U18919 ( .A(n18306), .B(n15451), .Z(n10603) );
  XOR U18920 ( .A(n18307), .B(n16522), .Z(n15451) );
  ANDN U18921 ( .B(n13743), .A(n14241), .Z(n18306) );
  IV U18922 ( .A(n13745), .Z(n14241) );
  XOR U18923 ( .A(n18308), .B(n18309), .Z(n13745) );
  XNOR U18924 ( .A(n18310), .B(n16008), .Z(n13743) );
  XNOR U18925 ( .A(n18311), .B(n15455), .Z(n12840) );
  XOR U18926 ( .A(n18312), .B(n16872), .Z(n15455) );
  NOR U18927 ( .A(n14238), .B(n13748), .Z(n18311) );
  XNOR U18928 ( .A(n18313), .B(n18314), .Z(n13748) );
  XOR U18929 ( .A(n18315), .B(n17024), .Z(n14238) );
  XOR U18930 ( .A(n18316), .B(n18317), .Z(n15059) );
  XOR U18931 ( .A(n9885), .B(n10737), .Z(n18317) );
  XNOR U18932 ( .A(n18318), .B(n17639), .Z(n10737) );
  IV U18933 ( .A(n14538), .Z(n17639) );
  XNOR U18934 ( .A(n18319), .B(n15339), .Z(n14538) );
  ANDN U18935 ( .B(n15552), .A(n14537), .Z(n18318) );
  XNOR U18936 ( .A(n18320), .B(n17740), .Z(n14537) );
  XNOR U18937 ( .A(n18321), .B(n18322), .Z(n15552) );
  XNOR U18938 ( .A(n18323), .B(n14524), .Z(n9885) );
  XNOR U18939 ( .A(n18324), .B(n16813), .Z(n14524) );
  ANDN U18940 ( .B(n15555), .A(n14523), .Z(n18323) );
  XOR U18941 ( .A(n18325), .B(n18326), .Z(n14523) );
  XOR U18942 ( .A(n18327), .B(n17306), .Z(n15555) );
  XNOR U18943 ( .A(n13417), .B(n18328), .Z(n18316) );
  XNOR U18944 ( .A(n12638), .B(n11336), .Z(n18328) );
  XNOR U18945 ( .A(n18329), .B(n14533), .Z(n11336) );
  XNOR U18946 ( .A(n18330), .B(n17586), .Z(n14533) );
  ANDN U18947 ( .B(n15563), .A(n15561), .Z(n18329) );
  XOR U18948 ( .A(n18331), .B(n18332), .Z(n15561) );
  XOR U18949 ( .A(n18333), .B(n16078), .Z(n15563) );
  XNOR U18950 ( .A(n18334), .B(n17615), .Z(n12638) );
  XOR U18951 ( .A(n18335), .B(n16744), .Z(n17615) );
  NOR U18952 ( .A(n16324), .B(n15565), .Z(n18334) );
  XNOR U18953 ( .A(n18336), .B(n18337), .Z(n15565) );
  IV U18954 ( .A(n15567), .Z(n16324) );
  XOR U18955 ( .A(n18338), .B(n17750), .Z(n15567) );
  XOR U18956 ( .A(n18339), .B(n14528), .Z(n13417) );
  XOR U18957 ( .A(n18340), .B(n17188), .Z(n14528) );
  NOR U18958 ( .A(n16320), .B(n14527), .Z(n18339) );
  XOR U18959 ( .A(n18341), .B(n14172), .Z(n14527) );
  XOR U18960 ( .A(n18342), .B(n18343), .Z(n14172) );
  IV U18961 ( .A(n15559), .Z(n16320) );
  XOR U18962 ( .A(n18344), .B(n14967), .Z(n15559) );
  XNOR U18963 ( .A(n18345), .B(n15448), .Z(n13741) );
  XOR U18964 ( .A(n18346), .B(n15899), .Z(n15448) );
  ANDN U18965 ( .B(n14253), .A(n14252), .Z(n18345) );
  XOR U18966 ( .A(n18347), .B(n17402), .Z(n14252) );
  IV U18967 ( .A(n17240), .Z(n17402) );
  XOR U18968 ( .A(n17026), .B(n18348), .Z(n14253) );
  XNOR U18969 ( .A(n17755), .B(n11902), .Z(n7672) );
  XOR U18970 ( .A(n18349), .B(n18350), .Z(n17755) );
  AND U18971 ( .A(n18351), .B(n18352), .Z(n18349) );
  XOR U18972 ( .A(n18353), .B(n18354), .Z(n5992) );
  XNOR U18973 ( .A(n1851), .B(n5228), .Z(n18354) );
  XOR U18974 ( .A(n18355), .B(n7731), .Z(n5228) );
  XOR U18975 ( .A(n17713), .B(n11688), .Z(n7731) );
  IV U18976 ( .A(n11221), .Z(n11688) );
  XNOR U18977 ( .A(n14982), .B(n12910), .Z(n11221) );
  XNOR U18978 ( .A(n18356), .B(n18357), .Z(n12910) );
  XOR U18979 ( .A(n11951), .B(n11551), .Z(n18357) );
  XOR U18980 ( .A(n18358), .B(n15728), .Z(n11551) );
  ANDN U18981 ( .B(n17719), .A(n18359), .Z(n18358) );
  XNOR U18982 ( .A(n15342), .B(n18360), .Z(n17719) );
  XNOR U18983 ( .A(n18361), .B(n15720), .Z(n11951) );
  ANDN U18984 ( .B(n17715), .A(n17716), .Z(n18361) );
  XNOR U18985 ( .A(n18362), .B(n17970), .Z(n17716) );
  XOR U18986 ( .A(n10760), .B(n18363), .Z(n18356) );
  XOR U18987 ( .A(n11974), .B(n11591), .Z(n18363) );
  XOR U18988 ( .A(n18364), .B(n15712), .Z(n11591) );
  AND U18989 ( .A(n18093), .B(n18365), .Z(n18364) );
  XNOR U18990 ( .A(n18366), .B(n15725), .Z(n11974) );
  ANDN U18991 ( .B(n17706), .A(n17707), .Z(n18366) );
  XNOR U18992 ( .A(n18368), .B(n15715), .Z(n10760) );
  ANDN U18993 ( .B(n17711), .A(n17709), .Z(n18368) );
  XOR U18994 ( .A(n18370), .B(n18371), .Z(n14982) );
  XOR U18995 ( .A(n9230), .B(n14153), .Z(n18371) );
  XOR U18996 ( .A(n18373), .B(n18374), .Z(n13255) );
  ANDN U18997 ( .B(n14140), .A(n14169), .Z(n18372) );
  XOR U18998 ( .A(n18375), .B(n15528), .Z(n14169) );
  XOR U18999 ( .A(n18376), .B(n15290), .Z(n14140) );
  XNOR U19000 ( .A(n18377), .B(n13267), .Z(n9230) );
  XOR U19001 ( .A(n18378), .B(n18379), .Z(n13267) );
  ANDN U19002 ( .B(n14164), .A(n14149), .Z(n18377) );
  XNOR U19003 ( .A(n18380), .B(n18381), .Z(n14149) );
  XOR U19004 ( .A(n16399), .B(n18382), .Z(n14164) );
  XOR U19005 ( .A(n10294), .B(n18383), .Z(n18370) );
  XOR U19006 ( .A(n9622), .B(n10270), .Z(n18383) );
  XNOR U19007 ( .A(n18384), .B(n13250), .Z(n10270) );
  XNOR U19008 ( .A(n18385), .B(n16105), .Z(n13250) );
  ANDN U19009 ( .B(n14142), .A(n15349), .Z(n18384) );
  IV U19010 ( .A(n14177), .Z(n15349) );
  XOR U19011 ( .A(n18386), .B(n18387), .Z(n14177) );
  XOR U19012 ( .A(n18388), .B(n16058), .Z(n14142) );
  XOR U19013 ( .A(n18389), .B(n13259), .Z(n9622) );
  XOR U19014 ( .A(n18390), .B(n14967), .Z(n13259) );
  NOR U19015 ( .A(n15334), .B(n14145), .Z(n18389) );
  XOR U19016 ( .A(n18391), .B(n17301), .Z(n14145) );
  XOR U19017 ( .A(n18392), .B(n14996), .Z(n15334) );
  IV U19018 ( .A(n16096), .Z(n14996) );
  XOR U19019 ( .A(n18393), .B(n18394), .Z(n16096) );
  XNOR U19020 ( .A(n18395), .B(n13263), .Z(n10294) );
  XOR U19021 ( .A(n18396), .B(n18397), .Z(n13263) );
  ANDN U19022 ( .B(n14147), .A(n15345), .Z(n18395) );
  XOR U19023 ( .A(n18398), .B(n16575), .Z(n15345) );
  XOR U19024 ( .A(n18399), .B(n18400), .Z(n14147) );
  XOR U19025 ( .A(n18401), .B(n18365), .Z(n17713) );
  ANDN U19026 ( .B(n15710), .A(n18093), .Z(n18401) );
  XOR U19027 ( .A(n16097), .B(n18402), .Z(n18093) );
  IV U19028 ( .A(n18403), .Z(n16097) );
  XOR U19029 ( .A(n18404), .B(n17788), .Z(n15710) );
  ANDN U19030 ( .B(n6907), .A(n7732), .Z(n18355) );
  XOR U19031 ( .A(n18405), .B(n10198), .Z(n7732) );
  XNOR U19032 ( .A(n18406), .B(n16179), .Z(n10198) );
  XNOR U19033 ( .A(n18407), .B(n18408), .Z(n16179) );
  XNOR U19034 ( .A(n12924), .B(n11931), .Z(n18408) );
  XOR U19035 ( .A(n18409), .B(n16386), .Z(n11931) );
  IV U19036 ( .A(n16414), .Z(n16386) );
  XNOR U19037 ( .A(n18410), .B(n16744), .Z(n16414) );
  ANDN U19038 ( .B(n15599), .A(n16413), .Z(n18409) );
  XNOR U19039 ( .A(n18411), .B(n14825), .Z(n12924) );
  XOR U19040 ( .A(n18412), .B(n18413), .Z(n14825) );
  AND U19041 ( .A(n15614), .B(n14826), .Z(n18411) );
  XNOR U19042 ( .A(n13038), .B(n18414), .Z(n18407) );
  XOR U19043 ( .A(n9444), .B(n9561), .Z(n18414) );
  XOR U19044 ( .A(n18415), .B(n15858), .Z(n9561) );
  XNOR U19045 ( .A(n18416), .B(n17294), .Z(n15858) );
  ANDN U19046 ( .B(n15859), .A(n15603), .Z(n18415) );
  XNOR U19047 ( .A(n18417), .B(n14818), .Z(n9444) );
  XOR U19048 ( .A(n18418), .B(n18419), .Z(n14818) );
  ANDN U19049 ( .B(n14819), .A(n15611), .Z(n18417) );
  XNOR U19050 ( .A(n18420), .B(n16373), .Z(n13038) );
  IV U19051 ( .A(n14814), .Z(n16373) );
  XOR U19052 ( .A(n18421), .B(n18422), .Z(n14814) );
  ANDN U19053 ( .B(n14815), .A(n15608), .Z(n18420) );
  XOR U19054 ( .A(n11637), .B(n13425), .Z(n6907) );
  XNOR U19055 ( .A(n18423), .B(n16849), .Z(n13425) );
  ANDN U19056 ( .B(n14027), .A(n16041), .Z(n18423) );
  IV U19057 ( .A(n14028), .Z(n16041) );
  XOR U19058 ( .A(n18424), .B(n16331), .Z(n14028) );
  XNOR U19059 ( .A(n13634), .B(n12817), .Z(n11637) );
  XOR U19060 ( .A(n18425), .B(n18426), .Z(n12817) );
  XNOR U19061 ( .A(n11795), .B(n9328), .Z(n18426) );
  XOR U19062 ( .A(n18427), .B(n14063), .Z(n9328) );
  XNOR U19063 ( .A(n18428), .B(n18429), .Z(n14063) );
  ANDN U19064 ( .B(n14064), .A(n15220), .Z(n18427) );
  XOR U19065 ( .A(n17180), .B(n18430), .Z(n14064) );
  XOR U19066 ( .A(n18431), .B(n14049), .Z(n11795) );
  XNOR U19067 ( .A(n18432), .B(n18433), .Z(n14050) );
  XOR U19068 ( .A(n10258), .B(n18434), .Z(n18425) );
  XOR U19069 ( .A(n11203), .B(n14044), .Z(n18434) );
  XNOR U19070 ( .A(n18435), .B(n14053), .Z(n14044) );
  IV U19071 ( .A(n15757), .Z(n14053) );
  XOR U19072 ( .A(n14158), .B(n18436), .Z(n15757) );
  ANDN U19073 ( .B(n15223), .A(n15222), .Z(n18435) );
  IV U19074 ( .A(n14054), .Z(n15222) );
  XOR U19075 ( .A(n18437), .B(n18438), .Z(n14054) );
  XNOR U19076 ( .A(n18439), .B(n15759), .Z(n11203) );
  IV U19077 ( .A(n14060), .Z(n15759) );
  XNOR U19078 ( .A(n18440), .B(n17589), .Z(n14060) );
  NOR U19079 ( .A(n15212), .B(n14059), .Z(n18439) );
  XNOR U19080 ( .A(n18441), .B(n18442), .Z(n14059) );
  XOR U19081 ( .A(n18443), .B(n15749), .Z(n10258) );
  XNOR U19082 ( .A(n18444), .B(n18445), .Z(n15749) );
  XOR U19083 ( .A(n16600), .B(n18446), .Z(n15214) );
  XOR U19084 ( .A(n18447), .B(n18448), .Z(n13634) );
  XOR U19085 ( .A(n10337), .B(n9971), .Z(n18448) );
  XOR U19086 ( .A(n18449), .B(n16042), .Z(n9971) );
  XOR U19087 ( .A(n18450), .B(n17506), .Z(n16042) );
  XOR U19088 ( .A(n18451), .B(n18452), .Z(n14027) );
  XOR U19089 ( .A(n15694), .B(n18453), .Z(n16849) );
  XOR U19090 ( .A(n18454), .B(n16038), .Z(n10337) );
  XNOR U19091 ( .A(n18455), .B(n18456), .Z(n16038) );
  NOR U19092 ( .A(n14034), .B(n14899), .Z(n18454) );
  XNOR U19093 ( .A(n18457), .B(n18458), .Z(n14899) );
  XOR U19094 ( .A(n18459), .B(n15269), .Z(n14034) );
  IV U19095 ( .A(n16154), .Z(n15269) );
  XOR U19096 ( .A(n11705), .B(n18462), .Z(n18447) );
  XOR U19097 ( .A(n10853), .B(n11695), .Z(n18462) );
  XNOR U19098 ( .A(n18463), .B(n16050), .Z(n11695) );
  XOR U19099 ( .A(n18464), .B(n18465), .Z(n16050) );
  ANDN U19100 ( .B(n13439), .A(n13437), .Z(n18463) );
  IV U19101 ( .A(n16853), .Z(n13437) );
  XNOR U19102 ( .A(n18466), .B(n17333), .Z(n16853) );
  XNOR U19103 ( .A(n18467), .B(n18468), .Z(n13439) );
  XNOR U19104 ( .A(n18469), .B(n16046), .Z(n10853) );
  XOR U19105 ( .A(n18470), .B(n17916), .Z(n16046) );
  NOR U19106 ( .A(n13427), .B(n13428), .Z(n18469) );
  XNOR U19107 ( .A(n18171), .B(n18471), .Z(n13428) );
  XOR U19108 ( .A(n18472), .B(n18473), .Z(n13427) );
  XOR U19109 ( .A(n18474), .B(n16033), .Z(n11705) );
  XOR U19110 ( .A(n17287), .B(n18475), .Z(n16033) );
  IV U19111 ( .A(n18476), .Z(n17287) );
  NOR U19112 ( .A(n13434), .B(n13433), .Z(n18474) );
  XOR U19113 ( .A(n18477), .B(n18478), .Z(n13433) );
  XNOR U19114 ( .A(n18479), .B(n18480), .Z(n13434) );
  XOR U19115 ( .A(n18481), .B(n7725), .Z(n1851) );
  XNOR U19116 ( .A(n9452), .B(n16536), .Z(n7725) );
  XNOR U19117 ( .A(n18482), .B(n14783), .Z(n16536) );
  NOR U19118 ( .A(n17775), .B(n18483), .Z(n18482) );
  IV U19119 ( .A(n14178), .Z(n9452) );
  XOR U19120 ( .A(n18059), .B(n18484), .Z(n14178) );
  XOR U19121 ( .A(n18485), .B(n18486), .Z(n18059) );
  XNOR U19122 ( .A(n11082), .B(n12021), .Z(n18486) );
  XNOR U19123 ( .A(n18487), .B(n15005), .Z(n12021) );
  XOR U19124 ( .A(n18488), .B(n17429), .Z(n15005) );
  NOR U19125 ( .A(n15004), .B(n17327), .Z(n18487) );
  XNOR U19126 ( .A(n18489), .B(n18203), .Z(n17327) );
  XOR U19127 ( .A(n18090), .B(n18490), .Z(n15004) );
  XNOR U19128 ( .A(n18491), .B(n16336), .Z(n11082) );
  XOR U19129 ( .A(n18492), .B(n17392), .Z(n16336) );
  XNOR U19130 ( .A(n18493), .B(n17432), .Z(n16880) );
  XOR U19131 ( .A(n18494), .B(n16074), .Z(n16337) );
  XOR U19132 ( .A(n11905), .B(n18495), .Z(n18485) );
  XNOR U19133 ( .A(n9120), .B(n10843), .Z(n18495) );
  XNOR U19134 ( .A(n18496), .B(n14796), .Z(n10843) );
  XNOR U19135 ( .A(n16809), .B(n18497), .Z(n14796) );
  ANDN U19136 ( .B(n14797), .A(n16870), .Z(n18496) );
  XNOR U19137 ( .A(n18498), .B(n17229), .Z(n16870) );
  XNOR U19138 ( .A(n16004), .B(n18499), .Z(n14797) );
  XNOR U19139 ( .A(n18500), .B(n16358), .Z(n9120) );
  XOR U19140 ( .A(n18501), .B(n18502), .Z(n16358) );
  ANDN U19141 ( .B(n14804), .A(n16866), .Z(n18500) );
  XOR U19142 ( .A(n17180), .B(n18503), .Z(n16866) );
  IV U19143 ( .A(n14970), .Z(n17180) );
  XOR U19144 ( .A(n18504), .B(n18237), .Z(n14804) );
  XOR U19145 ( .A(n18505), .B(n14792), .Z(n11905) );
  XOR U19146 ( .A(n18506), .B(n15351), .Z(n14792) );
  ANDN U19147 ( .B(n14793), .A(n16876), .Z(n18505) );
  IV U19148 ( .A(n17331), .Z(n16876) );
  XOR U19149 ( .A(n18507), .B(n18508), .Z(n17331) );
  XOR U19150 ( .A(n18509), .B(n18458), .Z(n14793) );
  ANDN U19151 ( .B(n6899), .A(n7726), .Z(n18481) );
  XNOR U19152 ( .A(n16015), .B(n12220), .Z(n7726) );
  XNOR U19153 ( .A(n18510), .B(n17721), .Z(n12220) );
  XNOR U19154 ( .A(n18511), .B(n18512), .Z(n17721) );
  XOR U19155 ( .A(n12643), .B(n12321), .Z(n18512) );
  XNOR U19156 ( .A(n18513), .B(n17675), .Z(n12321) );
  XOR U19157 ( .A(n18514), .B(n16813), .Z(n17675) );
  AND U19158 ( .A(n12451), .B(n12449), .Z(n18513) );
  XOR U19159 ( .A(n15875), .B(n18515), .Z(n12449) );
  XOR U19160 ( .A(n18516), .B(n18517), .Z(n12451) );
  XNOR U19161 ( .A(n18518), .B(n16138), .Z(n12643) );
  XOR U19162 ( .A(n18519), .B(n17699), .Z(n16138) );
  NOR U19163 ( .A(n13697), .B(n13698), .Z(n18518) );
  XOR U19164 ( .A(n18520), .B(n18521), .Z(n13698) );
  XOR U19165 ( .A(n18522), .B(n18523), .Z(n13697) );
  XOR U19166 ( .A(n11234), .B(n18524), .Z(n18511) );
  XNOR U19167 ( .A(n12669), .B(n12377), .Z(n18524) );
  XNOR U19168 ( .A(n18525), .B(n16125), .Z(n12377) );
  XNOR U19169 ( .A(n18526), .B(n16529), .Z(n16125) );
  AND U19170 ( .A(n17680), .B(n17723), .Z(n18525) );
  XNOR U19171 ( .A(n16600), .B(n18527), .Z(n17723) );
  XOR U19172 ( .A(n18528), .B(n18445), .Z(n17680) );
  XNOR U19173 ( .A(n18529), .B(n16135), .Z(n12669) );
  XOR U19174 ( .A(n18530), .B(n18531), .Z(n16135) );
  NOR U19175 ( .A(n14445), .B(n14446), .Z(n18529) );
  XNOR U19176 ( .A(n18532), .B(n16668), .Z(n14446) );
  IV U19177 ( .A(n17683), .Z(n14445) );
  XNOR U19178 ( .A(n18533), .B(n16579), .Z(n17683) );
  XNOR U19179 ( .A(n18534), .B(n16129), .Z(n11234) );
  XOR U19180 ( .A(n18535), .B(n18078), .Z(n16129) );
  ANDN U19181 ( .B(n12460), .A(n12461), .Z(n18534) );
  XOR U19182 ( .A(n18536), .B(n16504), .Z(n12461) );
  XNOR U19183 ( .A(n18537), .B(n16058), .Z(n12460) );
  XNOR U19184 ( .A(n18538), .B(n17694), .Z(n16015) );
  ANDN U19185 ( .B(n14555), .A(n14556), .Z(n18538) );
  XNOR U19186 ( .A(n18539), .B(n18540), .Z(n14556) );
  XNOR U19187 ( .A(n18541), .B(n9244), .Z(n6899) );
  XOR U19188 ( .A(n18542), .B(n16657), .Z(n9244) );
  XOR U19189 ( .A(n18543), .B(n18544), .Z(n16657) );
  XNOR U19190 ( .A(n14112), .B(n10644), .Z(n18544) );
  XNOR U19191 ( .A(n18545), .B(n18546), .Z(n10644) );
  ANDN U19192 ( .B(n17825), .A(n17823), .Z(n18545) );
  XOR U19193 ( .A(n18547), .B(n16998), .Z(n17825) );
  XNOR U19194 ( .A(n18548), .B(n14258), .Z(n14112) );
  ANDN U19195 ( .B(n17828), .A(n14257), .Z(n18548) );
  XOR U19196 ( .A(n18549), .B(n17861), .Z(n14257) );
  XNOR U19197 ( .A(n15196), .B(n18550), .Z(n17828) );
  XNOR U19198 ( .A(n10532), .B(n18553), .Z(n18543) );
  XOR U19199 ( .A(n10051), .B(n9779), .Z(n18553) );
  XOR U19200 ( .A(n18554), .B(n15099), .Z(n9779) );
  ANDN U19201 ( .B(n17831), .A(n15100), .Z(n18554) );
  XNOR U19202 ( .A(n18555), .B(n17898), .Z(n15100) );
  XNOR U19203 ( .A(n18556), .B(n18557), .Z(n17831) );
  XNOR U19204 ( .A(n18558), .B(n18559), .Z(n10051) );
  NOR U19205 ( .A(n17882), .B(n17818), .Z(n18558) );
  XOR U19206 ( .A(n18560), .B(n18561), .Z(n17882) );
  XOR U19207 ( .A(n18562), .B(n14119), .Z(n10532) );
  NOR U19208 ( .A(n17887), .B(n14120), .Z(n18562) );
  XOR U19209 ( .A(n18563), .B(n18564), .Z(n14120) );
  XOR U19210 ( .A(n18565), .B(n18150), .Z(n17887) );
  XOR U19211 ( .A(n4134), .B(n18566), .Z(n18353) );
  XOR U19212 ( .A(n7705), .B(n3636), .Z(n18566) );
  XOR U19213 ( .A(n18567), .B(n10091), .Z(n3636) );
  XOR U19214 ( .A(n13531), .B(n12169), .Z(n10091) );
  IV U19215 ( .A(n10759), .Z(n12169) );
  XNOR U19216 ( .A(n13074), .B(n18568), .Z(n10759) );
  XOR U19217 ( .A(n18569), .B(n18570), .Z(n13074) );
  XNOR U19218 ( .A(n11789), .B(n11956), .Z(n18570) );
  XOR U19219 ( .A(n18571), .B(n13843), .Z(n11956) );
  XNOR U19220 ( .A(n14158), .B(n18572), .Z(n13843) );
  ANDN U19221 ( .B(n13527), .A(n13526), .Z(n18571) );
  XNOR U19222 ( .A(n18573), .B(n17013), .Z(n13526) );
  XOR U19223 ( .A(n18574), .B(n17186), .Z(n13527) );
  XNOR U19224 ( .A(n18575), .B(n14209), .Z(n11789) );
  IV U19225 ( .A(n14762), .Z(n14209) );
  XOR U19226 ( .A(n18576), .B(n18577), .Z(n14762) );
  ANDN U19227 ( .B(n15279), .A(n14208), .Z(n18575) );
  XOR U19228 ( .A(n18578), .B(n18579), .Z(n14208) );
  XOR U19229 ( .A(n18580), .B(n18192), .Z(n15279) );
  XOR U19230 ( .A(n14201), .B(n18581), .Z(n18569) );
  XOR U19231 ( .A(n11450), .B(n10356), .Z(n18581) );
  XNOR U19232 ( .A(n18582), .B(n13579), .Z(n10356) );
  XNOR U19233 ( .A(n18583), .B(n18422), .Z(n13579) );
  NOR U19234 ( .A(n13533), .B(n13534), .Z(n18582) );
  XNOR U19235 ( .A(n15674), .B(n18584), .Z(n13534) );
  IV U19236 ( .A(n14213), .Z(n13533) );
  XOR U19237 ( .A(n18585), .B(n18586), .Z(n14213) );
  XOR U19238 ( .A(n18587), .B(n13585), .Z(n11450) );
  XNOR U19239 ( .A(n18588), .B(n15891), .Z(n13585) );
  NOR U19240 ( .A(n18160), .B(n14205), .Z(n18587) );
  IV U19241 ( .A(n18589), .Z(n18160) );
  XNOR U19242 ( .A(n18590), .B(n13587), .Z(n14201) );
  XOR U19243 ( .A(n18591), .B(n17516), .Z(n13587) );
  NOR U19244 ( .A(n13523), .B(n13522), .Z(n18590) );
  XOR U19245 ( .A(n18592), .B(n17958), .Z(n13522) );
  XOR U19246 ( .A(n15956), .B(n18593), .Z(n13523) );
  XNOR U19247 ( .A(n18594), .B(n14205), .Z(n13531) );
  XOR U19248 ( .A(n18595), .B(n15256), .Z(n14205) );
  NOR U19249 ( .A(n18589), .B(n13583), .Z(n18594) );
  XOR U19250 ( .A(n18596), .B(n18597), .Z(n13583) );
  XOR U19251 ( .A(n18598), .B(n18599), .Z(n18589) );
  NOR U19252 ( .A(n10126), .B(n6895), .Z(n18567) );
  XOR U19253 ( .A(n14093), .B(n9336), .Z(n6895) );
  XOR U19254 ( .A(n13912), .B(n13925), .Z(n9336) );
  XNOR U19255 ( .A(n18600), .B(n18601), .Z(n13925) );
  XNOR U19256 ( .A(n12184), .B(n13304), .Z(n18601) );
  XNOR U19257 ( .A(n18602), .B(n18603), .Z(n13304) );
  ANDN U19258 ( .B(n15828), .A(n14919), .Z(n18602) );
  XNOR U19259 ( .A(n18604), .B(n18468), .Z(n14919) );
  XNOR U19260 ( .A(n18605), .B(n17390), .Z(n15828) );
  IV U19261 ( .A(n16115), .Z(n17390) );
  XOR U19262 ( .A(n18606), .B(n18607), .Z(n16115) );
  XNOR U19263 ( .A(n18608), .B(n14914), .Z(n12184) );
  IV U19264 ( .A(n18609), .Z(n14914) );
  NOR U19265 ( .A(n16794), .B(n14913), .Z(n18608) );
  XNOR U19266 ( .A(n18610), .B(n18611), .Z(n14913) );
  XOR U19267 ( .A(n18612), .B(n18613), .Z(n16794) );
  XOR U19268 ( .A(n11090), .B(n18614), .Z(n18600) );
  XOR U19269 ( .A(n10867), .B(n11731), .Z(n18614) );
  XNOR U19270 ( .A(n18615), .B(n14909), .Z(n11731) );
  IV U19271 ( .A(n18616), .Z(n14909) );
  ANDN U19272 ( .B(n14910), .A(n15823), .Z(n18615) );
  XNOR U19273 ( .A(n18617), .B(n16045), .Z(n15823) );
  XOR U19274 ( .A(n18277), .B(n18618), .Z(n14910) );
  XNOR U19275 ( .A(n18619), .B(n14923), .Z(n10867) );
  ANDN U19276 ( .B(n14924), .A(n16799), .Z(n18619) );
  XOR U19277 ( .A(n18620), .B(n16149), .Z(n16799) );
  XNOR U19278 ( .A(n18621), .B(n18622), .Z(n14924) );
  XNOR U19279 ( .A(n18623), .B(n18624), .Z(n11090) );
  ANDN U19280 ( .B(n15819), .A(n16792), .Z(n18623) );
  XNOR U19281 ( .A(n18027), .B(n18625), .Z(n15819) );
  XOR U19282 ( .A(n18626), .B(n18627), .Z(n13912) );
  XOR U19283 ( .A(n9794), .B(n12791), .Z(n18627) );
  XNOR U19284 ( .A(n18628), .B(n14743), .Z(n12791) );
  IV U19285 ( .A(n15735), .Z(n14743) );
  XOR U19286 ( .A(n18629), .B(n17994), .Z(n15735) );
  NOR U19287 ( .A(n14108), .B(n14109), .Z(n18628) );
  XNOR U19288 ( .A(n18630), .B(n17613), .Z(n14108) );
  XNOR U19289 ( .A(n18631), .B(n14753), .Z(n9794) );
  XNOR U19290 ( .A(n18632), .B(n18177), .Z(n14753) );
  ANDN U19291 ( .B(n18633), .A(n15738), .Z(n18631) );
  XNOR U19292 ( .A(n14903), .B(n18634), .Z(n18626) );
  XNOR U19293 ( .A(n9814), .B(n12619), .Z(n18634) );
  XNOR U19294 ( .A(n18635), .B(n14747), .Z(n12619) );
  IV U19295 ( .A(n15744), .Z(n14747) );
  XOR U19296 ( .A(n15951), .B(n18636), .Z(n15744) );
  IV U19297 ( .A(n16399), .Z(n15951) );
  XNOR U19298 ( .A(n18637), .B(n18638), .Z(n16399) );
  NOR U19299 ( .A(n14104), .B(n14106), .Z(n18635) );
  XOR U19300 ( .A(n18639), .B(n18433), .Z(n14104) );
  XNOR U19301 ( .A(n18640), .B(n14739), .Z(n9814) );
  XOR U19302 ( .A(n18641), .B(n15671), .Z(n14739) );
  ANDN U19303 ( .B(n14100), .A(n14101), .Z(n18640) );
  XNOR U19304 ( .A(n18642), .B(n17009), .Z(n14100) );
  XNOR U19305 ( .A(n18643), .B(n14749), .Z(n14903) );
  XNOR U19306 ( .A(n18644), .B(n17630), .Z(n14749) );
  NOR U19307 ( .A(n14095), .B(n14097), .Z(n18643) );
  IV U19308 ( .A(n15742), .Z(n14095) );
  XNOR U19309 ( .A(n18645), .B(n18563), .Z(n15742) );
  XNOR U19310 ( .A(n18646), .B(n15738), .Z(n14093) );
  XOR U19311 ( .A(n18647), .B(n17982), .Z(n15738) );
  ANDN U19312 ( .B(n14752), .A(n18633), .Z(n18646) );
  XOR U19313 ( .A(n14123), .B(n10108), .Z(n10126) );
  XNOR U19314 ( .A(n18648), .B(n17889), .Z(n14123) );
  IV U19315 ( .A(n18649), .Z(n17889) );
  AND U19316 ( .A(n17823), .B(n18546), .Z(n18648) );
  XOR U19317 ( .A(n18650), .B(n17188), .Z(n17823) );
  XNOR U19318 ( .A(n18651), .B(n7723), .Z(n7705) );
  IV U19319 ( .A(n10081), .Z(n7723) );
  XOR U19320 ( .A(n16481), .B(n9783), .Z(n10081) );
  XNOR U19321 ( .A(n18652), .B(n15514), .Z(n16481) );
  ANDN U19322 ( .B(n18653), .A(n18654), .Z(n18652) );
  ANDN U19323 ( .B(n7666), .A(n6889), .Z(n18651) );
  XOR U19324 ( .A(n13928), .B(n10695), .Z(n6889) );
  XOR U19325 ( .A(n13305), .B(n17811), .Z(n10695) );
  XOR U19326 ( .A(n18655), .B(n18656), .Z(n17811) );
  XNOR U19327 ( .A(n18541), .B(n14260), .Z(n18656) );
  XNOR U19328 ( .A(n18657), .B(n16902), .Z(n14260) );
  IV U19329 ( .A(n18658), .Z(n16902) );
  ANDN U19330 ( .B(n14688), .A(n14687), .Z(n18657) );
  XOR U19331 ( .A(n18659), .B(n17977), .Z(n14688) );
  XNOR U19332 ( .A(n18660), .B(n13859), .Z(n18541) );
  ANDN U19333 ( .B(n16895), .A(n17218), .Z(n18660) );
  XNOR U19334 ( .A(n17145), .B(n18661), .Z(n16895) );
  XOR U19335 ( .A(n9243), .B(n18662), .Z(n18655) );
  XNOR U19336 ( .A(n10011), .B(n13550), .Z(n18662) );
  XNOR U19337 ( .A(n18663), .B(n13854), .Z(n13550) );
  XOR U19338 ( .A(n18664), .B(n17874), .Z(n14685) );
  XNOR U19339 ( .A(n18665), .B(n14196), .Z(n10011) );
  AND U19340 ( .A(n17833), .B(n16897), .Z(n18665) );
  XOR U19341 ( .A(n18666), .B(n17240), .Z(n16897) );
  XNOR U19342 ( .A(n18667), .B(n18668), .Z(n17240) );
  XNOR U19343 ( .A(n18669), .B(n13864), .Z(n9243) );
  ANDN U19344 ( .B(n15103), .A(n18670), .Z(n18669) );
  XOR U19345 ( .A(n16770), .B(n18671), .Z(n15103) );
  XNOR U19346 ( .A(n18672), .B(n18673), .Z(n13305) );
  XOR U19347 ( .A(n14763), .B(n18674), .Z(n18673) );
  XOR U19348 ( .A(n18675), .B(n15811), .Z(n14763) );
  NOR U19349 ( .A(n18676), .B(n13931), .Z(n18675) );
  XOR U19350 ( .A(n18677), .B(n18678), .Z(n13931) );
  XOR U19351 ( .A(n12189), .B(n18679), .Z(n18672) );
  XOR U19352 ( .A(n10268), .B(n13513), .Z(n18679) );
  XNOR U19353 ( .A(n18680), .B(n15815), .Z(n13513) );
  IV U19354 ( .A(n18681), .Z(n15815) );
  AND U19355 ( .A(n13938), .B(n13936), .Z(n18680) );
  XOR U19356 ( .A(n18682), .B(n18468), .Z(n13938) );
  IV U19357 ( .A(n18683), .Z(n18468) );
  XOR U19358 ( .A(n18684), .B(n15804), .Z(n10268) );
  ANDN U19359 ( .B(n13942), .A(n18685), .Z(n18684) );
  XNOR U19360 ( .A(n18686), .B(n16848), .Z(n13942) );
  IV U19361 ( .A(n18687), .Z(n16848) );
  XNOR U19362 ( .A(n18688), .B(n15801), .Z(n12189) );
  ANDN U19363 ( .B(n16806), .A(n18689), .Z(n18688) );
  XNOR U19364 ( .A(n4687), .B(n18691), .Z(n18690) );
  OR U19365 ( .A(n16806), .B(n15799), .Z(n18691) );
  XOR U19366 ( .A(n18692), .B(n18693), .Z(n15799) );
  XNOR U19367 ( .A(n17231), .B(n18694), .Z(n16806) );
  XNOR U19368 ( .A(n12329), .B(n18695), .Z(n7666) );
  XNOR U19369 ( .A(n12252), .B(n11975), .Z(n12329) );
  XOR U19370 ( .A(n18696), .B(n18697), .Z(n11975) );
  XNOR U19371 ( .A(n12129), .B(n13244), .Z(n18697) );
  XNOR U19372 ( .A(n18698), .B(n18097), .Z(n13244) );
  IV U19373 ( .A(n15729), .Z(n18097) );
  XOR U19374 ( .A(n18699), .B(n15541), .Z(n15729) );
  XNOR U19375 ( .A(n18700), .B(n18701), .Z(n15541) );
  NOR U19376 ( .A(n17718), .B(n15728), .Z(n18698) );
  XOR U19377 ( .A(n18702), .B(n18456), .Z(n15728) );
  IV U19378 ( .A(n18359), .Z(n17718) );
  XOR U19379 ( .A(n18703), .B(n17440), .Z(n18359) );
  XNOR U19380 ( .A(n18704), .B(n18089), .Z(n12129) );
  IV U19381 ( .A(n15721), .Z(n18089) );
  XOR U19382 ( .A(n18705), .B(n17744), .Z(n15721) );
  NOR U19383 ( .A(n17715), .B(n15720), .Z(n18704) );
  XOR U19384 ( .A(n18706), .B(n18707), .Z(n15720) );
  XOR U19385 ( .A(n18708), .B(n16507), .Z(n17715) );
  XNOR U19386 ( .A(n11602), .B(n18709), .Z(n18696) );
  XOR U19387 ( .A(n9792), .B(n12358), .Z(n18709) );
  XNOR U19388 ( .A(n18710), .B(n15711), .Z(n12358) );
  IV U19389 ( .A(n18094), .Z(n15711) );
  XNOR U19390 ( .A(n18711), .B(n18712), .Z(n18094) );
  NOR U19391 ( .A(n15712), .B(n18365), .Z(n18710) );
  XNOR U19392 ( .A(n17026), .B(n18713), .Z(n18365) );
  IV U19393 ( .A(n18714), .Z(n17026) );
  XOR U19394 ( .A(n18715), .B(n18064), .Z(n15712) );
  IV U19395 ( .A(n15653), .Z(n18064) );
  XNOR U19396 ( .A(n18716), .B(n15724), .Z(n9792) );
  XOR U19397 ( .A(n18717), .B(n18387), .Z(n15724) );
  ANDN U19398 ( .B(n15725), .A(n17706), .Z(n18716) );
  XNOR U19399 ( .A(n18171), .B(n18718), .Z(n17706) );
  XNOR U19400 ( .A(n18719), .B(n17249), .Z(n15725) );
  XOR U19401 ( .A(n18720), .B(n15716), .Z(n11602) );
  XOR U19402 ( .A(n17399), .B(n18721), .Z(n15716) );
  XOR U19403 ( .A(n18722), .B(n17024), .Z(n15715) );
  XOR U19404 ( .A(n18723), .B(n18521), .Z(n17709) );
  IV U19405 ( .A(n17546), .Z(n18521) );
  XOR U19406 ( .A(n18724), .B(n18725), .Z(n12252) );
  XOR U19407 ( .A(n15705), .B(n13017), .Z(n18725) );
  XOR U19408 ( .A(n18726), .B(n17166), .Z(n13017) );
  XOR U19409 ( .A(n18727), .B(n17918), .Z(n17166) );
  AND U19410 ( .A(n18728), .B(n17167), .Z(n18726) );
  XNOR U19411 ( .A(n18729), .B(n17156), .Z(n15705) );
  XOR U19412 ( .A(n18730), .B(n17574), .Z(n17156) );
  NOR U19413 ( .A(n17157), .B(n18731), .Z(n18729) );
  XOR U19414 ( .A(n10061), .B(n18732), .Z(n18724) );
  XOR U19415 ( .A(n9417), .B(n14440), .Z(n18732) );
  XOR U19416 ( .A(n18733), .B(n17152), .Z(n14440) );
  XOR U19417 ( .A(n18734), .B(n16529), .Z(n17152) );
  NOR U19418 ( .A(n18735), .B(n18736), .Z(n18733) );
  XOR U19419 ( .A(n18737), .B(n18084), .Z(n9417) );
  XOR U19420 ( .A(n18738), .B(n16967), .Z(n18084) );
  IV U19421 ( .A(n17503), .Z(n16967) );
  XOR U19422 ( .A(n18740), .B(n17163), .Z(n10061) );
  XNOR U19423 ( .A(n18706), .B(n18741), .Z(n17163) );
  ANDN U19424 ( .B(n18742), .A(n17162), .Z(n18740) );
  XOR U19425 ( .A(n16927), .B(n10185), .Z(n7734) );
  XNOR U19426 ( .A(n15965), .B(n12417), .Z(n10185) );
  XNOR U19427 ( .A(n18744), .B(n18745), .Z(n12417) );
  XNOR U19428 ( .A(n16702), .B(n11232), .Z(n18745) );
  XNOR U19429 ( .A(n18746), .B(n16434), .Z(n11232) );
  IV U19430 ( .A(n17424), .Z(n16434) );
  XOR U19431 ( .A(n18747), .B(n16516), .Z(n17424) );
  ANDN U19432 ( .B(n16933), .A(n16934), .Z(n18746) );
  XOR U19433 ( .A(n18748), .B(n17479), .Z(n16934) );
  XOR U19434 ( .A(n15654), .B(n18749), .Z(n16933) );
  IV U19435 ( .A(n16825), .Z(n15654) );
  XNOR U19436 ( .A(n18750), .B(n18751), .Z(n16825) );
  XNOR U19437 ( .A(n18752), .B(n16439), .Z(n16702) );
  XNOR U19438 ( .A(n18753), .B(n18458), .Z(n16439) );
  IV U19439 ( .A(n17059), .Z(n18458) );
  ANDN U19440 ( .B(n16929), .A(n16930), .Z(n18752) );
  XNOR U19441 ( .A(n18754), .B(n17333), .Z(n16930) );
  XOR U19442 ( .A(n18714), .B(n18755), .Z(n16929) );
  XOR U19443 ( .A(n18756), .B(n18757), .Z(n18714) );
  XNOR U19444 ( .A(n12901), .B(n18758), .Z(n18744) );
  XOR U19445 ( .A(n10713), .B(n17411), .Z(n18758) );
  XNOR U19446 ( .A(n18759), .B(n16422), .Z(n17411) );
  XOR U19447 ( .A(n18760), .B(n16527), .Z(n16422) );
  ANDN U19448 ( .B(n17946), .A(n18761), .Z(n18759) );
  XNOR U19449 ( .A(n18762), .B(n16426), .Z(n10713) );
  IV U19450 ( .A(n17416), .Z(n16426) );
  XOR U19451 ( .A(n18692), .B(n18763), .Z(n17416) );
  ANDN U19452 ( .B(n16922), .A(n16921), .Z(n18762) );
  XOR U19453 ( .A(n18764), .B(n17970), .Z(n16921) );
  XOR U19454 ( .A(n18765), .B(n18766), .Z(n16922) );
  XOR U19455 ( .A(n18767), .B(n17420), .Z(n12901) );
  XOR U19456 ( .A(n18768), .B(n17977), .Z(n17420) );
  ANDN U19457 ( .B(n16925), .A(n17419), .Z(n18767) );
  XOR U19458 ( .A(n18769), .B(n18770), .Z(n17419) );
  XNOR U19459 ( .A(n18771), .B(n18772), .Z(n16925) );
  XOR U19460 ( .A(n18773), .B(n18774), .Z(n15965) );
  XOR U19461 ( .A(n17071), .B(n12981), .Z(n18774) );
  XNOR U19462 ( .A(n18775), .B(n16759), .Z(n12981) );
  XNOR U19463 ( .A(n18776), .B(n18777), .Z(n16759) );
  ANDN U19464 ( .B(n15990), .A(n15991), .Z(n18775) );
  XNOR U19465 ( .A(n18778), .B(n17093), .Z(n15991) );
  XOR U19466 ( .A(n18779), .B(n16101), .Z(n15990) );
  XNOR U19467 ( .A(n18780), .B(n16764), .Z(n17071) );
  XOR U19468 ( .A(n18781), .B(n15347), .Z(n16764) );
  IV U19469 ( .A(n17788), .Z(n15347) );
  AND U19470 ( .A(n14387), .B(n14385), .Z(n18780) );
  XOR U19471 ( .A(n18171), .B(n18782), .Z(n14385) );
  XOR U19472 ( .A(n18783), .B(n18438), .Z(n14387) );
  XOR U19473 ( .A(n12494), .B(n18784), .Z(n18773) );
  XOR U19474 ( .A(n12576), .B(n11167), .Z(n18784) );
  XNOR U19475 ( .A(n18785), .B(n16772), .Z(n11167) );
  XOR U19476 ( .A(n18786), .B(n18787), .Z(n16772) );
  ANDN U19477 ( .B(n12858), .A(n12860), .Z(n18785) );
  XOR U19478 ( .A(n18788), .B(n18789), .Z(n12860) );
  XOR U19479 ( .A(n18790), .B(n18791), .Z(n12858) );
  XNOR U19480 ( .A(n18792), .B(n16768), .Z(n12576) );
  XOR U19481 ( .A(n18793), .B(n18078), .Z(n16768) );
  ANDN U19482 ( .B(n12866), .A(n17437), .Z(n18792) );
  IV U19483 ( .A(n12864), .Z(n17437) );
  XOR U19484 ( .A(n18794), .B(n18212), .Z(n12864) );
  XOR U19485 ( .A(n18795), .B(n16511), .Z(n12866) );
  XNOR U19486 ( .A(n18796), .B(n16755), .Z(n12494) );
  XOR U19487 ( .A(n18797), .B(n18798), .Z(n16755) );
  ANDN U19488 ( .B(n12868), .A(n12869), .Z(n18796) );
  XOR U19489 ( .A(n18692), .B(n18799), .Z(n12869) );
  XNOR U19490 ( .A(n18800), .B(n17586), .Z(n12868) );
  XNOR U19491 ( .A(n18801), .B(n18761), .Z(n16927) );
  IV U19492 ( .A(n17422), .Z(n18761) );
  XOR U19493 ( .A(n18802), .B(n16023), .Z(n17422) );
  NOR U19494 ( .A(n17946), .B(n16420), .Z(n18801) );
  XOR U19495 ( .A(n18803), .B(n18804), .Z(n16420) );
  XNOR U19496 ( .A(n18805), .B(n18806), .Z(n17946) );
  NOR U19497 ( .A(n7659), .B(n6885), .Z(n18743) );
  XOR U19498 ( .A(n15753), .B(n11754), .Z(n6885) );
  XNOR U19499 ( .A(n18807), .B(n12632), .Z(n11754) );
  XNOR U19500 ( .A(n18808), .B(n18809), .Z(n12632) );
  XNOR U19501 ( .A(n12984), .B(n11190), .Z(n18809) );
  XOR U19502 ( .A(n18810), .B(n15212), .Z(n11190) );
  XNOR U19503 ( .A(n18811), .B(n17592), .Z(n15212) );
  NOR U19504 ( .A(n14058), .B(n15211), .Z(n18810) );
  XOR U19505 ( .A(n18812), .B(n18813), .Z(n15211) );
  XOR U19506 ( .A(n18814), .B(n18815), .Z(n14058) );
  XOR U19507 ( .A(n18816), .B(n15216), .Z(n12984) );
  XOR U19508 ( .A(n18817), .B(n17740), .Z(n15216) );
  IV U19509 ( .A(n15671), .Z(n17740) );
  ANDN U19510 ( .B(n15748), .A(n15215), .Z(n18816) );
  XNOR U19511 ( .A(n18820), .B(n15351), .Z(n15215) );
  XOR U19512 ( .A(n18821), .B(n18822), .Z(n15748) );
  XOR U19513 ( .A(n15207), .B(n18823), .Z(n18808) );
  XNOR U19514 ( .A(n11935), .B(n11042), .Z(n18823) );
  XOR U19515 ( .A(n18824), .B(n15227), .Z(n11042) );
  XOR U19516 ( .A(n18825), .B(n18502), .Z(n15227) );
  ANDN U19517 ( .B(n14048), .A(n15226), .Z(n18824) );
  XNOR U19518 ( .A(n18826), .B(n15223), .Z(n11935) );
  XOR U19519 ( .A(n18827), .B(n18828), .Z(n15223) );
  XNOR U19520 ( .A(n18829), .B(n18830), .Z(n14052) );
  XNOR U19521 ( .A(n18692), .B(n18831), .Z(n15224) );
  XNOR U19522 ( .A(n18832), .B(n15220), .Z(n15207) );
  XOR U19523 ( .A(n18833), .B(n18834), .Z(n15220) );
  ANDN U19524 ( .B(n14062), .A(n15219), .Z(n18832) );
  XOR U19525 ( .A(n18835), .B(n18836), .Z(n15219) );
  XOR U19526 ( .A(n18837), .B(n18078), .Z(n14062) );
  IV U19527 ( .A(n18480), .Z(n18078) );
  XNOR U19528 ( .A(n18838), .B(n18839), .Z(n18606) );
  XOR U19529 ( .A(n18840), .B(n18841), .Z(n18839) );
  XOR U19530 ( .A(n14963), .B(n18842), .Z(n18838) );
  XOR U19531 ( .A(n18843), .B(n18267), .Z(n18842) );
  XNOR U19532 ( .A(n18844), .B(n18845), .Z(n18267) );
  ANDN U19533 ( .B(n18846), .A(n18847), .Z(n18844) );
  XNOR U19534 ( .A(n18848), .B(n18849), .Z(n14963) );
  XOR U19535 ( .A(n18853), .B(n15226), .Z(n15753) );
  XOR U19536 ( .A(n18854), .B(n18855), .Z(n15226) );
  NOR U19537 ( .A(n14048), .B(n14049), .Z(n18853) );
  XNOR U19538 ( .A(n18856), .B(n18857), .Z(n14049) );
  XNOR U19539 ( .A(n18858), .B(n18712), .Z(n14048) );
  XOR U19540 ( .A(n9966), .B(n13453), .Z(n7659) );
  XNOR U19541 ( .A(n18859), .B(n14889), .Z(n13453) );
  ANDN U19542 ( .B(n16564), .A(n16565), .Z(n18859) );
  XNOR U19543 ( .A(n18860), .B(n17699), .Z(n16565) );
  XNOR U19544 ( .A(n13373), .B(n13333), .Z(n9966) );
  XOR U19545 ( .A(n18861), .B(n18862), .Z(n13333) );
  XNOR U19546 ( .A(n9651), .B(n12622), .Z(n18862) );
  XNOR U19547 ( .A(n18863), .B(n14881), .Z(n12622) );
  XOR U19548 ( .A(n18864), .B(n18865), .Z(n14881) );
  ANDN U19549 ( .B(n13460), .A(n13461), .Z(n18863) );
  XOR U19550 ( .A(n18866), .B(n18177), .Z(n13461) );
  XOR U19551 ( .A(n18867), .B(n17500), .Z(n13460) );
  XNOR U19552 ( .A(n18868), .B(n14884), .Z(n9651) );
  XNOR U19553 ( .A(n18869), .B(n17140), .Z(n14884) );
  ANDN U19554 ( .B(n13446), .A(n16562), .Z(n18868) );
  IV U19555 ( .A(n13448), .Z(n16562) );
  XOR U19556 ( .A(n18870), .B(n16032), .Z(n13448) );
  XOR U19557 ( .A(n17635), .B(n18871), .Z(n13446) );
  XOR U19558 ( .A(n12390), .B(n18872), .Z(n18861) );
  XNOR U19559 ( .A(n9669), .B(n14089), .Z(n18872) );
  XOR U19560 ( .A(n18873), .B(n14892), .Z(n14089) );
  XOR U19561 ( .A(n18874), .B(n15904), .Z(n14892) );
  XOR U19562 ( .A(n17472), .B(n18875), .Z(n13450) );
  XOR U19563 ( .A(n18876), .B(n18877), .Z(n13452) );
  XOR U19564 ( .A(n18878), .B(n14888), .Z(n9669) );
  XNOR U19565 ( .A(n18879), .B(n16841), .Z(n14888) );
  ANDN U19566 ( .B(n14889), .A(n16564), .Z(n18878) );
  XOR U19567 ( .A(n18880), .B(n18248), .Z(n16564) );
  XNOR U19568 ( .A(n18881), .B(n15351), .Z(n14889) );
  XOR U19569 ( .A(n18882), .B(n14895), .Z(n12390) );
  XOR U19570 ( .A(n18100), .B(n18883), .Z(n14895) );
  XOR U19571 ( .A(n18884), .B(n15201), .Z(n13457) );
  XOR U19572 ( .A(n18885), .B(n16331), .Z(n13456) );
  XOR U19573 ( .A(n18886), .B(n18887), .Z(n13373) );
  XNOR U19574 ( .A(n12052), .B(n12958), .Z(n18887) );
  XOR U19575 ( .A(n18888), .B(n14106), .Z(n12958) );
  XOR U19576 ( .A(n18889), .B(n18890), .Z(n14106) );
  NOR U19577 ( .A(n14105), .B(n14746), .Z(n18888) );
  XOR U19578 ( .A(n18891), .B(n18260), .Z(n14746) );
  XOR U19579 ( .A(n18892), .B(n17451), .Z(n14105) );
  XNOR U19580 ( .A(n18893), .B(n14097), .Z(n12052) );
  XNOR U19581 ( .A(n17143), .B(n18894), .Z(n14097) );
  ANDN U19582 ( .B(n14750), .A(n14096), .Z(n18893) );
  XOR U19583 ( .A(n18895), .B(n15290), .Z(n14096) );
  IV U19584 ( .A(n18896), .Z(n15290) );
  XNOR U19585 ( .A(n18897), .B(n17699), .Z(n14750) );
  XNOR U19586 ( .A(n11742), .B(n18898), .Z(n18886) );
  XNOR U19587 ( .A(n11763), .B(n11594), .Z(n18898) );
  XOR U19588 ( .A(n18899), .B(n18633), .Z(n11594) );
  XOR U19589 ( .A(n18900), .B(n18473), .Z(n18633) );
  XNOR U19590 ( .A(n16374), .B(n18901), .Z(n14752) );
  XOR U19591 ( .A(n18902), .B(n17654), .Z(n14754) );
  XNOR U19592 ( .A(n18903), .B(n14101), .Z(n11763) );
  XOR U19593 ( .A(n18216), .B(n18904), .Z(n14101) );
  AND U19594 ( .A(n14740), .B(n14102), .Z(n18903) );
  XOR U19595 ( .A(n18905), .B(n18613), .Z(n14102) );
  XNOR U19596 ( .A(n18906), .B(n18804), .Z(n14740) );
  XNOR U19597 ( .A(n18907), .B(n14109), .Z(n11742) );
  XOR U19598 ( .A(n18908), .B(n17244), .Z(n14109) );
  ANDN U19599 ( .B(n14110), .A(n14742), .Z(n18907) );
  XOR U19600 ( .A(n14962), .B(n18840), .Z(n14742) );
  XOR U19601 ( .A(n18909), .B(n18910), .Z(n18840) );
  XOR U19602 ( .A(n18913), .B(n14168), .Z(n14110) );
  XOR U19603 ( .A(n18914), .B(n6863), .Z(n7669) );
  XNOR U19604 ( .A(n11698), .B(n14267), .Z(n6863) );
  XOR U19605 ( .A(n18915), .B(n14232), .Z(n14267) );
  ANDN U19606 ( .B(n17221), .A(n17242), .Z(n18915) );
  XOR U19607 ( .A(n18916), .B(n16668), .Z(n17221) );
  XOR U19608 ( .A(n18917), .B(n18918), .Z(n16668) );
  XOR U19609 ( .A(n17361), .B(n18568), .Z(n11698) );
  XNOR U19610 ( .A(n18919), .B(n18920), .Z(n18568) );
  XNOR U19611 ( .A(n9860), .B(n12759), .Z(n18920) );
  XNOR U19612 ( .A(n18921), .B(n13572), .Z(n12759) );
  XNOR U19613 ( .A(n18922), .B(n15891), .Z(n13572) );
  ANDN U19614 ( .B(n16861), .A(n14228), .Z(n18921) );
  XOR U19615 ( .A(n18923), .B(n18865), .Z(n14228) );
  XNOR U19616 ( .A(n18924), .B(n16892), .Z(n16861) );
  XNOR U19617 ( .A(n18927), .B(n13566), .Z(n9860) );
  XNOR U19618 ( .A(n18928), .B(n16613), .Z(n13566) );
  XOR U19619 ( .A(n15639), .B(n18929), .Z(n14225) );
  XOR U19620 ( .A(n18930), .B(n16086), .Z(n14275) );
  XOR U19621 ( .A(n12968), .B(n18931), .Z(n18919) );
  XNOR U19622 ( .A(n11889), .B(n9930), .Z(n18931) );
  XOR U19623 ( .A(n18932), .B(n14219), .Z(n9930) );
  XOR U19624 ( .A(n18933), .B(n17498), .Z(n14219) );
  AND U19625 ( .A(n14273), .B(n14220), .Z(n18932) );
  XNOR U19626 ( .A(n18934), .B(n17059), .Z(n14220) );
  XOR U19627 ( .A(n18935), .B(n18936), .Z(n17059) );
  XOR U19628 ( .A(n18937), .B(n17988), .Z(n14273) );
  IV U19629 ( .A(n18938), .Z(n17988) );
  XOR U19630 ( .A(n18939), .B(n14231), .Z(n11889) );
  XOR U19631 ( .A(n15645), .B(n18940), .Z(n14231) );
  XOR U19632 ( .A(n18941), .B(n18942), .Z(n17242) );
  XOR U19633 ( .A(n18943), .B(n18944), .Z(n14232) );
  XNOR U19634 ( .A(n18945), .B(n13562), .Z(n12968) );
  XOR U19635 ( .A(n18946), .B(n18167), .Z(n13562) );
  AND U19636 ( .A(n14671), .B(n14222), .Z(n18945) );
  XOR U19637 ( .A(n18947), .B(n17024), .Z(n14222) );
  XOR U19638 ( .A(n18948), .B(n18949), .Z(n14671) );
  XOR U19639 ( .A(n18950), .B(n18951), .Z(n17361) );
  XNOR U19640 ( .A(n14111), .B(n15104), .Z(n18951) );
  XNOR U19641 ( .A(n18952), .B(n15120), .Z(n15104) );
  IV U19642 ( .A(n16648), .Z(n15120) );
  XOR U19643 ( .A(n18953), .B(n17735), .Z(n16648) );
  IV U19644 ( .A(n16507), .Z(n17735) );
  XOR U19645 ( .A(n18954), .B(n18955), .Z(n16507) );
  ANDN U19646 ( .B(n14290), .A(n15119), .Z(n18952) );
  IV U19647 ( .A(n14289), .Z(n15119) );
  XNOR U19648 ( .A(n18956), .B(n17918), .Z(n14289) );
  XOR U19649 ( .A(n17143), .B(n18957), .Z(n14290) );
  XOR U19650 ( .A(n18958), .B(n15110), .Z(n14111) );
  XOR U19651 ( .A(n18959), .B(n18561), .Z(n15110) );
  ANDN U19652 ( .B(n14283), .A(n14284), .Z(n18958) );
  IV U19653 ( .A(n17991), .Z(n14284) );
  XOR U19654 ( .A(n18960), .B(n17982), .Z(n17991) );
  XOR U19655 ( .A(n17921), .B(n18961), .Z(n14283) );
  XOR U19656 ( .A(n14132), .B(n18962), .Z(n18950) );
  XOR U19657 ( .A(n12842), .B(n12121), .Z(n18962) );
  XOR U19658 ( .A(n18963), .B(n16624), .Z(n12121) );
  XOR U19659 ( .A(n18964), .B(n18965), .Z(n16624) );
  ANDN U19660 ( .B(n14279), .A(n14280), .Z(n18963) );
  XOR U19661 ( .A(n18966), .B(n17188), .Z(n14280) );
  IV U19662 ( .A(n18967), .Z(n17188) );
  XOR U19663 ( .A(n18539), .B(n18968), .Z(n14279) );
  XOR U19664 ( .A(n18969), .B(n15114), .Z(n12842) );
  XNOR U19665 ( .A(n18970), .B(n16608), .Z(n15114) );
  ANDN U19666 ( .B(n17364), .A(n15113), .Z(n18969) );
  XOR U19667 ( .A(n18971), .B(n17750), .Z(n15113) );
  XNOR U19668 ( .A(n17231), .B(n18972), .Z(n17364) );
  XNOR U19669 ( .A(n18973), .B(n15123), .Z(n14132) );
  XOR U19670 ( .A(n18974), .B(n17015), .Z(n15123) );
  ANDN U19671 ( .B(n14293), .A(n14294), .Z(n18973) );
  XNOR U19672 ( .A(n18975), .B(n17788), .Z(n14294) );
  XNOR U19673 ( .A(n18976), .B(n18977), .Z(n17788) );
  XNOR U19674 ( .A(n17233), .B(n18978), .Z(n14293) );
  NOR U19675 ( .A(n7569), .B(n9968), .Z(n18914) );
  XNOR U19676 ( .A(n9637), .B(n18979), .Z(n9968) );
  XNOR U19677 ( .A(n14357), .B(n10749), .Z(n7569) );
  XNOR U19678 ( .A(n18980), .B(n18981), .Z(n14357) );
  AND U19679 ( .A(n17538), .B(n12486), .Z(n18980) );
  XNOR U19680 ( .A(n18982), .B(n17564), .Z(n12486) );
  XOR U19681 ( .A(n18983), .B(n18984), .Z(n17564) );
  XOR U19682 ( .A(n1807), .B(n9265), .Z(n4105) );
  XNOR U19683 ( .A(n18985), .B(n9323), .Z(n9265) );
  ANDN U19684 ( .B(n6671), .A(n7132), .Z(n18985) );
  XOR U19685 ( .A(n9637), .B(n18986), .Z(n6671) );
  IV U19686 ( .A(n11808), .Z(n9637) );
  XNOR U19687 ( .A(n12670), .B(n14654), .Z(n11808) );
  XOR U19688 ( .A(n18987), .B(n18988), .Z(n14654) );
  XNOR U19689 ( .A(n16460), .B(n11944), .Z(n18988) );
  XOR U19690 ( .A(n18989), .B(n18653), .Z(n11944) );
  XNOR U19691 ( .A(n18990), .B(n16479), .Z(n16460) );
  NOR U19692 ( .A(n18991), .B(n16478), .Z(n18990) );
  XNOR U19693 ( .A(n10178), .B(n18992), .Z(n18987) );
  XOR U19694 ( .A(n9437), .B(n10877), .Z(n18992) );
  XOR U19695 ( .A(n18993), .B(n16484), .Z(n10877) );
  ANDN U19696 ( .B(n15517), .A(n16485), .Z(n18993) );
  XNOR U19697 ( .A(n18994), .B(n18995), .Z(n9437) );
  ANDN U19698 ( .B(n18996), .A(n15508), .Z(n18994) );
  XNOR U19699 ( .A(n18997), .B(n16488), .Z(n10178) );
  NOR U19700 ( .A(n15504), .B(n16487), .Z(n18997) );
  XOR U19701 ( .A(n18998), .B(n18999), .Z(n12670) );
  XOR U19702 ( .A(n12733), .B(n15388), .Z(n18999) );
  XNOR U19703 ( .A(n19000), .B(n15405), .Z(n15388) );
  XOR U19704 ( .A(n19001), .B(n17942), .Z(n15405) );
  IV U19705 ( .A(n16090), .Z(n17942) );
  ANDN U19706 ( .B(n15406), .A(n19002), .Z(n19000) );
  XNOR U19707 ( .A(n19003), .B(n15409), .Z(n12733) );
  XOR U19708 ( .A(n19004), .B(n16008), .Z(n15409) );
  ANDN U19709 ( .B(n15408), .A(n14586), .Z(n19003) );
  XOR U19710 ( .A(n12105), .B(n19005), .Z(n18998) );
  XOR U19711 ( .A(n10762), .B(n14481), .Z(n19005) );
  XOR U19712 ( .A(n19006), .B(n15397), .Z(n14481) );
  XNOR U19713 ( .A(n19007), .B(n18557), .Z(n15397) );
  XOR U19714 ( .A(n19009), .B(n15401), .Z(n10762) );
  XNOR U19715 ( .A(n19010), .B(n19011), .Z(n15401) );
  ANDN U19716 ( .B(n15402), .A(n13827), .Z(n19009) );
  XOR U19717 ( .A(n19012), .B(n15394), .Z(n12105) );
  XOR U19718 ( .A(n19013), .B(n16101), .Z(n15394) );
  XNOR U19719 ( .A(n19014), .B(n19015), .Z(n16101) );
  NOR U19720 ( .A(n19016), .B(n15393), .Z(n19012) );
  IV U19721 ( .A(n5201), .Z(n1807) );
  XNOR U19722 ( .A(n6641), .B(n6377), .Z(n5201) );
  XOR U19723 ( .A(n19017), .B(n19018), .Z(n6377) );
  XOR U19724 ( .A(n5951), .B(n4350), .Z(n19018) );
  XNOR U19725 ( .A(n19019), .B(n7227), .Z(n4350) );
  XOR U19726 ( .A(n16169), .B(n12325), .Z(n7227) );
  XOR U19727 ( .A(n16250), .B(n12125), .Z(n12325) );
  XOR U19728 ( .A(n19020), .B(n19021), .Z(n12125) );
  XOR U19729 ( .A(n11333), .B(n11182), .Z(n19021) );
  XOR U19730 ( .A(n19022), .B(n12542), .Z(n11182) );
  XNOR U19731 ( .A(n19023), .B(n16398), .Z(n12542) );
  IV U19732 ( .A(n15899), .Z(n16398) );
  NOR U19733 ( .A(n14344), .B(n14345), .Z(n19022) );
  XOR U19734 ( .A(n19024), .B(n19025), .Z(n14345) );
  IV U19735 ( .A(n12541), .Z(n14344) );
  XNOR U19736 ( .A(n19026), .B(n17744), .Z(n12541) );
  XNOR U19737 ( .A(n19027), .B(n12538), .Z(n11333) );
  XOR U19738 ( .A(n19028), .B(n18787), .Z(n12538) );
  NOR U19739 ( .A(n14338), .B(n14339), .Z(n19027) );
  XNOR U19740 ( .A(n19029), .B(n15891), .Z(n14339) );
  IV U19741 ( .A(n12537), .Z(n14338) );
  XOR U19742 ( .A(n17192), .B(n19030), .Z(n12537) );
  IV U19743 ( .A(n17272), .Z(n17192) );
  XNOR U19744 ( .A(n10328), .B(n19031), .Z(n19020) );
  XNOR U19745 ( .A(n11370), .B(n11156), .Z(n19031) );
  XNOR U19746 ( .A(n19032), .B(n12547), .Z(n11156) );
  XNOR U19747 ( .A(n19033), .B(n17479), .Z(n12547) );
  AND U19748 ( .A(n12546), .B(n14342), .Z(n19032) );
  XNOR U19749 ( .A(n19034), .B(n19035), .Z(n14342) );
  XOR U19750 ( .A(n19036), .B(n19037), .Z(n12546) );
  XNOR U19751 ( .A(n19038), .B(n12550), .Z(n11370) );
  XOR U19752 ( .A(n19039), .B(n18944), .Z(n12550) );
  IV U19753 ( .A(n18212), .Z(n18944) );
  ANDN U19754 ( .B(n14331), .A(n12551), .Z(n19038) );
  XOR U19755 ( .A(n19040), .B(n17001), .Z(n12551) );
  IV U19756 ( .A(n16608), .Z(n17001) );
  XOR U19757 ( .A(n19041), .B(n19042), .Z(n16608) );
  XOR U19758 ( .A(n16733), .B(n19043), .Z(n14331) );
  XOR U19759 ( .A(n19044), .B(n13603), .Z(n10328) );
  XOR U19760 ( .A(n19045), .B(n18221), .Z(n13603) );
  ANDN U19761 ( .B(n14335), .A(n14334), .Z(n19044) );
  IV U19762 ( .A(n12555), .Z(n14334) );
  XOR U19763 ( .A(n19046), .B(n17429), .Z(n12555) );
  IV U19764 ( .A(n18374), .Z(n17429) );
  XOR U19765 ( .A(n19047), .B(n19048), .Z(n18374) );
  XOR U19766 ( .A(n19049), .B(n18678), .Z(n14335) );
  IV U19767 ( .A(n18766), .Z(n18678) );
  XOR U19768 ( .A(n19050), .B(n19051), .Z(n16250) );
  XOR U19769 ( .A(n11694), .B(n10506), .Z(n19051) );
  XNOR U19770 ( .A(n19052), .B(n12565), .Z(n10506) );
  XOR U19771 ( .A(n19053), .B(n18212), .Z(n12565) );
  XOR U19772 ( .A(n19054), .B(n19055), .Z(n18212) );
  NOR U19773 ( .A(n12564), .B(n16171), .Z(n19052) );
  XOR U19774 ( .A(n19056), .B(n18309), .Z(n12564) );
  XNOR U19775 ( .A(n19057), .B(n13619), .Z(n11694) );
  IV U19776 ( .A(n13391), .Z(n13619) );
  XOR U19777 ( .A(n19058), .B(n16502), .Z(n13391) );
  ANDN U19778 ( .B(n13392), .A(n19059), .Z(n19057) );
  XOR U19779 ( .A(n19060), .B(n19061), .Z(n13392) );
  XOR U19780 ( .A(n9249), .B(n19062), .Z(n19050) );
  XOR U19781 ( .A(n12532), .B(n9803), .Z(n19062) );
  XNOR U19782 ( .A(n19063), .B(n13616), .Z(n9803) );
  IV U19783 ( .A(n12874), .Z(n13616) );
  XOR U19784 ( .A(n19064), .B(n15679), .Z(n12874) );
  NOR U19785 ( .A(n19065), .B(n12873), .Z(n19063) );
  XNOR U19786 ( .A(n19066), .B(n12569), .Z(n12532) );
  XNOR U19787 ( .A(n19067), .B(n17795), .Z(n12569) );
  ANDN U19788 ( .B(n16167), .A(n12568), .Z(n19066) );
  XOR U19789 ( .A(n19068), .B(n18227), .Z(n12568) );
  IV U19790 ( .A(n19069), .Z(n18227) );
  XNOR U19791 ( .A(n19070), .B(n13628), .Z(n9249) );
  XNOR U19792 ( .A(n19071), .B(n16404), .Z(n13628) );
  IV U19793 ( .A(n19072), .Z(n16404) );
  ANDN U19794 ( .B(n16164), .A(n13630), .Z(n19070) );
  XOR U19795 ( .A(n19073), .B(n15261), .Z(n13630) );
  XOR U19796 ( .A(n19074), .B(n12873), .Z(n16169) );
  XOR U19797 ( .A(n19075), .B(n17907), .Z(n12873) );
  ANDN U19798 ( .B(n19065), .A(n13615), .Z(n19074) );
  ANDN U19799 ( .B(n6714), .A(n6716), .Z(n19019) );
  XOR U19800 ( .A(n14916), .B(n10113), .Z(n6716) );
  XOR U19801 ( .A(n14735), .B(n19076), .Z(n10113) );
  XOR U19802 ( .A(n19077), .B(n19078), .Z(n14735) );
  XOR U19803 ( .A(n9890), .B(n13072), .Z(n19078) );
  XOR U19804 ( .A(n19079), .B(n15821), .Z(n13072) );
  XOR U19805 ( .A(n17321), .B(n19080), .Z(n15821) );
  XOR U19806 ( .A(n19082), .B(n18577), .Z(n15824) );
  IV U19807 ( .A(n17244), .Z(n18577) );
  ANDN U19808 ( .B(n14908), .A(n18616), .Z(n19081) );
  XNOR U19809 ( .A(n19083), .B(n18830), .Z(n18616) );
  XOR U19810 ( .A(n19084), .B(n17916), .Z(n14908) );
  XNOR U19811 ( .A(n19085), .B(n19086), .Z(n17916) );
  XOR U19812 ( .A(n15795), .B(n19087), .Z(n19077) );
  XOR U19813 ( .A(n9913), .B(n12789), .Z(n19087) );
  XNOR U19814 ( .A(n19088), .B(n15829), .Z(n12789) );
  XOR U19815 ( .A(n18016), .B(n19089), .Z(n15829) );
  ANDN U19816 ( .B(n15830), .A(n18603), .Z(n19088) );
  IV U19817 ( .A(n14920), .Z(n18603) );
  XOR U19818 ( .A(n19090), .B(n18400), .Z(n14920) );
  IV U19819 ( .A(n14918), .Z(n15830) );
  XOR U19820 ( .A(n19091), .B(n18836), .Z(n14918) );
  XOR U19821 ( .A(n19092), .B(n16800), .Z(n9913) );
  XNOR U19822 ( .A(n19093), .B(n17451), .Z(n16800) );
  XOR U19823 ( .A(n19094), .B(n19095), .Z(n17451) );
  ANDN U19824 ( .B(n14922), .A(n14923), .Z(n19092) );
  XNOR U19825 ( .A(n19096), .B(n17297), .Z(n14923) );
  XNOR U19826 ( .A(n19097), .B(n18309), .Z(n14922) );
  XNOR U19827 ( .A(n19098), .B(n15833), .Z(n15795) );
  XNOR U19828 ( .A(n16822), .B(n19099), .Z(n15833) );
  ANDN U19829 ( .B(n14912), .A(n18609), .Z(n19098) );
  XOR U19830 ( .A(n19100), .B(n16108), .Z(n18609) );
  XOR U19831 ( .A(n19101), .B(n19102), .Z(n14912) );
  XNOR U19832 ( .A(n19103), .B(n15820), .Z(n14916) );
  XOR U19833 ( .A(n19104), .B(n17622), .Z(n15820) );
  ANDN U19834 ( .B(n16792), .A(n18624), .Z(n19103) );
  XOR U19835 ( .A(n17231), .B(n19105), .Z(n18624) );
  XNOR U19836 ( .A(n19106), .B(n18804), .Z(n16792) );
  XNOR U19837 ( .A(n19107), .B(n11925), .Z(n6714) );
  XOR U19838 ( .A(n19108), .B(n7236), .Z(n5951) );
  XOR U19839 ( .A(n9263), .B(n18126), .Z(n7236) );
  XNOR U19840 ( .A(n19109), .B(n16711), .Z(n18126) );
  ANDN U19841 ( .B(n15914), .A(n19110), .Z(n19109) );
  IV U19842 ( .A(n12499), .Z(n9263) );
  XNOR U19843 ( .A(n12964), .B(n16205), .Z(n12499) );
  XOR U19844 ( .A(n19111), .B(n19112), .Z(n16205) );
  XNOR U19845 ( .A(n13786), .B(n14901), .Z(n19112) );
  XNOR U19846 ( .A(n19113), .B(n15916), .Z(n14901) );
  IV U19847 ( .A(n16712), .Z(n15916) );
  XOR U19848 ( .A(n19114), .B(n16008), .Z(n16712) );
  XNOR U19849 ( .A(n19115), .B(n19116), .Z(n16008) );
  XNOR U19850 ( .A(n18090), .B(n19117), .Z(n16711) );
  XOR U19851 ( .A(n19118), .B(n15924), .Z(n13786) );
  XOR U19852 ( .A(n19119), .B(n18804), .Z(n15924) );
  NOR U19853 ( .A(n18125), .B(n16715), .Z(n19118) );
  XOR U19854 ( .A(n19120), .B(n16992), .Z(n16715) );
  XNOR U19855 ( .A(n11351), .B(n19121), .Z(n19111) );
  XOR U19856 ( .A(n11238), .B(n15007), .Z(n19121) );
  XNOR U19857 ( .A(n19122), .B(n15920), .Z(n15007) );
  XNOR U19858 ( .A(n16957), .B(n19123), .Z(n15920) );
  ANDN U19859 ( .B(n18123), .A(n16717), .Z(n19122) );
  XOR U19860 ( .A(n16036), .B(n19124), .Z(n16717) );
  XNOR U19861 ( .A(n19125), .B(n15929), .Z(n11238) );
  IV U19862 ( .A(n16720), .Z(n15929) );
  XOR U19863 ( .A(n17522), .B(n19126), .Z(n16720) );
  NOR U19864 ( .A(n18129), .B(n16719), .Z(n19125) );
  XOR U19865 ( .A(n19127), .B(n18517), .Z(n16719) );
  XOR U19866 ( .A(n19128), .B(n16709), .Z(n11351) );
  IV U19867 ( .A(n15933), .Z(n16709) );
  XOR U19868 ( .A(n19129), .B(n17098), .Z(n15933) );
  NOR U19869 ( .A(n18131), .B(n16708), .Z(n19128) );
  XOR U19870 ( .A(n19130), .B(n18397), .Z(n16708) );
  XOR U19871 ( .A(n19131), .B(n19132), .Z(n12964) );
  XOR U19872 ( .A(n9953), .B(n11578), .Z(n19132) );
  XOR U19873 ( .A(n19133), .B(n15017), .Z(n11578) );
  ANDN U19874 ( .B(n15018), .A(n18135), .Z(n19133) );
  XOR U19875 ( .A(n19134), .B(n17994), .Z(n18135) );
  XNOR U19876 ( .A(n19137), .B(n16301), .Z(n15018) );
  XNOR U19877 ( .A(n19138), .B(n19139), .Z(n16301) );
  XNOR U19878 ( .A(n19140), .B(n15027), .Z(n9953) );
  ANDN U19879 ( .B(n16187), .A(n15028), .Z(n19140) );
  XNOR U19880 ( .A(n19141), .B(n19025), .Z(n15028) );
  XNOR U19881 ( .A(n19142), .B(n17578), .Z(n16187) );
  XOR U19882 ( .A(n10090), .B(n19143), .Z(n19131) );
  XNOR U19883 ( .A(n10937), .B(n10732), .Z(n19143) );
  XOR U19884 ( .A(n19144), .B(n19145), .Z(n10732) );
  ANDN U19885 ( .B(n16194), .A(n18140), .Z(n19144) );
  XNOR U19886 ( .A(n19146), .B(n16529), .Z(n16194) );
  XNOR U19887 ( .A(n19147), .B(n19148), .Z(n19095) );
  XOR U19888 ( .A(n14159), .B(n17611), .Z(n19148) );
  XOR U19889 ( .A(n19149), .B(n19150), .Z(n17611) );
  ANDN U19890 ( .B(n19151), .A(n19152), .Z(n19149) );
  XOR U19891 ( .A(n19153), .B(n19154), .Z(n14159) );
  ANDN U19892 ( .B(n19155), .A(n19156), .Z(n19153) );
  XNOR U19893 ( .A(n18436), .B(n19157), .Z(n19147) );
  XNOR U19894 ( .A(n19158), .B(n18572), .Z(n19157) );
  XNOR U19895 ( .A(n19159), .B(n19160), .Z(n18572) );
  ANDN U19896 ( .B(n19161), .A(n19162), .Z(n19159) );
  XNOR U19897 ( .A(n19163), .B(n19164), .Z(n18436) );
  NOR U19898 ( .A(n19165), .B(n19166), .Z(n19163) );
  XNOR U19899 ( .A(n19168), .B(n15013), .Z(n10937) );
  ANDN U19900 ( .B(n15014), .A(n16191), .Z(n19168) );
  XOR U19901 ( .A(n19169), .B(n19170), .Z(n16191) );
  XOR U19902 ( .A(n19171), .B(n15663), .Z(n15014) );
  XNOR U19903 ( .A(n19172), .B(n15023), .Z(n10090) );
  NOR U19904 ( .A(n18137), .B(n16183), .Z(n19172) );
  XNOR U19905 ( .A(n19173), .B(n18442), .Z(n16183) );
  IV U19906 ( .A(n15024), .Z(n18137) );
  XOR U19907 ( .A(n19174), .B(n17432), .Z(n15024) );
  ANDN U19908 ( .B(n6697), .A(n6698), .Z(n19108) );
  XOR U19909 ( .A(n14358), .B(n10749), .Z(n6698) );
  XOR U19910 ( .A(n12124), .B(n17702), .Z(n10749) );
  XNOR U19911 ( .A(n19175), .B(n19176), .Z(n17702) );
  XNOR U19912 ( .A(n11966), .B(n12908), .Z(n19176) );
  XOR U19913 ( .A(n19177), .B(n18742), .Z(n12908) );
  NOR U19914 ( .A(n17161), .B(n18108), .Z(n19177) );
  XOR U19915 ( .A(n19178), .B(n18611), .Z(n17161) );
  IV U19916 ( .A(n16023), .Z(n18611) );
  XOR U19917 ( .A(n19179), .B(n19180), .Z(n16023) );
  XOR U19918 ( .A(n19181), .B(n18728), .Z(n11966) );
  ANDN U19919 ( .B(n17165), .A(n19182), .Z(n19181) );
  XNOR U19920 ( .A(n19183), .B(n16086), .Z(n17165) );
  XOR U19921 ( .A(n11506), .B(n19184), .Z(n19175) );
  XOR U19922 ( .A(n9649), .B(n12192), .Z(n19184) );
  XNOR U19923 ( .A(n19185), .B(n18739), .Z(n12192) );
  ANDN U19924 ( .B(n18083), .A(n19186), .Z(n19185) );
  XNOR U19925 ( .A(n19187), .B(n17015), .Z(n18083) );
  XNOR U19926 ( .A(n19188), .B(n18736), .Z(n9649) );
  XOR U19927 ( .A(n19189), .B(n17203), .Z(n17151) );
  XNOR U19928 ( .A(n19190), .B(n18731), .Z(n11506) );
  XOR U19929 ( .A(n19191), .B(n15261), .Z(n17155) );
  XNOR U19930 ( .A(n19192), .B(n19193), .Z(n15261) );
  XOR U19931 ( .A(n19194), .B(n19195), .Z(n12124) );
  XOR U19932 ( .A(n14871), .B(n12712), .Z(n19195) );
  XNOR U19933 ( .A(n19196), .B(n19197), .Z(n12712) );
  AND U19934 ( .A(n14360), .B(n14361), .Z(n19196) );
  XNOR U19935 ( .A(n18070), .B(n19198), .Z(n14361) );
  XOR U19936 ( .A(n19199), .B(n17170), .Z(n14871) );
  ANDN U19937 ( .B(n14355), .A(n14353), .Z(n19199) );
  XOR U19938 ( .A(n19200), .B(n15698), .Z(n14355) );
  IV U19939 ( .A(n19201), .Z(n15698) );
  XOR U19940 ( .A(n15204), .B(n19202), .Z(n19194) );
  XNOR U19941 ( .A(n19203), .B(n13643), .Z(n19202) );
  XOR U19942 ( .A(n19204), .B(n12488), .Z(n13643) );
  ANDN U19943 ( .B(n18981), .A(n17538), .Z(n19204) );
  XOR U19944 ( .A(n19205), .B(n18275), .Z(n17538) );
  NOR U19945 ( .A(n19207), .B(n17529), .Z(n19206) );
  XNOR U19946 ( .A(n19208), .B(n19207), .Z(n14358) );
  IV U19947 ( .A(n19209), .Z(n19207) );
  ANDN U19948 ( .B(n17529), .A(n12472), .Z(n19208) );
  IV U19949 ( .A(n17530), .Z(n12472) );
  XOR U19950 ( .A(n19210), .B(n17626), .Z(n17530) );
  XOR U19951 ( .A(n14162), .B(n19211), .Z(n17529) );
  XOR U19952 ( .A(n16476), .B(n9783), .Z(n6697) );
  XOR U19953 ( .A(n19212), .B(n19213), .Z(n12895) );
  XOR U19954 ( .A(n12904), .B(n10304), .Z(n19213) );
  XOR U19955 ( .A(n19214), .B(n15519), .Z(n10304) );
  NOR U19956 ( .A(n16483), .B(n16484), .Z(n19214) );
  XOR U19957 ( .A(n19215), .B(n18938), .Z(n16484) );
  XOR U19958 ( .A(n19216), .B(n17654), .Z(n16483) );
  XNOR U19959 ( .A(n19217), .B(n15523), .Z(n12904) );
  AND U19960 ( .A(n15522), .B(n16479), .Z(n19217) );
  XOR U19961 ( .A(n17901), .B(n19218), .Z(n16479) );
  IV U19962 ( .A(n18216), .Z(n17901) );
  XNOR U19963 ( .A(n19219), .B(n19220), .Z(n18216) );
  XOR U19964 ( .A(n19221), .B(n18090), .Z(n15522) );
  XNOR U19965 ( .A(n12234), .B(n19222), .Z(n19212) );
  XOR U19966 ( .A(n10859), .B(n15500), .Z(n19222) );
  XNOR U19967 ( .A(n19223), .B(n15510), .Z(n15500) );
  ANDN U19968 ( .B(n18995), .A(n19224), .Z(n19223) );
  XOR U19969 ( .A(n19225), .B(n15515), .Z(n10859) );
  ANDN U19970 ( .B(n15514), .A(n18653), .Z(n19225) );
  XNOR U19971 ( .A(n19226), .B(n16509), .Z(n18653) );
  XOR U19972 ( .A(n19227), .B(n19228), .Z(n15514) );
  XOR U19973 ( .A(n19229), .B(n15505), .Z(n12234) );
  ANDN U19974 ( .B(n16488), .A(n15506), .Z(n19229) );
  XNOR U19975 ( .A(n19230), .B(n18412), .Z(n15506) );
  XOR U19976 ( .A(n19231), .B(n18221), .Z(n16488) );
  XOR U19977 ( .A(n19232), .B(n19233), .Z(n17492) );
  XOR U19978 ( .A(n9542), .B(n10314), .Z(n19233) );
  XOR U19979 ( .A(n19234), .B(n13226), .Z(n10314) );
  XOR U19980 ( .A(n17066), .B(n19235), .Z(n13226) );
  IV U19981 ( .A(n17197), .Z(n17066) );
  ANDN U19982 ( .B(n15538), .A(n14658), .Z(n19234) );
  XNOR U19983 ( .A(n19236), .B(n18712), .Z(n14658) );
  XNOR U19984 ( .A(n17268), .B(n19237), .Z(n15538) );
  XNOR U19985 ( .A(n19238), .B(n13218), .Z(n9542) );
  XOR U19986 ( .A(n19239), .B(n15351), .Z(n13218) );
  XNOR U19987 ( .A(n19240), .B(n19241), .Z(n15351) );
  ANDN U19988 ( .B(n14660), .A(n15542), .Z(n19238) );
  XOR U19989 ( .A(n15875), .B(n19242), .Z(n15542) );
  XOR U19990 ( .A(n19243), .B(n19244), .Z(n14660) );
  XOR U19991 ( .A(n10993), .B(n19245), .Z(n19232) );
  XNOR U19992 ( .A(n12587), .B(n12108), .Z(n19245) );
  XNOR U19993 ( .A(n19246), .B(n13222), .Z(n12108) );
  XNOR U19994 ( .A(n16390), .B(n19247), .Z(n13222) );
  ANDN U19995 ( .B(n15533), .A(n14663), .Z(n19246) );
  XOR U19996 ( .A(n19248), .B(n18186), .Z(n14663) );
  XOR U19997 ( .A(n18014), .B(n19249), .Z(n15533) );
  XOR U19998 ( .A(n19250), .B(n13239), .Z(n12587) );
  XOR U19999 ( .A(n19251), .B(n17297), .Z(n13239) );
  ANDN U20000 ( .B(n15529), .A(n14668), .Z(n19250) );
  IV U20001 ( .A(n16472), .Z(n14668) );
  XNOR U20002 ( .A(n17483), .B(n19252), .Z(n16472) );
  XNOR U20003 ( .A(n19253), .B(n18938), .Z(n15529) );
  XNOR U20004 ( .A(n19254), .B(n13214), .Z(n10993) );
  XOR U20005 ( .A(n19255), .B(n17015), .Z(n13214) );
  XNOR U20006 ( .A(n19256), .B(n19257), .Z(n17015) );
  AND U20007 ( .A(n15546), .B(n14665), .Z(n19254) );
  XOR U20008 ( .A(n19258), .B(n16509), .Z(n14665) );
  XOR U20009 ( .A(n19259), .B(n17028), .Z(n15546) );
  IV U20010 ( .A(n18283), .Z(n17028) );
  XNOR U20011 ( .A(n19260), .B(n15509), .Z(n16476) );
  IV U20012 ( .A(n19224), .Z(n15509) );
  XOR U20013 ( .A(n16082), .B(n19261), .Z(n19224) );
  NOR U20014 ( .A(n18996), .B(n18995), .Z(n19260) );
  XOR U20015 ( .A(n19262), .B(n19263), .Z(n18995) );
  XOR U20016 ( .A(n3748), .B(n19264), .Z(n19017) );
  XOR U20017 ( .A(n5496), .B(n2145), .Z(n19264) );
  XOR U20018 ( .A(n19265), .B(n7232), .Z(n2145) );
  XNOR U20019 ( .A(n9527), .B(n14398), .Z(n7232) );
  XNOR U20020 ( .A(n19266), .B(n14846), .Z(n14398) );
  NOR U20021 ( .A(n17803), .B(n19267), .Z(n19266) );
  XNOR U20022 ( .A(n13511), .B(n12306), .Z(n9527) );
  XOR U20023 ( .A(n19268), .B(n19269), .Z(n12306) );
  XNOR U20024 ( .A(n13472), .B(n13276), .Z(n19269) );
  XOR U20025 ( .A(n19270), .B(n14838), .Z(n13276) );
  XNOR U20026 ( .A(n19271), .B(n14958), .Z(n14838) );
  ANDN U20027 ( .B(n14409), .A(n14410), .Z(n19270) );
  XOR U20028 ( .A(n18814), .B(n19272), .Z(n14409) );
  XNOR U20029 ( .A(n19273), .B(n14842), .Z(n13472) );
  XNOR U20030 ( .A(n17483), .B(n19274), .Z(n14842) );
  NOR U20031 ( .A(n14401), .B(n14400), .Z(n19273) );
  XOR U20032 ( .A(n19275), .B(n18772), .Z(n14400) );
  XOR U20033 ( .A(n10854), .B(n19276), .Z(n19268) );
  XOR U20034 ( .A(n14831), .B(n11566), .Z(n19276) );
  XNOR U20035 ( .A(n19277), .B(n17779), .Z(n11566) );
  XOR U20036 ( .A(n19278), .B(n18706), .Z(n17779) );
  XOR U20037 ( .A(n19279), .B(n19280), .Z(n14405) );
  XNOR U20038 ( .A(n19281), .B(n14845), .Z(n14831) );
  XNOR U20039 ( .A(n18378), .B(n19282), .Z(n14845) );
  XOR U20040 ( .A(n19283), .B(n17647), .Z(n14846) );
  XNOR U20041 ( .A(n19284), .B(n14849), .Z(n10854) );
  XOR U20042 ( .A(n18530), .B(n19285), .Z(n14849) );
  ANDN U20043 ( .B(n14414), .A(n14413), .Z(n19284) );
  XOR U20044 ( .A(n18539), .B(n19286), .Z(n14413) );
  IV U20045 ( .A(n17474), .Z(n18539) );
  XOR U20046 ( .A(n19287), .B(n19288), .Z(n13511) );
  XNOR U20047 ( .A(n12070), .B(n15352), .Z(n19288) );
  XOR U20048 ( .A(n19289), .B(n15357), .Z(n15352) );
  XOR U20049 ( .A(n17926), .B(n19290), .Z(n15357) );
  ANDN U20050 ( .B(n14438), .A(n14435), .Z(n19289) );
  XOR U20051 ( .A(n16961), .B(n19291), .Z(n14435) );
  XOR U20052 ( .A(n19010), .B(n19292), .Z(n14438) );
  IV U20053 ( .A(n18814), .Z(n19010) );
  XOR U20054 ( .A(n19293), .B(n15370), .Z(n12070) );
  XNOR U20055 ( .A(n19294), .B(n15639), .Z(n15370) );
  NOR U20056 ( .A(n14419), .B(n14420), .Z(n19293) );
  XOR U20057 ( .A(n19295), .B(n19296), .Z(n14420) );
  XNOR U20058 ( .A(n19297), .B(n15645), .Z(n14419) );
  XOR U20059 ( .A(n19298), .B(n19299), .Z(n15645) );
  XOR U20060 ( .A(n11061), .B(n19300), .Z(n19287) );
  XOR U20061 ( .A(n13330), .B(n11510), .Z(n19300) );
  XNOR U20062 ( .A(n19301), .B(n15364), .Z(n11510) );
  XOR U20063 ( .A(n18476), .B(n19302), .Z(n15364) );
  ANDN U20064 ( .B(n14432), .A(n14433), .Z(n19301) );
  XOR U20065 ( .A(n19303), .B(n18161), .Z(n14433) );
  XNOR U20066 ( .A(n19304), .B(n18596), .Z(n14432) );
  XNOR U20067 ( .A(n19305), .B(n15367), .Z(n13330) );
  XOR U20068 ( .A(n16082), .B(n19306), .Z(n15367) );
  IV U20069 ( .A(n19307), .Z(n16082) );
  NOR U20070 ( .A(n14425), .B(n14423), .Z(n19305) );
  XNOR U20071 ( .A(n19308), .B(n18277), .Z(n14423) );
  XOR U20072 ( .A(n19310), .B(n19311), .Z(n15875) );
  XOR U20073 ( .A(n19312), .B(n15360), .Z(n11061) );
  XNOR U20074 ( .A(n19313), .B(n15674), .Z(n15360) );
  AND U20075 ( .A(n14428), .B(n14430), .Z(n19312) );
  XOR U20076 ( .A(n17143), .B(n19314), .Z(n14430) );
  XOR U20077 ( .A(n16390), .B(n19315), .Z(n14428) );
  ANDN U20078 ( .B(n6706), .A(n6707), .Z(n19265) );
  XOR U20079 ( .A(n15762), .B(n10496), .Z(n6707) );
  XNOR U20080 ( .A(n13971), .B(n18807), .Z(n10496) );
  XOR U20081 ( .A(n19316), .B(n19317), .Z(n18807) );
  XNOR U20082 ( .A(n14366), .B(n10213), .Z(n19317) );
  XNOR U20083 ( .A(n19318), .B(n15232), .Z(n10213) );
  XOR U20084 ( .A(n19319), .B(n17301), .Z(n15232) );
  ANDN U20085 ( .B(n15233), .A(n14077), .Z(n19318) );
  XOR U20086 ( .A(n19320), .B(n19321), .Z(n14077) );
  XOR U20087 ( .A(n19322), .B(n16502), .Z(n15233) );
  XNOR U20088 ( .A(n19323), .B(n15239), .Z(n14366) );
  XOR U20089 ( .A(n19324), .B(n19325), .Z(n15239) );
  AND U20090 ( .A(n14081), .B(n15240), .Z(n19323) );
  XOR U20091 ( .A(n18053), .B(n19326), .Z(n15240) );
  XNOR U20092 ( .A(n19327), .B(n17613), .Z(n14081) );
  XOR U20093 ( .A(n11237), .B(n19328), .Z(n19316) );
  XNOR U20094 ( .A(n9133), .B(n12127), .Z(n19328) );
  XNOR U20095 ( .A(n19329), .B(n15244), .Z(n12127) );
  XOR U20096 ( .A(n19330), .B(n16094), .Z(n15244) );
  NOR U20097 ( .A(n14068), .B(n15243), .Z(n19329) );
  XOR U20098 ( .A(n19331), .B(n19035), .Z(n15243) );
  XNOR U20099 ( .A(n19332), .B(n18830), .Z(n14068) );
  XNOR U20100 ( .A(n19333), .B(n17452), .Z(n9133) );
  XOR U20101 ( .A(n19334), .B(n17980), .Z(n17452) );
  NOR U20102 ( .A(n14072), .B(n15768), .Z(n19333) );
  XNOR U20103 ( .A(n18814), .B(n19335), .Z(n15768) );
  XOR U20104 ( .A(n18179), .B(n19336), .Z(n18814) );
  XOR U20105 ( .A(n19337), .B(n19338), .Z(n18179) );
  XOR U20106 ( .A(n16517), .B(n14966), .Z(n19338) );
  XOR U20107 ( .A(n19339), .B(n19340), .Z(n14966) );
  NOR U20108 ( .A(n19341), .B(n19342), .Z(n19339) );
  XNOR U20109 ( .A(n19343), .B(n19344), .Z(n16517) );
  NOR U20110 ( .A(n19345), .B(n19346), .Z(n19343) );
  XOR U20111 ( .A(n18344), .B(n19347), .Z(n19337) );
  XNOR U20112 ( .A(n18390), .B(n19348), .Z(n19347) );
  XNOR U20113 ( .A(n19349), .B(n19350), .Z(n18390) );
  NOR U20114 ( .A(n19351), .B(n19352), .Z(n19349) );
  XNOR U20115 ( .A(n19353), .B(n19354), .Z(n18344) );
  NOR U20116 ( .A(n19355), .B(n19356), .Z(n19353) );
  XOR U20117 ( .A(n19357), .B(n18419), .Z(n14072) );
  XNOR U20118 ( .A(n19358), .B(n15237), .Z(n11237) );
  XOR U20119 ( .A(n19359), .B(n17589), .Z(n15237) );
  ANDN U20120 ( .B(n14085), .A(n15236), .Z(n19358) );
  XOR U20121 ( .A(n19360), .B(n19361), .Z(n13971) );
  XNOR U20122 ( .A(n13593), .B(n11815), .Z(n19361) );
  XOR U20123 ( .A(n19362), .B(n14375), .Z(n11815) );
  XOR U20124 ( .A(n19363), .B(n19325), .Z(n14375) );
  ANDN U20125 ( .B(n13105), .A(n13107), .Z(n19362) );
  XNOR U20126 ( .A(n19364), .B(n16737), .Z(n13107) );
  XOR U20127 ( .A(n19365), .B(n18877), .Z(n13105) );
  XNOR U20128 ( .A(n19366), .B(n14380), .Z(n13593) );
  XOR U20129 ( .A(n19367), .B(n19228), .Z(n14380) );
  XOR U20130 ( .A(n19368), .B(n19369), .Z(n13969) );
  XOR U20131 ( .A(n19370), .B(n18683), .Z(n13968) );
  XNOR U20132 ( .A(n13005), .B(n19371), .Z(n19360) );
  XNOR U20133 ( .A(n10949), .B(n12982), .Z(n19371) );
  XOR U20134 ( .A(n19372), .B(n15772), .Z(n12982) );
  XOR U20135 ( .A(n19373), .B(n19374), .Z(n15772) );
  NOR U20136 ( .A(n17115), .B(n13100), .Z(n19372) );
  XNOR U20137 ( .A(n19375), .B(n18234), .Z(n13100) );
  IV U20138 ( .A(n13101), .Z(n17115) );
  XNOR U20139 ( .A(n19376), .B(n17105), .Z(n13101) );
  XOR U20140 ( .A(n19377), .B(n14372), .Z(n10949) );
  XOR U20141 ( .A(n19378), .B(n16809), .Z(n14372) );
  XOR U20142 ( .A(n19379), .B(n16830), .Z(n13110) );
  XOR U20143 ( .A(n19380), .B(n17907), .Z(n13109) );
  IV U20144 ( .A(n17548), .Z(n17907) );
  XNOR U20145 ( .A(n19381), .B(n17488), .Z(n13005) );
  XOR U20146 ( .A(n19382), .B(n18942), .Z(n17488) );
  XOR U20147 ( .A(n19383), .B(n16868), .Z(n13114) );
  XOR U20148 ( .A(n18100), .B(n19384), .Z(n13113) );
  XNOR U20149 ( .A(n19385), .B(n15236), .Z(n15762) );
  XNOR U20150 ( .A(n19386), .B(n16889), .Z(n15236) );
  XNOR U20151 ( .A(n18014), .B(n19387), .Z(n14085) );
  XOR U20152 ( .A(n19388), .B(n19389), .Z(n14087) );
  XNOR U20153 ( .A(n13831), .B(n10075), .Z(n6706) );
  XNOR U20154 ( .A(n17720), .B(n13207), .Z(n10075) );
  XNOR U20155 ( .A(n19390), .B(n19391), .Z(n13207) );
  XOR U20156 ( .A(n13654), .B(n12709), .Z(n19391) );
  XNOR U20157 ( .A(n19392), .B(n16487), .Z(n12709) );
  XNOR U20158 ( .A(n19393), .B(n18295), .Z(n16487) );
  ANDN U20159 ( .B(n15504), .A(n15505), .Z(n19392) );
  XOR U20160 ( .A(n19394), .B(n16996), .Z(n15505) );
  XOR U20161 ( .A(n19395), .B(n19396), .Z(n15504) );
  XOR U20162 ( .A(n19397), .B(n18996), .Z(n13654) );
  XOR U20163 ( .A(n19398), .B(n16367), .Z(n18996) );
  AND U20164 ( .A(n15508), .B(n15510), .Z(n19397) );
  XOR U20165 ( .A(n19399), .B(n19400), .Z(n15510) );
  XOR U20166 ( .A(n19401), .B(n18621), .Z(n15508) );
  XOR U20167 ( .A(n12788), .B(n19402), .Z(n19390) );
  XOR U20168 ( .A(n10342), .B(n14653), .Z(n19402) );
  XNOR U20169 ( .A(n19403), .B(n18654), .Z(n14653) );
  XOR U20170 ( .A(n19404), .B(n14970), .Z(n18654) );
  XNOR U20171 ( .A(n19405), .B(n19406), .Z(n18264) );
  XOR U20172 ( .A(n18797), .B(n19407), .Z(n19406) );
  XOR U20173 ( .A(n19408), .B(n19409), .Z(n18797) );
  ANDN U20174 ( .B(n19410), .A(n19411), .Z(n19408) );
  XNOR U20175 ( .A(n17540), .B(n19412), .Z(n19405) );
  XNOR U20176 ( .A(n19413), .B(n19414), .Z(n19412) );
  XNOR U20177 ( .A(n19415), .B(n19416), .Z(n17540) );
  NOR U20178 ( .A(n19417), .B(n19418), .Z(n19415) );
  ANDN U20179 ( .B(n15513), .A(n15515), .Z(n19403) );
  XNOR U20180 ( .A(n19420), .B(n16094), .Z(n15515) );
  XOR U20181 ( .A(n19421), .B(n19422), .Z(n16094) );
  XOR U20182 ( .A(n19423), .B(n17209), .Z(n15513) );
  IV U20183 ( .A(n18397), .Z(n17209) );
  XNOR U20184 ( .A(n19424), .B(n16485), .Z(n10342) );
  XNOR U20185 ( .A(n19425), .B(n17197), .Z(n16485) );
  XOR U20186 ( .A(n19426), .B(n19427), .Z(n17197) );
  ANDN U20187 ( .B(n15519), .A(n15517), .Z(n19424) );
  XOR U20188 ( .A(n19428), .B(n16088), .Z(n15517) );
  XNOR U20189 ( .A(n19429), .B(n16511), .Z(n15519) );
  IV U20190 ( .A(n18197), .Z(n16511) );
  XNOR U20191 ( .A(n19430), .B(n16478), .Z(n12788) );
  XNOR U20192 ( .A(n19431), .B(n19037), .Z(n16478) );
  ANDN U20193 ( .B(n15523), .A(n15521), .Z(n19430) );
  IV U20194 ( .A(n18991), .Z(n15521) );
  XOR U20195 ( .A(n19432), .B(n19035), .Z(n18991) );
  XOR U20196 ( .A(n19433), .B(n17632), .Z(n15523) );
  XOR U20197 ( .A(n19434), .B(n19435), .Z(n17720) );
  XNOR U20198 ( .A(n10828), .B(n18979), .Z(n19435) );
  XOR U20199 ( .A(n19436), .B(n15402), .Z(n18979) );
  XOR U20200 ( .A(n19437), .B(n18419), .Z(n15402) );
  AND U20201 ( .A(n13828), .B(n13827), .Z(n19436) );
  XOR U20202 ( .A(n16048), .B(n19439), .Z(n13828) );
  IV U20203 ( .A(n15299), .Z(n16048) );
  XNOR U20204 ( .A(n19440), .B(n15393), .Z(n10828) );
  XOR U20205 ( .A(n18621), .B(n19441), .Z(n15393) );
  IV U20206 ( .A(n19442), .Z(n18621) );
  NOR U20207 ( .A(n13837), .B(n13838), .Z(n19440) );
  XOR U20208 ( .A(n19443), .B(n19444), .Z(n13838) );
  IV U20209 ( .A(n19016), .Z(n13837) );
  XNOR U20210 ( .A(n19445), .B(n17861), .Z(n19016) );
  XOR U20211 ( .A(n11809), .B(n19446), .Z(n19434) );
  XOR U20212 ( .A(n9638), .B(n18986), .Z(n19446) );
  XNOR U20213 ( .A(n19447), .B(n15398), .Z(n18986) );
  XOR U20214 ( .A(n19295), .B(n19448), .Z(n15398) );
  ANDN U20215 ( .B(n17842), .A(n19008), .Z(n19447) );
  XNOR U20216 ( .A(n19449), .B(n15408), .Z(n9638) );
  XOR U20217 ( .A(n19450), .B(n19451), .Z(n15408) );
  XNOR U20218 ( .A(n19452), .B(n17186), .Z(n14588) );
  XOR U20219 ( .A(n19453), .B(n18248), .Z(n14586) );
  XOR U20220 ( .A(n19454), .B(n15406), .Z(n11809) );
  XOR U20221 ( .A(n19455), .B(n19456), .Z(n15406) );
  ANDN U20222 ( .B(n13835), .A(n13833), .Z(n19454) );
  IV U20223 ( .A(n19002), .Z(n13833) );
  XOR U20224 ( .A(n19457), .B(n19037), .Z(n19002) );
  IV U20225 ( .A(n18167), .Z(n19037) );
  XOR U20226 ( .A(n19458), .B(n19459), .Z(n18167) );
  XOR U20227 ( .A(n19460), .B(n18221), .Z(n13835) );
  XOR U20228 ( .A(n19461), .B(n19008), .Z(n13831) );
  XOR U20229 ( .A(n19462), .B(n16305), .Z(n19008) );
  NOR U20230 ( .A(n15396), .B(n17842), .Z(n19461) );
  XNOR U20231 ( .A(n19463), .B(n18561), .Z(n17842) );
  XOR U20232 ( .A(n19464), .B(n18613), .Z(n15396) );
  IV U20233 ( .A(n18517), .Z(n18613) );
  XNOR U20234 ( .A(n19467), .B(n9464), .Z(n5496) );
  IV U20235 ( .A(n9343), .Z(n9464) );
  XOR U20236 ( .A(n15153), .B(n9450), .Z(n9343) );
  XOR U20237 ( .A(n19468), .B(n19469), .Z(n14692) );
  XNOR U20238 ( .A(n9556), .B(n10055), .Z(n19469) );
  XNOR U20239 ( .A(n19470), .B(n19471), .Z(n10055) );
  ANDN U20240 ( .B(n15146), .A(n15145), .Z(n19470) );
  IV U20241 ( .A(n19472), .Z(n15146) );
  XOR U20242 ( .A(n19473), .B(n16693), .Z(n9556) );
  XOR U20243 ( .A(n19474), .B(n19475), .Z(n19468) );
  XOR U20244 ( .A(n12967), .B(n12892), .Z(n19475) );
  XOR U20245 ( .A(n19476), .B(n16686), .Z(n12892) );
  AND U20246 ( .A(n15156), .B(n15155), .Z(n19476) );
  XNOR U20247 ( .A(n19477), .B(n19478), .Z(n12967) );
  ANDN U20248 ( .B(n19479), .A(n19480), .Z(n19477) );
  XOR U20249 ( .A(n19481), .B(n19482), .Z(n17727) );
  XOR U20250 ( .A(n12626), .B(n9898), .Z(n19482) );
  XOR U20251 ( .A(n19483), .B(n16669), .Z(n9898) );
  ANDN U20252 ( .B(n15040), .A(n13344), .Z(n19483) );
  XOR U20253 ( .A(n19484), .B(n17098), .Z(n13344) );
  XNOR U20254 ( .A(n19485), .B(n16681), .Z(n12626) );
  NOR U20255 ( .A(n14484), .B(n15036), .Z(n19485) );
  XOR U20256 ( .A(n19486), .B(n16613), .Z(n14484) );
  XNOR U20257 ( .A(n16201), .B(n19487), .Z(n19481) );
  XNOR U20258 ( .A(n16553), .B(n9973), .Z(n19487) );
  XNOR U20259 ( .A(n19488), .B(n16677), .Z(n9973) );
  AND U20260 ( .A(n17725), .B(n13348), .Z(n19488) );
  XNOR U20261 ( .A(n17746), .B(n19489), .Z(n13348) );
  XOR U20262 ( .A(n19490), .B(n16675), .Z(n16553) );
  ANDN U20263 ( .B(n15034), .A(n14873), .Z(n19490) );
  XNOR U20264 ( .A(n19491), .B(n16841), .Z(n14873) );
  XNOR U20265 ( .A(n19492), .B(n16665), .Z(n16201) );
  ANDN U20266 ( .B(n15042), .A(n13338), .Z(n19492) );
  XNOR U20267 ( .A(n19493), .B(n16086), .Z(n13338) );
  XNOR U20268 ( .A(n19494), .B(n19480), .Z(n15153) );
  NOR U20269 ( .A(n19479), .B(n16696), .Z(n19494) );
  NOR U20270 ( .A(n9428), .B(n6710), .Z(n19467) );
  XOR U20271 ( .A(n12717), .B(n15020), .Z(n6710) );
  XNOR U20272 ( .A(n19495), .B(n16195), .Z(n15020) );
  ANDN U20273 ( .B(n18140), .A(n19145), .Z(n19495) );
  XOR U20274 ( .A(n19496), .B(n18877), .Z(n18140) );
  IV U20275 ( .A(n9459), .Z(n12717) );
  XOR U20276 ( .A(n13308), .B(n15910), .Z(n9459) );
  XNOR U20277 ( .A(n19497), .B(n19498), .Z(n15910) );
  XOR U20278 ( .A(n14582), .B(n15769), .Z(n19498) );
  XOR U20279 ( .A(n19499), .B(n16188), .Z(n15769) );
  XOR U20280 ( .A(n19500), .B(n17632), .Z(n16188) );
  ANDN U20281 ( .B(n15026), .A(n15027), .Z(n19499) );
  XOR U20282 ( .A(n19501), .B(n19389), .Z(n15027) );
  XNOR U20283 ( .A(n19502), .B(n15528), .Z(n15026) );
  XNOR U20284 ( .A(n19503), .B(n16192), .Z(n14582) );
  XOR U20285 ( .A(n19504), .B(n18791), .Z(n16192) );
  ANDN U20286 ( .B(n15012), .A(n15013), .Z(n19503) );
  XOR U20287 ( .A(n18302), .B(n19505), .Z(n15013) );
  XNOR U20288 ( .A(n19506), .B(n16078), .Z(n15012) );
  XOR U20289 ( .A(n11495), .B(n19507), .Z(n19497) );
  XOR U20290 ( .A(n11363), .B(n16178), .Z(n19507) );
  XNOR U20291 ( .A(n19508), .B(n18141), .Z(n16178) );
  XNOR U20292 ( .A(n15962), .B(n19509), .Z(n18141) );
  ANDN U20293 ( .B(n19145), .A(n16195), .Z(n19508) );
  XOR U20294 ( .A(n19510), .B(n19511), .Z(n16195) );
  XOR U20295 ( .A(n19512), .B(n16088), .Z(n19145) );
  XNOR U20296 ( .A(n19513), .B(n16199), .Z(n11363) );
  XNOR U20297 ( .A(n19514), .B(n16872), .Z(n16199) );
  IV U20298 ( .A(n18452), .Z(n16872) );
  XOR U20299 ( .A(n19515), .B(n19516), .Z(n18452) );
  NOR U20300 ( .A(n15016), .B(n15017), .Z(n19513) );
  XOR U20301 ( .A(n19517), .B(n18687), .Z(n15017) );
  IV U20302 ( .A(n16200), .Z(n15016) );
  XOR U20303 ( .A(n19442), .B(n19518), .Z(n16200) );
  XNOR U20304 ( .A(n19519), .B(n16185), .Z(n11495) );
  XOR U20305 ( .A(n19520), .B(n17601), .Z(n16185) );
  NOR U20306 ( .A(n15022), .B(n15023), .Z(n19519) );
  XNOR U20307 ( .A(n16855), .B(n19521), .Z(n15023) );
  IV U20308 ( .A(n14952), .Z(n16855) );
  XNOR U20309 ( .A(n19522), .B(n19047), .Z(n14952) );
  XNOR U20310 ( .A(n19523), .B(n19524), .Z(n19047) );
  XNOR U20311 ( .A(n19525), .B(n18194), .Z(n19524) );
  XNOR U20312 ( .A(n19526), .B(n19527), .Z(n18194) );
  ANDN U20313 ( .B(n19528), .A(n19529), .Z(n19526) );
  XOR U20314 ( .A(n19530), .B(n19531), .Z(n19523) );
  XNOR U20315 ( .A(n15531), .B(n18229), .Z(n19531) );
  XNOR U20316 ( .A(n19532), .B(n19533), .Z(n18229) );
  NOR U20317 ( .A(n19534), .B(n19535), .Z(n19532) );
  XNOR U20318 ( .A(n19536), .B(n19537), .Z(n15531) );
  NOR U20319 ( .A(n19538), .B(n19539), .Z(n19536) );
  IV U20320 ( .A(n16184), .Z(n15022) );
  XNOR U20321 ( .A(n19540), .B(n18186), .Z(n16184) );
  XOR U20322 ( .A(n19541), .B(n19542), .Z(n13308) );
  XOR U20323 ( .A(n18405), .B(n11717), .Z(n19542) );
  XOR U20324 ( .A(n19543), .B(n14826), .Z(n11717) );
  XOR U20325 ( .A(n19544), .B(n18502), .Z(n14826) );
  ANDN U20326 ( .B(n15615), .A(n15614), .Z(n19543) );
  XOR U20327 ( .A(n19545), .B(n19444), .Z(n15614) );
  XNOR U20328 ( .A(n17321), .B(n19546), .Z(n15615) );
  XOR U20329 ( .A(n19547), .B(n15859), .Z(n18405) );
  XOR U20330 ( .A(n18100), .B(n19548), .Z(n15859) );
  ANDN U20331 ( .B(n15603), .A(n16382), .Z(n19547) );
  XOR U20332 ( .A(n19549), .B(n15265), .Z(n16382) );
  XOR U20333 ( .A(n19550), .B(n19551), .Z(n15603) );
  XOR U20334 ( .A(n10197), .B(n19552), .Z(n19541) );
  XOR U20335 ( .A(n11880), .B(n11803), .Z(n19552) );
  XNOR U20336 ( .A(n19553), .B(n14819), .Z(n11803) );
  XOR U20337 ( .A(n19554), .B(n16509), .Z(n14819) );
  ANDN U20338 ( .B(n15611), .A(n15612), .Z(n19553) );
  XOR U20339 ( .A(n19555), .B(n17853), .Z(n15612) );
  XOR U20340 ( .A(n19559), .B(n16413), .Z(n11880) );
  XNOR U20341 ( .A(n17926), .B(n19560), .Z(n16413) );
  IV U20342 ( .A(n17619), .Z(n17926) );
  NOR U20343 ( .A(n16385), .B(n15599), .Z(n19559) );
  XOR U20344 ( .A(n19561), .B(n15688), .Z(n15599) );
  IV U20345 ( .A(n15600), .Z(n16385) );
  XOR U20346 ( .A(n19562), .B(n17533), .Z(n15600) );
  IV U20347 ( .A(n19025), .Z(n17533) );
  XOR U20348 ( .A(n19563), .B(n18552), .Z(n19025) );
  XNOR U20349 ( .A(n19564), .B(n19565), .Z(n18552) );
  XNOR U20350 ( .A(n18708), .B(n17726), .Z(n19565) );
  XNOR U20351 ( .A(n19566), .B(n19567), .Z(n17726) );
  ANDN U20352 ( .B(n19568), .A(n19569), .Z(n19566) );
  XNOR U20353 ( .A(n19570), .B(n19571), .Z(n18708) );
  XOR U20354 ( .A(n16506), .B(n19574), .Z(n19564) );
  XOR U20355 ( .A(n18953), .B(n17734), .Z(n19574) );
  XOR U20356 ( .A(n19575), .B(n19576), .Z(n17734) );
  ANDN U20357 ( .B(n19577), .A(n19578), .Z(n19575) );
  XOR U20358 ( .A(n19579), .B(n19580), .Z(n18953) );
  ANDN U20359 ( .B(n19581), .A(n19582), .Z(n19579) );
  XNOR U20360 ( .A(n19583), .B(n19584), .Z(n16506) );
  ANDN U20361 ( .B(n19585), .A(n19586), .Z(n19583) );
  XNOR U20362 ( .A(n19587), .B(n14815), .Z(n10197) );
  XOR U20363 ( .A(n16844), .B(n19588), .Z(n14815) );
  ANDN U20364 ( .B(n15608), .A(n16372), .Z(n19587) );
  XOR U20365 ( .A(n19589), .B(n18830), .Z(n16372) );
  XNOR U20366 ( .A(n19590), .B(n17578), .Z(n15608) );
  IV U20367 ( .A(n6711), .Z(n9428) );
  XNOR U20368 ( .A(n17603), .B(n10065), .Z(n6711) );
  XNOR U20369 ( .A(n19591), .B(n13964), .Z(n17603) );
  ANDN U20370 ( .B(n13153), .A(n15254), .Z(n19591) );
  IV U20371 ( .A(n19592), .Z(n15254) );
  XOR U20372 ( .A(n19593), .B(n16088), .Z(n13153) );
  XOR U20373 ( .A(n19594), .B(n19595), .Z(n16088) );
  XNOR U20374 ( .A(n19596), .B(n7224), .Z(n3748) );
  IV U20375 ( .A(n9347), .Z(n7224) );
  XOR U20376 ( .A(n17760), .B(n11902), .Z(n9347) );
  XNOR U20377 ( .A(n11836), .B(n11848), .Z(n11902) );
  XNOR U20378 ( .A(n19597), .B(n19598), .Z(n11848) );
  XNOR U20379 ( .A(n10994), .B(n11692), .Z(n19598) );
  XOR U20380 ( .A(n19599), .B(n16545), .Z(n11692) );
  NOR U20381 ( .A(n16544), .B(n14785), .Z(n19599) );
  XOR U20382 ( .A(n19600), .B(n19069), .Z(n14785) );
  XNOR U20383 ( .A(n19601), .B(n19451), .Z(n16544) );
  XOR U20384 ( .A(n19602), .B(n16569), .Z(n10994) );
  NOR U20385 ( .A(n16568), .B(n14777), .Z(n19602) );
  XOR U20386 ( .A(n18769), .B(n19603), .Z(n14777) );
  XOR U20387 ( .A(n15639), .B(n19604), .Z(n16568) );
  XNOR U20388 ( .A(n10740), .B(n19605), .Z(n19597) );
  XOR U20389 ( .A(n16175), .B(n11915), .Z(n19605) );
  XOR U20390 ( .A(n19606), .B(n18483), .Z(n11915) );
  ANDN U20391 ( .B(n17775), .A(n14781), .Z(n19606) );
  XOR U20392 ( .A(n19607), .B(n16575), .Z(n14781) );
  XNOR U20393 ( .A(n19608), .B(n18165), .Z(n17775) );
  XOR U20394 ( .A(n19609), .B(n16538), .Z(n16175) );
  ANDN U20395 ( .B(n16539), .A(n14768), .Z(n19609) );
  XOR U20396 ( .A(n15299), .B(n19610), .Z(n14768) );
  XOR U20397 ( .A(n19611), .B(n18949), .Z(n16539) );
  XNOR U20398 ( .A(n19612), .B(n16548), .Z(n10740) );
  XOR U20399 ( .A(n19613), .B(n15891), .Z(n14772) );
  XNOR U20400 ( .A(n18638), .B(n19614), .Z(n15891) );
  XOR U20401 ( .A(n19615), .B(n19616), .Z(n18638) );
  XNOR U20402 ( .A(n19462), .B(n19617), .Z(n19616) );
  XNOR U20403 ( .A(n19618), .B(n19619), .Z(n19462) );
  NOR U20404 ( .A(n19620), .B(n19621), .Z(n19618) );
  XOR U20405 ( .A(n19622), .B(n19623), .Z(n19615) );
  XOR U20406 ( .A(n16304), .B(n19624), .Z(n19623) );
  XNOR U20407 ( .A(n19625), .B(n19626), .Z(n16304) );
  NOR U20408 ( .A(n19627), .B(n19628), .Z(n19625) );
  XNOR U20409 ( .A(n19629), .B(n18400), .Z(n16549) );
  XOR U20410 ( .A(n19630), .B(n19631), .Z(n11836) );
  XOR U20411 ( .A(n16532), .B(n13943), .Z(n19631) );
  XNOR U20412 ( .A(n19632), .B(n17383), .Z(n13943) );
  ANDN U20413 ( .B(n17384), .A(n17762), .Z(n19632) );
  XNOR U20414 ( .A(n19633), .B(n18777), .Z(n17384) );
  XNOR U20415 ( .A(n19634), .B(n17380), .Z(n16532) );
  NOR U20416 ( .A(n17379), .B(n17758), .Z(n19634) );
  XOR U20417 ( .A(n19635), .B(n16465), .Z(n17379) );
  XOR U20418 ( .A(n12403), .B(n19636), .Z(n19630) );
  XOR U20419 ( .A(n13509), .B(n12116), .Z(n19636) );
  XOR U20420 ( .A(n19637), .B(n17370), .Z(n12116) );
  ANDN U20421 ( .B(n17371), .A(n19638), .Z(n19637) );
  XOR U20422 ( .A(n19639), .B(n19640), .Z(n13509) );
  NOR U20423 ( .A(n18352), .B(n18350), .Z(n19639) );
  XNOR U20424 ( .A(n19641), .B(n17375), .Z(n12403) );
  ANDN U20425 ( .B(n17376), .A(n17765), .Z(n19641) );
  XNOR U20426 ( .A(n19642), .B(n17630), .Z(n17376) );
  XOR U20427 ( .A(n19643), .B(n17371), .Z(n17760) );
  XOR U20428 ( .A(n19644), .B(n19321), .Z(n17371) );
  ANDN U20429 ( .B(n6701), .A(n6703), .Z(n19596) );
  XOR U20430 ( .A(n15176), .B(n11842), .Z(n6703) );
  XNOR U20431 ( .A(n19646), .B(n14627), .Z(n15176) );
  IV U20432 ( .A(n19647), .Z(n14627) );
  NOR U20433 ( .A(n16599), .B(n16490), .Z(n19646) );
  XOR U20434 ( .A(n19648), .B(n16575), .Z(n16490) );
  IV U20435 ( .A(n19649), .Z(n16575) );
  XOR U20436 ( .A(n9153), .B(n13311), .Z(n6701) );
  XOR U20437 ( .A(n19650), .B(n13882), .Z(n13311) );
  AND U20438 ( .A(n15620), .B(n15621), .Z(n19650) );
  XNOR U20439 ( .A(n19651), .B(n19228), .Z(n15621) );
  IV U20440 ( .A(n17215), .Z(n19228) );
  XOR U20441 ( .A(n19652), .B(n19653), .Z(n17215) );
  XNOR U20442 ( .A(n14185), .B(n18406), .Z(n9153) );
  XOR U20443 ( .A(n19654), .B(n19655), .Z(n18406) );
  XOR U20444 ( .A(n12211), .B(n12891), .Z(n19655) );
  XNOR U20445 ( .A(n19656), .B(n13886), .Z(n12891) );
  XOR U20446 ( .A(n19657), .B(n19069), .Z(n13886) );
  ANDN U20447 ( .B(n13321), .A(n13319), .Z(n19656) );
  XOR U20448 ( .A(n19658), .B(n19659), .Z(n13319) );
  XOR U20449 ( .A(n19660), .B(n18557), .Z(n13321) );
  XOR U20450 ( .A(n19661), .B(n13890), .Z(n12211) );
  XOR U20451 ( .A(n19662), .B(n15265), .Z(n13890) );
  ANDN U20452 ( .B(n14300), .A(n13889), .Z(n19661) );
  XNOR U20453 ( .A(n19663), .B(n19325), .Z(n13889) );
  IV U20454 ( .A(n19664), .Z(n19325) );
  XNOR U20455 ( .A(n18277), .B(n19665), .Z(n14300) );
  XNOR U20456 ( .A(n11038), .B(n19666), .Z(n19654) );
  XNOR U20457 ( .A(n13868), .B(n12989), .Z(n19666) );
  XNOR U20458 ( .A(n19667), .B(n13874), .Z(n12989) );
  XOR U20459 ( .A(n19668), .B(n18855), .Z(n13874) );
  ANDN U20460 ( .B(n13323), .A(n13324), .Z(n19667) );
  XNOR U20461 ( .A(n19670), .B(n19671), .Z(n16502) );
  XOR U20462 ( .A(n19672), .B(n18766), .Z(n13323) );
  XOR U20463 ( .A(n19673), .B(n13877), .Z(n13868) );
  XNOR U20464 ( .A(n18706), .B(n19674), .Z(n13877) );
  NOR U20465 ( .A(n13315), .B(n13316), .Z(n19673) );
  XOR U20466 ( .A(n19675), .B(n17506), .Z(n13316) );
  IV U20467 ( .A(n19444), .Z(n17506) );
  IV U20468 ( .A(n13878), .Z(n13315) );
  XOR U20469 ( .A(n17272), .B(n19678), .Z(n13878) );
  XNOR U20470 ( .A(n19679), .B(n13883), .Z(n11038) );
  NOR U20471 ( .A(n15620), .B(n13882), .Z(n19679) );
  XOR U20472 ( .A(n19681), .B(n18397), .Z(n13882) );
  XNOR U20473 ( .A(n19682), .B(n18954), .Z(n18397) );
  XOR U20474 ( .A(n19683), .B(n19684), .Z(n18954) );
  XOR U20475 ( .A(n19658), .B(n19685), .Z(n19684) );
  XOR U20476 ( .A(n19686), .B(n19687), .Z(n19658) );
  XOR U20477 ( .A(n19688), .B(n19689), .Z(n19683) );
  XNOR U20478 ( .A(n19550), .B(n19690), .Z(n19689) );
  XNOR U20479 ( .A(n19691), .B(n19692), .Z(n19550) );
  NOR U20480 ( .A(n19576), .B(n19577), .Z(n19691) );
  XOR U20481 ( .A(n19693), .B(n19694), .Z(n15620) );
  XOR U20482 ( .A(n19695), .B(n19696), .Z(n14185) );
  XOR U20483 ( .A(n19107), .B(n12089), .Z(n19696) );
  XNOR U20484 ( .A(n19697), .B(n15133), .Z(n12089) );
  NOR U20485 ( .A(n17251), .B(n17271), .Z(n19697) );
  XOR U20486 ( .A(n19698), .B(n16616), .Z(n17251) );
  XOR U20487 ( .A(n19699), .B(n15141), .Z(n19107) );
  AND U20488 ( .A(n14706), .B(n17256), .Z(n19699) );
  XOR U20489 ( .A(n19700), .B(n16992), .Z(n14706) );
  IV U20490 ( .A(n15644), .Z(n16992) );
  XOR U20491 ( .A(n12695), .B(n19703), .Z(n19695) );
  XOR U20492 ( .A(n19704), .B(n11924), .Z(n19703) );
  XNOR U20493 ( .A(n19705), .B(n15137), .Z(n11924) );
  AND U20494 ( .A(n14696), .B(n17267), .Z(n19705) );
  XNOR U20495 ( .A(n19706), .B(n17548), .Z(n14696) );
  XOR U20496 ( .A(n19707), .B(n19708), .Z(n17548) );
  XOR U20497 ( .A(n19709), .B(n15130), .Z(n12695) );
  ANDN U20498 ( .B(n17259), .A(n14710), .Z(n19709) );
  XOR U20499 ( .A(n19713), .B(n19714), .Z(n6641) );
  XNOR U20500 ( .A(n4907), .B(n4078), .Z(n19714) );
  XNOR U20501 ( .A(n19715), .B(n6677), .Z(n4078) );
  XOR U20502 ( .A(n15937), .B(n12381), .Z(n6677) );
  IV U20503 ( .A(n10833), .Z(n12381) );
  XOR U20504 ( .A(n14476), .B(n12244), .Z(n10833) );
  XNOR U20505 ( .A(n19716), .B(n19717), .Z(n12244) );
  XOR U20506 ( .A(n10266), .B(n11586), .Z(n19717) );
  XNOR U20507 ( .A(n19718), .B(n13186), .Z(n11586) );
  XOR U20508 ( .A(n19719), .B(n18282), .Z(n13186) );
  ANDN U20509 ( .B(n13668), .A(n13185), .Z(n19718) );
  XOR U20510 ( .A(n19720), .B(n18400), .Z(n13185) );
  XNOR U20511 ( .A(n19721), .B(n17136), .Z(n13668) );
  IV U20512 ( .A(n18429), .Z(n17136) );
  XNOR U20513 ( .A(n19722), .B(n13199), .Z(n10266) );
  IV U20514 ( .A(n18024), .Z(n13199) );
  XOR U20515 ( .A(n19723), .B(n17982), .Z(n18024) );
  XNOR U20516 ( .A(n19724), .B(n19725), .Z(n17982) );
  ANDN U20517 ( .B(n13665), .A(n13198), .Z(n19722) );
  XNOR U20518 ( .A(n9235), .B(n19726), .Z(n19716) );
  XOR U20519 ( .A(n9152), .B(n11438), .Z(n19726) );
  XNOR U20520 ( .A(n19727), .B(n13191), .Z(n11438) );
  IV U20521 ( .A(n18020), .Z(n13191) );
  XOR U20522 ( .A(n18843), .B(n14962), .Z(n18020) );
  IV U20523 ( .A(n18266), .Z(n14962) );
  XNOR U20524 ( .A(n19728), .B(n19729), .Z(n18843) );
  ANDN U20525 ( .B(n19730), .A(n19731), .Z(n19728) );
  ANDN U20526 ( .B(n13803), .A(n13190), .Z(n19727) );
  XOR U20527 ( .A(n19732), .B(n17098), .Z(n13190) );
  XOR U20528 ( .A(n19733), .B(n18203), .Z(n13803) );
  XOR U20529 ( .A(n19736), .B(n13195), .Z(n9152) );
  XOR U20530 ( .A(n19737), .B(n16737), .Z(n13195) );
  XOR U20531 ( .A(n17921), .B(n19738), .Z(n13194) );
  XOR U20532 ( .A(n19739), .B(n16061), .Z(n13660) );
  IV U20533 ( .A(n19740), .Z(n16061) );
  XOR U20534 ( .A(n19741), .B(n18010), .Z(n9235) );
  XNOR U20535 ( .A(n14158), .B(n19158), .Z(n18010) );
  XOR U20536 ( .A(n19742), .B(n19743), .Z(n19158) );
  AND U20537 ( .A(n15943), .B(n13789), .Z(n19741) );
  XOR U20538 ( .A(n19748), .B(n19749), .Z(n13789) );
  XOR U20539 ( .A(n19750), .B(n18248), .Z(n15943) );
  IV U20540 ( .A(n19751), .Z(n18248) );
  XOR U20541 ( .A(n19752), .B(n19753), .Z(n14476) );
  XOR U20542 ( .A(n14616), .B(n12223), .Z(n19753) );
  XOR U20543 ( .A(n19754), .B(n14648), .Z(n12223) );
  XOR U20544 ( .A(n18769), .B(n19755), .Z(n14648) );
  IV U20545 ( .A(n16727), .Z(n18769) );
  ANDN U20546 ( .B(n13686), .A(n13815), .Z(n19754) );
  XNOR U20547 ( .A(n19756), .B(n19757), .Z(n13815) );
  XOR U20548 ( .A(n18004), .B(n19758), .Z(n13686) );
  XNOR U20549 ( .A(n19759), .B(n14640), .Z(n14616) );
  XOR U20550 ( .A(n19760), .B(n18070), .Z(n14640) );
  NOR U20551 ( .A(n13682), .B(n14478), .Z(n19759) );
  XOR U20552 ( .A(n19761), .B(n16409), .Z(n14478) );
  XOR U20553 ( .A(n19510), .B(n19762), .Z(n13682) );
  IV U20554 ( .A(n16600), .Z(n19510) );
  XOR U20555 ( .A(n19763), .B(n19764), .Z(n16600) );
  XOR U20556 ( .A(n14584), .B(n19765), .Z(n19752) );
  XOR U20557 ( .A(n11491), .B(n10989), .Z(n19765) );
  XNOR U20558 ( .A(n19766), .B(n14646), .Z(n10989) );
  XNOR U20559 ( .A(n19767), .B(n16889), .Z(n14646) );
  AND U20560 ( .A(n13810), .B(n13677), .Z(n19766) );
  XNOR U20561 ( .A(n19768), .B(n19769), .Z(n13677) );
  XOR U20562 ( .A(n19770), .B(n17020), .Z(n13810) );
  XNOR U20563 ( .A(n19771), .B(n14643), .Z(n11491) );
  XNOR U20564 ( .A(n17467), .B(n19772), .Z(n14643) );
  IV U20565 ( .A(n15999), .Z(n17467) );
  XNOR U20566 ( .A(n19773), .B(n19774), .Z(n15999) );
  NOR U20567 ( .A(n13813), .B(n13690), .Z(n19771) );
  XOR U20568 ( .A(n19693), .B(n19775), .Z(n13690) );
  IV U20569 ( .A(n16844), .Z(n19693) );
  XOR U20570 ( .A(n19240), .B(n19776), .Z(n16844) );
  XOR U20571 ( .A(n19777), .B(n19778), .Z(n19240) );
  XNOR U20572 ( .A(n19779), .B(n19780), .Z(n19778) );
  XNOR U20573 ( .A(n19781), .B(n19782), .Z(n19777) );
  XNOR U20574 ( .A(n17869), .B(n19783), .Z(n19782) );
  XNOR U20575 ( .A(n19784), .B(n19785), .Z(n17869) );
  XNOR U20576 ( .A(n19787), .B(n16112), .Z(n13813) );
  XNOR U20577 ( .A(n19788), .B(n14650), .Z(n14584) );
  XOR U20578 ( .A(n18103), .B(n19789), .Z(n14650) );
  ANDN U20579 ( .B(n13817), .A(n13673), .Z(n19788) );
  IV U20580 ( .A(n13818), .Z(n13673) );
  XOR U20581 ( .A(n19790), .B(n18237), .Z(n13818) );
  XNOR U20582 ( .A(n19792), .B(n19793), .Z(n16036) );
  XOR U20583 ( .A(n19794), .B(n13198), .Z(n15937) );
  XOR U20584 ( .A(n19795), .B(n15296), .Z(n13198) );
  IV U20585 ( .A(n15883), .Z(n15296) );
  NOR U20586 ( .A(n13666), .B(n13665), .Z(n19794) );
  XOR U20587 ( .A(n19796), .B(n17520), .Z(n13665) );
  IV U20588 ( .A(n17301), .Z(n17520) );
  XOR U20589 ( .A(n19086), .B(n19797), .Z(n17301) );
  XNOR U20590 ( .A(n19798), .B(n19799), .Z(n19086) );
  XNOR U20591 ( .A(n15633), .B(n15540), .Z(n19799) );
  XNOR U20592 ( .A(n19800), .B(n19801), .Z(n15540) );
  NOR U20593 ( .A(n19802), .B(n19803), .Z(n19800) );
  XNOR U20594 ( .A(n19804), .B(n19805), .Z(n15633) );
  NOR U20595 ( .A(n19806), .B(n19807), .Z(n19804) );
  XOR U20596 ( .A(n16500), .B(n19808), .Z(n19798) );
  XOR U20597 ( .A(n16144), .B(n18699), .Z(n19808) );
  XNOR U20598 ( .A(n19809), .B(n19810), .Z(n18699) );
  NOR U20599 ( .A(n19811), .B(n19812), .Z(n19809) );
  XNOR U20600 ( .A(n19813), .B(n19814), .Z(n16144) );
  ANDN U20601 ( .B(n19815), .A(n19816), .Z(n19813) );
  XOR U20602 ( .A(n19817), .B(n19818), .Z(n16500) );
  ANDN U20603 ( .B(n19819), .A(n19820), .Z(n19817) );
  XNOR U20604 ( .A(n16733), .B(n19821), .Z(n13666) );
  IV U20605 ( .A(n14992), .Z(n16733) );
  XOR U20606 ( .A(n19822), .B(n19823), .Z(n14992) );
  ANDN U20607 ( .B(n9272), .A(n7135), .Z(n19715) );
  XNOR U20608 ( .A(n16978), .B(n9949), .Z(n7135) );
  XNOR U20609 ( .A(n18255), .B(n11833), .Z(n9949) );
  XNOR U20610 ( .A(n19824), .B(n19825), .Z(n11833) );
  XNOR U20611 ( .A(n15745), .B(n11555), .Z(n19825) );
  XOR U20612 ( .A(n19826), .B(n17765), .Z(n11555) );
  XOR U20613 ( .A(n19827), .B(n17918), .Z(n17765) );
  XNOR U20614 ( .A(n19828), .B(n19829), .Z(n17918) );
  ANDN U20615 ( .B(n17766), .A(n19830), .Z(n19826) );
  XNOR U20616 ( .A(n19831), .B(n19638), .Z(n15745) );
  XOR U20617 ( .A(n16822), .B(n19832), .Z(n19638) );
  ANDN U20618 ( .B(n19645), .A(n17369), .Z(n19831) );
  XOR U20619 ( .A(n11041), .B(n19833), .Z(n19824) );
  XNOR U20620 ( .A(n10879), .B(n17752), .Z(n19833) );
  XNOR U20621 ( .A(n19834), .B(n17758), .Z(n17752) );
  XNOR U20622 ( .A(n19835), .B(n18433), .Z(n17758) );
  ANDN U20623 ( .B(n17378), .A(n17757), .Z(n19834) );
  XNOR U20624 ( .A(n19836), .B(n17762), .Z(n10879) );
  XOR U20625 ( .A(n19837), .B(n16737), .Z(n17762) );
  ANDN U20626 ( .B(n17763), .A(n17382), .Z(n19836) );
  XNOR U20627 ( .A(n19840), .B(n18352), .Z(n11041) );
  XNOR U20628 ( .A(n19617), .B(n19841), .Z(n18352) );
  XOR U20629 ( .A(n19842), .B(n19843), .Z(n19617) );
  ANDN U20630 ( .B(n19844), .A(n19845), .Z(n19842) );
  ANDN U20631 ( .B(n19846), .A(n18351), .Z(n19840) );
  XOR U20632 ( .A(n19847), .B(n19848), .Z(n18255) );
  XNOR U20633 ( .A(n14591), .B(n13375), .Z(n19848) );
  XOR U20634 ( .A(n19849), .B(n14008), .Z(n13375) );
  XOR U20635 ( .A(n18027), .B(n19850), .Z(n14008) );
  NOR U20636 ( .A(n16980), .B(n14604), .Z(n19849) );
  XOR U20637 ( .A(n19851), .B(n18766), .Z(n14604) );
  XOR U20638 ( .A(n19426), .B(n19852), .Z(n18766) );
  XOR U20639 ( .A(n19853), .B(n19854), .Z(n19426) );
  XOR U20640 ( .A(n19083), .B(n19589), .Z(n19854) );
  XOR U20641 ( .A(n19855), .B(n19856), .Z(n19589) );
  XOR U20642 ( .A(n19859), .B(n19860), .Z(n19083) );
  ANDN U20643 ( .B(n19861), .A(n19862), .Z(n19859) );
  XNOR U20644 ( .A(n18829), .B(n19863), .Z(n19853) );
  XOR U20645 ( .A(n19332), .B(n19864), .Z(n19863) );
  XOR U20646 ( .A(n19865), .B(n19866), .Z(n19332) );
  ANDN U20647 ( .B(n19867), .A(n19868), .Z(n19865) );
  XOR U20648 ( .A(n19869), .B(n19870), .Z(n18829) );
  ANDN U20649 ( .B(n19871), .A(n19872), .Z(n19869) );
  XOR U20650 ( .A(n16071), .B(n19873), .Z(n16980) );
  XNOR U20651 ( .A(n19874), .B(n14601), .Z(n14591) );
  IV U20652 ( .A(n14019), .Z(n14601) );
  XOR U20653 ( .A(n19875), .B(n15635), .Z(n14019) );
  ANDN U20654 ( .B(n16976), .A(n14600), .Z(n19874) );
  IV U20655 ( .A(n16975), .Z(n14600) );
  XOR U20656 ( .A(n19876), .B(n16996), .Z(n16975) );
  IV U20657 ( .A(n16520), .Z(n16996) );
  XOR U20658 ( .A(n19877), .B(n18852), .Z(n16520) );
  XOR U20659 ( .A(n19878), .B(n19879), .Z(n18852) );
  XOR U20660 ( .A(n18755), .B(n17983), .Z(n19879) );
  XOR U20661 ( .A(n19880), .B(n19881), .Z(n17983) );
  ANDN U20662 ( .B(n19882), .A(n19883), .Z(n19880) );
  XNOR U20663 ( .A(n19884), .B(n19885), .Z(n18755) );
  ANDN U20664 ( .B(n19886), .A(n19887), .Z(n19884) );
  XOR U20665 ( .A(n18348), .B(n19888), .Z(n19878) );
  XOR U20666 ( .A(n17025), .B(n18713), .Z(n19888) );
  XNOR U20667 ( .A(n19889), .B(n19890), .Z(n18713) );
  AND U20668 ( .A(n19891), .B(n19892), .Z(n19889) );
  XOR U20669 ( .A(n19893), .B(n19894), .Z(n17025) );
  ANDN U20670 ( .B(n19895), .A(n19896), .Z(n19893) );
  XNOR U20671 ( .A(n19897), .B(n19898), .Z(n18348) );
  ANDN U20672 ( .B(n19899), .A(n19900), .Z(n19897) );
  XNOR U20673 ( .A(n19901), .B(n16331), .Z(n16976) );
  XNOR U20674 ( .A(n19902), .B(n19903), .Z(n18393) );
  XOR U20675 ( .A(n17455), .B(n19071), .Z(n19903) );
  XNOR U20676 ( .A(n19904), .B(n19905), .Z(n19071) );
  NOR U20677 ( .A(n19906), .B(n19907), .Z(n19904) );
  XNOR U20678 ( .A(n19908), .B(n19909), .Z(n17455) );
  XOR U20679 ( .A(n19912), .B(n19913), .Z(n19902) );
  XOR U20680 ( .A(n16403), .B(n19914), .Z(n19913) );
  XNOR U20681 ( .A(n19915), .B(n19916), .Z(n16403) );
  AND U20682 ( .A(n19917), .B(n19918), .Z(n19915) );
  XNOR U20683 ( .A(n19919), .B(n19920), .Z(n19557) );
  XOR U20684 ( .A(n19837), .B(n19737), .Z(n19920) );
  XOR U20685 ( .A(n19921), .B(n19922), .Z(n19737) );
  ANDN U20686 ( .B(n19923), .A(n19924), .Z(n19921) );
  XNOR U20687 ( .A(n19925), .B(n19926), .Z(n19837) );
  ANDN U20688 ( .B(n19927), .A(n19928), .Z(n19925) );
  XOR U20689 ( .A(n17283), .B(n19929), .Z(n19919) );
  XOR U20690 ( .A(n16736), .B(n19364), .Z(n19929) );
  XNOR U20691 ( .A(n19930), .B(n19931), .Z(n19364) );
  XNOR U20692 ( .A(n19934), .B(n19935), .Z(n16736) );
  AND U20693 ( .A(n19936), .B(n19937), .Z(n19934) );
  XNOR U20694 ( .A(n19938), .B(n19939), .Z(n17283) );
  ANDN U20695 ( .B(n19940), .A(n19941), .Z(n19938) );
  XOR U20696 ( .A(n12231), .B(n19942), .Z(n19847) );
  XOR U20697 ( .A(n13042), .B(n11954), .Z(n19942) );
  XNOR U20698 ( .A(n19943), .B(n14597), .Z(n11954) );
  XNOR U20699 ( .A(n19944), .B(n17980), .Z(n14597) );
  XNOR U20700 ( .A(n19945), .B(n14608), .Z(n13042) );
  IV U20701 ( .A(n14015), .Z(n14608) );
  XOR U20702 ( .A(n19946), .B(n17024), .Z(n14015) );
  XNOR U20703 ( .A(n19947), .B(n19948), .Z(n17024) );
  ANDN U20704 ( .B(n16973), .A(n14607), .Z(n19945) );
  XOR U20705 ( .A(n19949), .B(n15948), .Z(n14607) );
  XNOR U20706 ( .A(n19950), .B(n17626), .Z(n16973) );
  XOR U20707 ( .A(n19951), .B(n14005), .Z(n12231) );
  XOR U20708 ( .A(n18596), .B(n19952), .Z(n14005) );
  ANDN U20709 ( .B(n14611), .A(n17388), .Z(n19951) );
  IV U20710 ( .A(n16982), .Z(n17388) );
  XOR U20711 ( .A(n19953), .B(n17229), .Z(n16982) );
  XOR U20712 ( .A(n19954), .B(n15904), .Z(n14611) );
  IV U20713 ( .A(n16522), .Z(n15904) );
  XOR U20714 ( .A(n19955), .B(n19956), .Z(n16522) );
  XOR U20715 ( .A(n19957), .B(n14598), .Z(n16978) );
  XOR U20716 ( .A(n19958), .B(n18465), .Z(n14598) );
  IV U20717 ( .A(n18433), .Z(n18465) );
  XOR U20718 ( .A(n19959), .B(n19960), .Z(n18433) );
  ANDN U20719 ( .B(n17405), .A(n17404), .Z(n19957) );
  XNOR U20720 ( .A(n19961), .B(n17630), .Z(n17404) );
  XNOR U20721 ( .A(n17195), .B(n19962), .Z(n17405) );
  XOR U20722 ( .A(n19203), .B(n12713), .Z(n9272) );
  XOR U20723 ( .A(n11372), .B(n12909), .Z(n12713) );
  XOR U20724 ( .A(n19963), .B(n19964), .Z(n12909) );
  XNOR U20725 ( .A(n12330), .B(n10848), .Z(n19964) );
  XNOR U20726 ( .A(n19965), .B(n18085), .Z(n10848) );
  XOR U20727 ( .A(n19966), .B(n18772), .Z(n18085) );
  IV U20728 ( .A(n17249), .Z(n18772) );
  XOR U20729 ( .A(n19967), .B(n19839), .Z(n17249) );
  XOR U20730 ( .A(n19968), .B(n19969), .Z(n19839) );
  XOR U20731 ( .A(n19970), .B(n19100), .Z(n19969) );
  XOR U20732 ( .A(n19971), .B(n19972), .Z(n19100) );
  ANDN U20733 ( .B(n19932), .A(n19973), .Z(n19971) );
  XNOR U20734 ( .A(n16107), .B(n19974), .Z(n19968) );
  XNOR U20735 ( .A(n19680), .B(n17929), .Z(n19974) );
  XNOR U20736 ( .A(n19975), .B(n19976), .Z(n17929) );
  XNOR U20737 ( .A(n19977), .B(n19978), .Z(n19680) );
  ANDN U20738 ( .B(n19935), .A(n19937), .Z(n19977) );
  XNOR U20739 ( .A(n19979), .B(n19980), .Z(n16107) );
  ANDN U20740 ( .B(n19924), .A(n19922), .Z(n19979) );
  ANDN U20741 ( .B(n18739), .A(n18113), .Z(n19965) );
  IV U20742 ( .A(n19186), .Z(n18113) );
  XOR U20743 ( .A(n16961), .B(n19981), .Z(n19186) );
  IV U20744 ( .A(n17335), .Z(n16961) );
  XOR U20745 ( .A(n19982), .B(n19983), .Z(n17335) );
  XOR U20746 ( .A(n15694), .B(n19984), .Z(n18739) );
  XNOR U20747 ( .A(n19985), .B(n17157), .Z(n12330) );
  XOR U20748 ( .A(n19986), .B(n19987), .Z(n17157) );
  ANDN U20749 ( .B(n18731), .A(n18117), .Z(n19985) );
  XOR U20750 ( .A(n18283), .B(n19988), .Z(n18117) );
  XOR U20751 ( .A(n19989), .B(n19990), .Z(n18926) );
  XOR U20752 ( .A(n17868), .B(n18174), .Z(n19990) );
  XOR U20753 ( .A(n19991), .B(n19992), .Z(n18174) );
  ANDN U20754 ( .B(n19866), .A(n19993), .Z(n19991) );
  XNOR U20755 ( .A(n19994), .B(n19995), .Z(n17868) );
  ANDN U20756 ( .B(n19996), .A(n19856), .Z(n19994) );
  XOR U20757 ( .A(n18076), .B(n19997), .Z(n19989) );
  XOR U20758 ( .A(n19998), .B(n15303), .Z(n19997) );
  XNOR U20759 ( .A(n19999), .B(n20000), .Z(n15303) );
  XNOR U20760 ( .A(n20002), .B(n20003), .Z(n18076) );
  ANDN U20761 ( .B(n20004), .A(n20005), .Z(n20002) );
  XNOR U20762 ( .A(n20007), .B(n18282), .Z(n18731) );
  IV U20763 ( .A(n20008), .Z(n18282) );
  XOR U20764 ( .A(n13475), .B(n20009), .Z(n19963) );
  XOR U20765 ( .A(n9507), .B(n18695), .Z(n20009) );
  XNOR U20766 ( .A(n20010), .B(n18735), .Z(n18695) );
  IV U20767 ( .A(n17153), .Z(n18735) );
  XOR U20768 ( .A(n19748), .B(n20011), .Z(n17153) );
  IV U20769 ( .A(n17399), .Z(n19748) );
  XOR U20770 ( .A(n20012), .B(n20013), .Z(n17399) );
  ANDN U20771 ( .B(n18736), .A(n18115), .Z(n20010) );
  XOR U20772 ( .A(n20014), .B(n17958), .Z(n18115) );
  XOR U20773 ( .A(n20015), .B(n15201), .Z(n18736) );
  XNOR U20774 ( .A(n20016), .B(n20017), .Z(n15201) );
  XOR U20775 ( .A(n20018), .B(n17162), .Z(n9507) );
  XOR U20776 ( .A(n20019), .B(n18275), .Z(n17162) );
  ANDN U20777 ( .B(n18108), .A(n18742), .Z(n20018) );
  XOR U20778 ( .A(n19307), .B(n20020), .Z(n18742) );
  XOR U20779 ( .A(n19622), .B(n19841), .Z(n18108) );
  XNOR U20780 ( .A(n20021), .B(n20022), .Z(n19622) );
  XNOR U20781 ( .A(n20025), .B(n17167), .Z(n13475) );
  XNOR U20782 ( .A(n20026), .B(n19451), .Z(n17167) );
  NOR U20783 ( .A(n18110), .B(n18728), .Z(n20025) );
  XNOR U20784 ( .A(n20027), .B(n16613), .Z(n18728) );
  IV U20785 ( .A(n19182), .Z(n18110) );
  XOR U20786 ( .A(n19685), .B(n19659), .Z(n19182) );
  XOR U20787 ( .A(n20028), .B(n20029), .Z(n19685) );
  ANDN U20788 ( .B(n19584), .A(n19585), .Z(n20028) );
  XOR U20789 ( .A(n20030), .B(n20031), .Z(n11372) );
  XNOR U20790 ( .A(n11416), .B(n12251), .Z(n20031) );
  XNOR U20791 ( .A(n20032), .B(n12487), .Z(n12251) );
  XOR U20792 ( .A(n20033), .B(n17961), .Z(n12487) );
  ANDN U20793 ( .B(n12488), .A(n18981), .Z(n20032) );
  XOR U20794 ( .A(n20034), .B(n20008), .Z(n18981) );
  XOR U20795 ( .A(n20035), .B(n16112), .Z(n12488) );
  XOR U20796 ( .A(n20036), .B(n17169), .Z(n11416) );
  XNOR U20797 ( .A(n20037), .B(n18789), .Z(n17169) );
  XOR U20798 ( .A(n20038), .B(n20039), .Z(n14353) );
  XOR U20799 ( .A(n20040), .B(n18777), .Z(n17170) );
  XOR U20800 ( .A(n12132), .B(n20041), .Z(n20030) );
  XNOR U20801 ( .A(n11747), .B(n9941), .Z(n20041) );
  XOR U20802 ( .A(n20042), .B(n12483), .Z(n9941) );
  XOR U20803 ( .A(n20043), .B(n18938), .Z(n12483) );
  XOR U20804 ( .A(n20044), .B(n20045), .Z(n18938) );
  ANDN U20805 ( .B(n12484), .A(n14350), .Z(n20042) );
  IV U20806 ( .A(n20046), .Z(n14350) );
  XOR U20807 ( .A(n20047), .B(n12473), .Z(n11747) );
  XOR U20808 ( .A(n20048), .B(n18896), .Z(n12473) );
  XOR U20809 ( .A(n20049), .B(n19701), .Z(n18896) );
  XNOR U20810 ( .A(n20050), .B(n20051), .Z(n19701) );
  XNOR U20811 ( .A(n18149), .B(n20052), .Z(n20051) );
  XOR U20812 ( .A(n20053), .B(n20054), .Z(n18149) );
  NOR U20813 ( .A(n20055), .B(n20056), .Z(n20053) );
  XOR U20814 ( .A(n20057), .B(n20058), .Z(n20050) );
  XOR U20815 ( .A(n18565), .B(n16747), .Z(n20058) );
  XNOR U20816 ( .A(n20059), .B(n20060), .Z(n16747) );
  ANDN U20817 ( .B(n20061), .A(n20062), .Z(n20059) );
  XNOR U20818 ( .A(n20063), .B(n20064), .Z(n18565) );
  NOR U20819 ( .A(n20065), .B(n20066), .Z(n20063) );
  ANDN U20820 ( .B(n12474), .A(n19209), .Z(n20047) );
  XOR U20821 ( .A(n20067), .B(n17552), .Z(n19209) );
  XOR U20822 ( .A(n19690), .B(n19659), .Z(n12474) );
  IV U20823 ( .A(n19551), .Z(n19659) );
  XNOR U20824 ( .A(n20068), .B(n20069), .Z(n19690) );
  ANDN U20825 ( .B(n19582), .A(n19580), .Z(n20068) );
  IV U20826 ( .A(n20070), .Z(n19582) );
  XOR U20827 ( .A(n20071), .B(n12478), .Z(n12132) );
  XNOR U20828 ( .A(n18161), .B(n20072), .Z(n12478) );
  ANDN U20829 ( .B(n12477), .A(n14360), .Z(n20071) );
  XOR U20830 ( .A(n20073), .B(n20074), .Z(n14360) );
  IV U20831 ( .A(n19197), .Z(n12477) );
  XOR U20832 ( .A(n20075), .B(n17229), .Z(n19197) );
  XOR U20833 ( .A(n20076), .B(n20077), .Z(n17229) );
  XOR U20834 ( .A(n20078), .B(n12484), .Z(n19203) );
  XOR U20835 ( .A(n17483), .B(n20079), .Z(n12484) );
  ANDN U20836 ( .B(n14351), .A(n20046), .Z(n20078) );
  XOR U20837 ( .A(n20080), .B(n17958), .Z(n20046) );
  XOR U20838 ( .A(n20081), .B(n17646), .Z(n14351) );
  XOR U20839 ( .A(n20082), .B(n9337), .Z(n4907) );
  IV U20840 ( .A(n6690), .Z(n9337) );
  XOR U20841 ( .A(n9765), .B(n16002), .Z(n6690) );
  XNOR U20842 ( .A(n20083), .B(n13781), .Z(n16002) );
  ANDN U20843 ( .B(n14572), .A(n14573), .Z(n20083) );
  XOR U20844 ( .A(n20084), .B(n19649), .Z(n14573) );
  XOR U20845 ( .A(n20085), .B(n20086), .Z(n19649) );
  XNOR U20846 ( .A(n12136), .B(n18510), .Z(n9765) );
  XOR U20847 ( .A(n20087), .B(n20088), .Z(n18510) );
  XOR U20848 ( .A(n13271), .B(n11348), .Z(n20088) );
  XOR U20849 ( .A(n20089), .B(n16155), .Z(n11348) );
  XOR U20850 ( .A(n16753), .B(n20090), .Z(n16155) );
  NOR U20851 ( .A(n16017), .B(n14563), .Z(n20089) );
  XOR U20852 ( .A(n20091), .B(n16112), .Z(n14563) );
  XOR U20853 ( .A(n16603), .B(n20092), .Z(n16017) );
  IV U20854 ( .A(n18321), .Z(n16603) );
  XNOR U20855 ( .A(n20093), .B(n16145), .Z(n13271) );
  XOR U20856 ( .A(n20094), .B(n15193), .Z(n16145) );
  ANDN U20857 ( .B(n14559), .A(n16019), .Z(n20093) );
  XOR U20858 ( .A(n20095), .B(n18508), .Z(n16019) );
  XNOR U20859 ( .A(n20096), .B(n17333), .Z(n14559) );
  XNOR U20860 ( .A(n20098), .B(n20099), .Z(n19015) );
  XOR U20861 ( .A(n18974), .B(n19187), .Z(n20099) );
  XNOR U20862 ( .A(n20100), .B(n20101), .Z(n19187) );
  NOR U20863 ( .A(n20102), .B(n20103), .Z(n20100) );
  XNOR U20864 ( .A(n20104), .B(n20105), .Z(n18974) );
  ANDN U20865 ( .B(n20106), .A(n20107), .Z(n20104) );
  XOR U20866 ( .A(n17014), .B(n20108), .Z(n20098) );
  XNOR U20867 ( .A(n17913), .B(n19255), .Z(n20108) );
  XNOR U20868 ( .A(n20109), .B(n20110), .Z(n19255) );
  ANDN U20869 ( .B(n20111), .A(n20112), .Z(n20109) );
  XOR U20870 ( .A(n20113), .B(n20114), .Z(n17913) );
  AND U20871 ( .A(n20115), .B(n20116), .Z(n20113) );
  XNOR U20872 ( .A(n20117), .B(n20118), .Z(n17014) );
  ANDN U20873 ( .B(n20119), .A(n20120), .Z(n20117) );
  XNOR U20874 ( .A(n9923), .B(n20121), .Z(n20087) );
  XNOR U20875 ( .A(n9100), .B(n17670), .Z(n20121) );
  XNOR U20876 ( .A(n20122), .B(n16142), .Z(n17670) );
  XOR U20877 ( .A(n19998), .B(n15304), .Z(n16142) );
  XOR U20878 ( .A(n20123), .B(n20124), .Z(n15304) );
  XOR U20879 ( .A(n20125), .B(n20126), .Z(n19998) );
  ANDN U20880 ( .B(n20127), .A(n19870), .Z(n20125) );
  ANDN U20881 ( .B(n17694), .A(n14555), .Z(n20122) );
  XNOR U20882 ( .A(n20128), .B(n16516), .Z(n14555) );
  XOR U20883 ( .A(n20129), .B(n20130), .Z(n17694) );
  XNOR U20884 ( .A(n20131), .B(n16151), .Z(n9100) );
  XOR U20885 ( .A(n20132), .B(n15899), .Z(n16151) );
  XNOR U20886 ( .A(n20133), .B(n20134), .Z(n15899) );
  ANDN U20887 ( .B(n16013), .A(n14550), .Z(n20131) );
  XOR U20888 ( .A(n17746), .B(n20135), .Z(n14550) );
  XOR U20889 ( .A(n20136), .B(n17440), .Z(n16013) );
  XNOR U20890 ( .A(n20137), .B(n16158), .Z(n9923) );
  XOR U20891 ( .A(n18045), .B(n20138), .Z(n16158) );
  AND U20892 ( .A(n16366), .B(n14546), .Z(n20137) );
  XOR U20893 ( .A(n20139), .B(n18309), .Z(n14546) );
  IV U20894 ( .A(n19369), .Z(n18309) );
  XOR U20895 ( .A(n20140), .B(n20141), .Z(n19369) );
  XOR U20896 ( .A(n20142), .B(n20143), .Z(n16366) );
  XOR U20897 ( .A(n20144), .B(n20145), .Z(n12136) );
  XOR U20898 ( .A(n12172), .B(n13159), .Z(n20145) );
  XOR U20899 ( .A(n20146), .B(n13777), .Z(n13159) );
  XOR U20900 ( .A(n18053), .B(n20147), .Z(n13777) );
  XOR U20901 ( .A(n20148), .B(n18186), .Z(n13776) );
  XOR U20902 ( .A(n20149), .B(n18508), .Z(n14577) );
  XOR U20903 ( .A(n20150), .B(n13780), .Z(n12172) );
  XOR U20904 ( .A(n19307), .B(n20151), .Z(n13780) );
  XOR U20905 ( .A(n20152), .B(n20153), .Z(n19307) );
  ANDN U20906 ( .B(n13781), .A(n14572), .Z(n20150) );
  XOR U20907 ( .A(n20154), .B(n20155), .Z(n14572) );
  XOR U20908 ( .A(n20156), .B(n18260), .Z(n13781) );
  IV U20909 ( .A(n17795), .Z(n18260) );
  XNOR U20910 ( .A(n20157), .B(n20158), .Z(n20097) );
  XNOR U20911 ( .A(n16816), .B(n17277), .Z(n20158) );
  XNOR U20912 ( .A(n20159), .B(n19883), .Z(n17277) );
  ANDN U20913 ( .B(n20160), .A(n20161), .Z(n20159) );
  XNOR U20914 ( .A(n20162), .B(n19891), .Z(n16816) );
  ANDN U20915 ( .B(n20163), .A(n20164), .Z(n20162) );
  XNOR U20916 ( .A(n17736), .B(n20165), .Z(n20157) );
  XNOR U20917 ( .A(n20166), .B(n20167), .Z(n20165) );
  XOR U20918 ( .A(n20168), .B(n19900), .Z(n17736) );
  ANDN U20919 ( .B(n20169), .A(n20170), .Z(n20168) );
  XNOR U20920 ( .A(n20171), .B(n20172), .Z(n18343) );
  XNOR U20921 ( .A(n17648), .B(n19126), .Z(n20172) );
  XOR U20922 ( .A(n20173), .B(n19730), .Z(n19126) );
  ANDN U20923 ( .B(n20174), .A(n20175), .Z(n20173) );
  XNOR U20924 ( .A(n20176), .B(n18912), .Z(n17648) );
  NOR U20925 ( .A(n20177), .B(n20178), .Z(n20176) );
  XOR U20926 ( .A(n17523), .B(n20179), .Z(n20171) );
  XOR U20927 ( .A(n19283), .B(n20180), .Z(n20179) );
  XNOR U20928 ( .A(n20181), .B(n18847), .Z(n19283) );
  IV U20929 ( .A(n20182), .Z(n18847) );
  ANDN U20930 ( .B(n20183), .A(n20184), .Z(n20181) );
  XNOR U20931 ( .A(n20185), .B(n20186), .Z(n17523) );
  NOR U20932 ( .A(n20187), .B(n20188), .Z(n20185) );
  XOR U20933 ( .A(n11489), .B(n20189), .Z(n20144) );
  XNOR U20934 ( .A(n10330), .B(n12889), .Z(n20189) );
  XNOR U20935 ( .A(n20190), .B(n13771), .Z(n12889) );
  XNOR U20936 ( .A(n20191), .B(n18804), .Z(n13771) );
  XNOR U20937 ( .A(n20192), .B(n20193), .Z(n18804) );
  ANDN U20938 ( .B(n13772), .A(n16021), .Z(n20190) );
  XNOR U20939 ( .A(n20194), .B(n17294), .Z(n16021) );
  XNOR U20940 ( .A(n20195), .B(n17572), .Z(n13772) );
  IV U20941 ( .A(n18789), .Z(n17572) );
  XOR U20942 ( .A(n20196), .B(n13785), .Z(n10330) );
  XNOR U20943 ( .A(n20197), .B(n17586), .Z(n13785) );
  XOR U20944 ( .A(n20198), .B(n18607), .Z(n17586) );
  XNOR U20945 ( .A(n20199), .B(n20200), .Z(n18607) );
  XNOR U20946 ( .A(n19514), .B(n18451), .Z(n20200) );
  XNOR U20947 ( .A(n20201), .B(n20202), .Z(n18451) );
  NOR U20948 ( .A(n20203), .B(n20204), .Z(n20201) );
  XOR U20949 ( .A(n20205), .B(n20206), .Z(n19514) );
  NOR U20950 ( .A(n20207), .B(n20208), .Z(n20205) );
  XOR U20951 ( .A(n18312), .B(n20209), .Z(n20199) );
  XNOR U20952 ( .A(n16871), .B(n17796), .Z(n20209) );
  XNOR U20953 ( .A(n20210), .B(n20211), .Z(n17796) );
  XNOR U20954 ( .A(n20214), .B(n20215), .Z(n16871) );
  NOR U20955 ( .A(n20216), .B(n20217), .Z(n20214) );
  XNOR U20956 ( .A(n20218), .B(n20219), .Z(n18312) );
  ANDN U20957 ( .B(n20220), .A(n20221), .Z(n20218) );
  NOR U20958 ( .A(n14569), .B(n13784), .Z(n20196) );
  XOR U20959 ( .A(n15958), .B(n20222), .Z(n13784) );
  IV U20960 ( .A(n17659), .Z(n15958) );
  IV U20961 ( .A(n15998), .Z(n14569) );
  XOR U20962 ( .A(n20223), .B(n16516), .Z(n15998) );
  XNOR U20963 ( .A(n20224), .B(n13767), .Z(n11489) );
  XOR U20964 ( .A(n20225), .B(n18561), .Z(n13767) );
  IV U20965 ( .A(n15252), .Z(n18561) );
  XNOR U20966 ( .A(n19947), .B(n20226), .Z(n15252) );
  XOR U20967 ( .A(n20227), .B(n20228), .Z(n19947) );
  XNOR U20968 ( .A(n19452), .B(n18574), .Z(n20228) );
  XNOR U20969 ( .A(n20229), .B(n20230), .Z(n18574) );
  ANDN U20970 ( .B(n20231), .A(n20232), .Z(n20229) );
  XNOR U20971 ( .A(n20233), .B(n20234), .Z(n19452) );
  ANDN U20972 ( .B(n20235), .A(n20236), .Z(n20233) );
  XNOR U20973 ( .A(n20237), .B(n20238), .Z(n20227) );
  XOR U20974 ( .A(n17862), .B(n17185), .Z(n20238) );
  XNOR U20975 ( .A(n20239), .B(n20240), .Z(n17185) );
  ANDN U20976 ( .B(n20241), .A(n20242), .Z(n20239) );
  XNOR U20977 ( .A(n20243), .B(n20244), .Z(n17862) );
  ANDN U20978 ( .B(n20245), .A(n20246), .Z(n20243) );
  AND U20979 ( .A(n14580), .B(n13768), .Z(n20224) );
  XOR U20980 ( .A(n16523), .B(n20247), .Z(n13768) );
  IV U20981 ( .A(n17746), .Z(n16523) );
  XNOR U20982 ( .A(n20248), .B(n20249), .Z(n17746) );
  XOR U20983 ( .A(n20250), .B(n18400), .Z(n14580) );
  XNOR U20984 ( .A(n20251), .B(n20252), .Z(n18400) );
  NOR U20985 ( .A(n9268), .B(n7125), .Z(n20082) );
  XNOR U20986 ( .A(n16347), .B(n11437), .Z(n7125) );
  IV U20987 ( .A(n11210), .Z(n11437) );
  XOR U20988 ( .A(n11963), .B(n16862), .Z(n11210) );
  XNOR U20989 ( .A(n20253), .B(n20254), .Z(n16862) );
  XOR U20990 ( .A(n11559), .B(n10336), .Z(n20254) );
  XNOR U20991 ( .A(n20255), .B(n17349), .Z(n10336) );
  XOR U20992 ( .A(n20256), .B(n17944), .Z(n17349) );
  ANDN U20993 ( .B(n16349), .A(n12039), .Z(n20255) );
  XOR U20994 ( .A(n20257), .B(n18822), .Z(n12039) );
  IV U20995 ( .A(n16767), .Z(n18822) );
  XNOR U20996 ( .A(n20258), .B(n19116), .Z(n16767) );
  XNOR U20997 ( .A(n20259), .B(n20260), .Z(n19116) );
  XOR U20998 ( .A(n16953), .B(n17857), .Z(n20260) );
  XNOR U20999 ( .A(n20261), .B(n20262), .Z(n17857) );
  ANDN U21000 ( .B(n20263), .A(n20264), .Z(n20261) );
  XNOR U21001 ( .A(n20265), .B(n20266), .Z(n16953) );
  ANDN U21002 ( .B(n20267), .A(n20268), .Z(n20265) );
  XOR U21003 ( .A(n20269), .B(n20270), .Z(n20259) );
  XOR U21004 ( .A(n17668), .B(n20271), .Z(n20270) );
  XOR U21005 ( .A(n20272), .B(n20273), .Z(n17668) );
  ANDN U21006 ( .B(n20274), .A(n20275), .Z(n20272) );
  XNOR U21007 ( .A(n20276), .B(n17009), .Z(n16349) );
  XOR U21008 ( .A(n20278), .B(n20279), .Z(n19653) );
  XOR U21009 ( .A(n17947), .B(n18373), .Z(n20279) );
  XOR U21010 ( .A(n20280), .B(n19539), .Z(n18373) );
  ANDN U21011 ( .B(n19538), .A(n20281), .Z(n20280) );
  XNOR U21012 ( .A(n20282), .B(n19529), .Z(n17947) );
  NOR U21013 ( .A(n19785), .B(n19528), .Z(n20282) );
  XNOR U21014 ( .A(n17428), .B(n20283), .Z(n20278) );
  XNOR U21015 ( .A(n19046), .B(n18488), .Z(n20283) );
  XOR U21016 ( .A(n20284), .B(n19535), .Z(n18488) );
  ANDN U21017 ( .B(n19534), .A(n20285), .Z(n20284) );
  XNOR U21018 ( .A(n20286), .B(n20287), .Z(n19046) );
  AND U21019 ( .A(n20288), .B(n20289), .Z(n20286) );
  XNOR U21020 ( .A(n20290), .B(n20291), .Z(n17428) );
  NOR U21021 ( .A(n20292), .B(n20293), .Z(n20290) );
  XOR U21022 ( .A(n20294), .B(n17353), .Z(n11559) );
  XOR U21023 ( .A(n20295), .B(n16119), .Z(n17353) );
  IV U21024 ( .A(n18857), .Z(n16119) );
  XOR U21025 ( .A(n20296), .B(n20297), .Z(n18857) );
  ANDN U21026 ( .B(n12030), .A(n16351), .Z(n20294) );
  XOR U21027 ( .A(n20298), .B(n16868), .Z(n16351) );
  XNOR U21028 ( .A(n20299), .B(n17874), .Z(n12030) );
  XNOR U21029 ( .A(n12297), .B(n20300), .Z(n20253) );
  XNOR U21030 ( .A(n16159), .B(n9660), .Z(n20300) );
  XNOR U21031 ( .A(n20301), .B(n17346), .Z(n9660) );
  XOR U21032 ( .A(n20302), .B(n20303), .Z(n17346) );
  AND U21033 ( .A(n17345), .B(n12026), .Z(n20301) );
  XNOR U21034 ( .A(n20304), .B(n18072), .Z(n16159) );
  ANDN U21035 ( .B(n16341), .A(n12043), .Z(n20304) );
  IV U21036 ( .A(n16342), .Z(n12043) );
  XOR U21037 ( .A(n20306), .B(n15528), .Z(n16342) );
  IV U21038 ( .A(n17045), .Z(n15528) );
  XNOR U21039 ( .A(n19421), .B(n20307), .Z(n17045) );
  XOR U21040 ( .A(n20308), .B(n20309), .Z(n19421) );
  XOR U21041 ( .A(n20038), .B(n20310), .Z(n20309) );
  XNOR U21042 ( .A(n20311), .B(n20312), .Z(n20038) );
  XOR U21043 ( .A(n20314), .B(n20315), .Z(n20308) );
  XNOR U21044 ( .A(n18833), .B(n20316), .Z(n20315) );
  XOR U21045 ( .A(n20317), .B(n20318), .Z(n18833) );
  ANDN U21046 ( .B(n20319), .A(n19344), .Z(n20317) );
  XOR U21047 ( .A(n20320), .B(n18789), .Z(n16341) );
  XOR U21048 ( .A(n19220), .B(n19776), .Z(n18789) );
  XNOR U21049 ( .A(n20321), .B(n20322), .Z(n19776) );
  XNOR U21050 ( .A(n20323), .B(n18591), .Z(n20322) );
  ANDN U21051 ( .B(n20326), .A(n20327), .Z(n20324) );
  XNOR U21052 ( .A(n20328), .B(n20329), .Z(n20321) );
  XNOR U21053 ( .A(n17515), .B(n18181), .Z(n20329) );
  XNOR U21054 ( .A(n20330), .B(n20331), .Z(n18181) );
  ANDN U21055 ( .B(n20332), .A(n20333), .Z(n20330) );
  XOR U21056 ( .A(n20334), .B(n20335), .Z(n17515) );
  AND U21057 ( .A(n20336), .B(n20337), .Z(n20334) );
  XOR U21058 ( .A(n20338), .B(n20339), .Z(n19220) );
  XOR U21059 ( .A(n18324), .B(n17565), .Z(n20339) );
  XOR U21060 ( .A(n20340), .B(n20341), .Z(n17565) );
  ANDN U21061 ( .B(n20342), .A(n20343), .Z(n20340) );
  XNOR U21062 ( .A(n20344), .B(n20345), .Z(n18324) );
  ANDN U21063 ( .B(n20346), .A(n20347), .Z(n20344) );
  XOR U21064 ( .A(n18514), .B(n20348), .Z(n20338) );
  XNOR U21065 ( .A(n20349), .B(n16812), .Z(n20348) );
  XNOR U21066 ( .A(n20350), .B(n20351), .Z(n16812) );
  ANDN U21067 ( .B(n20352), .A(n20353), .Z(n20350) );
  XNOR U21068 ( .A(n20354), .B(n20355), .Z(n18514) );
  ANDN U21069 ( .B(n20356), .A(n20357), .Z(n20354) );
  XNOR U21070 ( .A(n20358), .B(n17351), .Z(n12297) );
  XOR U21071 ( .A(n18378), .B(n20359), .Z(n17351) );
  IV U21072 ( .A(n17284), .Z(n18378) );
  XNOR U21073 ( .A(n18756), .B(n20360), .Z(n17284) );
  XOR U21074 ( .A(n20361), .B(n20362), .Z(n18756) );
  XNOR U21075 ( .A(n20363), .B(n18325), .Z(n20362) );
  XNOR U21076 ( .A(n20364), .B(n20365), .Z(n18325) );
  NOR U21077 ( .A(n19899), .B(n19898), .Z(n20364) );
  XOR U21078 ( .A(n16464), .B(n20366), .Z(n20361) );
  XNOR U21079 ( .A(n19635), .B(n20367), .Z(n20366) );
  XNOR U21080 ( .A(n20368), .B(n20369), .Z(n19635) );
  NOR U21081 ( .A(n19892), .B(n19890), .Z(n20370) );
  ANDN U21082 ( .B(n12035), .A(n16344), .Z(n20358) );
  XOR U21083 ( .A(n20371), .B(n15688), .Z(n16344) );
  IV U21084 ( .A(n16585), .Z(n15688) );
  XOR U21085 ( .A(n20372), .B(n16739), .Z(n12035) );
  XOR U21086 ( .A(n20373), .B(n20374), .Z(n16739) );
  XOR U21087 ( .A(n20375), .B(n20376), .Z(n11963) );
  XOR U21088 ( .A(n10194), .B(n11246), .Z(n20376) );
  XOR U21089 ( .A(n20377), .B(n19065), .Z(n11246) );
  XNOR U21090 ( .A(n20378), .B(n17944), .Z(n19065) );
  IV U21091 ( .A(n18154), .Z(n17944) );
  ANDN U21092 ( .B(n13615), .A(n12872), .Z(n20377) );
  XNOR U21093 ( .A(n20381), .B(n14958), .Z(n12872) );
  IV U21094 ( .A(n15336), .Z(n14958) );
  XNOR U21095 ( .A(n20382), .B(n20383), .Z(n15336) );
  XNOR U21096 ( .A(n20384), .B(n18942), .Z(n13615) );
  IV U21097 ( .A(n17020), .Z(n18942) );
  XOR U21098 ( .A(n20385), .B(n20386), .Z(n17020) );
  XNOR U21099 ( .A(n20387), .B(n16173), .Z(n10194) );
  IV U21100 ( .A(n19059), .Z(n16173) );
  XNOR U21101 ( .A(n20388), .B(n17861), .Z(n19059) );
  ANDN U21102 ( .B(n13390), .A(n13618), .Z(n20387) );
  XNOR U21103 ( .A(n20389), .B(n17970), .Z(n13618) );
  XOR U21104 ( .A(n17321), .B(n20390), .Z(n13390) );
  XOR U21105 ( .A(n20391), .B(n20124), .Z(n17321) );
  XNOR U21106 ( .A(n20392), .B(n20393), .Z(n20124) );
  XNOR U21107 ( .A(n19463), .B(n15251), .Z(n20393) );
  XOR U21108 ( .A(n20394), .B(n19867), .Z(n15251) );
  ANDN U21109 ( .B(n19993), .A(n19992), .Z(n20394) );
  XOR U21110 ( .A(n20395), .B(n20396), .Z(n19463) );
  NOR U21111 ( .A(n19995), .B(n19996), .Z(n20395) );
  XOR U21112 ( .A(n20225), .B(n20397), .Z(n20392) );
  XOR U21113 ( .A(n18560), .B(n18959), .Z(n20397) );
  XNOR U21114 ( .A(n20398), .B(n19861), .Z(n18959) );
  NOR U21115 ( .A(n20000), .B(n20001), .Z(n20398) );
  XOR U21116 ( .A(n20399), .B(n19872), .Z(n18560) );
  ANDN U21117 ( .B(n20126), .A(n20127), .Z(n20399) );
  XNOR U21118 ( .A(n20400), .B(n20401), .Z(n20225) );
  ANDN U21119 ( .B(n20003), .A(n20004), .Z(n20400) );
  XOR U21120 ( .A(n11863), .B(n20402), .Z(n20375) );
  XOR U21121 ( .A(n11057), .B(n11204), .Z(n20402) );
  XNOR U21122 ( .A(n20403), .B(n16167), .Z(n11204) );
  XNOR U21123 ( .A(n20404), .B(n18806), .Z(n16167) );
  ANDN U21124 ( .B(n12567), .A(n13622), .Z(n20403) );
  XNOR U21125 ( .A(n20405), .B(n15265), .Z(n13622) );
  XNOR U21126 ( .A(n20406), .B(n20407), .Z(n19746) );
  XNOR U21127 ( .A(n18604), .B(n20408), .Z(n20407) );
  XOR U21128 ( .A(n20409), .B(n20410), .Z(n18604) );
  NOR U21129 ( .A(n19160), .B(n19161), .Z(n20409) );
  XOR U21130 ( .A(n18682), .B(n20411), .Z(n20406) );
  XNOR U21131 ( .A(n19370), .B(n18467), .Z(n20411) );
  XNOR U21132 ( .A(n20412), .B(n20413), .Z(n18467) );
  ANDN U21133 ( .B(n19166), .A(n19164), .Z(n20412) );
  NOR U21134 ( .A(n20416), .B(n19155), .Z(n20414) );
  XOR U21135 ( .A(n20417), .B(n20418), .Z(n18682) );
  XOR U21136 ( .A(n20419), .B(n20420), .Z(n19823) );
  XOR U21137 ( .A(n17968), .B(n16062), .Z(n20420) );
  XNOR U21138 ( .A(n20421), .B(n20422), .Z(n16062) );
  ANDN U21139 ( .B(n20423), .A(n20424), .Z(n20421) );
  XOR U21140 ( .A(n20425), .B(n20426), .Z(n17968) );
  ANDN U21141 ( .B(n20427), .A(n20428), .Z(n20425) );
  XOR U21142 ( .A(n20372), .B(n20429), .Z(n20419) );
  XOR U21143 ( .A(n17356), .B(n16738), .Z(n20429) );
  XNOR U21144 ( .A(n20430), .B(n20431), .Z(n16738) );
  AND U21145 ( .A(n20432), .B(n20433), .Z(n20430) );
  XNOR U21146 ( .A(n20434), .B(n20435), .Z(n17356) );
  ANDN U21147 ( .B(n20436), .A(n20437), .Z(n20434) );
  XNOR U21148 ( .A(n20438), .B(n20439), .Z(n20372) );
  ANDN U21149 ( .B(n20440), .A(n20441), .Z(n20438) );
  XOR U21150 ( .A(n20442), .B(n18192), .Z(n12567) );
  IV U21151 ( .A(n17282), .Z(n18192) );
  XOR U21152 ( .A(n20443), .B(n16171), .Z(n11057) );
  XOR U21153 ( .A(n20444), .B(n17102), .Z(n16171) );
  IV U21154 ( .A(n17980), .Z(n17102) );
  XOR U21155 ( .A(n19298), .B(n20445), .Z(n17980) );
  XOR U21156 ( .A(n20446), .B(n20447), .Z(n19298) );
  XNOR U21157 ( .A(n20448), .B(n18778), .Z(n20447) );
  XNOR U21158 ( .A(n20449), .B(n20450), .Z(n18778) );
  ANDN U21159 ( .B(n20451), .A(n20452), .Z(n20449) );
  XNOR U21160 ( .A(n17289), .B(n20453), .Z(n20446) );
  XNOR U21161 ( .A(n20454), .B(n17092), .Z(n20453) );
  XNOR U21162 ( .A(n20455), .B(n20456), .Z(n17092) );
  ANDN U21163 ( .B(n20457), .A(n20458), .Z(n20455) );
  XNOR U21164 ( .A(n20459), .B(n20460), .Z(n17289) );
  ANDN U21165 ( .B(n20461), .A(n20462), .Z(n20459) );
  ANDN U21166 ( .B(n12563), .A(n13624), .Z(n20443) );
  XOR U21167 ( .A(n20237), .B(n17186), .Z(n13624) );
  XNOR U21168 ( .A(n20463), .B(n20464), .Z(n19852) );
  XOR U21169 ( .A(n20465), .B(n20466), .Z(n20464) );
  XOR U21170 ( .A(n17975), .B(n20467), .Z(n20463) );
  XOR U21171 ( .A(n19398), .B(n16368), .Z(n20467) );
  XNOR U21172 ( .A(n20468), .B(n20469), .Z(n16368) );
  AND U21173 ( .A(n20470), .B(n20471), .Z(n20468) );
  XNOR U21174 ( .A(n20472), .B(n20473), .Z(n19398) );
  ANDN U21175 ( .B(n20236), .A(n20234), .Z(n20472) );
  XNOR U21176 ( .A(n20474), .B(n20475), .Z(n17975) );
  NOR U21177 ( .A(n20241), .B(n20240), .Z(n20474) );
  XNOR U21178 ( .A(n20477), .B(n20470), .Z(n20237) );
  ANDN U21179 ( .B(n20478), .A(n20471), .Z(n20477) );
  XNOR U21180 ( .A(n20479), .B(n17589), .Z(n12563) );
  XNOR U21181 ( .A(n20482), .B(n16164), .Z(n11863) );
  XOR U21182 ( .A(n20483), .B(n17294), .Z(n16164) );
  XOR U21183 ( .A(n20484), .B(n20485), .Z(n17294) );
  ANDN U21184 ( .B(n13627), .A(n16165), .Z(n20482) );
  XOR U21185 ( .A(n20486), .B(n16613), .Z(n16165) );
  XOR U21186 ( .A(n20489), .B(n18787), .Z(n13627) );
  XNOR U21187 ( .A(n20490), .B(n17345), .Z(n16347) );
  XOR U21188 ( .A(n19914), .B(n19072), .Z(n17345) );
  XNOR U21189 ( .A(n20491), .B(n20492), .Z(n19914) );
  ANDN U21190 ( .B(n20493), .A(n20494), .Z(n20491) );
  NOR U21191 ( .A(n12027), .B(n12026), .Z(n20490) );
  XOR U21192 ( .A(n20495), .B(n16878), .Z(n12026) );
  XOR U21193 ( .A(n18014), .B(n20496), .Z(n12027) );
  XNOR U21194 ( .A(n19299), .B(n20497), .Z(n18014) );
  XOR U21195 ( .A(n20498), .B(n20499), .Z(n19299) );
  XOR U21196 ( .A(n19668), .B(n18854), .Z(n20499) );
  XNOR U21197 ( .A(n20500), .B(n20501), .Z(n18854) );
  NOR U21198 ( .A(n20502), .B(n20503), .Z(n20500) );
  XOR U21199 ( .A(n20504), .B(n20505), .Z(n19668) );
  AND U21200 ( .A(n20506), .B(n20507), .Z(n20504) );
  XOR U21201 ( .A(n20508), .B(n20509), .Z(n20498) );
  XNOR U21202 ( .A(n18294), .B(n19393), .Z(n20509) );
  XNOR U21203 ( .A(n20510), .B(n20511), .Z(n19393) );
  XOR U21204 ( .A(n20514), .B(n20515), .Z(n18294) );
  ANDN U21205 ( .B(n19409), .A(n20516), .Z(n20514) );
  XOR U21206 ( .A(n18674), .B(n10269), .Z(n9268) );
  XNOR U21207 ( .A(n18542), .B(n19076), .Z(n10269) );
  XNOR U21208 ( .A(n20517), .B(n20518), .Z(n19076) );
  XNOR U21209 ( .A(n12334), .B(n13846), .Z(n20518) );
  XNOR U21210 ( .A(n20519), .B(n15807), .Z(n13846) );
  XOR U21211 ( .A(n18045), .B(n20520), .Z(n15807) );
  IV U21212 ( .A(n16004), .Z(n18045) );
  XOR U21213 ( .A(n20521), .B(n20487), .Z(n16004) );
  XNOR U21214 ( .A(n20522), .B(n20523), .Z(n20487) );
  XOR U21215 ( .A(n20007), .B(n19719), .Z(n20523) );
  XOR U21216 ( .A(n20524), .B(n20525), .Z(n19719) );
  ANDN U21217 ( .B(n20526), .A(n20527), .Z(n20524) );
  XNOR U21218 ( .A(n20528), .B(n20529), .Z(n20007) );
  AND U21219 ( .A(n20530), .B(n20531), .Z(n20528) );
  XOR U21220 ( .A(n18281), .B(n20532), .Z(n20522) );
  XNOR U21221 ( .A(n20034), .B(n20533), .Z(n20532) );
  XNOR U21222 ( .A(n20534), .B(n20535), .Z(n20034) );
  ANDN U21223 ( .B(n20536), .A(n20537), .Z(n20534) );
  XNOR U21224 ( .A(n20538), .B(n20539), .Z(n18281) );
  ANDN U21225 ( .B(n20540), .A(n20541), .Z(n20538) );
  NOR U21226 ( .A(n20542), .B(n15808), .Z(n20519) );
  XOR U21227 ( .A(n20543), .B(n15803), .Z(n12334) );
  XOR U21228 ( .A(n20544), .B(n16527), .Z(n15803) );
  XOR U21229 ( .A(n20545), .B(n20546), .Z(n16527) );
  ANDN U21230 ( .B(n15804), .A(n13940), .Z(n20543) );
  IV U21231 ( .A(n18685), .Z(n13940) );
  XOR U21232 ( .A(n19442), .B(n20547), .Z(n18685) );
  XNOR U21233 ( .A(n20548), .B(n20379), .Z(n19442) );
  XNOR U21234 ( .A(n20549), .B(n20550), .Z(n20379) );
  XOR U21235 ( .A(n17510), .B(n18288), .Z(n20550) );
  XOR U21236 ( .A(n20551), .B(n20552), .Z(n18288) );
  ANDN U21237 ( .B(n20553), .A(n20554), .Z(n20551) );
  XOR U21238 ( .A(n20555), .B(n20556), .Z(n17510) );
  XOR U21239 ( .A(n20559), .B(n20560), .Z(n20549) );
  XNOR U21240 ( .A(n16102), .B(n17299), .Z(n20560) );
  XNOR U21241 ( .A(n20561), .B(n20562), .Z(n17299) );
  ANDN U21242 ( .B(n20563), .A(n20564), .Z(n20561) );
  XNOR U21243 ( .A(n20565), .B(n20566), .Z(n16102) );
  NOR U21244 ( .A(n20567), .B(n20568), .Z(n20565) );
  XOR U21245 ( .A(n20569), .B(n17440), .Z(n15804) );
  XNOR U21246 ( .A(n20571), .B(n20572), .Z(n19427) );
  XOR U21247 ( .A(n20095), .B(n18218), .Z(n20572) );
  XNOR U21248 ( .A(n20573), .B(n20574), .Z(n18218) );
  AND U21249 ( .A(n20575), .B(n20576), .Z(n20573) );
  XNOR U21250 ( .A(n20577), .B(n20578), .Z(n20095) );
  ANDN U21251 ( .B(n20579), .A(n20580), .Z(n20577) );
  XNOR U21252 ( .A(n18507), .B(n20581), .Z(n20571) );
  XOR U21253 ( .A(n20149), .B(n20582), .Z(n20581) );
  XNOR U21254 ( .A(n20583), .B(n20584), .Z(n20149) );
  ANDN U21255 ( .B(n20585), .A(n20586), .Z(n20583) );
  XOR U21256 ( .A(n20587), .B(n20588), .Z(n18507) );
  ANDN U21257 ( .B(n20589), .A(n20590), .Z(n20587) );
  XOR U21258 ( .A(n11218), .B(n20591), .Z(n20517) );
  XOR U21259 ( .A(n10984), .B(n12079), .Z(n20591) );
  XNOR U21260 ( .A(n20592), .B(n15800), .Z(n12079) );
  XNOR U21261 ( .A(n20593), .B(n19664), .Z(n15800) );
  XOR U21262 ( .A(n20595), .B(n18438), .Z(n18689) );
  IV U21263 ( .A(n17500), .Z(n18438) );
  XNOR U21264 ( .A(n20596), .B(n20597), .Z(n17500) );
  XNOR U21265 ( .A(n20598), .B(n15814), .Z(n10984) );
  XNOR U21266 ( .A(n20599), .B(n17013), .Z(n15814) );
  NOR U21267 ( .A(n18681), .B(n13936), .Z(n20598) );
  XOR U21268 ( .A(n20600), .B(n18523), .Z(n13936) );
  IV U21269 ( .A(n16412), .Z(n18523) );
  XOR U21270 ( .A(n20601), .B(n20602), .Z(n16412) );
  XOR U21271 ( .A(n19243), .B(n20603), .Z(n18681) );
  XNOR U21272 ( .A(n20604), .B(n15812), .Z(n11218) );
  XOR U21273 ( .A(n17921), .B(n20605), .Z(n15812) );
  NOR U21274 ( .A(n13930), .B(n15811), .Z(n20604) );
  XOR U21275 ( .A(n20606), .B(n16149), .Z(n15811) );
  IV U21276 ( .A(n18791), .Z(n16149) );
  XOR U21277 ( .A(n20607), .B(n18918), .Z(n18791) );
  XNOR U21278 ( .A(n20608), .B(n20609), .Z(n18918) );
  XOR U21279 ( .A(n16680), .B(n16024), .Z(n20609) );
  XOR U21280 ( .A(n20610), .B(n20611), .Z(n16024) );
  NOR U21281 ( .A(n20612), .B(n20613), .Z(n20610) );
  XOR U21282 ( .A(n20614), .B(n20615), .Z(n16680) );
  ANDN U21283 ( .B(n20616), .A(n20617), .Z(n20614) );
  XOR U21284 ( .A(n16104), .B(n20618), .Z(n20608) );
  XNOR U21285 ( .A(n20619), .B(n18385), .Z(n20618) );
  XNOR U21286 ( .A(n20620), .B(n20621), .Z(n18385) );
  ANDN U21287 ( .B(n20622), .A(n20623), .Z(n20620) );
  XNOR U21288 ( .A(n20624), .B(n20625), .Z(n16104) );
  NOR U21289 ( .A(n20626), .B(n20627), .Z(n20624) );
  IV U21290 ( .A(n18676), .Z(n13930) );
  XOR U21291 ( .A(n20628), .B(n19757), .Z(n18676) );
  XOR U21292 ( .A(n20629), .B(n20630), .Z(n18542) );
  XNOR U21293 ( .A(n10117), .B(n10826), .Z(n20630) );
  XNOR U21294 ( .A(n20631), .B(n16899), .Z(n10826) );
  XNOR U21295 ( .A(n20632), .B(n16596), .Z(n16899) );
  ANDN U21296 ( .B(n14687), .A(n18658), .Z(n20631) );
  XNOR U21297 ( .A(n20633), .B(n18777), .Z(n18658) );
  XOR U21298 ( .A(n18476), .B(n20634), .Z(n14687) );
  XNOR U21299 ( .A(n13860), .B(n20635), .Z(n10117) );
  XOR U21300 ( .A(n20636), .B(n4694), .Z(n20635) );
  AND U21301 ( .A(n17218), .B(n13859), .Z(n20636) );
  XNOR U21302 ( .A(n17921), .B(n20637), .Z(n13859) );
  XNOR U21303 ( .A(n19773), .B(n20638), .Z(n17921) );
  XOR U21304 ( .A(n20639), .B(n20640), .Z(n19773) );
  XNOR U21305 ( .A(n18753), .B(n18509), .Z(n20640) );
  XNOR U21306 ( .A(n20641), .B(n20642), .Z(n18509) );
  AND U21307 ( .A(n20643), .B(n20644), .Z(n20641) );
  XNOR U21308 ( .A(n20645), .B(n20646), .Z(n18753) );
  XNOR U21309 ( .A(n18934), .B(n20649), .Z(n20639) );
  XOR U21310 ( .A(n18457), .B(n17058), .Z(n20649) );
  XNOR U21311 ( .A(n20650), .B(n20651), .Z(n17058) );
  NOR U21312 ( .A(n20652), .B(n20653), .Z(n20650) );
  XNOR U21313 ( .A(n20654), .B(n20655), .Z(n18457) );
  AND U21314 ( .A(n20656), .B(n20657), .Z(n20654) );
  XOR U21315 ( .A(n20658), .B(n20659), .Z(n18934) );
  AND U21316 ( .A(n20660), .B(n20661), .Z(n20658) );
  XOR U21317 ( .A(n18207), .B(n20662), .Z(n17218) );
  IV U21318 ( .A(n16757), .Z(n18207) );
  XOR U21319 ( .A(n20665), .B(n17613), .Z(n13860) );
  XNOR U21320 ( .A(n20666), .B(n20667), .Z(n17613) );
  XNOR U21321 ( .A(n9925), .B(n20668), .Z(n20629) );
  XOR U21322 ( .A(n12595), .B(n10298), .Z(n20668) );
  XOR U21323 ( .A(n20669), .B(n13853), .Z(n10298) );
  XOR U21324 ( .A(n20670), .B(n19451), .Z(n13853) );
  ANDN U21325 ( .B(n13854), .A(n14684), .Z(n20669) );
  XOR U21326 ( .A(n20671), .B(n16868), .Z(n14684) );
  XNOR U21327 ( .A(n20673), .B(n20674), .Z(n19595) );
  XNOR U21328 ( .A(n15200), .B(n18098), .Z(n20674) );
  XOR U21329 ( .A(n20675), .B(n20676), .Z(n18098) );
  NOR U21330 ( .A(n20677), .B(n20678), .Z(n20675) );
  XNOR U21331 ( .A(n20679), .B(n20680), .Z(n15200) );
  ANDN U21332 ( .B(n20681), .A(n20682), .Z(n20679) );
  XOR U21333 ( .A(n17407), .B(n20683), .Z(n20673) );
  XNOR U21334 ( .A(n18884), .B(n20015), .Z(n20683) );
  XNOR U21335 ( .A(n20684), .B(n20685), .Z(n20015) );
  NOR U21336 ( .A(n20686), .B(n20687), .Z(n20684) );
  XNOR U21337 ( .A(n20688), .B(n20689), .Z(n18884) );
  XNOR U21338 ( .A(n20692), .B(n20693), .Z(n17407) );
  ANDN U21339 ( .B(n20694), .A(n20695), .Z(n20692) );
  XOR U21340 ( .A(n19780), .B(n20696), .Z(n13854) );
  XOR U21341 ( .A(n20697), .B(n20293), .Z(n19780) );
  AND U21342 ( .A(n20698), .B(n20699), .Z(n20697) );
  XOR U21343 ( .A(n20700), .B(n14195), .Z(n12595) );
  XNOR U21344 ( .A(n20701), .B(n18557), .Z(n14195) );
  ANDN U21345 ( .B(n14196), .A(n17833), .Z(n20700) );
  XOR U21346 ( .A(n20702), .B(n15702), .Z(n17833) );
  IV U21347 ( .A(n17646), .Z(n15702) );
  XOR U21348 ( .A(n20705), .B(n18429), .Z(n14196) );
  XOR U21349 ( .A(n20706), .B(n13863), .Z(n9925) );
  XOR U21350 ( .A(n19243), .B(n20707), .Z(n13863) );
  IV U21351 ( .A(n18412), .Z(n19243) );
  XOR U21352 ( .A(n18751), .B(n19055), .Z(n18412) );
  XNOR U21353 ( .A(n20708), .B(n20709), .Z(n19055) );
  XOR U21354 ( .A(n18307), .B(n19954), .Z(n20709) );
  XNOR U21355 ( .A(n20710), .B(n20711), .Z(n19954) );
  ANDN U21356 ( .B(n20712), .A(n20713), .Z(n20710) );
  XNOR U21357 ( .A(n20714), .B(n20715), .Z(n18307) );
  ANDN U21358 ( .B(n20716), .A(n20717), .Z(n20714) );
  XNOR U21359 ( .A(n15903), .B(n20718), .Z(n20708) );
  XOR U21360 ( .A(n16521), .B(n18874), .Z(n20718) );
  XNOR U21361 ( .A(n20719), .B(n20720), .Z(n18874) );
  ANDN U21362 ( .B(n20721), .A(n20722), .Z(n20719) );
  XNOR U21363 ( .A(n20723), .B(n20724), .Z(n16521) );
  XNOR U21364 ( .A(n20727), .B(n20728), .Z(n15903) );
  XOR U21365 ( .A(n20731), .B(n20732), .Z(n18751) );
  XNOR U21366 ( .A(n20733), .B(n19373), .Z(n20732) );
  XNOR U21367 ( .A(n20734), .B(n20735), .Z(n19373) );
  ANDN U21368 ( .B(n20736), .A(n20737), .Z(n20734) );
  XOR U21369 ( .A(n19104), .B(n20738), .Z(n20731) );
  XOR U21370 ( .A(n20739), .B(n17621), .Z(n20738) );
  XNOR U21371 ( .A(n20740), .B(n20741), .Z(n17621) );
  NOR U21372 ( .A(n20742), .B(n20743), .Z(n20740) );
  XNOR U21373 ( .A(n20744), .B(n20745), .Z(n19104) );
  ANDN U21374 ( .B(n20746), .A(n20556), .Z(n20744) );
  ANDN U21375 ( .B(n13864), .A(n15102), .Z(n20706) );
  IV U21376 ( .A(n18670), .Z(n15102) );
  XOR U21377 ( .A(n18266), .B(n18841), .Z(n18670) );
  XNOR U21378 ( .A(n20747), .B(n20748), .Z(n18841) );
  XNOR U21379 ( .A(n20750), .B(n20751), .Z(n18757) );
  XNOR U21380 ( .A(n17588), .B(n19359), .Z(n20751) );
  XNOR U21381 ( .A(n20752), .B(n20753), .Z(n19359) );
  ANDN U21382 ( .B(n18849), .A(n18851), .Z(n20752) );
  XOR U21383 ( .A(n20754), .B(n20187), .Z(n17588) );
  NOR U21384 ( .A(n20749), .B(n20748), .Z(n20754) );
  XOR U21385 ( .A(n17848), .B(n20755), .Z(n20750) );
  XOR U21386 ( .A(n20479), .B(n18440), .Z(n20755) );
  XOR U21387 ( .A(n20756), .B(n20177), .Z(n18440) );
  AND U21388 ( .A(n18911), .B(n18910), .Z(n20756) );
  XNOR U21389 ( .A(n20757), .B(n20183), .Z(n20479) );
  ANDN U21390 ( .B(n18845), .A(n18846), .Z(n20757) );
  IV U21391 ( .A(n20758), .Z(n18846) );
  XNOR U21392 ( .A(n20759), .B(n20174), .Z(n17848) );
  ANDN U21393 ( .B(n19731), .A(n19729), .Z(n20759) );
  XOR U21394 ( .A(n20760), .B(n20761), .Z(n19516) );
  XNOR U21395 ( .A(n20762), .B(n18536), .Z(n20761) );
  XOR U21396 ( .A(n20763), .B(n20764), .Z(n18536) );
  ANDN U21397 ( .B(n20211), .A(n20213), .Z(n20763) );
  XOR U21398 ( .A(n20765), .B(n20766), .Z(n20760) );
  XNOR U21399 ( .A(n20073), .B(n16503), .Z(n20766) );
  XOR U21400 ( .A(n20767), .B(n20768), .Z(n16503) );
  ANDN U21401 ( .B(n20219), .A(n20769), .Z(n20767) );
  XOR U21402 ( .A(n20770), .B(n20771), .Z(n20073) );
  AND U21403 ( .A(n20215), .B(n20216), .Z(n20770) );
  XOR U21404 ( .A(n20772), .B(n18502), .Z(n13864) );
  XNOR U21405 ( .A(n20773), .B(n20545), .Z(n18502) );
  XOR U21406 ( .A(n20774), .B(n20775), .Z(n20545) );
  XNOR U21407 ( .A(n17610), .B(n17925), .Z(n20775) );
  XNOR U21408 ( .A(n20776), .B(n20494), .Z(n17925) );
  NOR U21409 ( .A(n20493), .B(n20777), .Z(n20776) );
  XNOR U21410 ( .A(n20778), .B(n19910), .Z(n17610) );
  NOR U21411 ( .A(n19911), .B(n20779), .Z(n20778) );
  XNOR U21412 ( .A(n14995), .B(n20780), .Z(n20774) );
  XNOR U21413 ( .A(n16095), .B(n18392), .Z(n20780) );
  XOR U21414 ( .A(n20781), .B(n19906), .Z(n18392) );
  ANDN U21415 ( .B(n19907), .A(n20782), .Z(n20781) );
  XNOR U21416 ( .A(n20783), .B(n19917), .Z(n16095) );
  NOR U21417 ( .A(n20784), .B(n19918), .Z(n20783) );
  XNOR U21418 ( .A(n20785), .B(n20786), .Z(n14995) );
  ANDN U21419 ( .B(n20787), .A(n20788), .Z(n20785) );
  XOR U21420 ( .A(n20789), .B(n15808), .Z(n18674) );
  XOR U21421 ( .A(n20790), .B(n18429), .Z(n15808) );
  XOR U21422 ( .A(n19682), .B(n20791), .Z(n18429) );
  XOR U21423 ( .A(n20792), .B(n20793), .Z(n19682) );
  XNOR U21424 ( .A(n20794), .B(n18540), .Z(n20793) );
  XOR U21425 ( .A(n20795), .B(n20796), .Z(n18540) );
  ANDN U21426 ( .B(n20797), .A(n20798), .Z(n20795) );
  XOR U21427 ( .A(n18968), .B(n20799), .Z(n20792) );
  XOR U21428 ( .A(n19286), .B(n17475), .Z(n20799) );
  XNOR U21429 ( .A(n20800), .B(n20801), .Z(n17475) );
  NOR U21430 ( .A(n20802), .B(n20803), .Z(n20800) );
  XOR U21431 ( .A(n20804), .B(n20805), .Z(n19286) );
  NOR U21432 ( .A(n20806), .B(n20807), .Z(n20804) );
  XNOR U21433 ( .A(n20808), .B(n20809), .Z(n18968) );
  NOR U21434 ( .A(n20810), .B(n20811), .Z(n20808) );
  NOR U21435 ( .A(n15497), .B(n15498), .Z(n20789) );
  XNOR U21436 ( .A(n20812), .B(n15193), .Z(n15498) );
  IV U21437 ( .A(n19769), .Z(n15193) );
  IV U21438 ( .A(n20542), .Z(n15497) );
  XOR U21439 ( .A(n20762), .B(n20074), .Z(n20542) );
  XOR U21440 ( .A(n20813), .B(n20814), .Z(n20762) );
  AND U21441 ( .A(n20204), .B(n20202), .Z(n20813) );
  XOR U21442 ( .A(n2566), .B(n20815), .Z(n19713) );
  XNOR U21443 ( .A(n3531), .B(n9317), .Z(n20815) );
  XNOR U21444 ( .A(n20816), .B(n6686), .Z(n9317) );
  IV U21445 ( .A(n9333), .Z(n6686) );
  XNOR U21446 ( .A(n12352), .B(n10521), .Z(n9333) );
  XNOR U21447 ( .A(n13972), .B(n15181), .Z(n10521) );
  XNOR U21448 ( .A(n20817), .B(n20818), .Z(n15181) );
  XOR U21449 ( .A(n10817), .B(n11948), .Z(n20818) );
  XNOR U21450 ( .A(n20819), .B(n14858), .Z(n11948) );
  XOR U21451 ( .A(n18403), .B(n20820), .Z(n14858) );
  ANDN U21452 ( .B(n15660), .A(n15661), .Z(n20819) );
  IV U21453 ( .A(n14307), .Z(n15661) );
  XOR U21454 ( .A(n19970), .B(n16108), .Z(n14307) );
  XNOR U21455 ( .A(n19959), .B(n20821), .Z(n16108) );
  XOR U21456 ( .A(n20822), .B(n20823), .Z(n19959) );
  XNOR U21457 ( .A(n20824), .B(n20825), .Z(n20823) );
  XOR U21458 ( .A(n18287), .B(n20826), .Z(n20822) );
  XOR U21459 ( .A(n18049), .B(n20827), .Z(n20826) );
  XNOR U21460 ( .A(n20828), .B(n20788), .Z(n18049) );
  NOR U21461 ( .A(n20829), .B(n20830), .Z(n20828) );
  XOR U21462 ( .A(n20831), .B(n20779), .Z(n18287) );
  ANDN U21463 ( .B(n20832), .A(n19909), .Z(n20831) );
  IV U21464 ( .A(n20833), .Z(n19909) );
  XNOR U21465 ( .A(n20834), .B(n20835), .Z(n19970) );
  XOR U21466 ( .A(n18563), .B(n20836), .Z(n15660) );
  XNOR U21467 ( .A(n20837), .B(n14865), .Z(n10817) );
  ANDN U21468 ( .B(n15665), .A(n15666), .Z(n20837) );
  XNOR U21469 ( .A(n20839), .B(n16889), .Z(n15666) );
  XNOR U21470 ( .A(n20328), .B(n18182), .Z(n15665) );
  XOR U21471 ( .A(n20840), .B(n20841), .Z(n20328) );
  ANDN U21472 ( .B(n20842), .A(n20843), .Z(n20840) );
  XOR U21473 ( .A(n9769), .B(n20844), .Z(n20817) );
  XOR U21474 ( .A(n9279), .B(n11308), .Z(n20844) );
  XNOR U21475 ( .A(n20845), .B(n14862), .Z(n11308) );
  XNOR U21476 ( .A(n20846), .B(n19987), .Z(n14862) );
  IV U21477 ( .A(n19389), .Z(n19987) );
  ANDN U21478 ( .B(n14312), .A(n16955), .Z(n20845) );
  XOR U21479 ( .A(n19060), .B(n20847), .Z(n16955) );
  IV U21480 ( .A(n20302), .Z(n19060) );
  XOR U21481 ( .A(n20848), .B(n20849), .Z(n14312) );
  XNOR U21482 ( .A(n20850), .B(n14856), .Z(n9279) );
  XNOR U21483 ( .A(n20851), .B(n16090), .Z(n14856) );
  XOR U21484 ( .A(n20852), .B(n18955), .Z(n16090) );
  XNOR U21485 ( .A(n20853), .B(n20854), .Z(n18955) );
  XNOR U21486 ( .A(n20855), .B(n20856), .Z(n20854) );
  XOR U21487 ( .A(n20857), .B(n20858), .Z(n20853) );
  XOR U21488 ( .A(n20859), .B(n17303), .Z(n20858) );
  XNOR U21489 ( .A(n20860), .B(n20861), .Z(n17303) );
  ANDN U21490 ( .B(n20862), .A(n20863), .Z(n20860) );
  XOR U21491 ( .A(n18476), .B(n20864), .Z(n15673) );
  XNOR U21492 ( .A(n20865), .B(n19054), .Z(n18476) );
  XOR U21493 ( .A(n20866), .B(n20867), .Z(n19054) );
  XOR U21494 ( .A(n17447), .B(n20868), .Z(n20867) );
  XNOR U21495 ( .A(n20869), .B(n20870), .Z(n17447) );
  ANDN U21496 ( .B(n20871), .A(n20872), .Z(n20869) );
  XNOR U21497 ( .A(n15255), .B(n20873), .Z(n20866) );
  XOR U21498 ( .A(n20874), .B(n18595), .Z(n20873) );
  XNOR U21499 ( .A(n20875), .B(n20876), .Z(n18595) );
  ANDN U21500 ( .B(n20877), .A(n20878), .Z(n20875) );
  XNOR U21501 ( .A(n20879), .B(n20880), .Z(n15255) );
  XOR U21502 ( .A(n20883), .B(n18177), .Z(n14316) );
  IV U21503 ( .A(n18586), .Z(n18177) );
  XNOR U21504 ( .A(n20884), .B(n18700), .Z(n18586) );
  XOR U21505 ( .A(n20885), .B(n20886), .Z(n18700) );
  XNOR U21506 ( .A(n18693), .B(n18799), .Z(n20886) );
  XNOR U21507 ( .A(n20887), .B(n20888), .Z(n18799) );
  ANDN U21508 ( .B(n19807), .A(n19805), .Z(n20887) );
  XNOR U21509 ( .A(n20889), .B(n20890), .Z(n18693) );
  ANDN U21510 ( .B(n19816), .A(n20891), .Z(n20889) );
  XNOR U21511 ( .A(n18763), .B(n20892), .Z(n20885) );
  XNOR U21512 ( .A(n20893), .B(n18831), .Z(n20892) );
  XOR U21513 ( .A(n20894), .B(n20895), .Z(n18831) );
  ANDN U21514 ( .B(n19803), .A(n20896), .Z(n20894) );
  XOR U21515 ( .A(n20897), .B(n20898), .Z(n18763) );
  ANDN U21516 ( .B(n19812), .A(n19810), .Z(n20897) );
  XNOR U21517 ( .A(n20899), .B(n14868), .Z(n9769) );
  XNOR U21518 ( .A(n20900), .B(n15883), .Z(n14868) );
  XOR U21519 ( .A(n20901), .B(n20902), .Z(n15883) );
  ANDN U21520 ( .B(n14320), .A(n15677), .Z(n20899) );
  XOR U21521 ( .A(n20903), .B(n18337), .Z(n15677) );
  XNOR U21522 ( .A(n18016), .B(n20904), .Z(n14320) );
  XOR U21523 ( .A(n20905), .B(n20906), .Z(n13972) );
  XNOR U21524 ( .A(n16938), .B(n12490), .Z(n20906) );
  XNOR U21525 ( .A(n20907), .B(n15793), .Z(n12490) );
  XOR U21526 ( .A(n20908), .B(n20302), .Z(n15793) );
  NOR U21527 ( .A(n12355), .B(n12354), .Z(n20907) );
  XNOR U21528 ( .A(n17483), .B(n20909), .Z(n12354) );
  XOR U21529 ( .A(n19515), .B(n20910), .Z(n17483) );
  XOR U21530 ( .A(n20911), .B(n20912), .Z(n19515) );
  XNOR U21531 ( .A(n16153), .B(n17663), .Z(n20912) );
  XNOR U21532 ( .A(n20913), .B(n20914), .Z(n17663) );
  NOR U21533 ( .A(n20915), .B(n20916), .Z(n20913) );
  XNOR U21534 ( .A(n20917), .B(n20918), .Z(n16153) );
  NOR U21535 ( .A(n20919), .B(n20920), .Z(n20917) );
  XNOR U21536 ( .A(n15268), .B(n20921), .Z(n20911) );
  XNOR U21537 ( .A(n17593), .B(n18459), .Z(n20921) );
  XOR U21538 ( .A(n20922), .B(n20923), .Z(n18459) );
  NOR U21539 ( .A(n20924), .B(n20925), .Z(n20922) );
  XNOR U21540 ( .A(n20926), .B(n20927), .Z(n17593) );
  NOR U21541 ( .A(n20928), .B(n20929), .Z(n20926) );
  XOR U21542 ( .A(n20930), .B(n20931), .Z(n15268) );
  ANDN U21543 ( .B(n20932), .A(n20933), .Z(n20930) );
  XOR U21544 ( .A(n17302), .B(n20855), .Z(n12355) );
  XNOR U21545 ( .A(n20934), .B(n20935), .Z(n20855) );
  NOR U21546 ( .A(n20936), .B(n20937), .Z(n20934) );
  XNOR U21547 ( .A(n20938), .B(n16947), .Z(n16938) );
  XNOR U21548 ( .A(n20939), .B(n16841), .Z(n16947) );
  XOR U21549 ( .A(n20940), .B(n19822), .Z(n16841) );
  XOR U21550 ( .A(n20941), .B(n20942), .Z(n19822) );
  XNOR U21551 ( .A(n17202), .B(n17652), .Z(n20942) );
  XNOR U21552 ( .A(n20943), .B(n20944), .Z(n17652) );
  XNOR U21553 ( .A(n20947), .B(n20948), .Z(n17202) );
  XOR U21554 ( .A(n20951), .B(n20952), .Z(n20941) );
  XNOR U21555 ( .A(n17937), .B(n19189), .Z(n20952) );
  XNOR U21556 ( .A(n20953), .B(n20954), .Z(n19189) );
  ANDN U21557 ( .B(n20955), .A(n20956), .Z(n20953) );
  XOR U21558 ( .A(n20957), .B(n20958), .Z(n17937) );
  NOR U21559 ( .A(n17128), .B(n12347), .Z(n20938) );
  XNOR U21560 ( .A(n18321), .B(n20961), .Z(n12347) );
  XOR U21561 ( .A(n20962), .B(n20664), .Z(n18321) );
  XOR U21562 ( .A(n20963), .B(n20964), .Z(n20664) );
  XOR U21563 ( .A(n16746), .B(n18310), .Z(n20964) );
  XNOR U21564 ( .A(n20965), .B(n20966), .Z(n18310) );
  NOR U21565 ( .A(n20967), .B(n20651), .Z(n20965) );
  XNOR U21566 ( .A(n20968), .B(n20969), .Z(n16746) );
  ANDN U21567 ( .B(n20655), .A(n20970), .Z(n20968) );
  XOR U21568 ( .A(n16007), .B(n20971), .Z(n20963) );
  XOR U21569 ( .A(n19004), .B(n19114), .Z(n20971) );
  XOR U21570 ( .A(n20972), .B(n20973), .Z(n19114) );
  ANDN U21571 ( .B(n20642), .A(n20974), .Z(n20972) );
  XNOR U21572 ( .A(n20975), .B(n20976), .Z(n19004) );
  NOR U21573 ( .A(n20659), .B(n20977), .Z(n20975) );
  XNOR U21574 ( .A(n20978), .B(n20979), .Z(n16007) );
  NOR U21575 ( .A(n20646), .B(n20980), .Z(n20978) );
  IV U21576 ( .A(n20981), .Z(n20646) );
  XOR U21577 ( .A(n20310), .B(n18834), .Z(n17128) );
  XNOR U21578 ( .A(n20982), .B(n20983), .Z(n20310) );
  ANDN U21579 ( .B(n20984), .A(n20985), .Z(n20982) );
  XNOR U21580 ( .A(n12502), .B(n20986), .Z(n20905) );
  XOR U21581 ( .A(n11354), .B(n10849), .Z(n20986) );
  XNOR U21582 ( .A(n20987), .B(n15782), .Z(n10849) );
  XNOR U21583 ( .A(n20349), .B(n16813), .Z(n15782) );
  XOR U21584 ( .A(n20990), .B(n20991), .Z(n20349) );
  NOR U21585 ( .A(n20992), .B(n20993), .Z(n20990) );
  NOR U21586 ( .A(n17134), .B(n16944), .Z(n20987) );
  XNOR U21587 ( .A(n20994), .B(n15789), .Z(n11354) );
  XNOR U21588 ( .A(n18187), .B(n20995), .Z(n15789) );
  ANDN U21589 ( .B(n15275), .A(n17138), .Z(n20994) );
  IV U21590 ( .A(n15277), .Z(n17138) );
  XOR U21591 ( .A(n20996), .B(n16579), .Z(n15277) );
  XNOR U21592 ( .A(n20997), .B(n20998), .Z(n16579) );
  XNOR U21593 ( .A(n18563), .B(n20999), .Z(n15275) );
  XNOR U21594 ( .A(n21000), .B(n15778), .Z(n12502) );
  XOR U21595 ( .A(n18048), .B(n20827), .Z(n15778) );
  XNOR U21596 ( .A(n21001), .B(n20784), .Z(n20827) );
  NOR U21597 ( .A(n21002), .B(n19916), .Z(n21001) );
  ANDN U21598 ( .B(n12429), .A(n12430), .Z(n21000) );
  XOR U21599 ( .A(n21003), .B(n17503), .Z(n12430) );
  XNOR U21600 ( .A(n20307), .B(n20297), .Z(n17503) );
  XNOR U21601 ( .A(n21004), .B(n21005), .Z(n20297) );
  XOR U21602 ( .A(n18528), .B(n18477), .Z(n21005) );
  XNOR U21603 ( .A(n21006), .B(n21007), .Z(n18477) );
  ANDN U21604 ( .B(n21008), .A(n21009), .Z(n21006) );
  XNOR U21605 ( .A(n21010), .B(n21011), .Z(n18528) );
  NOR U21606 ( .A(n21012), .B(n21013), .Z(n21010) );
  XOR U21607 ( .A(n18444), .B(n21014), .Z(n21004) );
  XOR U21608 ( .A(n21015), .B(n21016), .Z(n21014) );
  XNOR U21609 ( .A(n21017), .B(n21018), .Z(n18444) );
  ANDN U21610 ( .B(n21019), .A(n21020), .Z(n21017) );
  XNOR U21611 ( .A(n21021), .B(n21022), .Z(n20307) );
  XNOR U21612 ( .A(n21023), .B(n17339), .Z(n21022) );
  XNOR U21613 ( .A(n21024), .B(n21025), .Z(n17339) );
  AND U21614 ( .A(n21026), .B(n21027), .Z(n21024) );
  XOR U21615 ( .A(n18231), .B(n21028), .Z(n21021) );
  XOR U21616 ( .A(n18278), .B(n21029), .Z(n21028) );
  XNOR U21617 ( .A(n21030), .B(n21031), .Z(n18278) );
  ANDN U21618 ( .B(n21032), .A(n21033), .Z(n21030) );
  XNOR U21619 ( .A(n21034), .B(n21035), .Z(n18231) );
  NOR U21620 ( .A(n21036), .B(n21037), .Z(n21034) );
  XOR U21621 ( .A(n21038), .B(n16531), .Z(n12429) );
  XNOR U21622 ( .A(n21039), .B(n16944), .Z(n12352) );
  XNOR U21623 ( .A(n19407), .B(n17541), .Z(n16944) );
  IV U21624 ( .A(n18798), .Z(n17541) );
  XOR U21625 ( .A(n21040), .B(n20507), .Z(n19407) );
  ANDN U21626 ( .B(n21041), .A(n21042), .Z(n21040) );
  AND U21627 ( .A(n15780), .B(n17134), .Z(n21039) );
  XOR U21628 ( .A(n21043), .B(n16110), .Z(n17134) );
  IV U21629 ( .A(n16620), .Z(n16110) );
  XOR U21630 ( .A(n20485), .B(n19614), .Z(n16620) );
  XNOR U21631 ( .A(n21044), .B(n21045), .Z(n19614) );
  XOR U21632 ( .A(n19124), .B(n19791), .Z(n21045) );
  XOR U21633 ( .A(n21046), .B(n21047), .Z(n19791) );
  ANDN U21634 ( .B(n21048), .A(n21049), .Z(n21046) );
  XNOR U21635 ( .A(n21050), .B(n21051), .Z(n19124) );
  ANDN U21636 ( .B(n21052), .A(n21053), .Z(n21050) );
  XNOR U21637 ( .A(n16037), .B(n21054), .Z(n21044) );
  XOR U21638 ( .A(n18021), .B(n17696), .Z(n21054) );
  XNOR U21639 ( .A(n21055), .B(n21056), .Z(n17696) );
  ANDN U21640 ( .B(n21057), .A(n21058), .Z(n21055) );
  XNOR U21641 ( .A(n21059), .B(n21060), .Z(n18021) );
  NOR U21642 ( .A(n21061), .B(n21062), .Z(n21059) );
  XOR U21643 ( .A(n21063), .B(n21064), .Z(n16037) );
  ANDN U21644 ( .B(n21065), .A(n21066), .Z(n21063) );
  XNOR U21645 ( .A(n21067), .B(n21068), .Z(n20485) );
  XOR U21646 ( .A(n19388), .B(n19986), .Z(n21068) );
  XNOR U21647 ( .A(n21069), .B(n21070), .Z(n19986) );
  AND U21648 ( .A(n21071), .B(n21072), .Z(n21069) );
  XOR U21649 ( .A(n21073), .B(n21074), .Z(n19388) );
  ANDN U21650 ( .B(n21075), .A(n21076), .Z(n21073) );
  XOR U21651 ( .A(n21077), .B(n21078), .Z(n21067) );
  XNOR U21652 ( .A(n19501), .B(n20846), .Z(n21078) );
  XNOR U21653 ( .A(n21079), .B(n21080), .Z(n20846) );
  NOR U21654 ( .A(n21081), .B(n21082), .Z(n21079) );
  XNOR U21655 ( .A(n21083), .B(n21084), .Z(n19501) );
  AND U21656 ( .A(n21085), .B(n21086), .Z(n21083) );
  XOR U21657 ( .A(n19530), .B(n15532), .Z(n15780) );
  IV U21658 ( .A(n18195), .Z(n15532) );
  XNOR U21659 ( .A(n21087), .B(n20699), .Z(n19530) );
  ANDN U21660 ( .B(n20292), .A(n20291), .Z(n21087) );
  NOR U21661 ( .A(n7127), .B(n9262), .Z(n20816) );
  XNOR U21662 ( .A(n14943), .B(n11448), .Z(n9262) );
  IV U21663 ( .A(n9870), .Z(n11448) );
  XOR U21664 ( .A(n13117), .B(n12756), .Z(n9870) );
  XNOR U21665 ( .A(n21088), .B(n21089), .Z(n12756) );
  XNOR U21666 ( .A(n12884), .B(n11785), .Z(n21089) );
  XNOR U21667 ( .A(n21090), .B(n15202), .Z(n11785) );
  XOR U21668 ( .A(n15299), .B(n21091), .Z(n15202) );
  ANDN U21669 ( .B(n14941), .A(n12833), .Z(n21090) );
  XOR U21670 ( .A(n21094), .B(n15679), .Z(n12833) );
  IV U21671 ( .A(n21095), .Z(n15679) );
  XNOR U21672 ( .A(n21097), .B(n19763), .Z(n18100) );
  XNOR U21673 ( .A(n21098), .B(n21099), .Z(n19763) );
  XNOR U21674 ( .A(n18297), .B(n16958), .Z(n21099) );
  XOR U21675 ( .A(n21100), .B(n19620), .Z(n16958) );
  ANDN U21676 ( .B(n21101), .A(n21102), .Z(n21100) );
  XNOR U21677 ( .A(n21103), .B(n21104), .Z(n18297) );
  NOR U21678 ( .A(n21105), .B(n21106), .Z(n21103) );
  XOR U21679 ( .A(n19123), .B(n21107), .Z(n21098) );
  XOR U21680 ( .A(n21108), .B(n21109), .Z(n21107) );
  XNOR U21681 ( .A(n21110), .B(n20024), .Z(n19123) );
  ANDN U21682 ( .B(n21111), .A(n21112), .Z(n21110) );
  XNOR U21683 ( .A(n21113), .B(n15187), .Z(n12884) );
  XNOR U21684 ( .A(n15962), .B(n21114), .Z(n15187) );
  ANDN U21685 ( .B(n12822), .A(n14945), .Z(n21113) );
  XOR U21686 ( .A(n19348), .B(n14967), .Z(n14945) );
  XNOR U21687 ( .A(n21115), .B(n20133), .Z(n14967) );
  XNOR U21688 ( .A(n21116), .B(n21117), .Z(n20133) );
  XOR U21689 ( .A(n18191), .B(n20442), .Z(n21117) );
  XOR U21690 ( .A(n21118), .B(n21119), .Z(n20442) );
  AND U21691 ( .A(n21084), .B(n21120), .Z(n21118) );
  XNOR U21692 ( .A(n21121), .B(n21122), .Z(n18191) );
  ANDN U21693 ( .B(n21070), .A(n21123), .Z(n21121) );
  XOR U21694 ( .A(n18580), .B(n21124), .Z(n21116) );
  XNOR U21695 ( .A(n21125), .B(n17281), .Z(n21124) );
  XNOR U21696 ( .A(n21126), .B(n21127), .Z(n17281) );
  XNOR U21697 ( .A(n21129), .B(n21130), .Z(n18580) );
  AND U21698 ( .A(n21131), .B(n21132), .Z(n21129) );
  XOR U21699 ( .A(n21133), .B(n20984), .Z(n19348) );
  NOR U21700 ( .A(n21134), .B(n21135), .Z(n21133) );
  XOR U21701 ( .A(n21136), .B(n16664), .Z(n12822) );
  XOR U21702 ( .A(n11921), .B(n21137), .Z(n21088) );
  XOR U21703 ( .A(n9564), .B(n10384), .Z(n21137) );
  XNOR U21704 ( .A(n21138), .B(n15684), .Z(n10384) );
  IV U21705 ( .A(n15189), .Z(n15684) );
  XOR U21706 ( .A(n17276), .B(n20167), .Z(n15189) );
  XOR U21707 ( .A(n21139), .B(n19896), .Z(n20167) );
  IV U21708 ( .A(n21140), .Z(n19896) );
  NOR U21709 ( .A(n21141), .B(n20369), .Z(n21139) );
  ANDN U21710 ( .B(n15685), .A(n14828), .Z(n21138) );
  IV U21711 ( .A(n21142), .Z(n14828) );
  XOR U21712 ( .A(n21143), .B(n15198), .Z(n9564) );
  XOR U21713 ( .A(n21144), .B(n15653), .Z(n15198) );
  XOR U21714 ( .A(n21145), .B(n18578), .Z(n12826) );
  XNOR U21715 ( .A(n21108), .B(n16957), .Z(n14947) );
  XNOR U21716 ( .A(n21146), .B(n19844), .Z(n21108) );
  NOR U21717 ( .A(n21147), .B(n21148), .Z(n21146) );
  XNOR U21718 ( .A(n21149), .B(n15194), .Z(n11921) );
  XOR U21719 ( .A(n21150), .B(n18403), .Z(n15194) );
  XOR U21720 ( .A(n19670), .B(n20484), .Z(n18403) );
  XNOR U21721 ( .A(n21151), .B(n21152), .Z(n20484) );
  XNOR U21722 ( .A(n17047), .B(n18178), .Z(n21152) );
  XNOR U21723 ( .A(n21153), .B(n19355), .Z(n18178) );
  ANDN U21724 ( .B(n19356), .A(n21154), .Z(n21153) );
  XNOR U21725 ( .A(n21155), .B(n21134), .Z(n17047) );
  AND U21726 ( .A(n20983), .B(n21135), .Z(n21155) );
  XOR U21727 ( .A(n17211), .B(n21156), .Z(n21151) );
  XNOR U21728 ( .A(n18081), .B(n17408), .Z(n21156) );
  XNOR U21729 ( .A(n21157), .B(n19345), .Z(n17408) );
  ANDN U21730 ( .B(n19346), .A(n20318), .Z(n21157) );
  IV U21731 ( .A(n21158), .Z(n20318) );
  XNOR U21732 ( .A(n21159), .B(n19351), .Z(n18081) );
  AND U21733 ( .A(n21160), .B(n19352), .Z(n21159) );
  XNOR U21734 ( .A(n21161), .B(n19342), .Z(n17211) );
  AND U21735 ( .A(n19341), .B(n20312), .Z(n21161) );
  XOR U21736 ( .A(n21162), .B(n21163), .Z(n19670) );
  XNOR U21737 ( .A(n19011), .B(n18815), .Z(n21163) );
  XNOR U21738 ( .A(n21164), .B(n21165), .Z(n18815) );
  AND U21739 ( .A(n21166), .B(n21167), .Z(n21164) );
  XOR U21740 ( .A(n21168), .B(n21169), .Z(n19011) );
  XNOR U21741 ( .A(n19335), .B(n21171), .Z(n21162) );
  XNOR U21742 ( .A(n19292), .B(n19272), .Z(n21171) );
  XNOR U21743 ( .A(n21172), .B(n21173), .Z(n19272) );
  ANDN U21744 ( .B(n21174), .A(n21025), .Z(n21172) );
  IV U21745 ( .A(n21175), .Z(n21025) );
  XNOR U21746 ( .A(n21176), .B(n21177), .Z(n19292) );
  ANDN U21747 ( .B(n21178), .A(n21035), .Z(n21176) );
  XNOR U21748 ( .A(n21179), .B(n21180), .Z(n19335) );
  ANDN U21749 ( .B(n21181), .A(n21182), .Z(n21179) );
  ANDN U21750 ( .B(n14938), .A(n14937), .Z(n21149) );
  XOR U21751 ( .A(n17195), .B(n21183), .Z(n14937) );
  XOR U21752 ( .A(n21184), .B(n21185), .Z(n17195) );
  XOR U21753 ( .A(n20951), .B(n17203), .Z(n14938) );
  XNOR U21754 ( .A(n21186), .B(n21187), .Z(n20373) );
  XOR U21755 ( .A(n21188), .B(n20091), .Z(n21187) );
  XOR U21756 ( .A(n21189), .B(n21190), .Z(n20091) );
  NOR U21757 ( .A(n21191), .B(n20440), .Z(n21189) );
  XOR U21758 ( .A(n16111), .B(n21192), .Z(n21186) );
  XOR U21759 ( .A(n19787), .B(n20035), .Z(n21192) );
  XNOR U21760 ( .A(n21193), .B(n21194), .Z(n20035) );
  NOR U21761 ( .A(n21195), .B(n20436), .Z(n21193) );
  XNOR U21762 ( .A(n21196), .B(n21197), .Z(n19787) );
  ANDN U21763 ( .B(n20422), .A(n21198), .Z(n21196) );
  XNOR U21764 ( .A(n21199), .B(n21200), .Z(n16111) );
  ANDN U21765 ( .B(n20428), .A(n20426), .Z(n21199) );
  XNOR U21766 ( .A(n21202), .B(n21203), .Z(n20951) );
  ANDN U21767 ( .B(n21204), .A(n21205), .Z(n21202) );
  XOR U21768 ( .A(n21206), .B(n21207), .Z(n13117) );
  XNOR U21769 ( .A(n10160), .B(n11903), .Z(n21207) );
  XNOR U21770 ( .A(n21208), .B(n13167), .Z(n11903) );
  XOR U21771 ( .A(n20166), .B(n16815), .Z(n13167) );
  IV U21772 ( .A(n17276), .Z(n16815) );
  XNOR U21773 ( .A(n21209), .B(n19256), .Z(n17276) );
  XNOR U21774 ( .A(n21210), .B(n21211), .Z(n19256) );
  XNOR U21775 ( .A(n18793), .B(n18837), .Z(n21211) );
  XOR U21776 ( .A(n21212), .B(n19895), .Z(n18837) );
  XOR U21777 ( .A(n21213), .B(n21214), .Z(n19895) );
  ANDN U21778 ( .B(n21141), .A(n21140), .Z(n21212) );
  XNOR U21779 ( .A(n21215), .B(n21216), .Z(n21140) );
  XNOR U21780 ( .A(n21217), .B(n19892), .Z(n18793) );
  XOR U21781 ( .A(n21218), .B(n21219), .Z(n19892) );
  XOR U21782 ( .A(n21220), .B(n21221), .Z(n19891) );
  XOR U21783 ( .A(n18535), .B(n21222), .Z(n21210) );
  XNOR U21784 ( .A(n18077), .B(n18479), .Z(n21222) );
  XNOR U21785 ( .A(n21223), .B(n19899), .Z(n18479) );
  XNOR U21786 ( .A(n21224), .B(n21225), .Z(n19899) );
  ANDN U21787 ( .B(n19900), .A(n20169), .Z(n21223) );
  XOR U21788 ( .A(n21226), .B(n21227), .Z(n19900) );
  XNOR U21789 ( .A(n21228), .B(n19882), .Z(n18077) );
  ANDN U21790 ( .B(n19883), .A(n20160), .Z(n21228) );
  XNOR U21791 ( .A(n21229), .B(n21230), .Z(n19883) );
  XNOR U21792 ( .A(n21231), .B(n21232), .Z(n18535) );
  NOR U21793 ( .A(n21233), .B(n19886), .Z(n21231) );
  XNOR U21794 ( .A(n21234), .B(n19886), .Z(n20166) );
  XOR U21795 ( .A(n21235), .B(n21236), .Z(n19886) );
  AND U21796 ( .A(n21237), .B(n21233), .Z(n21234) );
  AND U21797 ( .A(n13291), .B(n14951), .Z(n21208) );
  XNOR U21798 ( .A(n16770), .B(n21238), .Z(n14951) );
  XNOR U21799 ( .A(n21239), .B(n19069), .Z(n13291) );
  XNOR U21800 ( .A(n21240), .B(n21241), .Z(n20017) );
  XNOR U21801 ( .A(n19061), .B(n20847), .Z(n21241) );
  XNOR U21802 ( .A(n21242), .B(n21243), .Z(n20847) );
  ANDN U21803 ( .B(n20695), .A(n20693), .Z(n21242) );
  IV U21804 ( .A(n21244), .Z(n20693) );
  XOR U21805 ( .A(n21245), .B(n21246), .Z(n19061) );
  AND U21806 ( .A(n20686), .B(n20685), .Z(n21245) );
  XOR U21807 ( .A(n21247), .B(n21248), .Z(n21240) );
  XOR U21808 ( .A(n20908), .B(n20303), .Z(n21248) );
  XOR U21809 ( .A(n21249), .B(n21250), .Z(n20303) );
  AND U21810 ( .A(n20678), .B(n20676), .Z(n21249) );
  XOR U21811 ( .A(n21251), .B(n21252), .Z(n20908) );
  AND U21812 ( .A(n20689), .B(n20690), .Z(n21251) );
  XNOR U21813 ( .A(n21254), .B(n12941), .Z(n10160) );
  XOR U21814 ( .A(n21255), .B(n17635), .Z(n12941) );
  IV U21815 ( .A(n17233), .Z(n17635) );
  XOR U21816 ( .A(n19219), .B(n21256), .Z(n17233) );
  XOR U21817 ( .A(n21257), .B(n21258), .Z(n19219) );
  XOR U21818 ( .A(n19375), .B(n21259), .Z(n21258) );
  XOR U21819 ( .A(n21260), .B(n21261), .Z(n19375) );
  ANDN U21820 ( .B(n21262), .A(n21263), .Z(n21260) );
  XOR U21821 ( .A(n21264), .B(n21265), .Z(n21257) );
  XNOR U21822 ( .A(n21266), .B(n18233), .Z(n21265) );
  XOR U21823 ( .A(n21267), .B(n21268), .Z(n18233) );
  ANDN U21824 ( .B(n21269), .A(n21270), .Z(n21267) );
  ANDN U21825 ( .B(n14955), .A(n13177), .Z(n21254) );
  IV U21826 ( .A(n14956), .Z(n13177) );
  XOR U21827 ( .A(n21271), .B(n18712), .Z(n14956) );
  XOR U21828 ( .A(n20859), .B(n17302), .Z(n14955) );
  IV U21829 ( .A(n21272), .Z(n17302) );
  XNOR U21830 ( .A(n21273), .B(n21274), .Z(n20859) );
  NOR U21831 ( .A(n21275), .B(n21276), .Z(n21273) );
  XOR U21832 ( .A(n11452), .B(n21277), .Z(n21206) );
  XOR U21833 ( .A(n15934), .B(n15627), .Z(n21277) );
  XNOR U21834 ( .A(n21278), .B(n12937), .Z(n15627) );
  XNOR U21835 ( .A(n21279), .B(n16071), .Z(n12937) );
  XOR U21836 ( .A(n21280), .B(n15650), .Z(n13173) );
  XNOR U21837 ( .A(n21281), .B(n20386), .Z(n15650) );
  XNOR U21838 ( .A(n21282), .B(n21283), .Z(n20386) );
  XNOR U21839 ( .A(n17624), .B(n17457), .Z(n21283) );
  XNOR U21840 ( .A(n21284), .B(n21285), .Z(n17457) );
  NOR U21841 ( .A(n21286), .B(n21287), .Z(n21284) );
  XNOR U21842 ( .A(n21288), .B(n21289), .Z(n17624) );
  AND U21843 ( .A(n21290), .B(n21291), .Z(n21288) );
  XNOR U21844 ( .A(n17269), .B(n21292), .Z(n21282) );
  XOR U21845 ( .A(n19237), .B(n21293), .Z(n21292) );
  XNOR U21846 ( .A(n21294), .B(n21295), .Z(n19237) );
  NOR U21847 ( .A(n21296), .B(n21297), .Z(n21294) );
  XOR U21848 ( .A(n21298), .B(n21299), .Z(n17269) );
  ANDN U21849 ( .B(n21300), .A(n21301), .Z(n21298) );
  XNOR U21850 ( .A(n17231), .B(n21302), .Z(n14961) );
  XOR U21851 ( .A(n19115), .B(n19797), .Z(n17231) );
  XNOR U21852 ( .A(n21303), .B(n21304), .Z(n19797) );
  XOR U21853 ( .A(n17911), .B(n19608), .Z(n21304) );
  XOR U21854 ( .A(n21305), .B(n21306), .Z(n19608) );
  NOR U21855 ( .A(n21307), .B(n21308), .Z(n21305) );
  XNOR U21856 ( .A(n21309), .B(n21310), .Z(n17911) );
  XOR U21857 ( .A(n18164), .B(n21313), .Z(n21303) );
  XOR U21858 ( .A(n17657), .B(n21314), .Z(n21313) );
  XNOR U21859 ( .A(n21315), .B(n21316), .Z(n17657) );
  ANDN U21860 ( .B(n21317), .A(n21318), .Z(n21315) );
  XOR U21861 ( .A(n21319), .B(n21320), .Z(n18164) );
  NOR U21862 ( .A(n21321), .B(n21322), .Z(n21319) );
  XOR U21863 ( .A(n21323), .B(n21324), .Z(n19115) );
  XNOR U21864 ( .A(n21325), .B(n21326), .Z(n21324) );
  XOR U21865 ( .A(n18235), .B(n21327), .Z(n21323) );
  XOR U21866 ( .A(n19376), .B(n17104), .Z(n21327) );
  XNOR U21867 ( .A(n21328), .B(n20648), .Z(n17104) );
  ANDN U21868 ( .B(n20980), .A(n20979), .Z(n21328) );
  IV U21869 ( .A(n21329), .Z(n20979) );
  XNOR U21870 ( .A(n21330), .B(n20652), .Z(n19376) );
  IV U21871 ( .A(n21331), .Z(n20652) );
  ANDN U21872 ( .B(n20967), .A(n20966), .Z(n21330) );
  XNOR U21873 ( .A(n21332), .B(n20644), .Z(n18235) );
  AND U21874 ( .A(n20974), .B(n20973), .Z(n21332) );
  XOR U21875 ( .A(n21333), .B(n12945), .Z(n15934) );
  XOR U21876 ( .A(n18171), .B(n21334), .Z(n12945) );
  XOR U21877 ( .A(n21335), .B(n21336), .Z(n18171) );
  AND U21878 ( .A(n13273), .B(n14965), .Z(n21333) );
  XNOR U21879 ( .A(n19781), .B(n20696), .Z(n14965) );
  XOR U21880 ( .A(n21337), .B(n20289), .Z(n19781) );
  AND U21881 ( .A(n21338), .B(n21339), .Z(n21337) );
  XNOR U21882 ( .A(n20533), .B(n20008), .Z(n13273) );
  XOR U21883 ( .A(n21340), .B(n21341), .Z(n20008) );
  XOR U21884 ( .A(n21342), .B(n21343), .Z(n20533) );
  ANDN U21885 ( .B(n21344), .A(n21345), .Z(n21342) );
  XOR U21886 ( .A(n21346), .B(n12933), .Z(n11452) );
  XNOR U21887 ( .A(n21347), .B(n19201), .Z(n12933) );
  XOR U21888 ( .A(n21348), .B(n19702), .Z(n19201) );
  XOR U21889 ( .A(n21349), .B(n21350), .Z(n19702) );
  XNOR U21890 ( .A(n20520), .B(n20138), .Z(n21350) );
  XNOR U21891 ( .A(n21351), .B(n20536), .Z(n20138) );
  ANDN U21892 ( .B(n20537), .A(n21352), .Z(n21351) );
  XNOR U21893 ( .A(n21353), .B(n21344), .Z(n20520) );
  XOR U21894 ( .A(n16005), .B(n21355), .Z(n21349) );
  XNOR U21895 ( .A(n18046), .B(n18499), .Z(n21355) );
  XNOR U21896 ( .A(n21356), .B(n20526), .Z(n18499) );
  ANDN U21897 ( .B(n21357), .A(n21358), .Z(n21356) );
  XNOR U21898 ( .A(n21359), .B(n20540), .Z(n18046) );
  XNOR U21899 ( .A(n21361), .B(n20531), .Z(n16005) );
  ANDN U21900 ( .B(n21362), .A(n20530), .Z(n21361) );
  XNOR U21901 ( .A(n20408), .B(n18683), .Z(n13179) );
  XNOR U21902 ( .A(n21363), .B(n21364), .Z(n20374) );
  XOR U21903 ( .A(n19030), .B(n19678), .Z(n21364) );
  XNOR U21904 ( .A(n21365), .B(n21366), .Z(n19678) );
  ANDN U21905 ( .B(n19164), .A(n20413), .Z(n21365) );
  XNOR U21906 ( .A(n21367), .B(n21368), .Z(n19164) );
  XNOR U21907 ( .A(n21369), .B(n21370), .Z(n19030) );
  ANDN U21908 ( .B(n20416), .A(n20415), .Z(n21369) );
  IV U21909 ( .A(n19154), .Z(n20416) );
  XOR U21910 ( .A(n21371), .B(n21372), .Z(n19154) );
  XOR U21911 ( .A(n21373), .B(n21374), .Z(n21363) );
  XNOR U21912 ( .A(n17273), .B(n17193), .Z(n21374) );
  XNOR U21913 ( .A(n21375), .B(n21376), .Z(n17193) );
  ANDN U21914 ( .B(n21377), .A(n21378), .Z(n21375) );
  XOR U21915 ( .A(n21379), .B(n21380), .Z(n17273) );
  XOR U21916 ( .A(n21381), .B(n21382), .Z(n19160) );
  XNOR U21917 ( .A(n21384), .B(n21378), .Z(n20408) );
  NOR U21918 ( .A(n21377), .B(n19151), .Z(n21384) );
  IV U21919 ( .A(n19150), .Z(n21377) );
  XOR U21920 ( .A(n21385), .B(n21386), .Z(n19150) );
  XOR U21921 ( .A(n21387), .B(n18387), .Z(n14969) );
  IV U21922 ( .A(n18890), .Z(n18387) );
  XNOR U21923 ( .A(n21388), .B(n15685), .Z(n14943) );
  XNOR U21924 ( .A(n21389), .B(n18197), .Z(n15685) );
  XNOR U21925 ( .A(n21390), .B(n21391), .Z(n18197) );
  ANDN U21926 ( .B(n14829), .A(n21142), .Z(n21388) );
  XOR U21927 ( .A(n21392), .B(n18813), .Z(n21142) );
  IV U21928 ( .A(n15638), .Z(n18813) );
  XOR U21929 ( .A(n21393), .B(n17244), .Z(n14829) );
  XNOR U21930 ( .A(n21394), .B(n21395), .Z(n17244) );
  XOR U21931 ( .A(n19704), .B(n11925), .Z(n7127) );
  IV U21932 ( .A(n12090), .Z(n11925) );
  XNOR U21933 ( .A(n21396), .B(n21397), .Z(n12366) );
  XOR U21934 ( .A(n12393), .B(n9799), .Z(n21397) );
  XNOR U21935 ( .A(n21398), .B(n15151), .Z(n9799) );
  XOR U21936 ( .A(n20323), .B(n18182), .Z(n15151) );
  IV U21937 ( .A(n17516), .Z(n18182) );
  XOR U21938 ( .A(n21399), .B(n20989), .Z(n17516) );
  XNOR U21939 ( .A(n21400), .B(n21401), .Z(n20989) );
  XNOR U21940 ( .A(n17076), .B(n17688), .Z(n21401) );
  XNOR U21941 ( .A(n21402), .B(n21403), .Z(n17688) );
  ANDN U21942 ( .B(n20993), .A(n20991), .Z(n21402) );
  XOR U21943 ( .A(n21404), .B(n21405), .Z(n17076) );
  ANDN U21944 ( .B(n20345), .A(n21406), .Z(n21404) );
  XNOR U21945 ( .A(n15260), .B(n21407), .Z(n21400) );
  XNOR U21946 ( .A(n19191), .B(n19073), .Z(n21407) );
  XNOR U21947 ( .A(n21408), .B(n21409), .Z(n19073) );
  ANDN U21948 ( .B(n20341), .A(n21410), .Z(n21408) );
  XOR U21949 ( .A(n21411), .B(n21412), .Z(n19191) );
  NOR U21950 ( .A(n20351), .B(n20352), .Z(n21411) );
  XNOR U21951 ( .A(n21413), .B(n21414), .Z(n15260) );
  NOR U21952 ( .A(n20355), .B(n20356), .Z(n21413) );
  XNOR U21953 ( .A(n21415), .B(n21416), .Z(n20323) );
  ANDN U21954 ( .B(n21417), .A(n21418), .Z(n21415) );
  ANDN U21955 ( .B(n15150), .A(n16694), .Z(n21398) );
  XNOR U21956 ( .A(n21419), .B(n16078), .Z(n15150) );
  XNOR U21957 ( .A(n21340), .B(n19180), .Z(n16078) );
  XNOR U21958 ( .A(n21420), .B(n21421), .Z(n19180) );
  XOR U21959 ( .A(n18923), .B(n18057), .Z(n21421) );
  XNOR U21960 ( .A(n21422), .B(n21423), .Z(n18057) );
  NOR U21961 ( .A(n21424), .B(n21425), .Z(n21422) );
  XNOR U21962 ( .A(n21426), .B(n21427), .Z(n18923) );
  NOR U21963 ( .A(n21428), .B(n21429), .Z(n21426) );
  XOR U21964 ( .A(n18864), .B(n21430), .Z(n21420) );
  XOR U21965 ( .A(n21431), .B(n21432), .Z(n21430) );
  XNOR U21966 ( .A(n21433), .B(n21434), .Z(n18864) );
  ANDN U21967 ( .B(n21435), .A(n21436), .Z(n21433) );
  XOR U21968 ( .A(n21437), .B(n21438), .Z(n21340) );
  XNOR U21969 ( .A(n21439), .B(n17873), .Z(n21438) );
  XOR U21970 ( .A(n21440), .B(n21441), .Z(n17873) );
  AND U21971 ( .A(n21442), .B(n20064), .Z(n21440) );
  XOR U21972 ( .A(n20299), .B(n21443), .Z(n21437) );
  XOR U21973 ( .A(n18664), .B(n20129), .Z(n21443) );
  XNOR U21974 ( .A(n21444), .B(n21445), .Z(n20129) );
  AND U21975 ( .A(n21446), .B(n20060), .Z(n21444) );
  XOR U21976 ( .A(n21447), .B(n21448), .Z(n18664) );
  ANDN U21977 ( .B(n21449), .A(n21450), .Z(n21447) );
  XNOR U21978 ( .A(n21451), .B(n21452), .Z(n20299) );
  AND U21979 ( .A(n21453), .B(n21454), .Z(n21451) );
  XNOR U21980 ( .A(n21455), .B(n15160), .Z(n12393) );
  ANDN U21981 ( .B(n16690), .A(n15161), .Z(n21455) );
  XOR U21982 ( .A(n21456), .B(n17592), .Z(n15161) );
  IV U21983 ( .A(n16732), .Z(n17592) );
  XOR U21984 ( .A(n21457), .B(n21458), .Z(n16732) );
  XNOR U21985 ( .A(n15029), .B(n21459), .Z(n21396) );
  XNOR U21986 ( .A(n14615), .B(n9906), .Z(n21459) );
  XNOR U21987 ( .A(n21460), .B(n19479), .Z(n9906) );
  XOR U21988 ( .A(n19624), .B(n16305), .Z(n19479) );
  IV U21989 ( .A(n19841), .Z(n16305) );
  XOR U21990 ( .A(n19793), .B(n21461), .Z(n19841) );
  XNOR U21991 ( .A(n21462), .B(n21463), .Z(n19793) );
  XOR U21992 ( .A(n17228), .B(n20075), .Z(n21463) );
  XNOR U21993 ( .A(n21464), .B(n21465), .Z(n20075) );
  ANDN U21994 ( .B(n19628), .A(n19626), .Z(n21464) );
  XOR U21995 ( .A(n21466), .B(n21101), .Z(n17228) );
  ANDN U21996 ( .B(n19621), .A(n19619), .Z(n21466) );
  XOR U21997 ( .A(n17992), .B(n21467), .Z(n21462) );
  XNOR U21998 ( .A(n18498), .B(n19953), .Z(n21467) );
  XNOR U21999 ( .A(n21468), .B(n21148), .Z(n19953) );
  ANDN U22000 ( .B(n19845), .A(n19843), .Z(n21468) );
  XNOR U22001 ( .A(n21469), .B(n21105), .Z(n18498) );
  IV U22002 ( .A(n21470), .Z(n21105) );
  ANDN U22003 ( .B(n21471), .A(n21472), .Z(n21469) );
  XOR U22004 ( .A(n21473), .B(n21111), .Z(n17992) );
  ANDN U22005 ( .B(n20022), .A(n20023), .Z(n21473) );
  XNOR U22006 ( .A(n21474), .B(n21472), .Z(n19624) );
  NOR U22007 ( .A(n21471), .B(n21104), .Z(n21474) );
  ANDN U22008 ( .B(n16696), .A(n16697), .Z(n21460) );
  XOR U22009 ( .A(n21475), .B(n19769), .Z(n16696) );
  XNOR U22010 ( .A(n21476), .B(n19829), .Z(n19769) );
  XNOR U22011 ( .A(n21477), .B(n21478), .Z(n19829) );
  XNOR U22012 ( .A(n19239), .B(n18506), .Z(n21478) );
  XOR U22013 ( .A(n21479), .B(n21480), .Z(n18506) );
  ANDN U22014 ( .B(n21481), .A(n21482), .Z(n21479) );
  XNOR U22015 ( .A(n21483), .B(n21484), .Z(n19239) );
  NOR U22016 ( .A(n21485), .B(n21486), .Z(n21483) );
  XOR U22017 ( .A(n15350), .B(n21487), .Z(n21477) );
  XOR U22018 ( .A(n18820), .B(n18881), .Z(n21487) );
  XNOR U22019 ( .A(n21488), .B(n21489), .Z(n18881) );
  NOR U22020 ( .A(n21490), .B(n21491), .Z(n21488) );
  XNOR U22021 ( .A(n21492), .B(n21493), .Z(n18820) );
  NOR U22022 ( .A(n21494), .B(n21495), .Z(n21492) );
  XNOR U22023 ( .A(n21496), .B(n21497), .Z(n15350) );
  NOR U22024 ( .A(n21498), .B(n21499), .Z(n21496) );
  XNOR U22025 ( .A(n21500), .B(n15156), .Z(n14615) );
  XOR U22026 ( .A(n21501), .B(n17306), .Z(n15156) );
  ANDN U22027 ( .B(n15157), .A(n16687), .Z(n21500) );
  XOR U22028 ( .A(n21502), .B(n17552), .Z(n15157) );
  IV U22029 ( .A(n17131), .Z(n17552) );
  XNOR U22030 ( .A(n21503), .B(n21504), .Z(n17131) );
  XOR U22031 ( .A(n21505), .B(n19472), .Z(n15029) );
  XNOR U22032 ( .A(n21506), .B(n17654), .Z(n19472) );
  XNOR U22033 ( .A(n21185), .B(n21507), .Z(n17654) );
  XOR U22034 ( .A(n21508), .B(n21509), .Z(n21185) );
  XNOR U22035 ( .A(n18933), .B(n21510), .Z(n21509) );
  XOR U22036 ( .A(n21511), .B(n21512), .Z(n18933) );
  NOR U22037 ( .A(n21513), .B(n21514), .Z(n21511) );
  XOR U22038 ( .A(n18029), .B(n21515), .Z(n21508) );
  XOR U22039 ( .A(n17497), .B(n21516), .Z(n21515) );
  XOR U22040 ( .A(n21517), .B(n21518), .Z(n17497) );
  ANDN U22041 ( .B(n21519), .A(n21520), .Z(n21517) );
  XNOR U22042 ( .A(n21521), .B(n21522), .Z(n18029) );
  AND U22043 ( .A(n21523), .B(n21524), .Z(n21521) );
  ANDN U22044 ( .B(n15147), .A(n16700), .Z(n21505) );
  XOR U22045 ( .A(n21266), .B(n18234), .Z(n15147) );
  XNOR U22046 ( .A(n21525), .B(n21526), .Z(n21266) );
  ANDN U22047 ( .B(n21527), .A(n21528), .Z(n21525) );
  XOR U22048 ( .A(n21529), .B(n21530), .Z(n13869) );
  XOR U22049 ( .A(n9253), .B(n12775), .Z(n21530) );
  XNOR U22050 ( .A(n21531), .B(n14701), .Z(n12775) );
  XOR U22051 ( .A(n21532), .B(n21533), .Z(n14701) );
  ANDN U22052 ( .B(n15139), .A(n17264), .Z(n21531) );
  XOR U22053 ( .A(n21534), .B(n14711), .Z(n9253) );
  XNOR U22054 ( .A(n18706), .B(n21535), .Z(n14711) );
  XNOR U22055 ( .A(n20901), .B(n20997), .Z(n18706) );
  XOR U22056 ( .A(n21536), .B(n21537), .Z(n20997) );
  XNOR U22057 ( .A(n21538), .B(n17513), .Z(n21537) );
  XNOR U22058 ( .A(n21539), .B(n21540), .Z(n17513) );
  ANDN U22059 ( .B(n21541), .A(n21542), .Z(n21539) );
  XOR U22060 ( .A(n18421), .B(n21543), .Z(n21536) );
  XNOR U22061 ( .A(n18583), .B(n17693), .Z(n21543) );
  XNOR U22062 ( .A(n21544), .B(n21545), .Z(n17693) );
  ANDN U22063 ( .B(n21546), .A(n21547), .Z(n21544) );
  XNOR U22064 ( .A(n21548), .B(n21549), .Z(n18583) );
  AND U22065 ( .A(n21550), .B(n21551), .Z(n21548) );
  XNOR U22066 ( .A(n21552), .B(n21275), .Z(n18421) );
  IV U22067 ( .A(n21553), .Z(n21275) );
  XOR U22068 ( .A(n21556), .B(n21557), .Z(n20901) );
  XNOR U22069 ( .A(n20191), .B(n18906), .Z(n21557) );
  XNOR U22070 ( .A(n21558), .B(n21559), .Z(n18906) );
  ANDN U22071 ( .B(n21560), .A(n21561), .Z(n21558) );
  XOR U22072 ( .A(n21562), .B(n21563), .Z(n20191) );
  XOR U22073 ( .A(n19119), .B(n21566), .Z(n21556) );
  XNOR U22074 ( .A(n18803), .B(n19106), .Z(n21566) );
  XOR U22075 ( .A(n21567), .B(n21568), .Z(n19106) );
  XOR U22076 ( .A(n21571), .B(n21572), .Z(n18803) );
  ANDN U22077 ( .B(n21573), .A(n21574), .Z(n21571) );
  XNOR U22078 ( .A(n21575), .B(n21576), .Z(n19119) );
  ANDN U22079 ( .B(n21577), .A(n21578), .Z(n21575) );
  ANDN U22080 ( .B(n15130), .A(n17259), .Z(n21534) );
  XNOR U22081 ( .A(n21579), .B(n18473), .Z(n17259) );
  IV U22082 ( .A(n18442), .Z(n18473) );
  XNOR U22083 ( .A(n21580), .B(n21581), .Z(n20226) );
  XOR U22084 ( .A(n18765), .B(n19049), .Z(n21581) );
  XOR U22085 ( .A(n21582), .B(n19862), .Z(n19049) );
  XOR U22086 ( .A(n21585), .B(n21586), .Z(n20000) );
  XOR U22087 ( .A(n21587), .B(n21588), .Z(n18765) );
  NOR U22088 ( .A(n20003), .B(n20401), .Z(n21587) );
  XNOR U22089 ( .A(n21589), .B(n21590), .Z(n20003) );
  XOR U22090 ( .A(n18677), .B(n21591), .Z(n21580) );
  XOR U22091 ( .A(n19851), .B(n19672), .Z(n21591) );
  XNOR U22092 ( .A(n21592), .B(n19858), .Z(n19672) );
  ANDN U22093 ( .B(n19995), .A(n19857), .Z(n21592) );
  IV U22094 ( .A(n20396), .Z(n19857) );
  XNOR U22095 ( .A(n21593), .B(n21594), .Z(n20396) );
  XOR U22096 ( .A(n21595), .B(n21596), .Z(n19995) );
  XOR U22097 ( .A(n21597), .B(n19871), .Z(n19851) );
  ANDN U22098 ( .B(n19872), .A(n20126), .Z(n21597) );
  XOR U22099 ( .A(n21598), .B(n21599), .Z(n20126) );
  XOR U22100 ( .A(n21600), .B(n21601), .Z(n19872) );
  XNOR U22101 ( .A(n21602), .B(n19868), .Z(n18677) );
  ANDN U22102 ( .B(n19992), .A(n19867), .Z(n21602) );
  XOR U22103 ( .A(n21603), .B(n21604), .Z(n19867) );
  XOR U22104 ( .A(n21605), .B(n21606), .Z(n19992) );
  XOR U22105 ( .A(n21607), .B(n21608), .Z(n20086) );
  XNOR U22106 ( .A(n17198), .B(n19235), .Z(n21608) );
  XNOR U22107 ( .A(n21609), .B(n20585), .Z(n19235) );
  XOR U22108 ( .A(n21611), .B(n20589), .Z(n17198) );
  XOR U22109 ( .A(n17536), .B(n21613), .Z(n21607) );
  XNOR U22110 ( .A(n19425), .B(n17067), .Z(n21613) );
  XNOR U22111 ( .A(n21614), .B(n21615), .Z(n17067) );
  AND U22112 ( .A(n21616), .B(n21617), .Z(n21614) );
  XOR U22113 ( .A(n21618), .B(n20580), .Z(n19425) );
  NOR U22114 ( .A(n21619), .B(n20579), .Z(n21618) );
  XNOR U22115 ( .A(n21620), .B(n20576), .Z(n17536) );
  ANDN U22116 ( .B(n21621), .A(n20575), .Z(n21620) );
  XOR U22117 ( .A(n19399), .B(n21622), .Z(n15130) );
  XOR U22118 ( .A(n15126), .B(n21623), .Z(n21529) );
  XNOR U22119 ( .A(n9454), .B(n12668), .Z(n21623) );
  XOR U22120 ( .A(n21624), .B(n14698), .Z(n12668) );
  XOR U22121 ( .A(n21625), .B(n18777), .Z(n14698) );
  XNOR U22122 ( .A(n19458), .B(n20006), .Z(n18777) );
  XNOR U22123 ( .A(n21626), .B(n21627), .Z(n20006) );
  XNOR U22124 ( .A(n21628), .B(n19663), .Z(n21627) );
  XNOR U22125 ( .A(n21629), .B(n20235), .Z(n19663) );
  ANDN U22126 ( .B(n21630), .A(n21631), .Z(n21629) );
  XOR U22127 ( .A(n19363), .B(n21632), .Z(n21626) );
  XOR U22128 ( .A(n20593), .B(n19324), .Z(n21632) );
  XNOR U22129 ( .A(n21633), .B(n20245), .Z(n19324) );
  NOR U22130 ( .A(n21634), .B(n21635), .Z(n21633) );
  XOR U22131 ( .A(n21636), .B(n20242), .Z(n20593) );
  ANDN U22132 ( .B(n21637), .A(n21638), .Z(n21636) );
  XNOR U22133 ( .A(n21639), .B(n20231), .Z(n19363) );
  ANDN U22134 ( .B(n21640), .A(n21641), .Z(n21639) );
  XOR U22135 ( .A(n21642), .B(n21643), .Z(n19458) );
  XNOR U22136 ( .A(n15876), .B(n19242), .Z(n21643) );
  XNOR U22137 ( .A(n21644), .B(n21645), .Z(n19242) );
  ANDN U22138 ( .B(n21646), .A(n21647), .Z(n21644) );
  XNOR U22139 ( .A(n21648), .B(n21649), .Z(n15876) );
  NOR U22140 ( .A(n21650), .B(n21651), .Z(n21648) );
  XNOR U22141 ( .A(n17935), .B(n21652), .Z(n21642) );
  XOR U22142 ( .A(n19309), .B(n18515), .Z(n21652) );
  XOR U22143 ( .A(n21653), .B(n21654), .Z(n18515) );
  ANDN U22144 ( .B(n21655), .A(n21656), .Z(n21653) );
  XNOR U22145 ( .A(n21657), .B(n21658), .Z(n19309) );
  ANDN U22146 ( .B(n21659), .A(n21660), .Z(n21657) );
  XNOR U22147 ( .A(n21661), .B(n21662), .Z(n17935) );
  ANDN U22148 ( .B(n21663), .A(n21664), .Z(n21661) );
  NOR U22149 ( .A(n15137), .B(n17267), .Z(n21624) );
  XNOR U22150 ( .A(n21665), .B(n16998), .Z(n17267) );
  XNOR U22151 ( .A(n21667), .B(n21668), .Z(n21458) );
  XNOR U22152 ( .A(n18475), .B(n20864), .Z(n21668) );
  XNOR U22153 ( .A(n21669), .B(n20881), .Z(n20864) );
  NOR U22154 ( .A(n20882), .B(n21670), .Z(n21669) );
  XNOR U22155 ( .A(n21671), .B(n21672), .Z(n18475) );
  ANDN U22156 ( .B(n21673), .A(n21674), .Z(n21671) );
  XOR U22157 ( .A(n20634), .B(n21675), .Z(n21667) );
  XOR U22158 ( .A(n19302), .B(n17288), .Z(n21675) );
  XOR U22159 ( .A(n21676), .B(n20877), .Z(n17288) );
  ANDN U22160 ( .B(n20878), .A(n21677), .Z(n21676) );
  XOR U22161 ( .A(n21678), .B(n21679), .Z(n19302) );
  NOR U22162 ( .A(n21680), .B(n21681), .Z(n21678) );
  XOR U22163 ( .A(n21682), .B(n20871), .Z(n20634) );
  NOR U22164 ( .A(n21683), .B(n21684), .Z(n21682) );
  XOR U22165 ( .A(n21685), .B(n16852), .Z(n15137) );
  XNOR U22166 ( .A(n14707), .B(n21686), .Z(n9454) );
  XOR U22167 ( .A(n21687), .B(n21688), .Z(n21686) );
  XOR U22168 ( .A(n19525), .B(n18195), .Z(n17256) );
  XNOR U22169 ( .A(n21476), .B(n20140), .Z(n18195) );
  XOR U22170 ( .A(n21689), .B(n21690), .Z(n20140) );
  XNOR U22171 ( .A(n18788), .B(n20195), .Z(n21690) );
  XOR U22172 ( .A(n21691), .B(n20336), .Z(n20195) );
  ANDN U22173 ( .B(n21692), .A(n20337), .Z(n21691) );
  XNOR U22174 ( .A(n21693), .B(n20327), .Z(n18788) );
  ANDN U22175 ( .B(n21694), .A(n20326), .Z(n21693) );
  XOR U22176 ( .A(n17571), .B(n21695), .Z(n21689) );
  XOR U22177 ( .A(n20037), .B(n20320), .Z(n21695) );
  XOR U22178 ( .A(n21696), .B(n20332), .Z(n20320) );
  ANDN U22179 ( .B(n20333), .A(n21697), .Z(n21696) );
  XNOR U22180 ( .A(n21698), .B(n21417), .Z(n20037) );
  XNOR U22181 ( .A(n21700), .B(n20842), .Z(n17571) );
  IV U22182 ( .A(n21701), .Z(n20842) );
  ANDN U22183 ( .B(n21702), .A(n21703), .Z(n21700) );
  XOR U22184 ( .A(n21704), .B(n21705), .Z(n21476) );
  XNOR U22185 ( .A(n19588), .B(n16845), .Z(n21705) );
  XOR U22186 ( .A(n21706), .B(n21339), .Z(n16845) );
  ANDN U22187 ( .B(n20287), .A(n21338), .Z(n21706) );
  XNOR U22188 ( .A(n21707), .B(n21708), .Z(n19588) );
  ANDN U22189 ( .B(n19539), .A(n19537), .Z(n21707) );
  XOR U22190 ( .A(n21709), .B(n21710), .Z(n19539) );
  XOR U22191 ( .A(n19775), .B(n21711), .Z(n21704) );
  XOR U22192 ( .A(n18019), .B(n19694), .Z(n21711) );
  XOR U22193 ( .A(n21712), .B(n20698), .Z(n19694) );
  ANDN U22194 ( .B(n20291), .A(n20699), .Z(n21712) );
  XOR U22195 ( .A(n21713), .B(n21714), .Z(n20699) );
  XNOR U22196 ( .A(n21715), .B(n21716), .Z(n20291) );
  XOR U22197 ( .A(n21717), .B(n19786), .Z(n18019) );
  ANDN U22198 ( .B(n19529), .A(n19527), .Z(n21717) );
  XOR U22199 ( .A(n21718), .B(n21719), .Z(n19527) );
  XOR U22200 ( .A(n21720), .B(n21721), .Z(n19529) );
  XOR U22201 ( .A(n21722), .B(n21723), .Z(n19775) );
  ANDN U22202 ( .B(n19535), .A(n19533), .Z(n21722) );
  XOR U22203 ( .A(n21724), .B(n21725), .Z(n19535) );
  XNOR U22204 ( .A(n21726), .B(n21338), .Z(n19525) );
  XOR U22205 ( .A(n21727), .B(n21728), .Z(n21338) );
  NOR U22206 ( .A(n20288), .B(n20287), .Z(n21726) );
  XOR U22207 ( .A(n21729), .B(n21730), .Z(n20287) );
  XOR U22208 ( .A(n21731), .B(n16409), .Z(n15141) );
  IV U22209 ( .A(n18828), .Z(n16409) );
  XOR U22210 ( .A(n21732), .B(n18186), .Z(n14707) );
  XOR U22211 ( .A(n21733), .B(n21734), .Z(n18186) );
  XNOR U22212 ( .A(n21735), .B(n15134), .Z(n15126) );
  XNOR U22213 ( .A(n17145), .B(n21736), .Z(n15134) );
  IV U22214 ( .A(n17472), .Z(n17145) );
  XOR U22215 ( .A(n19014), .B(n20476), .Z(n17472) );
  XOR U22216 ( .A(n21737), .B(n21738), .Z(n20476) );
  XNOR U22217 ( .A(n17989), .B(n18319), .Z(n21738) );
  XOR U22218 ( .A(n21739), .B(n21651), .Z(n18319) );
  ANDN U22219 ( .B(n21740), .A(n21741), .Z(n21739) );
  XNOR U22220 ( .A(n21742), .B(n21656), .Z(n17989) );
  AND U22221 ( .A(n21743), .B(n21744), .Z(n21742) );
  XOR U22222 ( .A(n15338), .B(n21745), .Z(n21737) );
  XOR U22223 ( .A(n21746), .B(n16989), .Z(n21745) );
  XNOR U22224 ( .A(n21747), .B(n21646), .Z(n16989) );
  ANDN U22225 ( .B(n21748), .A(n21749), .Z(n21747) );
  XNOR U22226 ( .A(n21750), .B(n21659), .Z(n15338) );
  AND U22227 ( .A(n21751), .B(n21752), .Z(n21750) );
  XOR U22228 ( .A(n21753), .B(n21754), .Z(n19014) );
  XNOR U22229 ( .A(n16673), .B(n17895), .Z(n21754) );
  XOR U22230 ( .A(n21755), .B(n21756), .Z(n17895) );
  ANDN U22231 ( .B(n21757), .A(n21758), .Z(n21755) );
  XNOR U22232 ( .A(n21759), .B(n21760), .Z(n16673) );
  XOR U22233 ( .A(n21763), .B(n21764), .Z(n21753) );
  XOR U22234 ( .A(n18369), .B(n16883), .Z(n21764) );
  XNOR U22235 ( .A(n21765), .B(n21766), .Z(n16883) );
  ANDN U22236 ( .B(n21767), .A(n21768), .Z(n21765) );
  ANDN U22237 ( .B(n21771), .A(n21772), .Z(n21769) );
  IV U22238 ( .A(n21773), .Z(n21772) );
  AND U22239 ( .A(n15133), .B(n17271), .Z(n21735) );
  XNOR U22240 ( .A(n21774), .B(n19456), .Z(n17271) );
  IV U22241 ( .A(n17750), .Z(n19456) );
  XNOR U22242 ( .A(n21775), .B(n21776), .Z(n20602) );
  XOR U22243 ( .A(n19489), .B(n20135), .Z(n21776) );
  XNOR U22244 ( .A(n21777), .B(n21514), .Z(n20135) );
  AND U22245 ( .A(n21778), .B(n21779), .Z(n21777) );
  XNOR U22246 ( .A(n21780), .B(n21781), .Z(n19489) );
  ANDN U22247 ( .B(n21782), .A(n21783), .Z(n21780) );
  XOR U22248 ( .A(n20247), .B(n21784), .Z(n21775) );
  XOR U22249 ( .A(n17745), .B(n16524), .Z(n21784) );
  XNOR U22250 ( .A(n21785), .B(n21520), .Z(n16524) );
  ANDN U22251 ( .B(n21786), .A(n21787), .Z(n21785) );
  XOR U22252 ( .A(n21788), .B(n21524), .Z(n17745) );
  ANDN U22253 ( .B(n21789), .A(n21790), .Z(n21788) );
  XOR U22254 ( .A(n21791), .B(n21792), .Z(n20247) );
  XNOR U22255 ( .A(n21795), .B(n21796), .Z(n20902) );
  XNOR U22256 ( .A(n18593), .B(n17086), .Z(n21796) );
  XNOR U22257 ( .A(n21797), .B(n21798), .Z(n17086) );
  AND U22258 ( .A(n21799), .B(n21800), .Z(n21797) );
  XNOR U22259 ( .A(n21801), .B(n21802), .Z(n18593) );
  AND U22260 ( .A(n21803), .B(n20611), .Z(n21801) );
  XNOR U22261 ( .A(n21804), .B(n21805), .Z(n21795) );
  XNOR U22262 ( .A(n15955), .B(n17525), .Z(n21805) );
  XOR U22263 ( .A(n21806), .B(n21807), .Z(n17525) );
  XNOR U22264 ( .A(n21809), .B(n21810), .Z(n15955) );
  ANDN U22265 ( .B(n21811), .A(n20615), .Z(n21809) );
  XOR U22266 ( .A(n21812), .B(n15635), .Z(n15133) );
  XOR U22267 ( .A(n21814), .B(n21815), .Z(n21341) );
  XOR U22268 ( .A(n18705), .B(n18002), .Z(n21815) );
  XNOR U22269 ( .A(n21816), .B(n21817), .Z(n18002) );
  ANDN U22270 ( .B(n20525), .A(n20526), .Z(n21816) );
  XNOR U22271 ( .A(n21818), .B(n21819), .Z(n20526) );
  XNOR U22272 ( .A(n21820), .B(n21821), .Z(n18705) );
  NOR U22273 ( .A(n20529), .B(n20531), .Z(n21820) );
  XNOR U22274 ( .A(n21822), .B(n21823), .Z(n20531) );
  XNOR U22275 ( .A(n19026), .B(n21824), .Z(n21814) );
  XOR U22276 ( .A(n17743), .B(n21825), .Z(n21824) );
  XNOR U22277 ( .A(n21826), .B(n21827), .Z(n17743) );
  NOR U22278 ( .A(n20536), .B(n20535), .Z(n21826) );
  XNOR U22279 ( .A(n21828), .B(n21829), .Z(n20536) );
  XNOR U22280 ( .A(n21830), .B(n21831), .Z(n19026) );
  ANDN U22281 ( .B(n20539), .A(n20540), .Z(n21830) );
  XOR U22282 ( .A(n21832), .B(n21833), .Z(n20540) );
  XNOR U22283 ( .A(n21834), .B(n15139), .Z(n19704) );
  XOR U22284 ( .A(n20508), .B(n18295), .Z(n15139) );
  IV U22285 ( .A(n18855), .Z(n18295) );
  XNOR U22286 ( .A(n19982), .B(n21835), .Z(n18855) );
  XOR U22287 ( .A(n21836), .B(n21837), .Z(n19982) );
  XOR U22288 ( .A(n19770), .B(n17019), .Z(n21837) );
  XNOR U22289 ( .A(n21838), .B(n21839), .Z(n17019) );
  ANDN U22290 ( .B(n21297), .A(n21840), .Z(n21838) );
  XNOR U22291 ( .A(n21841), .B(n21842), .Z(n19770) );
  ANDN U22292 ( .B(n21843), .A(n21300), .Z(n21841) );
  XOR U22293 ( .A(n19382), .B(n21844), .Z(n21836) );
  XOR U22294 ( .A(n18941), .B(n20384), .Z(n21844) );
  XNOR U22295 ( .A(n21845), .B(n21290), .Z(n20384) );
  NOR U22296 ( .A(n21846), .B(n21291), .Z(n21845) );
  XOR U22297 ( .A(n21847), .B(n21286), .Z(n18941) );
  ANDN U22298 ( .B(n21287), .A(n21848), .Z(n21847) );
  XNOR U22299 ( .A(n21849), .B(n21850), .Z(n19382) );
  ANDN U22300 ( .B(n21851), .A(n21852), .Z(n21849) );
  XNOR U22301 ( .A(n21853), .B(n21854), .Z(n20508) );
  NOR U22302 ( .A(n19416), .B(n21855), .Z(n21853) );
  ANDN U22303 ( .B(n17264), .A(n14700), .Z(n21834) );
  XOR U22304 ( .A(n18016), .B(n21856), .Z(n14700) );
  IV U22305 ( .A(n20154), .Z(n18016) );
  XNOR U22306 ( .A(n19652), .B(n20076), .Z(n20154) );
  XOR U22307 ( .A(n21857), .B(n21858), .Z(n20076) );
  XNOR U22308 ( .A(n19262), .B(n21859), .Z(n21858) );
  XNOR U22309 ( .A(n21860), .B(n21861), .Z(n19262) );
  ANDN U22310 ( .B(n21862), .A(n21863), .Z(n21860) );
  XOR U22311 ( .A(n18702), .B(n21864), .Z(n21857) );
  XOR U22312 ( .A(n18455), .B(n21865), .Z(n21864) );
  XNOR U22313 ( .A(n21866), .B(n21867), .Z(n18455) );
  XOR U22314 ( .A(n21870), .B(n21871), .Z(n18702) );
  NOR U22315 ( .A(n21872), .B(n21873), .Z(n21870) );
  XOR U22316 ( .A(n21874), .B(n21875), .Z(n19652) );
  XNOR U22317 ( .A(n16856), .B(n14953), .Z(n21875) );
  XNOR U22318 ( .A(n21876), .B(n21486), .Z(n14953) );
  NOR U22319 ( .A(n21877), .B(n21878), .Z(n21876) );
  XNOR U22320 ( .A(n21879), .B(n21490), .Z(n16856) );
  IV U22321 ( .A(n21880), .Z(n21490) );
  NOR U22322 ( .A(n21881), .B(n21882), .Z(n21879) );
  XNOR U22323 ( .A(n16377), .B(n21883), .Z(n21874) );
  XOR U22324 ( .A(n18025), .B(n19521), .Z(n21883) );
  XNOR U22325 ( .A(n21884), .B(n21495), .Z(n19521) );
  NOR U22326 ( .A(n21885), .B(n21886), .Z(n21884) );
  XOR U22327 ( .A(n21887), .B(n21481), .Z(n18025) );
  ANDN U22328 ( .B(n21888), .A(n21889), .Z(n21887) );
  XNOR U22329 ( .A(n21890), .B(n21499), .Z(n16377) );
  NOR U22330 ( .A(n21891), .B(n21892), .Z(n21890) );
  XNOR U22331 ( .A(n21893), .B(n17626), .Z(n17264) );
  XNOR U22332 ( .A(n21894), .B(n21895), .Z(n17626) );
  XOR U22333 ( .A(n21896), .B(n9330), .Z(n3531) );
  IV U22334 ( .A(n6682), .Z(n9330) );
  XNOR U22335 ( .A(n14121), .B(n10108), .Z(n6682) );
  XNOR U22336 ( .A(n12920), .B(n16884), .Z(n10108) );
  XNOR U22337 ( .A(n21897), .B(n21898), .Z(n16884) );
  XNOR U22338 ( .A(n10225), .B(n10929), .Z(n21898) );
  XOR U22339 ( .A(n21899), .B(n17830), .Z(n10929) );
  XOR U22340 ( .A(n21900), .B(n21023), .Z(n17830) );
  XNOR U22341 ( .A(n21901), .B(n21182), .Z(n21023) );
  NOR U22342 ( .A(n15098), .B(n15099), .Z(n21899) );
  XOR U22343 ( .A(n21904), .B(n15638), .Z(n15099) );
  XNOR U22344 ( .A(n21905), .B(n18984), .Z(n15638) );
  XNOR U22345 ( .A(n21906), .B(n21907), .Z(n18984) );
  XNOR U22346 ( .A(n19365), .B(n18876), .Z(n21907) );
  XNOR U22347 ( .A(n21908), .B(n21909), .Z(n18876) );
  ANDN U22348 ( .B(n21910), .A(n21911), .Z(n21908) );
  XNOR U22349 ( .A(n21912), .B(n21913), .Z(n19365) );
  ANDN U22350 ( .B(n21914), .A(n21915), .Z(n21912) );
  XOR U22351 ( .A(n17226), .B(n21916), .Z(n21906) );
  XNOR U22352 ( .A(n19496), .B(n21917), .Z(n21916) );
  XNOR U22353 ( .A(n21918), .B(n21919), .Z(n19496) );
  NOR U22354 ( .A(n21920), .B(n21921), .Z(n21918) );
  XNOR U22355 ( .A(n21922), .B(n21923), .Z(n17226) );
  IV U22356 ( .A(n17891), .Z(n15098) );
  XOR U22357 ( .A(n21926), .B(n17574), .Z(n17891) );
  XNOR U22358 ( .A(n17816), .B(n21927), .Z(n10225) );
  XOR U22359 ( .A(n21928), .B(n21688), .Z(n21927) );
  ANDN U22360 ( .B(n14118), .A(n14119), .Z(n21928) );
  XNOR U22361 ( .A(n21325), .B(n17105), .Z(n14119) );
  XNOR U22362 ( .A(n21929), .B(n20661), .Z(n21325) );
  ANDN U22363 ( .B(n20977), .A(n20976), .Z(n21929) );
  XOR U22364 ( .A(n21930), .B(n18051), .Z(n14118) );
  IV U22365 ( .A(n17977), .Z(n18051) );
  XNOR U22366 ( .A(n19138), .B(n20962), .Z(n17977) );
  XOR U22367 ( .A(n21931), .B(n21932), .Z(n20962) );
  XNOR U22368 ( .A(n20257), .B(n16766), .Z(n21932) );
  ANDN U22369 ( .B(n21934), .A(n20263), .Z(n21933) );
  XNOR U22370 ( .A(n21935), .B(n20275), .Z(n20257) );
  ANDN U22371 ( .B(n21936), .A(n20274), .Z(n21935) );
  XOR U22372 ( .A(n18006), .B(n21937), .Z(n21931) );
  XOR U22373 ( .A(n18821), .B(n18271), .Z(n21937) );
  XNOR U22374 ( .A(n21938), .B(n21939), .Z(n18271) );
  XNOR U22375 ( .A(n21942), .B(n20267), .Z(n18821) );
  ANDN U22376 ( .B(n20268), .A(n21943), .Z(n21942) );
  IV U22377 ( .A(n21944), .Z(n20268) );
  XNOR U22378 ( .A(n21945), .B(n21946), .Z(n18006) );
  NOR U22379 ( .A(n21947), .B(n21948), .Z(n21945) );
  XOR U22380 ( .A(n21949), .B(n21950), .Z(n19138) );
  XNOR U22381 ( .A(n15675), .B(n17290), .Z(n21950) );
  XNOR U22382 ( .A(n21951), .B(n21952), .Z(n17290) );
  NOR U22383 ( .A(n21953), .B(n21954), .Z(n21951) );
  XNOR U22384 ( .A(n21955), .B(n21956), .Z(n15675) );
  NOR U22385 ( .A(n21957), .B(n21958), .Z(n21955) );
  XOR U22386 ( .A(n21959), .B(n21960), .Z(n21949) );
  XNOR U22387 ( .A(n19313), .B(n18584), .Z(n21960) );
  XNOR U22388 ( .A(n21961), .B(n21962), .Z(n18584) );
  ANDN U22389 ( .B(n21963), .A(n21964), .Z(n21961) );
  XOR U22390 ( .A(n21965), .B(n21966), .Z(n19313) );
  NOR U22391 ( .A(n21967), .B(n21968), .Z(n21965) );
  XOR U22392 ( .A(n20733), .B(n19374), .Z(n17816) );
  XNOR U22393 ( .A(n21969), .B(n21970), .Z(n20733) );
  XNOR U22394 ( .A(n4549), .B(n21971), .Z(n21970) );
  NANDN U22395 ( .A(n21972), .B(n20562), .Z(n21971) );
  XOR U22396 ( .A(n17876), .B(n21973), .Z(n21897) );
  XOR U22397 ( .A(n12688), .B(n10398), .Z(n21973) );
  XOR U22398 ( .A(n21974), .B(n17827), .Z(n10398) );
  XNOR U22399 ( .A(n21976), .B(n21977), .Z(n20910) );
  XOR U22400 ( .A(n17308), .B(n20632), .Z(n21977) );
  XNOR U22401 ( .A(n21978), .B(n21019), .Z(n20632) );
  ANDN U22402 ( .B(n21979), .A(n21980), .Z(n21978) );
  XNOR U22403 ( .A(n21981), .B(n21012), .Z(n17308) );
  ANDN U22404 ( .B(n21982), .A(n21983), .Z(n21981) );
  XNOR U22405 ( .A(n16595), .B(n21984), .Z(n21976) );
  XOR U22406 ( .A(n21985), .B(n16588), .Z(n21984) );
  XOR U22407 ( .A(n21986), .B(n21987), .Z(n16588) );
  ANDN U22408 ( .B(n21988), .A(n21989), .Z(n21986) );
  XNOR U22409 ( .A(n21990), .B(n21009), .Z(n16595) );
  ANDN U22410 ( .B(n21991), .A(n21992), .Z(n21990) );
  XNOR U22411 ( .A(n21993), .B(n21994), .Z(n19336) );
  XNOR U22412 ( .A(n17469), .B(n21685), .Z(n21994) );
  XOR U22413 ( .A(n21995), .B(n21037), .Z(n21685) );
  NOR U22414 ( .A(n21177), .B(n21178), .Z(n21995) );
  XNOR U22415 ( .A(n21996), .B(n21903), .Z(n17469) );
  NOR U22416 ( .A(n21181), .B(n21180), .Z(n21996) );
  XOR U22417 ( .A(n16851), .B(n21997), .Z(n21993) );
  XOR U22418 ( .A(n17561), .B(n21998), .Z(n21997) );
  XNOR U22419 ( .A(n21999), .B(n22000), .Z(n17561) );
  NOR U22420 ( .A(n21165), .B(n21166), .Z(n21999) );
  XNOR U22421 ( .A(n22001), .B(n21033), .Z(n16851) );
  ANDN U22422 ( .B(n21169), .A(n21170), .Z(n22001) );
  ANDN U22423 ( .B(n14258), .A(n14256), .Z(n21974) );
  IV U22424 ( .A(n17880), .Z(n14256) );
  XOR U22425 ( .A(n22002), .B(n19751), .Z(n17880) );
  XOR U22426 ( .A(n22003), .B(n19048), .Z(n19751) );
  XNOR U22427 ( .A(n22004), .B(n22005), .Z(n19048) );
  XOR U22428 ( .A(n18308), .B(n19056), .Z(n22005) );
  XOR U22429 ( .A(n22006), .B(n20333), .Z(n19056) );
  XOR U22430 ( .A(n22007), .B(n22008), .Z(n20333) );
  ANDN U22431 ( .B(n21697), .A(n22009), .Z(n22006) );
  XNOR U22432 ( .A(n22010), .B(n20326), .Z(n18308) );
  XOR U22433 ( .A(n22011), .B(n22012), .Z(n20326) );
  ANDN U22434 ( .B(n22013), .A(n21694), .Z(n22010) );
  XOR U22435 ( .A(n20139), .B(n22014), .Z(n22004) );
  XNOR U22436 ( .A(n19368), .B(n19097), .Z(n22014) );
  XOR U22437 ( .A(n22015), .B(n21418), .Z(n19097) );
  XOR U22438 ( .A(n22016), .B(n22017), .Z(n21418) );
  ANDN U22439 ( .B(n22018), .A(n21699), .Z(n22015) );
  XNOR U22440 ( .A(n22019), .B(n20337), .Z(n19368) );
  XOR U22441 ( .A(n22020), .B(n22021), .Z(n20337) );
  ANDN U22442 ( .B(n22022), .A(n21692), .Z(n22019) );
  XNOR U22443 ( .A(n22023), .B(n21703), .Z(n20139) );
  IV U22444 ( .A(n20843), .Z(n21703) );
  XOR U22445 ( .A(n22024), .B(n22025), .Z(n20843) );
  NOR U22446 ( .A(n22026), .B(n21702), .Z(n22023) );
  XOR U22447 ( .A(n20302), .B(n21247), .Z(n14258) );
  XOR U22448 ( .A(n22027), .B(n22028), .Z(n21247) );
  ANDN U22449 ( .B(n20680), .A(n22029), .Z(n22027) );
  XOR U22450 ( .A(n22030), .B(n22031), .Z(n20302) );
  XOR U22451 ( .A(n22032), .B(n17824), .Z(n12688) );
  XNOR U22452 ( .A(n19399), .B(n22033), .Z(n17824) );
  NOR U22453 ( .A(n18649), .B(n18546), .Z(n22032) );
  XNOR U22454 ( .A(n19395), .B(n22034), .Z(n18546) );
  IV U22455 ( .A(n15694), .Z(n19395) );
  XNOR U22456 ( .A(n22035), .B(n22036), .Z(n20884) );
  XNOR U22457 ( .A(n17239), .B(n17401), .Z(n22036) );
  XNOR U22458 ( .A(n22037), .B(n22038), .Z(n17401) );
  ANDN U22459 ( .B(n22039), .A(n22040), .Z(n22037) );
  XNOR U22460 ( .A(n22041), .B(n22042), .Z(n17239) );
  ANDN U22461 ( .B(n22043), .A(n22044), .Z(n22041) );
  XNOR U22462 ( .A(n18213), .B(n22045), .Z(n22035) );
  XOR U22463 ( .A(n18347), .B(n18666), .Z(n22045) );
  XOR U22464 ( .A(n22046), .B(n22047), .Z(n18666) );
  XNOR U22465 ( .A(n22050), .B(n22051), .Z(n18347) );
  XOR U22466 ( .A(n22054), .B(n22055), .Z(n18213) );
  XOR U22467 ( .A(n22058), .B(n22059), .Z(n21256) );
  XNOR U22468 ( .A(n14163), .B(n19448), .Z(n22059) );
  XNOR U22469 ( .A(n22060), .B(n22061), .Z(n19448) );
  ANDN U22470 ( .B(n22062), .A(n22063), .Z(n22060) );
  XOR U22471 ( .A(n22064), .B(n22065), .Z(n14163) );
  ANDN U22472 ( .B(n22066), .A(n22067), .Z(n22064) );
  XOR U22473 ( .A(n19211), .B(n22068), .Z(n22058) );
  XOR U22474 ( .A(n19296), .B(n22069), .Z(n22068) );
  XOR U22475 ( .A(n22070), .B(n22071), .Z(n19296) );
  ANDN U22476 ( .B(n22072), .A(n22073), .Z(n22070) );
  XOR U22477 ( .A(n22074), .B(n22075), .Z(n19211) );
  ANDN U22478 ( .B(n22076), .A(n22077), .Z(n22074) );
  XNOR U22479 ( .A(n22078), .B(n16889), .Z(n18649) );
  XOR U22480 ( .A(n22079), .B(n21733), .Z(n16889) );
  XNOR U22481 ( .A(n22080), .B(n22081), .Z(n21733) );
  XOR U22482 ( .A(n16578), .B(n18533), .Z(n22081) );
  XNOR U22483 ( .A(n22082), .B(n19573), .Z(n18533) );
  NOR U22484 ( .A(n22083), .B(n22084), .Z(n22082) );
  XNOR U22485 ( .A(n22085), .B(n22086), .Z(n16578) );
  NOR U22486 ( .A(n22087), .B(n20029), .Z(n22085) );
  XOR U22487 ( .A(n20996), .B(n22088), .Z(n22080) );
  XOR U22488 ( .A(n17964), .B(n17799), .Z(n22088) );
  XNOR U22489 ( .A(n22089), .B(n19581), .Z(n17799) );
  NOR U22490 ( .A(n22090), .B(n20069), .Z(n22089) );
  XNOR U22491 ( .A(n22091), .B(n22092), .Z(n17964) );
  NOR U22492 ( .A(n22093), .B(n22094), .Z(n22091) );
  XNOR U22493 ( .A(n22095), .B(n19568), .Z(n20996) );
  NOR U22494 ( .A(n22096), .B(n19687), .Z(n22095) );
  XNOR U22495 ( .A(n22097), .B(n17884), .Z(n17876) );
  XOR U22496 ( .A(n22098), .B(n17835), .Z(n17884) );
  XNOR U22497 ( .A(n19711), .B(n18983), .Z(n17835) );
  XNOR U22498 ( .A(n22099), .B(n22100), .Z(n18983) );
  XNOR U22499 ( .A(n17629), .B(n19642), .Z(n22100) );
  XOR U22500 ( .A(n22101), .B(n21681), .Z(n19642) );
  ANDN U22501 ( .B(n22102), .A(n22103), .Z(n22101) );
  XNOR U22502 ( .A(n22104), .B(n21684), .Z(n17629) );
  ANDN U22503 ( .B(n20870), .A(n22105), .Z(n22104) );
  XOR U22504 ( .A(n18644), .B(n22106), .Z(n22099) );
  XNOR U22505 ( .A(n22107), .B(n19961), .Z(n22106) );
  XNOR U22506 ( .A(n22108), .B(n21677), .Z(n19961) );
  ANDN U22507 ( .B(n20876), .A(n22109), .Z(n22108) );
  XNOR U22508 ( .A(n22110), .B(n21670), .Z(n18644) );
  ANDN U22509 ( .B(n20880), .A(n22111), .Z(n22110) );
  XOR U22510 ( .A(n22112), .B(n22113), .Z(n19711) );
  XNOR U22511 ( .A(n16314), .B(n17069), .Z(n22113) );
  XNOR U22512 ( .A(n22114), .B(n22115), .Z(n17069) );
  ANDN U22513 ( .B(n22116), .A(n20728), .Z(n22114) );
  XNOR U22514 ( .A(n22117), .B(n22118), .Z(n16314) );
  NOR U22515 ( .A(n20724), .B(n22119), .Z(n22117) );
  XOR U22516 ( .A(n16804), .B(n22120), .Z(n22112) );
  XNOR U22517 ( .A(n22121), .B(n17141), .Z(n22120) );
  XOR U22518 ( .A(n22122), .B(n22123), .Z(n17141) );
  XNOR U22519 ( .A(n22126), .B(n22127), .Z(n16804) );
  ANDN U22520 ( .B(n20715), .A(n22128), .Z(n22126) );
  AND U22521 ( .A(n18559), .B(n17883), .Z(n22097) );
  XOR U22522 ( .A(n22129), .B(n22130), .Z(n12920) );
  XNOR U22523 ( .A(n10155), .B(n11781), .Z(n22130) );
  XOR U22524 ( .A(n22131), .B(n16276), .Z(n11781) );
  XNOR U22525 ( .A(n22132), .B(n18712), .Z(n16276) );
  XNOR U22526 ( .A(n19725), .B(n21394), .Z(n18712) );
  XNOR U22527 ( .A(n22133), .B(n22134), .Z(n21394) );
  XOR U22528 ( .A(n18966), .B(n22135), .Z(n22134) );
  XOR U22529 ( .A(n22136), .B(n19811), .Z(n18966) );
  XOR U22530 ( .A(n17187), .B(n22138), .Z(n22133) );
  XOR U22531 ( .A(n18340), .B(n18650), .Z(n22138) );
  XNOR U22532 ( .A(n22139), .B(n19802), .Z(n18650) );
  AND U22533 ( .A(n22140), .B(n20895), .Z(n22139) );
  XNOR U22534 ( .A(n22141), .B(n19806), .Z(n18340) );
  XNOR U22535 ( .A(n22143), .B(n19815), .Z(n17187) );
  ANDN U22536 ( .B(n20890), .A(n22144), .Z(n22143) );
  XOR U22537 ( .A(n22145), .B(n22146), .Z(n19725) );
  XNOR U22538 ( .A(n20151), .B(n19261), .Z(n22146) );
  XNOR U22539 ( .A(n22147), .B(n22148), .Z(n19261) );
  ANDN U22540 ( .B(n22149), .A(n22047), .Z(n22147) );
  XNOR U22541 ( .A(n22150), .B(n22151), .Z(n20151) );
  ANDN U22542 ( .B(n22152), .A(n22055), .Z(n22150) );
  XOR U22543 ( .A(n20020), .B(n22153), .Z(n22145) );
  XOR U22544 ( .A(n19306), .B(n16083), .Z(n22153) );
  XOR U22545 ( .A(n22154), .B(n22155), .Z(n16083) );
  XOR U22546 ( .A(n22157), .B(n22158), .Z(n19306) );
  NOR U22547 ( .A(n22051), .B(n22159), .Z(n22157) );
  IV U22548 ( .A(n22160), .Z(n22051) );
  XOR U22549 ( .A(n22161), .B(n22162), .Z(n20020) );
  AND U22550 ( .A(n22163), .B(n22042), .Z(n22161) );
  XOR U22551 ( .A(n21314), .B(n18165), .Z(n16235) );
  IV U22552 ( .A(n17658), .Z(n18165) );
  XOR U22553 ( .A(n18701), .B(n22164), .Z(n17658) );
  XNOR U22554 ( .A(n22165), .B(n22166), .Z(n18701) );
  XNOR U22555 ( .A(n16987), .B(n16000), .Z(n22166) );
  XNOR U22556 ( .A(n22167), .B(n22168), .Z(n16000) );
  AND U22557 ( .A(n21310), .B(n21311), .Z(n22167) );
  XNOR U22558 ( .A(n22169), .B(n22170), .Z(n16987) );
  NOR U22559 ( .A(n22171), .B(n21306), .Z(n22169) );
  XNOR U22560 ( .A(n18272), .B(n22172), .Z(n22165) );
  XNOR U22561 ( .A(n19772), .B(n17468), .Z(n22172) );
  XNOR U22562 ( .A(n22173), .B(n22174), .Z(n17468) );
  AND U22563 ( .A(n21318), .B(n21316), .Z(n22173) );
  XOR U22564 ( .A(n22175), .B(n22176), .Z(n19772) );
  ANDN U22565 ( .B(n22177), .A(n22178), .Z(n22175) );
  XOR U22566 ( .A(n22179), .B(n22180), .Z(n18272) );
  NOR U22567 ( .A(n22181), .B(n21320), .Z(n22179) );
  XNOR U22568 ( .A(n22182), .B(n22177), .Z(n21314) );
  ANDN U22569 ( .B(n22178), .A(n22183), .Z(n22182) );
  XOR U22570 ( .A(n22184), .B(n17306), .Z(n16237) );
  IV U22571 ( .A(n18314), .Z(n17306) );
  XOR U22572 ( .A(n19967), .B(n22185), .Z(n18314) );
  XOR U22573 ( .A(n22186), .B(n22187), .Z(n19967) );
  XNOR U22574 ( .A(n16847), .B(n17355), .Z(n22187) );
  XNOR U22575 ( .A(n22188), .B(n22189), .Z(n17355) );
  ANDN U22576 ( .B(n22190), .A(n22191), .Z(n22188) );
  XNOR U22577 ( .A(n22192), .B(n22193), .Z(n16847) );
  ANDN U22578 ( .B(n22194), .A(n22195), .Z(n22192) );
  XOR U22579 ( .A(n18686), .B(n22196), .Z(n22186) );
  XNOR U22580 ( .A(n19517), .B(n22197), .Z(n22196) );
  XNOR U22581 ( .A(n22198), .B(n22199), .Z(n19517) );
  AND U22582 ( .A(n22200), .B(n22201), .Z(n22198) );
  XOR U22583 ( .A(n22202), .B(n22203), .Z(n18686) );
  ANDN U22584 ( .B(n22204), .A(n22205), .Z(n22202) );
  XOR U22585 ( .A(n22206), .B(n16279), .Z(n10155) );
  XOR U22586 ( .A(n22207), .B(n19757), .Z(n16279) );
  ANDN U22587 ( .B(n16232), .A(n16230), .Z(n22206) );
  XNOR U22588 ( .A(n22208), .B(n17601), .Z(n16230) );
  XOR U22589 ( .A(n21503), .B(n22031), .Z(n17601) );
  XNOR U22590 ( .A(n22209), .B(n22210), .Z(n22031) );
  XOR U22591 ( .A(n17556), .B(n18202), .Z(n22210) );
  XNOR U22592 ( .A(n22211), .B(n22212), .Z(n18202) );
  ANDN U22593 ( .B(n21243), .A(n21244), .Z(n22211) );
  XOR U22594 ( .A(n22213), .B(n22214), .Z(n21244) );
  XOR U22595 ( .A(n22215), .B(n22216), .Z(n17556) );
  ANDN U22596 ( .B(n21246), .A(n20685), .Z(n22215) );
  XOR U22597 ( .A(n22217), .B(n22218), .Z(n20685) );
  XNOR U22598 ( .A(n18489), .B(n22219), .Z(n22209) );
  XOR U22599 ( .A(n17260), .B(n19733), .Z(n22219) );
  XNOR U22600 ( .A(n22220), .B(n22221), .Z(n19733) );
  NOR U22601 ( .A(n20689), .B(n21252), .Z(n22220) );
  XNOR U22602 ( .A(n22224), .B(n22225), .Z(n17260) );
  ANDN U22603 ( .B(n21250), .A(n20676), .Z(n22224) );
  XOR U22604 ( .A(n22226), .B(n22227), .Z(n20676) );
  XNOR U22605 ( .A(n22228), .B(n22229), .Z(n18489) );
  ANDN U22606 ( .B(n22028), .A(n20680), .Z(n22228) );
  XOR U22607 ( .A(n22230), .B(n22231), .Z(n20680) );
  XOR U22608 ( .A(n22232), .B(n22233), .Z(n21503) );
  XOR U22609 ( .A(n17858), .B(n17844), .Z(n22233) );
  XOR U22610 ( .A(n22234), .B(n22235), .Z(n17844) );
  NOR U22611 ( .A(n22236), .B(n22237), .Z(n22234) );
  XNOR U22612 ( .A(n22238), .B(n22239), .Z(n17858) );
  ANDN U22613 ( .B(n22240), .A(n22241), .Z(n22238) );
  XOR U22614 ( .A(n17798), .B(n22242), .Z(n22232) );
  XNOR U22615 ( .A(n17107), .B(n22243), .Z(n22242) );
  XOR U22616 ( .A(n22244), .B(n22245), .Z(n17107) );
  ANDN U22617 ( .B(n22246), .A(n22247), .Z(n22244) );
  XNOR U22618 ( .A(n22248), .B(n22249), .Z(n17798) );
  ANDN U22619 ( .B(n22250), .A(n22251), .Z(n22248) );
  XOR U22620 ( .A(n16367), .B(n20465), .Z(n16232) );
  XNOR U22621 ( .A(n22252), .B(n21635), .Z(n20465) );
  ANDN U22622 ( .B(n20244), .A(n22253), .Z(n22252) );
  XOR U22623 ( .A(n9878), .B(n22254), .Z(n22129) );
  XOR U22624 ( .A(n14925), .B(n10652), .Z(n22254) );
  XOR U22625 ( .A(n22255), .B(n17070), .Z(n10652) );
  XOR U22626 ( .A(n18187), .B(n22256), .Z(n17070) );
  ANDN U22627 ( .B(n16228), .A(n16226), .Z(n22255) );
  XOR U22628 ( .A(n22257), .B(n19102), .Z(n16226) );
  IV U22629 ( .A(n16664), .Z(n19102) );
  XNOR U22630 ( .A(n22259), .B(n22260), .Z(n20045) );
  XOR U22631 ( .A(n18754), .B(n18466), .Z(n22260) );
  XNOR U22632 ( .A(n22261), .B(n20111), .Z(n18466) );
  AND U22633 ( .A(n20112), .B(n22262), .Z(n22261) );
  XOR U22634 ( .A(n22263), .B(n20102), .Z(n18754) );
  IV U22635 ( .A(n22264), .Z(n20102) );
  ANDN U22636 ( .B(n20103), .A(n22265), .Z(n22263) );
  XOR U22637 ( .A(n20096), .B(n22266), .Z(n22259) );
  XNOR U22638 ( .A(n17332), .B(n17665), .Z(n22266) );
  XNOR U22639 ( .A(n22267), .B(n20120), .Z(n17665) );
  IV U22640 ( .A(n22268), .Z(n20120) );
  ANDN U22641 ( .B(n22269), .A(n20119), .Z(n22267) );
  XNOR U22642 ( .A(n22270), .B(n20106), .Z(n17332) );
  ANDN U22643 ( .B(n22271), .A(n22272), .Z(n22270) );
  XOR U22644 ( .A(n22273), .B(n20115), .Z(n20096) );
  NOR U22645 ( .A(n22274), .B(n20116), .Z(n22273) );
  XOR U22646 ( .A(n21431), .B(n18865), .Z(n16228) );
  XOR U22647 ( .A(n22275), .B(n22276), .Z(n21431) );
  ANDN U22648 ( .B(n22277), .A(n22278), .Z(n22275) );
  XNOR U22649 ( .A(n22279), .B(n16272), .Z(n14925) );
  XNOR U22650 ( .A(n22280), .B(n21095), .Z(n16272) );
  XNOR U22651 ( .A(n22281), .B(n22282), .Z(n21095) );
  ANDN U22652 ( .B(n16241), .A(n16239), .Z(n22279) );
  XOR U22653 ( .A(n22283), .B(n18221), .Z(n16239) );
  XNOR U22654 ( .A(n20391), .B(n19179), .Z(n18221) );
  XOR U22655 ( .A(n22284), .B(n22285), .Z(n19179) );
  XNOR U22656 ( .A(n18398), .B(n20084), .Z(n22285) );
  XNOR U22657 ( .A(n22286), .B(n22287), .Z(n20084) );
  NOR U22658 ( .A(n22288), .B(n22289), .Z(n22286) );
  XOR U22659 ( .A(n22290), .B(n22291), .Z(n18398) );
  NOR U22660 ( .A(n22292), .B(n22293), .Z(n22290) );
  XOR U22661 ( .A(n19648), .B(n22294), .Z(n22284) );
  XOR U22662 ( .A(n19607), .B(n16574), .Z(n22294) );
  XOR U22663 ( .A(n22295), .B(n22296), .Z(n16574) );
  AND U22664 ( .A(n22297), .B(n22298), .Z(n22295) );
  XOR U22665 ( .A(n22299), .B(n22300), .Z(n19607) );
  ANDN U22666 ( .B(n22301), .A(n22302), .Z(n22299) );
  XNOR U22667 ( .A(n22303), .B(n22304), .Z(n19648) );
  NOR U22668 ( .A(n22305), .B(n22306), .Z(n22303) );
  XOR U22669 ( .A(n22307), .B(n22308), .Z(n20391) );
  XNOR U22670 ( .A(n21579), .B(n19173), .Z(n22308) );
  XOR U22671 ( .A(n22309), .B(n20579), .Z(n19173) );
  XOR U22672 ( .A(n22310), .B(n21833), .Z(n20579) );
  ANDN U22673 ( .B(n21619), .A(n22311), .Z(n22309) );
  XOR U22674 ( .A(n22312), .B(n20590), .Z(n21579) );
  XOR U22675 ( .A(n22313), .B(n22314), .Z(n20590) );
  ANDN U22676 ( .B(n21612), .A(n22315), .Z(n22312) );
  XOR U22677 ( .A(n18441), .B(n22316), .Z(n22307) );
  XOR U22678 ( .A(n18900), .B(n18472), .Z(n22316) );
  XOR U22679 ( .A(n22317), .B(n20586), .Z(n18472) );
  XNOR U22680 ( .A(n22318), .B(n22319), .Z(n20586) );
  NOR U22681 ( .A(n21610), .B(n22320), .Z(n22317) );
  XOR U22682 ( .A(n22321), .B(n21616), .Z(n18900) );
  NOR U22683 ( .A(n22322), .B(n21617), .Z(n22321) );
  XNOR U22684 ( .A(n22323), .B(n20575), .Z(n18441) );
  XOR U22685 ( .A(n22324), .B(n21596), .Z(n20575) );
  IV U22686 ( .A(n22325), .Z(n21596) );
  NOR U22687 ( .A(n22326), .B(n21621), .Z(n22323) );
  XOR U22688 ( .A(n21272), .B(n20856), .Z(n16241) );
  XNOR U22689 ( .A(n22327), .B(n22328), .Z(n20856) );
  ANDN U22690 ( .B(n22329), .A(n21549), .Z(n22327) );
  IV U22691 ( .A(n22330), .Z(n21549) );
  XNOR U22692 ( .A(n22331), .B(n16269), .Z(n9878) );
  XNOR U22693 ( .A(n16071), .B(n22332), .Z(n16269) );
  XOR U22694 ( .A(n20773), .B(n22333), .Z(n16071) );
  XOR U22695 ( .A(n22334), .B(n22335), .Z(n20773) );
  XOR U22696 ( .A(n19901), .B(n18424), .Z(n22335) );
  XOR U22697 ( .A(n22336), .B(n19924), .Z(n18424) );
  XOR U22698 ( .A(n22337), .B(n22338), .Z(n19924) );
  NOR U22699 ( .A(n22339), .B(n19923), .Z(n22336) );
  XNOR U22700 ( .A(n22340), .B(n19928), .Z(n19901) );
  XOR U22701 ( .A(n22341), .B(n22342), .Z(n19928) );
  NOR U22702 ( .A(n22343), .B(n19927), .Z(n22340) );
  XOR U22703 ( .A(n18885), .B(n22344), .Z(n22334) );
  XOR U22704 ( .A(n17312), .B(n16330), .Z(n22344) );
  XNOR U22705 ( .A(n22345), .B(n19932), .Z(n16330) );
  XNOR U22706 ( .A(n22346), .B(n22347), .Z(n19932) );
  NOR U22707 ( .A(n19933), .B(n22348), .Z(n22345) );
  XOR U22708 ( .A(n22349), .B(n19937), .Z(n17312) );
  XOR U22709 ( .A(n22350), .B(n21728), .Z(n19937) );
  ANDN U22710 ( .B(n22351), .A(n19936), .Z(n22349) );
  XNOR U22711 ( .A(n22352), .B(n19941), .Z(n18885) );
  XOR U22712 ( .A(n22353), .B(n22354), .Z(n19941) );
  ANDN U22713 ( .B(n22355), .A(n19940), .Z(n22352) );
  IV U22714 ( .A(n22356), .Z(n19940) );
  ANDN U22715 ( .B(n16245), .A(n16243), .Z(n22331) );
  XNOR U22716 ( .A(n20454), .B(n17093), .Z(n16243) );
  XNOR U22717 ( .A(n22357), .B(n22358), .Z(n20454) );
  ANDN U22718 ( .B(n22359), .A(n22360), .Z(n22357) );
  XNOR U22719 ( .A(n19279), .B(n22361), .Z(n16245) );
  IV U22720 ( .A(n19399), .Z(n19279) );
  XNOR U22721 ( .A(n18750), .B(n22362), .Z(n19399) );
  XOR U22722 ( .A(n22363), .B(n22364), .Z(n18750) );
  XNOR U22723 ( .A(n17182), .B(n17965), .Z(n22364) );
  XNOR U22724 ( .A(n22365), .B(n22366), .Z(n17965) );
  ANDN U22725 ( .B(n22367), .A(n22368), .Z(n22365) );
  XOR U22726 ( .A(n22369), .B(n22370), .Z(n17182) );
  ANDN U22727 ( .B(n22371), .A(n22372), .Z(n22369) );
  XOR U22728 ( .A(n20495), .B(n22373), .Z(n22363) );
  XOR U22729 ( .A(n16877), .B(n22374), .Z(n22373) );
  XNOR U22730 ( .A(n22375), .B(n22376), .Z(n16877) );
  ANDN U22731 ( .B(n22377), .A(n22378), .Z(n22375) );
  XNOR U22732 ( .A(n22379), .B(n22380), .Z(n20495) );
  AND U22733 ( .A(n22381), .B(n22382), .Z(n22379) );
  XNOR U22734 ( .A(n22383), .B(n17883), .Z(n14121) );
  XOR U22735 ( .A(n19912), .B(n19072), .Z(n17883) );
  XNOR U22736 ( .A(n19838), .B(n22384), .Z(n19072) );
  XNOR U22737 ( .A(n22385), .B(n22386), .Z(n19838) );
  XNOR U22738 ( .A(n18639), .B(n19958), .Z(n22386) );
  XNOR U22739 ( .A(n22387), .B(n22388), .Z(n19958) );
  ANDN U22740 ( .B(n19906), .A(n22389), .Z(n22387) );
  XOR U22741 ( .A(n22390), .B(n22391), .Z(n19906) );
  XOR U22742 ( .A(n22392), .B(n20832), .Z(n18639) );
  ANDN U22743 ( .B(n19910), .A(n20833), .Z(n22392) );
  XOR U22744 ( .A(n22393), .B(n22394), .Z(n20833) );
  XNOR U22745 ( .A(n22395), .B(n22396), .Z(n19910) );
  XNOR U22746 ( .A(n18432), .B(n22397), .Z(n22385) );
  XNOR U22747 ( .A(n18464), .B(n19835), .Z(n22397) );
  XNOR U22748 ( .A(n22398), .B(n22399), .Z(n19835) );
  XOR U22749 ( .A(n22400), .B(n22401), .Z(n20494) );
  XNOR U22750 ( .A(n22402), .B(n21002), .Z(n18464) );
  ANDN U22751 ( .B(n19916), .A(n19917), .Z(n22402) );
  XOR U22752 ( .A(n22403), .B(n22404), .Z(n19917) );
  XNOR U22753 ( .A(n22405), .B(n22406), .Z(n19916) );
  XNOR U22754 ( .A(n22407), .B(n20830), .Z(n18432) );
  ANDN U22755 ( .B(n20829), .A(n20786), .Z(n22407) );
  XNOR U22756 ( .A(n22408), .B(n20829), .Z(n19912) );
  XOR U22757 ( .A(n22409), .B(n22410), .Z(n20829) );
  ANDN U22758 ( .B(n20786), .A(n20787), .Z(n22408) );
  XNOR U22759 ( .A(n22411), .B(n22412), .Z(n20786) );
  ANDN U22760 ( .B(n17818), .A(n18559), .Z(n22383) );
  XOR U22761 ( .A(n18027), .B(n22413), .Z(n18559) );
  XNOR U22762 ( .A(n20296), .B(n18342), .Z(n18027) );
  XNOR U22763 ( .A(n22414), .B(n22415), .Z(n18342) );
  XNOR U22764 ( .A(n22416), .B(n17486), .Z(n22415) );
  XOR U22765 ( .A(n22417), .B(n20217), .Z(n17486) );
  ANDN U22766 ( .B(n20771), .A(n22418), .Z(n22417) );
  XOR U22767 ( .A(n19331), .B(n22419), .Z(n22414) );
  XOR U22768 ( .A(n19034), .B(n19432), .Z(n22419) );
  XNOR U22769 ( .A(n22420), .B(n20208), .Z(n19432) );
  AND U22770 ( .A(n22421), .B(n22422), .Z(n22420) );
  XNOR U22771 ( .A(n22423), .B(n20212), .Z(n19034) );
  XNOR U22772 ( .A(n22425), .B(n22426), .Z(n19331) );
  ANDN U22773 ( .B(n20814), .A(n22427), .Z(n22425) );
  XOR U22774 ( .A(n22428), .B(n22429), .Z(n20296) );
  XOR U22775 ( .A(n19450), .B(n20670), .Z(n22429) );
  XNOR U22776 ( .A(n22430), .B(n22431), .Z(n20670) );
  NOR U22777 ( .A(n22432), .B(n22433), .Z(n22430) );
  XNOR U22778 ( .A(n22434), .B(n22435), .Z(n19450) );
  NOR U22779 ( .A(n22436), .B(n20927), .Z(n22434) );
  XOR U22780 ( .A(n19601), .B(n22437), .Z(n22428) );
  XOR U22781 ( .A(n20026), .B(n22438), .Z(n22437) );
  XNOR U22782 ( .A(n22439), .B(n22440), .Z(n20026) );
  NOR U22783 ( .A(n22441), .B(n20914), .Z(n22439) );
  XOR U22784 ( .A(n22442), .B(n22443), .Z(n19601) );
  XOR U22785 ( .A(n22445), .B(n17098), .Z(n17818) );
  XNOR U22786 ( .A(n20672), .B(n19708), .Z(n17098) );
  XNOR U22787 ( .A(n22446), .B(n22447), .Z(n19708) );
  XNOR U22788 ( .A(n20090), .B(n18531), .Z(n22447) );
  XOR U22789 ( .A(n22448), .B(n22449), .Z(n18531) );
  AND U22790 ( .A(n22450), .B(n22451), .Z(n22448) );
  XOR U22791 ( .A(n22452), .B(n22453), .Z(n20090) );
  ANDN U22792 ( .B(n22454), .A(n22455), .Z(n22452) );
  XOR U22793 ( .A(n22456), .B(n22457), .Z(n22446) );
  XOR U22794 ( .A(n19285), .B(n16754), .Z(n22457) );
  XNOR U22795 ( .A(n22458), .B(n22459), .Z(n16754) );
  AND U22796 ( .A(n22460), .B(n22461), .Z(n22458) );
  XOR U22797 ( .A(n22462), .B(n22463), .Z(n19285) );
  ANDN U22798 ( .B(n22464), .A(n22465), .Z(n22462) );
  XOR U22799 ( .A(n22466), .B(n22467), .Z(n20672) );
  XOR U22800 ( .A(n19068), .B(n18226), .Z(n22467) );
  XOR U22801 ( .A(n22468), .B(n22237), .Z(n18226) );
  ANDN U22802 ( .B(n22469), .A(n22470), .Z(n22468) );
  XNOR U22803 ( .A(n22471), .B(n22247), .Z(n19068) );
  ANDN U22804 ( .B(n22472), .A(n22473), .Z(n22471) );
  XOR U22805 ( .A(n19600), .B(n22474), .Z(n22466) );
  XNOR U22806 ( .A(n19657), .B(n21239), .Z(n22474) );
  XOR U22807 ( .A(n22475), .B(n22476), .Z(n21239) );
  NOR U22808 ( .A(n22477), .B(n22478), .Z(n22475) );
  XNOR U22809 ( .A(n22479), .B(n22241), .Z(n19657) );
  ANDN U22810 ( .B(n22480), .A(n22481), .Z(n22479) );
  XNOR U22811 ( .A(n22482), .B(n22251), .Z(n19600) );
  NOR U22812 ( .A(n9258), .B(n9257), .Z(n21896) );
  XNOR U22813 ( .A(n10200), .B(n17367), .Z(n9257) );
  XOR U22814 ( .A(n22485), .B(n19846), .Z(n17367) );
  ANDN U22815 ( .B(n18350), .A(n19640), .Z(n22485) );
  XNOR U22816 ( .A(n22486), .B(n18033), .Z(n18350) );
  IV U22817 ( .A(n10690), .Z(n10200) );
  XOR U22818 ( .A(n22487), .B(n22488), .Z(n16969) );
  XNOR U22819 ( .A(n11767), .B(n11831), .Z(n22488) );
  XOR U22820 ( .A(n20765), .B(n16504), .Z(n17766) );
  IV U22821 ( .A(n20074), .Z(n16504) );
  XNOR U22822 ( .A(n22490), .B(n22491), .Z(n20480) );
  XNOR U22823 ( .A(n22413), .B(n18625), .Z(n22491) );
  XNOR U22824 ( .A(n22492), .B(n22427), .Z(n18625) );
  NOR U22825 ( .A(n20814), .B(n20202), .Z(n22492) );
  XNOR U22826 ( .A(n22493), .B(n22494), .Z(n20202) );
  XNOR U22827 ( .A(n22495), .B(n22496), .Z(n20814) );
  XOR U22828 ( .A(n22497), .B(n22498), .Z(n22413) );
  ANDN U22829 ( .B(n20768), .A(n20219), .Z(n22497) );
  XNOR U22830 ( .A(n22499), .B(n22500), .Z(n20219) );
  XOR U22831 ( .A(n19850), .B(n22501), .Z(n22490) );
  XOR U22832 ( .A(n18037), .B(n18028), .Z(n22501) );
  XNOR U22833 ( .A(n22502), .B(n22418), .Z(n18028) );
  NOR U22834 ( .A(n20215), .B(n20771), .Z(n22502) );
  XNOR U22835 ( .A(n22503), .B(n22504), .Z(n20771) );
  XNOR U22836 ( .A(n22505), .B(n22506), .Z(n20215) );
  XOR U22837 ( .A(n22507), .B(n22421), .Z(n18037) );
  NOR U22838 ( .A(n22508), .B(n22422), .Z(n22507) );
  XNOR U22839 ( .A(n22509), .B(n22424), .Z(n19850) );
  ANDN U22840 ( .B(n20764), .A(n20211), .Z(n22509) );
  XNOR U22841 ( .A(n22510), .B(n21829), .Z(n20211) );
  XNOR U22842 ( .A(n22511), .B(n22512), .Z(n20764) );
  XNOR U22843 ( .A(n22513), .B(n22514), .Z(n18460) );
  XNOR U22844 ( .A(n18856), .B(n16380), .Z(n22514) );
  XOR U22845 ( .A(n22515), .B(n22444), .Z(n16380) );
  NOR U22846 ( .A(n20931), .B(n20932), .Z(n22515) );
  XOR U22847 ( .A(n22516), .B(n22517), .Z(n20931) );
  XNOR U22848 ( .A(n22518), .B(n22433), .Z(n18856) );
  ANDN U22849 ( .B(n22432), .A(n22519), .Z(n22518) );
  IV U22850 ( .A(n20923), .Z(n22432) );
  XNOR U22851 ( .A(n22520), .B(n22521), .Z(n20923) );
  XOR U22852 ( .A(n17638), .B(n22522), .Z(n22513) );
  XOR U22853 ( .A(n20295), .B(n16118), .Z(n22522) );
  XOR U22854 ( .A(n22523), .B(n22524), .Z(n16118) );
  XOR U22855 ( .A(n22525), .B(n22526), .Z(n20927) );
  XOR U22856 ( .A(n22527), .B(n22528), .Z(n20295) );
  AND U22857 ( .A(n20916), .B(n20914), .Z(n22527) );
  XOR U22858 ( .A(n22511), .B(n22529), .Z(n20914) );
  XNOR U22859 ( .A(n22530), .B(n22531), .Z(n17638) );
  ANDN U22860 ( .B(n20919), .A(n20918), .Z(n22530) );
  XNOR U22861 ( .A(n22532), .B(n22422), .Z(n20765) );
  XNOR U22862 ( .A(n22533), .B(n22534), .Z(n22422) );
  ANDN U22863 ( .B(n20207), .A(n20206), .Z(n22532) );
  IV U22864 ( .A(n22508), .Z(n20206) );
  XOR U22865 ( .A(n22535), .B(n22536), .Z(n22508) );
  NOR U22866 ( .A(n17374), .B(n17375), .Z(n22489) );
  XOR U22867 ( .A(n19041), .B(n18819), .Z(n15639) );
  XOR U22868 ( .A(n22538), .B(n22539), .Z(n18819) );
  XNOR U22869 ( .A(n19590), .B(n17577), .Z(n22539) );
  XOR U22870 ( .A(n22540), .B(n22541), .Z(n17577) );
  ANDN U22871 ( .B(n21203), .A(n22542), .Z(n22540) );
  XNOR U22872 ( .A(n22543), .B(n22544), .Z(n19590) );
  ANDN U22873 ( .B(n20948), .A(n22545), .Z(n22543) );
  XOR U22874 ( .A(n18080), .B(n22546), .Z(n22538) );
  XOR U22875 ( .A(n19142), .B(n22547), .Z(n22546) );
  XNOR U22876 ( .A(n22548), .B(n22549), .Z(n19142) );
  ANDN U22877 ( .B(n22550), .A(n20944), .Z(n22548) );
  XOR U22878 ( .A(n22551), .B(n22552), .Z(n18080) );
  ANDN U22879 ( .B(n20954), .A(n22553), .Z(n22551) );
  XOR U22880 ( .A(n22554), .B(n22555), .Z(n19041) );
  XOR U22881 ( .A(n19271), .B(n14957), .Z(n22555) );
  XNOR U22882 ( .A(n22556), .B(n22557), .Z(n14957) );
  NOR U22883 ( .A(n22558), .B(n22559), .Z(n22556) );
  XOR U22884 ( .A(n22560), .B(n22561), .Z(n19271) );
  NOR U22885 ( .A(n22562), .B(n22563), .Z(n22560) );
  XOR U22886 ( .A(n15335), .B(n22564), .Z(n22554) );
  XNOR U22887 ( .A(n20381), .B(n16069), .Z(n22564) );
  XOR U22888 ( .A(n22565), .B(n22566), .Z(n16069) );
  NOR U22889 ( .A(n22567), .B(n22568), .Z(n22565) );
  XNOR U22890 ( .A(n22569), .B(n22570), .Z(n20381) );
  NOR U22891 ( .A(n22571), .B(n22572), .Z(n22569) );
  XNOR U22892 ( .A(n22573), .B(n22574), .Z(n15335) );
  NOR U22893 ( .A(n22575), .B(n22576), .Z(n22573) );
  IV U22894 ( .A(n19830), .Z(n17374) );
  XOR U22895 ( .A(n22577), .B(n16585), .Z(n19830) );
  XNOR U22896 ( .A(n22578), .B(n22579), .Z(n16585) );
  XNOR U22897 ( .A(n22580), .B(n17763), .Z(n11767) );
  XOR U22898 ( .A(n22581), .B(n22582), .Z(n17763) );
  XOR U22899 ( .A(n22583), .B(n19757), .Z(n17383) );
  XOR U22900 ( .A(n22584), .B(n19740), .Z(n17382) );
  XOR U22901 ( .A(n22586), .B(n22587), .Z(n19042) );
  XNOR U22902 ( .A(n22588), .B(n19379), .Z(n22587) );
  XOR U22903 ( .A(n22589), .B(n22590), .Z(n19379) );
  XNOR U22904 ( .A(n22593), .B(n22594), .Z(n22586) );
  XNOR U22905 ( .A(n16829), .B(n17030), .Z(n22594) );
  XNOR U22906 ( .A(n22595), .B(n22596), .Z(n17030) );
  AND U22907 ( .A(n22597), .B(n22598), .Z(n22595) );
  XNOR U22908 ( .A(n22599), .B(n22600), .Z(n16829) );
  ANDN U22909 ( .B(n22601), .A(n22602), .Z(n22599) );
  XOR U22910 ( .A(n9873), .B(n22603), .Z(n22487) );
  XOR U22911 ( .A(n10781), .B(n10594), .Z(n22603) );
  XOR U22912 ( .A(n22604), .B(n18351), .Z(n10594) );
  XNOR U22913 ( .A(n22135), .B(n18967), .Z(n18351) );
  XNOR U22914 ( .A(n20152), .B(n20663), .Z(n18967) );
  XNOR U22915 ( .A(n22605), .B(n22606), .Z(n20663) );
  XNOR U22916 ( .A(n19105), .B(n17232), .Z(n22606) );
  XOR U22917 ( .A(n22607), .B(n21318), .Z(n17232) );
  XOR U22918 ( .A(n22608), .B(n22609), .Z(n21318) );
  ANDN U22919 ( .B(n22610), .A(n21317), .Z(n22607) );
  XNOR U22920 ( .A(n22611), .B(n22178), .Z(n19105) );
  XOR U22921 ( .A(n22612), .B(n22613), .Z(n22178) );
  ANDN U22922 ( .B(n22183), .A(n22614), .Z(n22611) );
  XOR U22923 ( .A(n18972), .B(n22615), .Z(n22605) );
  XOR U22924 ( .A(n21302), .B(n18694), .Z(n22615) );
  XNOR U22925 ( .A(n22616), .B(n21307), .Z(n18694) );
  IV U22926 ( .A(n22171), .Z(n21307) );
  XOR U22927 ( .A(n22617), .B(n21214), .Z(n22171) );
  ANDN U22928 ( .B(n21308), .A(n22618), .Z(n22616) );
  XNOR U22929 ( .A(n22619), .B(n22181), .Z(n21302) );
  IV U22930 ( .A(n21321), .Z(n22181) );
  XOR U22931 ( .A(n22620), .B(n22621), .Z(n21321) );
  ANDN U22932 ( .B(n21322), .A(n22622), .Z(n22619) );
  XNOR U22933 ( .A(n22623), .B(n21311), .Z(n18972) );
  XOR U22934 ( .A(n22624), .B(n22625), .Z(n21311) );
  ANDN U22935 ( .B(n21312), .A(n22626), .Z(n22623) );
  XOR U22936 ( .A(n22627), .B(n22628), .Z(n20152) );
  XOR U22937 ( .A(n19319), .B(n18391), .Z(n22628) );
  XNOR U22938 ( .A(n22629), .B(n19812), .Z(n18391) );
  XOR U22939 ( .A(n22630), .B(n22631), .Z(n19812) );
  ANDN U22940 ( .B(n19811), .A(n22137), .Z(n22629) );
  XOR U22941 ( .A(n22632), .B(n22346), .Z(n19811) );
  XNOR U22942 ( .A(n22633), .B(n19807), .Z(n19319) );
  XNOR U22943 ( .A(n22634), .B(n22635), .Z(n19807) );
  ANDN U22944 ( .B(n19806), .A(n22142), .Z(n22633) );
  XOR U22945 ( .A(n22636), .B(n22637), .Z(n19806) );
  XOR U22946 ( .A(n17519), .B(n22638), .Z(n22627) );
  XNOR U22947 ( .A(n19796), .B(n17300), .Z(n22638) );
  XNOR U22948 ( .A(n22639), .B(n19816), .Z(n17300) );
  XOR U22949 ( .A(n22640), .B(n22641), .Z(n19816) );
  ANDN U22950 ( .B(n22144), .A(n19815), .Z(n22639) );
  XOR U22951 ( .A(n22642), .B(n22643), .Z(n19815) );
  XNOR U22952 ( .A(n22644), .B(n19803), .Z(n19796) );
  XOR U22953 ( .A(n22645), .B(n22646), .Z(n19803) );
  ANDN U22954 ( .B(n19802), .A(n22140), .Z(n22644) );
  XOR U22955 ( .A(n22647), .B(n22648), .Z(n19802) );
  XNOR U22956 ( .A(n22649), .B(n19820), .Z(n17519) );
  IV U22957 ( .A(n22650), .Z(n19820) );
  NOR U22958 ( .A(n22651), .B(n19819), .Z(n22649) );
  XOR U22959 ( .A(n22652), .B(n19819), .Z(n22135) );
  XOR U22960 ( .A(n22653), .B(n22654), .Z(n19819) );
  ANDN U22961 ( .B(n22655), .A(n22656), .Z(n22652) );
  ANDN U22962 ( .B(n19640), .A(n19846), .Z(n22604) );
  XOR U22963 ( .A(n18103), .B(n22657), .Z(n19846) );
  XNOR U22964 ( .A(n21746), .B(n15339), .Z(n19640) );
  XNOR U22965 ( .A(n22660), .B(n22661), .Z(n21746) );
  AND U22966 ( .A(n22662), .B(n22663), .Z(n22660) );
  XOR U22967 ( .A(n22664), .B(n19645), .Z(n10781) );
  XOR U22968 ( .A(n22665), .B(n22666), .Z(n19645) );
  XNOR U22969 ( .A(n22667), .B(n17479), .Z(n17370) );
  XOR U22970 ( .A(n22668), .B(n22669), .Z(n21281) );
  XNOR U22971 ( .A(n17605), .B(n18262), .Z(n22669) );
  XOR U22972 ( .A(n22670), .B(n19418), .Z(n18262) );
  ANDN U22973 ( .B(n19417), .A(n21854), .Z(n22670) );
  XNOR U22974 ( .A(n22671), .B(n22672), .Z(n17605) );
  NOR U22975 ( .A(n22673), .B(n20511), .Z(n22671) );
  XOR U22976 ( .A(n17054), .B(n22674), .Z(n22668) );
  XNOR U22977 ( .A(n17083), .B(n18225), .Z(n22674) );
  XNOR U22978 ( .A(n22675), .B(n19411), .Z(n18225) );
  NOR U22979 ( .A(n19410), .B(n20515), .Z(n22675) );
  XNOR U22980 ( .A(n22676), .B(n21041), .Z(n17083) );
  NOR U22981 ( .A(n22677), .B(n20505), .Z(n22676) );
  XNOR U22982 ( .A(n22678), .B(n22679), .Z(n17054) );
  NOR U22983 ( .A(n22680), .B(n20501), .Z(n22678) );
  XNOR U22984 ( .A(n22681), .B(n22682), .Z(n19139) );
  XOR U22985 ( .A(n18430), .B(n17181), .Z(n22682) );
  XNOR U22986 ( .A(n22683), .B(n22684), .Z(n17181) );
  ANDN U22987 ( .B(n22685), .A(n22358), .Z(n22683) );
  XNOR U22988 ( .A(n22686), .B(n22687), .Z(n18430) );
  ANDN U22989 ( .B(n22688), .A(n20460), .Z(n22686) );
  XOR U22990 ( .A(n14971), .B(n22689), .Z(n22681) );
  XOR U22991 ( .A(n19404), .B(n18503), .Z(n22689) );
  XNOR U22992 ( .A(n22690), .B(n22691), .Z(n18503) );
  ANDN U22993 ( .B(n22692), .A(n22693), .Z(n22690) );
  XNOR U22994 ( .A(n22694), .B(n22695), .Z(n19404) );
  ANDN U22995 ( .B(n20456), .A(n22696), .Z(n22694) );
  XNOR U22996 ( .A(n22697), .B(n22698), .Z(n14971) );
  ANDN U22997 ( .B(n20450), .A(n22699), .Z(n22697) );
  XNOR U22998 ( .A(n20269), .B(n16954), .Z(n17369) );
  XOR U22999 ( .A(n22700), .B(n22701), .Z(n20269) );
  ANDN U23000 ( .B(n21948), .A(n22702), .Z(n22700) );
  XOR U23001 ( .A(n22703), .B(n17757), .Z(n9873) );
  XOR U23002 ( .A(n22704), .B(n18890), .Z(n17757) );
  XOR U23003 ( .A(n21813), .B(n19735), .Z(n18890) );
  XOR U23004 ( .A(n22705), .B(n22706), .Z(n19735) );
  XNOR U23005 ( .A(n17560), .B(n21094), .Z(n22706) );
  XOR U23006 ( .A(n22707), .B(n22708), .Z(n21094) );
  NOR U23007 ( .A(n22709), .B(n22710), .Z(n22707) );
  XNOR U23008 ( .A(n22711), .B(n22712), .Z(n17560) );
  ANDN U23009 ( .B(n22713), .A(n22714), .Z(n22711) );
  XNOR U23010 ( .A(n22280), .B(n22715), .Z(n22705) );
  XOR U23011 ( .A(n19064), .B(n15678), .Z(n22715) );
  XNOR U23012 ( .A(n22716), .B(n22717), .Z(n15678) );
  NOR U23013 ( .A(n22718), .B(n22719), .Z(n22716) );
  XNOR U23014 ( .A(n22720), .B(n22721), .Z(n19064) );
  NOR U23015 ( .A(n22722), .B(n22723), .Z(n22720) );
  XNOR U23016 ( .A(n22724), .B(n22725), .Z(n22280) );
  NOR U23017 ( .A(n22726), .B(n22727), .Z(n22724) );
  XOR U23018 ( .A(n22728), .B(n22729), .Z(n21813) );
  XNOR U23019 ( .A(n16391), .B(n22730), .Z(n22729) );
  XNOR U23020 ( .A(n22731), .B(n22732), .Z(n16391) );
  ANDN U23021 ( .B(n22733), .A(n22734), .Z(n22731) );
  XOR U23022 ( .A(n19247), .B(n22735), .Z(n22728) );
  XNOR U23023 ( .A(n19315), .B(n17496), .Z(n22735) );
  XNOR U23024 ( .A(n22736), .B(n22737), .Z(n17496) );
  XNOR U23025 ( .A(n22740), .B(n22741), .Z(n19315) );
  ANDN U23026 ( .B(n22742), .A(n22743), .Z(n22740) );
  XNOR U23027 ( .A(n22744), .B(n22745), .Z(n19247) );
  AND U23028 ( .A(n22746), .B(n22747), .Z(n22744) );
  NOR U23029 ( .A(n17380), .B(n17378), .Z(n22703) );
  XNOR U23030 ( .A(n21125), .B(n17282), .Z(n17378) );
  XOR U23031 ( .A(n21097), .B(n19422), .Z(n17282) );
  XNOR U23032 ( .A(n22748), .B(n22749), .Z(n19422) );
  XNOR U23033 ( .A(n20222), .B(n22750), .Z(n22749) );
  XNOR U23034 ( .A(n22751), .B(n21085), .Z(n20222) );
  NOR U23035 ( .A(n21119), .B(n21120), .Z(n22751) );
  XOR U23036 ( .A(n17660), .B(n22752), .Z(n22748) );
  XOR U23037 ( .A(n18031), .B(n15959), .Z(n22752) );
  XOR U23038 ( .A(n22753), .B(n21081), .Z(n15959) );
  ANDN U23039 ( .B(n21127), .A(n21128), .Z(n22753) );
  XNOR U23040 ( .A(n22754), .B(n21071), .Z(n18031) );
  ANDN U23041 ( .B(n21122), .A(n22755), .Z(n22754) );
  XNOR U23042 ( .A(n22756), .B(n22757), .Z(n17660) );
  XOR U23043 ( .A(n22758), .B(n22759), .Z(n21097) );
  XNOR U23044 ( .A(n17866), .B(n19950), .Z(n22759) );
  XOR U23045 ( .A(n22760), .B(n21062), .Z(n19950) );
  ANDN U23046 ( .B(n22761), .A(n22762), .Z(n22760) );
  XOR U23047 ( .A(n22763), .B(n21048), .Z(n17866) );
  ANDN U23048 ( .B(n22764), .A(n22765), .Z(n22763) );
  XOR U23049 ( .A(n19210), .B(n22766), .Z(n22758) );
  XOR U23050 ( .A(n17625), .B(n21893), .Z(n22766) );
  XNOR U23051 ( .A(n22767), .B(n21053), .Z(n21893) );
  IV U23052 ( .A(n22768), .Z(n21053) );
  NOR U23053 ( .A(n22769), .B(n22770), .Z(n22767) );
  XNOR U23054 ( .A(n22771), .B(n21058), .Z(n17625) );
  XNOR U23055 ( .A(n22774), .B(n22775), .Z(n19210) );
  ANDN U23056 ( .B(n22776), .A(n22777), .Z(n22774) );
  XOR U23057 ( .A(n22778), .B(n22779), .Z(n21125) );
  ANDN U23058 ( .B(n21074), .A(n22780), .Z(n22778) );
  XOR U23059 ( .A(n22781), .B(n16056), .Z(n17380) );
  XNOR U23060 ( .A(n22782), .B(n22783), .Z(n18484) );
  XOR U23061 ( .A(n14188), .B(n14764), .Z(n22783) );
  XOR U23062 ( .A(n22784), .B(n14778), .Z(n14764) );
  XNOR U23063 ( .A(n21985), .B(n16589), .Z(n14778) );
  IV U23064 ( .A(n16596), .Z(n16589) );
  XOR U23065 ( .A(n22785), .B(n18461), .Z(n16596) );
  XNOR U23066 ( .A(n22786), .B(n22787), .Z(n18461) );
  XNOR U23067 ( .A(n17786), .B(n16966), .Z(n22787) );
  XNOR U23068 ( .A(n22788), .B(n21008), .Z(n16966) );
  ANDN U23069 ( .B(n21009), .A(n21991), .Z(n22788) );
  XNOR U23070 ( .A(n22789), .B(n22790), .Z(n21009) );
  XNOR U23071 ( .A(n22791), .B(n21013), .Z(n17786) );
  XOR U23072 ( .A(n22792), .B(n22793), .Z(n21012) );
  XOR U23073 ( .A(n17502), .B(n22794), .Z(n22786) );
  XOR U23074 ( .A(n18738), .B(n21003), .Z(n22794) );
  XOR U23075 ( .A(n22795), .B(n21020), .Z(n21003) );
  NOR U23076 ( .A(n21019), .B(n21979), .Z(n22795) );
  XOR U23077 ( .A(n22796), .B(n21219), .Z(n21019) );
  ANDN U23078 ( .B(n22799), .A(n22800), .Z(n22797) );
  XNOR U23079 ( .A(n22801), .B(n22802), .Z(n17502) );
  ANDN U23080 ( .B(n21989), .A(n22803), .Z(n22801) );
  XNOR U23081 ( .A(n22804), .B(n22799), .Z(n21985) );
  AND U23082 ( .A(n22805), .B(n22800), .Z(n22804) );
  XNOR U23083 ( .A(n22806), .B(n17574), .Z(n14779) );
  XNOR U23084 ( .A(n18286), .B(n20825), .Z(n16569) );
  XOR U23085 ( .A(n22807), .B(n20777), .Z(n20825) );
  XNOR U23086 ( .A(n22808), .B(n22809), .Z(n20492) );
  XOR U23087 ( .A(n22811), .B(n14999), .Z(n14782) );
  IV U23088 ( .A(n18332), .Z(n14999) );
  XNOR U23089 ( .A(n22812), .B(n22813), .Z(n20360) );
  XOR U23090 ( .A(n19101), .B(n16663), .Z(n22813) );
  XOR U23091 ( .A(n22815), .B(n22816), .Z(n20119) );
  NOR U23092 ( .A(n22817), .B(n22269), .Z(n22814) );
  XNOR U23093 ( .A(n22818), .B(n20103), .Z(n19101) );
  XNOR U23094 ( .A(n22819), .B(n22820), .Z(n20103) );
  ANDN U23095 ( .B(n22265), .A(n22821), .Z(n22818) );
  XOR U23096 ( .A(n16964), .B(n22822), .Z(n22812) );
  XOR U23097 ( .A(n22257), .B(n21136), .Z(n22822) );
  XOR U23098 ( .A(n22823), .B(n20116), .Z(n21136) );
  XOR U23099 ( .A(n22824), .B(n22825), .Z(n20116) );
  NOR U23100 ( .A(n22826), .B(n22827), .Z(n22823) );
  XNOR U23101 ( .A(n22828), .B(n22272), .Z(n22257) );
  IV U23102 ( .A(n20107), .Z(n22272) );
  XOR U23103 ( .A(n22829), .B(n22830), .Z(n20107) );
  NOR U23104 ( .A(n22831), .B(n22271), .Z(n22828) );
  XNOR U23105 ( .A(n22832), .B(n20112), .Z(n16964) );
  XOR U23106 ( .A(n22833), .B(n22834), .Z(n20112) );
  ANDN U23107 ( .B(n22835), .A(n22262), .Z(n22832) );
  XOR U23108 ( .A(n22836), .B(n22837), .Z(n19311) );
  XNOR U23109 ( .A(n20043), .B(n19215), .Z(n22837) );
  XNOR U23110 ( .A(n22838), .B(n21767), .Z(n19215) );
  ANDN U23111 ( .B(n22839), .A(n22840), .Z(n22838) );
  XOR U23112 ( .A(n22841), .B(n22842), .Z(n20043) );
  XOR U23113 ( .A(n17987), .B(n22845), .Z(n22836) );
  XNOR U23114 ( .A(n18937), .B(n19253), .Z(n22845) );
  XOR U23115 ( .A(n22846), .B(n21761), .Z(n19253) );
  XNOR U23116 ( .A(n22849), .B(n21773), .Z(n18937) );
  ANDN U23117 ( .B(n22850), .A(n22851), .Z(n22849) );
  XNOR U23118 ( .A(n22852), .B(n21757), .Z(n17987) );
  ANDN U23119 ( .B(n22853), .A(n22854), .Z(n22852) );
  ANDN U23120 ( .B(n18483), .A(n14783), .Z(n22810) );
  XOR U23121 ( .A(n22855), .B(n18237), .Z(n14783) );
  IV U23122 ( .A(n18965), .Z(n18237) );
  XOR U23123 ( .A(n22856), .B(n20667), .Z(n18965) );
  XNOR U23124 ( .A(n22857), .B(n22858), .Z(n20667) );
  XNOR U23125 ( .A(n18749), .B(n16394), .Z(n22858) );
  XNOR U23126 ( .A(n22859), .B(n22367), .Z(n16394) );
  AND U23127 ( .A(n22368), .B(n22860), .Z(n22859) );
  XNOR U23128 ( .A(n22861), .B(n22382), .Z(n18749) );
  ANDN U23129 ( .B(n22862), .A(n22381), .Z(n22861) );
  XOR U23130 ( .A(n15655), .B(n22863), .Z(n22857) );
  XOR U23131 ( .A(n18242), .B(n16826), .Z(n22863) );
  XNOR U23132 ( .A(n22864), .B(n22371), .Z(n16826) );
  AND U23133 ( .A(n22865), .B(n22372), .Z(n22864) );
  XNOR U23134 ( .A(n22866), .B(n22867), .Z(n18242) );
  ANDN U23135 ( .B(n22868), .A(n22869), .Z(n22866) );
  XNOR U23136 ( .A(n22870), .B(n22377), .Z(n15655) );
  NOR U23137 ( .A(n22871), .B(n22872), .Z(n22870) );
  XOR U23138 ( .A(n21859), .B(n19263), .Z(n18483) );
  XOR U23139 ( .A(n22873), .B(n22874), .Z(n21859) );
  ANDN U23140 ( .B(n22875), .A(n22876), .Z(n22873) );
  XNOR U23141 ( .A(n12248), .B(n22877), .Z(n22782) );
  XNOR U23142 ( .A(n12593), .B(n12635), .Z(n22877) );
  XOR U23143 ( .A(n22878), .B(n14786), .Z(n12635) );
  XNOR U23144 ( .A(n22879), .B(n16074), .Z(n14786) );
  IV U23145 ( .A(n16117), .Z(n16074) );
  XNOR U23146 ( .A(n19094), .B(n22880), .Z(n16117) );
  XOR U23147 ( .A(n22881), .B(n22882), .Z(n19094) );
  XOR U23148 ( .A(n20405), .B(n19549), .Z(n22882) );
  XOR U23149 ( .A(n22883), .B(n20432), .Z(n19549) );
  ANDN U23150 ( .B(n22884), .A(n20433), .Z(n22883) );
  XNOR U23151 ( .A(n22885), .B(n20428), .Z(n20405) );
  XOR U23152 ( .A(n22886), .B(n22887), .Z(n20428) );
  ANDN U23153 ( .B(n22888), .A(n20427), .Z(n22885) );
  XNOR U23154 ( .A(n15264), .B(n22889), .Z(n22881) );
  XOR U23155 ( .A(n15286), .B(n19662), .Z(n22889) );
  XOR U23156 ( .A(n22890), .B(n20424), .Z(n19662) );
  IV U23157 ( .A(n21198), .Z(n20424) );
  XNOR U23158 ( .A(n22891), .B(n22892), .Z(n21198) );
  NOR U23159 ( .A(n22893), .B(n20423), .Z(n22890) );
  XNOR U23160 ( .A(n22894), .B(n20436), .Z(n15286) );
  XOR U23161 ( .A(n22895), .B(n22325), .Z(n20436) );
  XNOR U23162 ( .A(n22897), .B(n20440), .Z(n15264) );
  XNOR U23163 ( .A(n22898), .B(n22899), .Z(n20440) );
  ANDN U23164 ( .B(n16545), .A(n16543), .Z(n22878) );
  XOR U23165 ( .A(n22901), .B(n22902), .Z(n16543) );
  XOR U23166 ( .A(n22903), .B(n17970), .Z(n16545) );
  XNOR U23167 ( .A(n22904), .B(n22905), .Z(n17970) );
  XNOR U23168 ( .A(n22906), .B(n14774), .Z(n12593) );
  IV U23169 ( .A(n17771), .Z(n14774) );
  XOR U23170 ( .A(n20052), .B(n18150), .Z(n17771) );
  XOR U23171 ( .A(n22907), .B(n21450), .Z(n20052) );
  NOR U23172 ( .A(n14773), .B(n16548), .Z(n22906) );
  XOR U23173 ( .A(n22910), .B(n19321), .Z(n16548) );
  IV U23174 ( .A(n18836), .Z(n19321) );
  XOR U23175 ( .A(n22911), .B(n20546), .Z(n18836) );
  XNOR U23176 ( .A(n22912), .B(n22913), .Z(n20546) );
  XNOR U23177 ( .A(n22914), .B(n18492), .Z(n22913) );
  XOR U23178 ( .A(n22915), .B(n22916), .Z(n18492) );
  ANDN U23179 ( .B(n22917), .A(n22918), .Z(n22915) );
  XOR U23180 ( .A(n17391), .B(n22919), .Z(n22912) );
  XOR U23181 ( .A(n19171), .B(n15662), .Z(n22919) );
  XNOR U23182 ( .A(n22920), .B(n22921), .Z(n15662) );
  NOR U23183 ( .A(n22922), .B(n22923), .Z(n22920) );
  XNOR U23184 ( .A(n22924), .B(n22925), .Z(n19171) );
  NOR U23185 ( .A(n22926), .B(n22927), .Z(n22924) );
  XNOR U23186 ( .A(n22928), .B(n22929), .Z(n17391) );
  ANDN U23187 ( .B(n22930), .A(n22931), .Z(n22928) );
  IV U23188 ( .A(n16547), .Z(n14773) );
  XOR U23189 ( .A(n17522), .B(n20180), .Z(n16547) );
  XOR U23190 ( .A(n22932), .B(n18850), .Z(n20180) );
  ANDN U23191 ( .B(n20753), .A(n22933), .Z(n22932) );
  IV U23192 ( .A(n17647), .Z(n17522) );
  XNOR U23193 ( .A(n21209), .B(n22934), .Z(n17647) );
  XOR U23194 ( .A(n22935), .B(n22936), .Z(n21209) );
  XNOR U23195 ( .A(n17690), .B(n18605), .Z(n22936) );
  XNOR U23196 ( .A(n22937), .B(n18911), .Z(n18605) );
  XOR U23197 ( .A(n22938), .B(n21606), .Z(n18911) );
  ANDN U23198 ( .B(n20178), .A(n18912), .Z(n22937) );
  XOR U23199 ( .A(n22939), .B(n22940), .Z(n18912) );
  XNOR U23200 ( .A(n22941), .B(n20758), .Z(n17690) );
  XNOR U23201 ( .A(n22942), .B(n22943), .Z(n20758) );
  ANDN U23202 ( .B(n20184), .A(n20182), .Z(n22941) );
  XOR U23203 ( .A(n22944), .B(n22945), .Z(n20182) );
  XNOR U23204 ( .A(n17389), .B(n22946), .Z(n22935) );
  XOR U23205 ( .A(n17555), .B(n16114), .Z(n22946) );
  XNOR U23206 ( .A(n22947), .B(n20749), .Z(n16114) );
  XOR U23207 ( .A(n22948), .B(n22949), .Z(n20749) );
  ANDN U23208 ( .B(n20188), .A(n20186), .Z(n22947) );
  XOR U23209 ( .A(n22950), .B(n22951), .Z(n20186) );
  XNOR U23210 ( .A(n22952), .B(n18851), .Z(n17555) );
  XOR U23211 ( .A(n22953), .B(n22954), .Z(n18851) );
  XNOR U23212 ( .A(n22955), .B(n22534), .Z(n18850) );
  XNOR U23213 ( .A(n22956), .B(n19731), .Z(n17389) );
  XOR U23214 ( .A(n22957), .B(n22958), .Z(n19731) );
  ANDN U23215 ( .B(n20175), .A(n19730), .Z(n22956) );
  XOR U23216 ( .A(n22959), .B(n22960), .Z(n19730) );
  XOR U23217 ( .A(n22961), .B(n14769), .Z(n12248) );
  XOR U23218 ( .A(n19413), .B(n18798), .Z(n14769) );
  XNOR U23219 ( .A(n22962), .B(n22963), .Z(n19413) );
  AND U23220 ( .A(n22680), .B(n22679), .Z(n22962) );
  ANDN U23221 ( .B(n14770), .A(n16538), .Z(n22961) );
  XOR U23222 ( .A(n22197), .B(n18687), .Z(n16538) );
  XNOR U23223 ( .A(n20821), .B(n21905), .Z(n18687) );
  XNOR U23224 ( .A(n22964), .B(n22965), .Z(n21905) );
  XNOR U23225 ( .A(n15907), .B(n17649), .Z(n22965) );
  XNOR U23226 ( .A(n22966), .B(n22967), .Z(n17649) );
  XNOR U23227 ( .A(n22968), .B(n22969), .Z(n15907) );
  ANDN U23228 ( .B(n22970), .A(n22971), .Z(n22968) );
  XOR U23229 ( .A(n17641), .B(n22972), .Z(n22964) );
  XOR U23230 ( .A(n22973), .B(n15880), .Z(n22972) );
  XNOR U23231 ( .A(n22974), .B(n22975), .Z(n15880) );
  ANDN U23232 ( .B(n22189), .A(n22190), .Z(n22974) );
  XNOR U23233 ( .A(n22976), .B(n22977), .Z(n17641) );
  ANDN U23234 ( .B(n22199), .A(n22200), .Z(n22976) );
  XOR U23235 ( .A(n22978), .B(n22979), .Z(n20821) );
  XNOR U23236 ( .A(n18781), .B(n18975), .Z(n22979) );
  XNOR U23237 ( .A(n22980), .B(n22343), .Z(n18975) );
  ANDN U23238 ( .B(n19926), .A(n19976), .Z(n22980) );
  XNOR U23239 ( .A(n22981), .B(n22982), .Z(n19926) );
  XNOR U23240 ( .A(n22983), .B(n22355), .Z(n18781) );
  ANDN U23241 ( .B(n20835), .A(n19939), .Z(n22983) );
  XOR U23242 ( .A(n22984), .B(n22521), .Z(n19939) );
  XNOR U23243 ( .A(n15346), .B(n22985), .Z(n22978) );
  XNOR U23244 ( .A(n17787), .B(n18404), .Z(n22985) );
  XOR U23245 ( .A(n22986), .B(n22351), .Z(n18404) );
  NOR U23246 ( .A(n19978), .B(n19935), .Z(n22986) );
  XOR U23247 ( .A(n22987), .B(n22988), .Z(n19935) );
  XNOR U23248 ( .A(n22989), .B(n22348), .Z(n17787) );
  IV U23249 ( .A(n19931), .Z(n19973) );
  XOR U23250 ( .A(n22990), .B(n22991), .Z(n19931) );
  XOR U23251 ( .A(n22992), .B(n22993), .Z(n15346) );
  ANDN U23252 ( .B(n19922), .A(n19980), .Z(n22992) );
  XOR U23253 ( .A(n22645), .B(n22994), .Z(n19922) );
  XNOR U23254 ( .A(n22995), .B(n22970), .Z(n22197) );
  ANDN U23255 ( .B(n22971), .A(n22996), .Z(n22995) );
  XOR U23256 ( .A(n16809), .B(n22997), .Z(n14770) );
  IV U23257 ( .A(n17462), .Z(n16809) );
  XNOR U23258 ( .A(n22998), .B(n22999), .Z(n17462) );
  XOR U23259 ( .A(n17597), .B(n10065), .Z(n9258) );
  XNOR U23260 ( .A(n16253), .B(n17088), .Z(n10065) );
  XNOR U23261 ( .A(n23000), .B(n23001), .Z(n17088) );
  XNOR U23262 ( .A(n13009), .B(n12917), .Z(n23001) );
  XOR U23263 ( .A(n23002), .B(n13155), .Z(n12917) );
  XOR U23264 ( .A(n23003), .B(n15653), .Z(n13155) );
  XNOR U23265 ( .A(n23004), .B(n23005), .Z(n15653) );
  ANDN U23266 ( .B(n13964), .A(n19592), .Z(n23002) );
  XOR U23267 ( .A(n21326), .B(n17105), .Z(n19592) );
  XNOR U23268 ( .A(n23006), .B(n22164), .Z(n17105) );
  XNOR U23269 ( .A(n23007), .B(n23008), .Z(n22164) );
  XOR U23270 ( .A(n20637), .B(n18961), .Z(n23008) );
  XOR U23271 ( .A(n23009), .B(n20656), .Z(n18961) );
  NOR U23272 ( .A(n20969), .B(n20657), .Z(n23009) );
  IV U23273 ( .A(n23010), .Z(n20969) );
  XNOR U23274 ( .A(n23011), .B(n20643), .Z(n20637) );
  NOR U23275 ( .A(n20644), .B(n20973), .Z(n23011) );
  XOR U23276 ( .A(n23012), .B(n23013), .Z(n20973) );
  XOR U23277 ( .A(n23014), .B(n23015), .Z(n20644) );
  XOR U23278 ( .A(n17922), .B(n23016), .Z(n23007) );
  XOR U23279 ( .A(n19738), .B(n20605), .Z(n23016) );
  XNOR U23280 ( .A(n23017), .B(n20653), .Z(n20605) );
  ANDN U23281 ( .B(n20966), .A(n21331), .Z(n23017) );
  XOR U23282 ( .A(n23018), .B(n23019), .Z(n21331) );
  XNOR U23283 ( .A(n23020), .B(n23021), .Z(n20966) );
  XNOR U23284 ( .A(n23022), .B(n20660), .Z(n19738) );
  ANDN U23285 ( .B(n20976), .A(n20661), .Z(n23022) );
  XNOR U23286 ( .A(n23023), .B(n23024), .Z(n20661) );
  XOR U23287 ( .A(n23025), .B(n23026), .Z(n20976) );
  XOR U23288 ( .A(n23027), .B(n20647), .Z(n17922) );
  ANDN U23289 ( .B(n20648), .A(n21329), .Z(n23027) );
  XOR U23290 ( .A(n23028), .B(n23029), .Z(n21329) );
  XOR U23291 ( .A(n23030), .B(n23031), .Z(n20648) );
  XOR U23292 ( .A(n23032), .B(n20657), .Z(n21326) );
  XOR U23293 ( .A(n23033), .B(n23034), .Z(n20657) );
  ANDN U23294 ( .B(n20970), .A(n23010), .Z(n23032) );
  XOR U23295 ( .A(n23035), .B(n23036), .Z(n23010) );
  XNOR U23296 ( .A(n21015), .B(n18478), .Z(n13964) );
  XNOR U23297 ( .A(n23037), .B(n23038), .Z(n21015) );
  ANDN U23298 ( .B(n22798), .A(n22799), .Z(n23037) );
  XNOR U23299 ( .A(n23039), .B(n23040), .Z(n22799) );
  XNOR U23300 ( .A(n23041), .B(n13151), .Z(n13009) );
  XOR U23301 ( .A(n22416), .B(n19035), .Z(n13151) );
  IV U23302 ( .A(n17487), .Z(n19035) );
  XNOR U23303 ( .A(n22934), .B(n23042), .Z(n17487) );
  XOR U23304 ( .A(n23043), .B(n23044), .Z(n22934) );
  XNOR U23305 ( .A(n20197), .B(n18330), .Z(n23044) );
  XOR U23306 ( .A(n23045), .B(n20216), .Z(n18330) );
  XOR U23307 ( .A(n23046), .B(n22943), .Z(n20216) );
  AND U23308 ( .A(n22418), .B(n20217), .Z(n23045) );
  XOR U23309 ( .A(n23047), .B(n23048), .Z(n20217) );
  XOR U23310 ( .A(n23049), .B(n23050), .Z(n22418) );
  XOR U23311 ( .A(n23051), .B(n20769), .Z(n20197) );
  IV U23312 ( .A(n20221), .Z(n20769) );
  XOR U23313 ( .A(n23052), .B(n23053), .Z(n20221) );
  ANDN U23314 ( .B(n22498), .A(n20220), .Z(n23051) );
  XOR U23315 ( .A(n17585), .B(n23054), .Z(n23043) );
  XOR U23316 ( .A(n18800), .B(n17661), .Z(n23054) );
  XOR U23317 ( .A(n23055), .B(n20204), .Z(n17661) );
  XOR U23318 ( .A(n23056), .B(n23057), .Z(n20204) );
  ANDN U23319 ( .B(n22427), .A(n22426), .Z(n23055) );
  IV U23320 ( .A(n20203), .Z(n22426) );
  XNOR U23321 ( .A(n23058), .B(n23059), .Z(n20203) );
  XNOR U23322 ( .A(n21603), .B(n23060), .Z(n22427) );
  XNOR U23323 ( .A(n23061), .B(n20213), .Z(n18800) );
  XOR U23324 ( .A(n23062), .B(n23063), .Z(n20213) );
  ANDN U23325 ( .B(n20212), .A(n22424), .Z(n23061) );
  XOR U23326 ( .A(n23064), .B(n23065), .Z(n22424) );
  XNOR U23327 ( .A(n23066), .B(n23067), .Z(n20212) );
  XNOR U23328 ( .A(n23068), .B(n20207), .Z(n17585) );
  XOR U23329 ( .A(n23069), .B(n21584), .Z(n20207) );
  ANDN U23330 ( .B(n20208), .A(n22421), .Z(n23068) );
  XOR U23331 ( .A(n23070), .B(n22521), .Z(n22421) );
  XNOR U23332 ( .A(n23071), .B(n23072), .Z(n20208) );
  XOR U23333 ( .A(n23074), .B(n23075), .Z(n20220) );
  NOR U23334 ( .A(n20768), .B(n22498), .Z(n23073) );
  XOR U23335 ( .A(n23076), .B(n23077), .Z(n22498) );
  XOR U23336 ( .A(n23078), .B(n23079), .Z(n20768) );
  ANDN U23337 ( .B(n13960), .A(n15267), .Z(n23041) );
  XOR U23338 ( .A(n21510), .B(n23080), .Z(n15267) );
  XNOR U23339 ( .A(n23081), .B(n23082), .Z(n21510) );
  ANDN U23340 ( .B(n23083), .A(n21781), .Z(n23081) );
  XNOR U23341 ( .A(n23084), .B(n17958), .Z(n13960) );
  XNOR U23342 ( .A(n22333), .B(n21666), .Z(n17958) );
  XNOR U23343 ( .A(n23085), .B(n23086), .Z(n21666) );
  XNOR U23344 ( .A(n16823), .B(n22902), .Z(n23086) );
  XNOR U23345 ( .A(n23087), .B(n23088), .Z(n22902) );
  ANDN U23346 ( .B(n23089), .A(n21919), .Z(n23087) );
  IV U23347 ( .A(n23090), .Z(n21919) );
  XNOR U23348 ( .A(n23091), .B(n23092), .Z(n16823) );
  ANDN U23349 ( .B(n21913), .A(n23093), .Z(n23091) );
  XOR U23350 ( .A(n19832), .B(n23094), .Z(n23085) );
  XOR U23351 ( .A(n19099), .B(n23095), .Z(n23094) );
  XNOR U23352 ( .A(n23096), .B(n23097), .Z(n19099) );
  NOR U23353 ( .A(n23098), .B(n23099), .Z(n23096) );
  XOR U23354 ( .A(n23100), .B(n23101), .Z(n19832) );
  NOR U23355 ( .A(n21923), .B(n23102), .Z(n23100) );
  XOR U23356 ( .A(n23103), .B(n23104), .Z(n22333) );
  XOR U23357 ( .A(n17144), .B(n18894), .Z(n23104) );
  XNOR U23358 ( .A(n23105), .B(n22201), .Z(n18894) );
  ANDN U23359 ( .B(n23106), .A(n22977), .Z(n23105) );
  XNOR U23360 ( .A(n23107), .B(n23108), .Z(n17144) );
  AND U23361 ( .A(n23109), .B(n23110), .Z(n23107) );
  XOR U23362 ( .A(n18957), .B(n23111), .Z(n23103) );
  XOR U23363 ( .A(n19314), .B(n19556), .Z(n23111) );
  XNOR U23364 ( .A(n23112), .B(n23113), .Z(n19556) );
  NOR U23365 ( .A(n22975), .B(n23114), .Z(n23112) );
  IV U23366 ( .A(n23115), .Z(n22975) );
  XNOR U23367 ( .A(n23116), .B(n22204), .Z(n19314) );
  NOR U23368 ( .A(n23117), .B(n22967), .Z(n23116) );
  XOR U23369 ( .A(n23118), .B(n22996), .Z(n18957) );
  XNOR U23370 ( .A(n10755), .B(n23120), .Z(n23000) );
  XNOR U23371 ( .A(n11431), .B(n13948), .Z(n23120) );
  XNOR U23372 ( .A(n23121), .B(n13141), .Z(n13948) );
  XOR U23373 ( .A(n21763), .B(n16674), .Z(n13141) );
  XOR U23374 ( .A(n19257), .B(n22658), .Z(n16674) );
  XNOR U23375 ( .A(n23122), .B(n23123), .Z(n22658) );
  XOR U23376 ( .A(n20836), .B(n18564), .Z(n23123) );
  XNOR U23377 ( .A(n23124), .B(n22850), .Z(n18564) );
  ANDN U23378 ( .B(n21770), .A(n21771), .Z(n23124) );
  XOR U23379 ( .A(n23125), .B(n22853), .Z(n20836) );
  AND U23380 ( .A(n21758), .B(n21756), .Z(n23125) );
  XOR U23381 ( .A(n20999), .B(n23126), .Z(n23122) );
  XOR U23382 ( .A(n18645), .B(n23127), .Z(n23126) );
  XNOR U23383 ( .A(n23128), .B(n22844), .Z(n18645) );
  ANDN U23384 ( .B(n23129), .A(n23130), .Z(n23128) );
  XNOR U23385 ( .A(n23131), .B(n22839), .Z(n20999) );
  AND U23386 ( .A(n21768), .B(n21766), .Z(n23131) );
  XOR U23387 ( .A(n23132), .B(n23133), .Z(n19257) );
  XNOR U23388 ( .A(n16995), .B(n16519), .Z(n23133) );
  XOR U23389 ( .A(n23134), .B(n22827), .Z(n16519) );
  NOR U23390 ( .A(n20115), .B(n20114), .Z(n23134) );
  XOR U23391 ( .A(n23135), .B(n23136), .Z(n20115) );
  XNOR U23392 ( .A(n23137), .B(n22817), .Z(n16995) );
  NOR U23393 ( .A(n22268), .B(n20118), .Z(n23137) );
  XNOR U23394 ( .A(n23138), .B(n23139), .Z(n22268) );
  XOR U23395 ( .A(n19394), .B(n23140), .Z(n23132) );
  XNOR U23396 ( .A(n19876), .B(n17575), .Z(n23140) );
  XNOR U23397 ( .A(n23141), .B(n22831), .Z(n17575) );
  NOR U23398 ( .A(n20105), .B(n20106), .Z(n23141) );
  XNOR U23399 ( .A(n23142), .B(n23143), .Z(n20106) );
  XOR U23400 ( .A(n23144), .B(n22835), .Z(n19876) );
  NOR U23401 ( .A(n20111), .B(n20110), .Z(n23144) );
  XNOR U23402 ( .A(n23145), .B(n23146), .Z(n20111) );
  XNOR U23403 ( .A(n23147), .B(n22821), .Z(n19394) );
  ANDN U23404 ( .B(n23148), .A(n22264), .Z(n23147) );
  XOR U23405 ( .A(n23149), .B(n23150), .Z(n22264) );
  XOR U23406 ( .A(n23151), .B(n23130), .Z(n21763) );
  NOR U23407 ( .A(n23129), .B(n22842), .Z(n23151) );
  ANDN U23408 ( .B(n13953), .A(n15259), .Z(n23121) );
  IV U23409 ( .A(n23152), .Z(n15259) );
  XNOR U23410 ( .A(n23153), .B(n13146), .Z(n11431) );
  XOR U23411 ( .A(n19688), .B(n19551), .Z(n13146) );
  XNOR U23412 ( .A(n23156), .B(n22083), .Z(n19688) );
  NOR U23413 ( .A(n19571), .B(n19572), .Z(n23156) );
  NOR U23414 ( .A(n15250), .B(n13962), .Z(n23153) );
  XNOR U23415 ( .A(n23157), .B(n18557), .Z(n13962) );
  XNOR U23416 ( .A(n23158), .B(n23159), .Z(n21507) );
  XOR U23417 ( .A(n18897), .B(n18519), .Z(n23159) );
  XNOR U23418 ( .A(n23160), .B(n23161), .Z(n18519) );
  ANDN U23419 ( .B(n23162), .A(n23163), .Z(n23160) );
  XOR U23420 ( .A(n23164), .B(n23165), .Z(n18897) );
  ANDN U23421 ( .B(n23166), .A(n23167), .Z(n23164) );
  XNOR U23422 ( .A(n23168), .B(n23169), .Z(n23158) );
  XNOR U23423 ( .A(n18860), .B(n17698), .Z(n23169) );
  XOR U23424 ( .A(n23170), .B(n23171), .Z(n17698) );
  ANDN U23425 ( .B(n23172), .A(n23173), .Z(n23170) );
  NOR U23426 ( .A(n23176), .B(n23177), .Z(n23174) );
  IV U23427 ( .A(n23178), .Z(n23176) );
  IV U23428 ( .A(n17599), .Z(n15250) );
  XOR U23429 ( .A(n23180), .B(n17546), .Z(n17599) );
  XNOR U23430 ( .A(n23181), .B(n13956), .Z(n10755) );
  IV U23431 ( .A(n14513), .Z(n13956) );
  XNOR U23432 ( .A(n23182), .B(n16516), .Z(n14513) );
  XOR U23433 ( .A(n22579), .B(n19960), .Z(n16516) );
  XNOR U23434 ( .A(n23183), .B(n23184), .Z(n19960) );
  XOR U23435 ( .A(n19380), .B(n17547), .Z(n23184) );
  XNOR U23436 ( .A(n23185), .B(n22927), .Z(n17547) );
  ANDN U23437 ( .B(n23186), .A(n23187), .Z(n23185) );
  XNOR U23438 ( .A(n23188), .B(n23189), .Z(n19380) );
  ANDN U23439 ( .B(n23190), .A(n23191), .Z(n23188) );
  XNOR U23440 ( .A(n17906), .B(n23192), .Z(n23183) );
  XNOR U23441 ( .A(n19706), .B(n19075), .Z(n23192) );
  XNOR U23442 ( .A(n23193), .B(n22918), .Z(n19075) );
  NOR U23443 ( .A(n23194), .B(n23195), .Z(n23193) );
  XNOR U23444 ( .A(n23196), .B(n22923), .Z(n19706) );
  ANDN U23445 ( .B(n23197), .A(n23198), .Z(n23196) );
  XNOR U23446 ( .A(n23199), .B(n23200), .Z(n17906) );
  ANDN U23447 ( .B(n23201), .A(n23202), .Z(n23199) );
  XNOR U23448 ( .A(n23203), .B(n23204), .Z(n22579) );
  XOR U23449 ( .A(n19732), .B(n22445), .Z(n23204) );
  XOR U23450 ( .A(n23205), .B(n23206), .Z(n22445) );
  XNOR U23451 ( .A(n23209), .B(n22464), .Z(n19732) );
  AND U23452 ( .A(n22465), .B(n23210), .Z(n23209) );
  XOR U23453 ( .A(n17097), .B(n23211), .Z(n23203) );
  XNOR U23454 ( .A(n19484), .B(n19129), .Z(n23211) );
  XOR U23455 ( .A(n23212), .B(n22450), .Z(n19129) );
  ANDN U23456 ( .B(n23213), .A(n22451), .Z(n23212) );
  XOR U23457 ( .A(n23214), .B(n22454), .Z(n19484) );
  IV U23458 ( .A(n23216), .Z(n22455) );
  XOR U23459 ( .A(n23217), .B(n22460), .Z(n17097) );
  ANDN U23460 ( .B(n23218), .A(n22461), .Z(n23217) );
  AND U23461 ( .A(n15263), .B(n13957), .Z(n23181) );
  XNOR U23462 ( .A(n18053), .B(n23219), .Z(n13957) );
  IV U23463 ( .A(n17237), .Z(n18053) );
  XNOR U23464 ( .A(n23220), .B(n19563), .Z(n17237) );
  XNOR U23465 ( .A(n23221), .B(n23222), .Z(n19563) );
  XOR U23466 ( .A(n19423), .B(n19681), .Z(n23222) );
  XNOR U23467 ( .A(n23223), .B(n20802), .Z(n19681) );
  IV U23468 ( .A(n23224), .Z(n20802) );
  ANDN U23469 ( .B(n20803), .A(n23225), .Z(n23223) );
  XNOR U23470 ( .A(n23226), .B(n23227), .Z(n19423) );
  ANDN U23471 ( .B(n23228), .A(n23229), .Z(n23226) );
  XOR U23472 ( .A(n19130), .B(n23230), .Z(n23221) );
  XOR U23473 ( .A(n17208), .B(n18396), .Z(n23230) );
  XNOR U23474 ( .A(n23231), .B(n20806), .Z(n18396) );
  IV U23475 ( .A(n23232), .Z(n20806) );
  ANDN U23476 ( .B(n20807), .A(n23233), .Z(n23231) );
  XNOR U23477 ( .A(n23234), .B(n20810), .Z(n17208) );
  ANDN U23478 ( .B(n20811), .A(n23235), .Z(n23234) );
  XNOR U23479 ( .A(n23236), .B(n20798), .Z(n19130) );
  IV U23480 ( .A(n23237), .Z(n20798) );
  ANDN U23481 ( .B(n23238), .A(n20797), .Z(n23236) );
  XOR U23482 ( .A(n20739), .B(n17622), .Z(n15263) );
  IV U23483 ( .A(n19374), .Z(n17622) );
  XNOR U23484 ( .A(n19955), .B(n23239), .Z(n19374) );
  XOR U23485 ( .A(n23240), .B(n23241), .Z(n19955) );
  XOR U23486 ( .A(n17834), .B(n22098), .Z(n23241) );
  XOR U23487 ( .A(n23242), .B(n22116), .Z(n22098) );
  AND U23488 ( .A(n20728), .B(n20729), .Z(n23242) );
  XOR U23489 ( .A(n23243), .B(n23244), .Z(n20728) );
  XNOR U23490 ( .A(n23245), .B(n23246), .Z(n17834) );
  ANDN U23491 ( .B(n20713), .A(n20711), .Z(n23245) );
  XNOR U23492 ( .A(n17509), .B(n23247), .Z(n23240) );
  XOR U23493 ( .A(n16402), .B(n15536), .Z(n23247) );
  XNOR U23494 ( .A(n23248), .B(n22119), .Z(n15536) );
  ANDN U23495 ( .B(n20724), .A(n20726), .Z(n23248) );
  XNOR U23496 ( .A(n23249), .B(n23250), .Z(n20724) );
  XNOR U23497 ( .A(n23251), .B(n22128), .Z(n16402) );
  ANDN U23498 ( .B(n20717), .A(n20715), .Z(n23251) );
  XOR U23499 ( .A(n23252), .B(n23253), .Z(n20715) );
  XOR U23500 ( .A(n23254), .B(n22125), .Z(n17509) );
  ANDN U23501 ( .B(n20722), .A(n22124), .Z(n23254) );
  IV U23502 ( .A(n20720), .Z(n22124) );
  XNOR U23503 ( .A(n23255), .B(n22790), .Z(n20720) );
  XNOR U23504 ( .A(n23256), .B(n23257), .Z(n20739) );
  ANDN U23505 ( .B(n20552), .A(n23258), .Z(n23256) );
  XOR U23506 ( .A(n23259), .B(n23260), .Z(n16253) );
  XOR U23507 ( .A(n11718), .B(n14395), .Z(n23260) );
  XOR U23508 ( .A(n23261), .B(n14401), .Z(n14395) );
  XOR U23509 ( .A(n18302), .B(n23262), .Z(n14401) );
  IV U23510 ( .A(n18004), .Z(n18302) );
  XOR U23511 ( .A(n20601), .B(n19466), .Z(n18004) );
  XOR U23512 ( .A(n23263), .B(n23264), .Z(n19466) );
  XNOR U23513 ( .A(n20595), .B(n18437), .Z(n23264) );
  XNOR U23514 ( .A(n23265), .B(n23266), .Z(n18437) );
  NOR U23515 ( .A(n23267), .B(n23268), .Z(n23265) );
  XNOR U23516 ( .A(n23269), .B(n23270), .Z(n20595) );
  XOR U23517 ( .A(n23271), .B(n23272), .Z(n23270) );
  NAND U23518 ( .A(n23273), .B(n23274), .Z(n23272) );
  ANDN U23519 ( .B(n11417), .A(rc_i[1]), .Z(n23271) );
  XOR U23520 ( .A(n18867), .B(n23275), .Z(n23263) );
  XOR U23521 ( .A(n18783), .B(n17499), .Z(n23275) );
  XNOR U23522 ( .A(n23276), .B(n23277), .Z(n17499) );
  ANDN U23523 ( .B(n23278), .A(n23279), .Z(n23276) );
  XNOR U23524 ( .A(n23280), .B(n23281), .Z(n18783) );
  AND U23525 ( .A(n23282), .B(n23283), .Z(n23280) );
  XNOR U23526 ( .A(n23284), .B(n23285), .Z(n18867) );
  ANDN U23527 ( .B(n23286), .A(n23287), .Z(n23284) );
  XOR U23528 ( .A(n23288), .B(n23289), .Z(n20601) );
  XNOR U23529 ( .A(n23290), .B(n18948), .Z(n23289) );
  XOR U23530 ( .A(n23291), .B(n23172), .Z(n18948) );
  ANDN U23531 ( .B(n23292), .A(n23293), .Z(n23291) );
  XOR U23532 ( .A(n19611), .B(n23294), .Z(n23288) );
  XNOR U23533 ( .A(n22486), .B(n18032), .Z(n23294) );
  XOR U23534 ( .A(n23295), .B(n23167), .Z(n18032) );
  ANDN U23535 ( .B(n23296), .A(n23297), .Z(n23295) );
  XOR U23536 ( .A(n23298), .B(n23178), .Z(n22486) );
  ANDN U23537 ( .B(n23299), .A(n23300), .Z(n23298) );
  XNOR U23538 ( .A(n23301), .B(n23162), .Z(n19611) );
  ANDN U23539 ( .B(n14841), .A(n17807), .Z(n23261) );
  XOR U23540 ( .A(n19414), .B(n18798), .Z(n17807) );
  XOR U23541 ( .A(n19676), .B(n22585), .Z(n18798) );
  XNOR U23542 ( .A(n23304), .B(n23305), .Z(n22585) );
  XNOR U23543 ( .A(n17394), .B(n23306), .Z(n23305) );
  XOR U23544 ( .A(n23307), .B(n21851), .Z(n17394) );
  ANDN U23545 ( .B(n23308), .A(n23309), .Z(n23307) );
  XOR U23546 ( .A(n18201), .B(n23310), .Z(n23304) );
  XOR U23547 ( .A(n18290), .B(n23311), .Z(n23310) );
  XNOR U23548 ( .A(n23312), .B(n21848), .Z(n18290) );
  ANDN U23549 ( .B(n21285), .A(n23313), .Z(n23312) );
  XNOR U23550 ( .A(n23314), .B(n21846), .Z(n18201) );
  NOR U23551 ( .A(n21289), .B(n23315), .Z(n23314) );
  IV U23552 ( .A(n23316), .Z(n21289) );
  XOR U23553 ( .A(n23317), .B(n23318), .Z(n19676) );
  XNOR U23554 ( .A(n19387), .B(n18152), .Z(n23318) );
  XNOR U23555 ( .A(n23319), .B(n20503), .Z(n18152) );
  NOR U23556 ( .A(n22963), .B(n22679), .Z(n23319) );
  XNOR U23557 ( .A(n23320), .B(n23321), .Z(n22679) );
  IV U23558 ( .A(n20502), .Z(n22963) );
  XOR U23559 ( .A(n23322), .B(n23323), .Z(n20502) );
  XNOR U23560 ( .A(n23324), .B(n21855), .Z(n19387) );
  AND U23561 ( .A(n19416), .B(n19418), .Z(n23324) );
  XNOR U23562 ( .A(n23325), .B(n21368), .Z(n19418) );
  XOR U23563 ( .A(n23326), .B(n23327), .Z(n19416) );
  XNOR U23564 ( .A(n20496), .B(n23328), .Z(n23317) );
  XOR U23565 ( .A(n18015), .B(n19249), .Z(n23328) );
  XNOR U23566 ( .A(n23329), .B(n20512), .Z(n19249) );
  ANDN U23567 ( .B(n22672), .A(n20513), .Z(n23329) );
  XOR U23568 ( .A(n23330), .B(n20506), .Z(n18015) );
  NOR U23569 ( .A(n20507), .B(n21041), .Z(n23330) );
  XNOR U23570 ( .A(n23331), .B(n21833), .Z(n21041) );
  XOR U23571 ( .A(n23332), .B(n23333), .Z(n20507) );
  XNOR U23572 ( .A(n23334), .B(n20516), .Z(n20496) );
  ANDN U23573 ( .B(n19411), .A(n19409), .Z(n23334) );
  XOR U23574 ( .A(n23335), .B(n23336), .Z(n19409) );
  XNOR U23575 ( .A(n22217), .B(n23337), .Z(n19411) );
  XOR U23576 ( .A(n23338), .B(n20513), .Z(n19414) );
  XOR U23577 ( .A(n23339), .B(n22391), .Z(n20513) );
  ANDN U23578 ( .B(n22673), .A(n22672), .Z(n23338) );
  XOR U23579 ( .A(n23340), .B(n22504), .Z(n22672) );
  XNOR U23580 ( .A(n21016), .B(n18445), .Z(n14841) );
  IV U23581 ( .A(n18478), .Z(n18445) );
  XOR U23582 ( .A(n23341), .B(n23342), .Z(n18478) );
  XOR U23583 ( .A(n23343), .B(n23344), .Z(n21016) );
  NOR U23584 ( .A(n21987), .B(n22802), .Z(n23343) );
  IV U23585 ( .A(n22803), .Z(n21987) );
  XOR U23586 ( .A(n23345), .B(n23346), .Z(n22803) );
  XNOR U23587 ( .A(n23347), .B(n19267), .Z(n11718) );
  XNOR U23588 ( .A(n18596), .B(n23348), .Z(n19267) );
  IV U23589 ( .A(n22581), .Z(n18596) );
  XNOR U23590 ( .A(n20385), .B(n20940), .Z(n22581) );
  XOR U23591 ( .A(n23349), .B(n23350), .Z(n20940) );
  XNOR U23592 ( .A(n19174), .B(n17431), .Z(n23350) );
  XOR U23593 ( .A(n23351), .B(n22576), .Z(n17431) );
  ANDN U23594 ( .B(n23352), .A(n23353), .Z(n23351) );
  XOR U23595 ( .A(n23354), .B(n22558), .Z(n19174) );
  ANDN U23596 ( .B(n23355), .A(n23356), .Z(n23354) );
  XOR U23597 ( .A(n18493), .B(n23357), .Z(n23349) );
  XNOR U23598 ( .A(n23358), .B(n23359), .Z(n23357) );
  XOR U23599 ( .A(n23360), .B(n22563), .Z(n18493) );
  ANDN U23600 ( .B(n23361), .A(n23362), .Z(n23360) );
  XOR U23601 ( .A(n23363), .B(n23364), .Z(n20385) );
  XOR U23602 ( .A(n23003), .B(n21144), .Z(n23364) );
  XOR U23603 ( .A(n23365), .B(n23366), .Z(n21144) );
  ANDN U23604 ( .B(n23367), .A(n23368), .Z(n23365) );
  XOR U23605 ( .A(n23369), .B(n22601), .Z(n23003) );
  ANDN U23606 ( .B(n23370), .A(n23371), .Z(n23369) );
  XOR U23607 ( .A(n18715), .B(n23372), .Z(n23363) );
  XNOR U23608 ( .A(n18063), .B(n15652), .Z(n23372) );
  XOR U23609 ( .A(n23373), .B(n22598), .Z(n15652) );
  ANDN U23610 ( .B(n23374), .A(n23375), .Z(n23373) );
  XNOR U23611 ( .A(n23376), .B(n22591), .Z(n18063) );
  IV U23612 ( .A(n23377), .Z(n22591) );
  ANDN U23613 ( .B(n23378), .A(n23379), .Z(n23376) );
  XNOR U23614 ( .A(n23380), .B(n23381), .Z(n18715) );
  ANDN U23615 ( .B(n17803), .A(n14844), .Z(n23347) );
  XNOR U23616 ( .A(n23384), .B(n17546), .Z(n14844) );
  XOR U23617 ( .A(n23385), .B(n23386), .Z(n17546) );
  XNOR U23618 ( .A(n15674), .B(n21959), .Z(n17803) );
  XNOR U23619 ( .A(n23387), .B(n23388), .Z(n21959) );
  ANDN U23620 ( .B(n23389), .A(n23390), .Z(n23387) );
  XOR U23621 ( .A(n20258), .B(n19419), .Z(n15674) );
  XOR U23622 ( .A(n23391), .B(n23392), .Z(n19419) );
  XNOR U23623 ( .A(n19545), .B(n18450), .Z(n23392) );
  XOR U23624 ( .A(n23393), .B(n22360), .Z(n18450) );
  ANDN U23625 ( .B(n23394), .A(n22685), .Z(n23393) );
  XNOR U23626 ( .A(n23395), .B(n20452), .Z(n19545) );
  AND U23627 ( .A(n22699), .B(n22698), .Z(n23395) );
  XOR U23628 ( .A(n19675), .B(n23396), .Z(n23391) );
  XOR U23629 ( .A(n17505), .B(n19443), .Z(n23396) );
  XNOR U23630 ( .A(n23397), .B(n23398), .Z(n19443) );
  XNOR U23631 ( .A(n23399), .B(n23400), .Z(n17505) );
  XNOR U23632 ( .A(n23401), .B(n20462), .Z(n19675) );
  IV U23633 ( .A(n23402), .Z(n20462) );
  NOR U23634 ( .A(n22687), .B(n22688), .Z(n23401) );
  XOR U23635 ( .A(n23403), .B(n23404), .Z(n20258) );
  XOR U23636 ( .A(n23405), .B(n17934), .Z(n23404) );
  XNOR U23637 ( .A(n23406), .B(n23407), .Z(n17934) );
  ANDN U23638 ( .B(n21967), .A(n21966), .Z(n23406) );
  XOR U23639 ( .A(n17897), .B(n23408), .Z(n23403) );
  XNOR U23640 ( .A(n18555), .B(n16762), .Z(n23408) );
  XNOR U23641 ( .A(n23409), .B(n23410), .Z(n16762) );
  XNOR U23642 ( .A(n23411), .B(n23412), .Z(n18555) );
  ANDN U23643 ( .B(n21957), .A(n23413), .Z(n23411) );
  XNOR U23644 ( .A(n23414), .B(n23415), .Z(n17897) );
  ANDN U23645 ( .B(n21964), .A(n23416), .Z(n23414) );
  XOR U23646 ( .A(n10970), .B(n23417), .Z(n23259) );
  XOR U23647 ( .A(n12966), .B(n11367), .Z(n23417) );
  XNOR U23648 ( .A(n23418), .B(n14414), .Z(n11367) );
  XNOR U23649 ( .A(n16313), .B(n22121), .Z(n14414) );
  XOR U23650 ( .A(n23419), .B(n23420), .Z(n22121) );
  ANDN U23651 ( .B(n20711), .A(n23246), .Z(n23419) );
  IV U23652 ( .A(n23421), .Z(n23246) );
  XOR U23653 ( .A(n23422), .B(n23423), .Z(n20711) );
  XNOR U23654 ( .A(n23424), .B(n20380), .Z(n16313) );
  XOR U23655 ( .A(n23425), .B(n23426), .Z(n20380) );
  XOR U23656 ( .A(n18811), .B(n21456), .Z(n23426) );
  XNOR U23657 ( .A(n23427), .B(n20725), .Z(n21456) );
  ANDN U23658 ( .B(n22119), .A(n22118), .Z(n23427) );
  XNOR U23659 ( .A(n23428), .B(n23429), .Z(n22119) );
  XNOR U23660 ( .A(n23430), .B(n20716), .Z(n18811) );
  ANDN U23661 ( .B(n22128), .A(n22127), .Z(n23430) );
  XNOR U23662 ( .A(n23431), .B(n23432), .Z(n22128) );
  XNOR U23663 ( .A(n17591), .B(n23433), .Z(n23425) );
  XOR U23664 ( .A(n16731), .B(n18200), .Z(n23433) );
  XNOR U23665 ( .A(n23434), .B(n20730), .Z(n18200) );
  ANDN U23666 ( .B(n22115), .A(n22116), .Z(n23434) );
  XOR U23667 ( .A(n23435), .B(n23436), .Z(n22116) );
  XNOR U23668 ( .A(n23437), .B(n20712), .Z(n16731) );
  NOR U23669 ( .A(n23421), .B(n23420), .Z(n23437) );
  XOR U23670 ( .A(n23438), .B(n23439), .Z(n23421) );
  XNOR U23671 ( .A(n23440), .B(n20721), .Z(n17591) );
  ANDN U23672 ( .B(n22123), .A(n22125), .Z(n23440) );
  XOR U23673 ( .A(n23441), .B(n23442), .Z(n22125) );
  AND U23674 ( .A(n14848), .B(n14415), .Z(n23418) );
  XOR U23675 ( .A(n17395), .B(n23311), .Z(n14415) );
  XNOR U23676 ( .A(n23443), .B(n21840), .Z(n23311) );
  ANDN U23677 ( .B(n23444), .A(n21295), .Z(n23443) );
  XOR U23678 ( .A(n17272), .B(n21373), .Z(n14848) );
  XNOR U23679 ( .A(n23445), .B(n23446), .Z(n21373) );
  NOR U23680 ( .A(n19743), .B(n20418), .Z(n23445) );
  XOR U23681 ( .A(n23447), .B(n21710), .Z(n19743) );
  XNOR U23682 ( .A(n23220), .B(n23448), .Z(n17272) );
  XOR U23683 ( .A(n23449), .B(n23450), .Z(n23220) );
  XNOR U23684 ( .A(n20790), .B(n19721), .Z(n23450) );
  XNOR U23685 ( .A(n23451), .B(n23452), .Z(n19721) );
  XNOR U23686 ( .A(n23455), .B(n23456), .Z(n20790) );
  ANDN U23687 ( .B(n23457), .A(n23458), .Z(n23455) );
  XOR U23688 ( .A(n20705), .B(n23459), .Z(n23449) );
  XOR U23689 ( .A(n17135), .B(n18428), .Z(n23459) );
  XOR U23690 ( .A(n23460), .B(n23461), .Z(n18428) );
  NOR U23691 ( .A(n23462), .B(n23463), .Z(n23460) );
  XNOR U23692 ( .A(n23464), .B(n23465), .Z(n17135) );
  AND U23693 ( .A(n23466), .B(n23467), .Z(n23464) );
  XNOR U23694 ( .A(n23468), .B(n23469), .Z(n20705) );
  ANDN U23695 ( .B(n23470), .A(n23471), .Z(n23468) );
  XNOR U23696 ( .A(n23472), .B(n14407), .Z(n12966) );
  XOR U23697 ( .A(n19295), .B(n22069), .Z(n14407) );
  XOR U23698 ( .A(n23473), .B(n23474), .Z(n22069) );
  ANDN U23699 ( .B(n23475), .A(n23476), .Z(n23473) );
  IV U23700 ( .A(n14162), .Z(n19295) );
  XOR U23701 ( .A(n18667), .B(n23477), .Z(n14162) );
  XOR U23702 ( .A(n23478), .B(n23479), .Z(n18667) );
  XOR U23703 ( .A(n18858), .B(n18711), .Z(n23479) );
  XOR U23704 ( .A(n23480), .B(n22163), .Z(n18711) );
  NOR U23705 ( .A(n22043), .B(n22042), .Z(n23480) );
  XOR U23706 ( .A(n23481), .B(n23482), .Z(n22042) );
  XNOR U23707 ( .A(n23483), .B(n22159), .Z(n18858) );
  NOR U23708 ( .A(n22160), .B(n22052), .Z(n23483) );
  XOR U23709 ( .A(n23484), .B(n23485), .Z(n22160) );
  XOR U23710 ( .A(n19236), .B(n23486), .Z(n23478) );
  XOR U23711 ( .A(n21271), .B(n22132), .Z(n23486) );
  XNOR U23712 ( .A(n23487), .B(n22152), .Z(n22132) );
  XOR U23713 ( .A(n23488), .B(n23489), .Z(n22055) );
  XNOR U23714 ( .A(n23490), .B(n22149), .Z(n21271) );
  ANDN U23715 ( .B(n22047), .A(n22049), .Z(n23490) );
  XOR U23716 ( .A(n23491), .B(n21368), .Z(n22047) );
  XNOR U23717 ( .A(n23492), .B(n22156), .Z(n19236) );
  ANDN U23718 ( .B(n22040), .A(n22038), .Z(n23492) );
  XOR U23719 ( .A(n23493), .B(n23494), .Z(n22038) );
  NOR U23720 ( .A(n17778), .B(n14406), .Z(n23472) );
  XOR U23721 ( .A(n17063), .B(n23495), .Z(n14406) );
  XNOR U23722 ( .A(n17974), .B(n20466), .Z(n17778) );
  XNOR U23723 ( .A(n23496), .B(n21640), .Z(n20466) );
  IV U23724 ( .A(n16367), .Z(n17974) );
  XOR U23725 ( .A(n23497), .B(n22659), .Z(n16367) );
  XNOR U23726 ( .A(n23498), .B(n23499), .Z(n22659) );
  XNOR U23727 ( .A(n19431), .B(n18946), .Z(n23499) );
  XNOR U23728 ( .A(n23500), .B(n23501), .Z(n18946) );
  NOR U23729 ( .A(n21659), .B(n21752), .Z(n23500) );
  XOR U23730 ( .A(n23502), .B(n23503), .Z(n21659) );
  XOR U23731 ( .A(n23504), .B(n21647), .Z(n19431) );
  ANDN U23732 ( .B(n21749), .A(n21646), .Z(n23504) );
  XOR U23733 ( .A(n23505), .B(n23506), .Z(n21646) );
  XOR U23734 ( .A(n19036), .B(n23507), .Z(n23498) );
  XNOR U23735 ( .A(n19457), .B(n18166), .Z(n23507) );
  XNOR U23736 ( .A(n23508), .B(n21663), .Z(n18166) );
  NOR U23737 ( .A(n22661), .B(n22663), .Z(n23508) );
  IV U23738 ( .A(n21664), .Z(n22661) );
  XNOR U23739 ( .A(n23509), .B(n23510), .Z(n21664) );
  XOR U23740 ( .A(n23511), .B(n21650), .Z(n19457) );
  ANDN U23741 ( .B(n21651), .A(n21740), .Z(n23511) );
  XOR U23742 ( .A(n23512), .B(n23513), .Z(n21651) );
  XNOR U23743 ( .A(n23514), .B(n21655), .Z(n19036) );
  XOR U23744 ( .A(n23515), .B(n23516), .Z(n21656) );
  XNOR U23745 ( .A(n23517), .B(n14410), .Z(n10970) );
  XOR U23746 ( .A(n18187), .B(n23518), .Z(n14410) );
  NOR U23747 ( .A(n17810), .B(n14837), .Z(n23517) );
  XNOR U23748 ( .A(n21917), .B(n18877), .Z(n14837) );
  IV U23749 ( .A(n17227), .Z(n18877) );
  XOR U23750 ( .A(n23519), .B(n23520), .Z(n17227) );
  XNOR U23751 ( .A(n23521), .B(n23098), .Z(n21917) );
  ANDN U23752 ( .B(n23522), .A(n23523), .Z(n23521) );
  IV U23753 ( .A(n14411), .Z(n17810) );
  XOR U23754 ( .A(n23524), .B(n16509), .Z(n14411) );
  XNOR U23755 ( .A(n22030), .B(n20488), .Z(n16509) );
  XNOR U23756 ( .A(n23525), .B(n23526), .Z(n20488) );
  XOR U23757 ( .A(n18230), .B(n19875), .Z(n23526) );
  XOR U23758 ( .A(n23527), .B(n22733), .Z(n19875) );
  AND U23759 ( .A(n22734), .B(n23528), .Z(n23527) );
  XNOR U23760 ( .A(n23529), .B(n23530), .Z(n18230) );
  ANDN U23761 ( .B(n23531), .A(n23532), .Z(n23529) );
  XOR U23762 ( .A(n21812), .B(n23533), .Z(n23525) );
  XOR U23763 ( .A(n20594), .B(n15634), .Z(n23533) );
  XOR U23764 ( .A(n23534), .B(n22743), .Z(n15634) );
  ANDN U23765 ( .B(n23535), .A(n22742), .Z(n23534) );
  XNOR U23766 ( .A(n23536), .B(n22746), .Z(n20594) );
  ANDN U23767 ( .B(n23537), .A(n22747), .Z(n23536) );
  XNOR U23768 ( .A(n23538), .B(n22738), .Z(n21812) );
  ANDN U23769 ( .B(n23539), .A(n22739), .Z(n23538) );
  XOR U23770 ( .A(n23540), .B(n23541), .Z(n22030) );
  XOR U23771 ( .A(n21387), .B(n18386), .Z(n23541) );
  XOR U23772 ( .A(n23542), .B(n22723), .Z(n18386) );
  XOR U23773 ( .A(n23544), .B(n22726), .Z(n21387) );
  AND U23774 ( .A(n23545), .B(n22727), .Z(n23544) );
  XOR U23775 ( .A(n22704), .B(n23546), .Z(n23540) );
  XNOR U23776 ( .A(n18889), .B(n18717), .Z(n23546) );
  XOR U23777 ( .A(n23547), .B(n22714), .Z(n18717) );
  ANDN U23778 ( .B(n23548), .A(n22713), .Z(n23547) );
  XNOR U23779 ( .A(n23549), .B(n22718), .Z(n18889) );
  AND U23780 ( .A(n22719), .B(n23550), .Z(n23549) );
  XNOR U23781 ( .A(n23551), .B(n23552), .Z(n22704) );
  ANDN U23782 ( .B(n22710), .A(n23553), .Z(n23551) );
  XNOR U23783 ( .A(n23554), .B(n13953), .Z(n17597) );
  XOR U23784 ( .A(n20367), .B(n16465), .Z(n13953) );
  IV U23785 ( .A(n18326), .Z(n16465) );
  XNOR U23786 ( .A(n23555), .B(n23556), .Z(n20367) );
  ANDN U23787 ( .B(n19881), .A(n19882), .Z(n23555) );
  XOR U23788 ( .A(n23557), .B(n23558), .Z(n19882) );
  ANDN U23789 ( .B(n13140), .A(n23152), .Z(n23554) );
  XOR U23790 ( .A(n17395), .B(n23306), .Z(n23152) );
  XNOR U23791 ( .A(n23559), .B(n21843), .Z(n23306) );
  NOR U23792 ( .A(n21299), .B(n23560), .Z(n23559) );
  XOR U23793 ( .A(n20497), .B(n23561), .Z(n17395) );
  XNOR U23794 ( .A(n23562), .B(n23563), .Z(n20497) );
  XOR U23795 ( .A(n17594), .B(n16962), .Z(n23563) );
  XNOR U23796 ( .A(n23564), .B(n21300), .Z(n16962) );
  XNOR U23797 ( .A(n23565), .B(n23566), .Z(n21300) );
  ANDN U23798 ( .B(n23560), .A(n21843), .Z(n23564) );
  XOR U23799 ( .A(n23567), .B(n23568), .Z(n21843) );
  XNOR U23800 ( .A(n23569), .B(n21291), .Z(n17594) );
  XOR U23801 ( .A(n23570), .B(n23571), .Z(n21291) );
  AND U23802 ( .A(n21846), .B(n23315), .Z(n23569) );
  XOR U23803 ( .A(n23572), .B(n23573), .Z(n21846) );
  XOR U23804 ( .A(n19981), .B(n23574), .Z(n23562) );
  XNOR U23805 ( .A(n19291), .B(n17336), .Z(n23574) );
  XNOR U23806 ( .A(n23575), .B(n21287), .Z(n17336) );
  XNOR U23807 ( .A(n23576), .B(n23577), .Z(n21287) );
  AND U23808 ( .A(n23313), .B(n21848), .Z(n23575) );
  XNOR U23809 ( .A(n23035), .B(n23578), .Z(n21848) );
  XOR U23810 ( .A(n21297), .B(n23579), .Z(n19291) );
  XOR U23811 ( .A(n23580), .B(n4407), .Z(n23579) );
  ANDN U23812 ( .B(n21840), .A(n23444), .Z(n23580) );
  XOR U23813 ( .A(n23581), .B(n23582), .Z(n21840) );
  XNOR U23814 ( .A(n23583), .B(n23584), .Z(n21297) );
  XNOR U23815 ( .A(n23585), .B(n21852), .Z(n19981) );
  NOR U23816 ( .A(n23308), .B(n21851), .Z(n23585) );
  XOR U23817 ( .A(n23586), .B(n23587), .Z(n21851) );
  XNOR U23818 ( .A(n18187), .B(n23588), .Z(n13140) );
  XNOR U23819 ( .A(n18935), .B(n21093), .Z(n18187) );
  XOR U23820 ( .A(n23589), .B(n23590), .Z(n21093) );
  XNOR U23821 ( .A(n19137), .B(n16300), .Z(n23590) );
  XNOR U23822 ( .A(n23591), .B(n21957), .Z(n16300) );
  XOR U23823 ( .A(n23592), .B(n23593), .Z(n21957) );
  ANDN U23824 ( .B(n21958), .A(n23594), .Z(n23591) );
  XNOR U23825 ( .A(n23595), .B(n21967), .Z(n19137) );
  XNOR U23826 ( .A(n23596), .B(n23597), .Z(n21967) );
  ANDN U23827 ( .B(n21968), .A(n23598), .Z(n23595) );
  XOR U23828 ( .A(n16383), .B(n23599), .Z(n23589) );
  XOR U23829 ( .A(n16473), .B(n17875), .Z(n23599) );
  XNOR U23830 ( .A(n23600), .B(n23389), .Z(n17875) );
  XNOR U23831 ( .A(n23601), .B(n23602), .Z(n23389) );
  ANDN U23832 ( .B(n23603), .A(n23604), .Z(n23600) );
  XNOR U23833 ( .A(n23605), .B(n21953), .Z(n16473) );
  AND U23834 ( .A(n23606), .B(n21954), .Z(n23605) );
  XNOR U23835 ( .A(n23607), .B(n21964), .Z(n16383) );
  XOR U23836 ( .A(n23608), .B(n22954), .Z(n21964) );
  NOR U23837 ( .A(n23609), .B(n21963), .Z(n23607) );
  XOR U23838 ( .A(n23610), .B(n23611), .Z(n18935) );
  XOR U23839 ( .A(n18050), .B(n17976), .Z(n23611) );
  XNOR U23840 ( .A(n23612), .B(n21944), .Z(n17976) );
  XNOR U23841 ( .A(n23613), .B(n22231), .Z(n21944) );
  NOR U23842 ( .A(n23614), .B(n23615), .Z(n23612) );
  XNOR U23843 ( .A(n23616), .B(n21948), .Z(n18050) );
  XOR U23844 ( .A(n23617), .B(n21710), .Z(n21948) );
  ANDN U23845 ( .B(n21947), .A(n23618), .Z(n23616) );
  XOR U23846 ( .A(n21930), .B(n23619), .Z(n23610) );
  XOR U23847 ( .A(n18659), .B(n18768), .Z(n23619) );
  XNOR U23848 ( .A(n23620), .B(n20263), .Z(n18768) );
  XOR U23849 ( .A(n23621), .B(n23013), .Z(n20263) );
  NOR U23850 ( .A(n23622), .B(n21934), .Z(n23620) );
  XNOR U23851 ( .A(n23623), .B(n21940), .Z(n18659) );
  NOR U23852 ( .A(n21941), .B(n23624), .Z(n23623) );
  XNOR U23853 ( .A(n23625), .B(n20274), .Z(n21930) );
  XOR U23854 ( .A(n23626), .B(n23627), .Z(n20274) );
  NOR U23855 ( .A(n23628), .B(n21936), .Z(n23625) );
  XNOR U23856 ( .A(n23629), .B(n6673), .Z(n2566) );
  XOR U23857 ( .A(n19474), .B(n9557), .Z(n6673) );
  IV U23858 ( .A(n12893), .Z(n9557) );
  XNOR U23859 ( .A(n16554), .B(n17252), .Z(n12893) );
  XNOR U23860 ( .A(n23630), .B(n23631), .Z(n17252) );
  XOR U23861 ( .A(n12523), .B(n13701), .Z(n23631) );
  XNOR U23862 ( .A(n23632), .B(n16690), .Z(n13701) );
  XNOR U23863 ( .A(n18070), .B(n23633), .Z(n16690) );
  IV U23864 ( .A(n18598), .Z(n18070) );
  XNOR U23865 ( .A(n20251), .B(n19594), .Z(n18598) );
  XNOR U23866 ( .A(n23634), .B(n23635), .Z(n19594) );
  XNOR U23867 ( .A(n23636), .B(n18276), .Z(n23635) );
  XNOR U23868 ( .A(n23637), .B(n23550), .Z(n18276) );
  ANDN U23869 ( .B(n23638), .A(n22717), .Z(n23637) );
  XNOR U23870 ( .A(n19665), .B(n23639), .Z(n23634) );
  XOR U23871 ( .A(n19308), .B(n18618), .Z(n23639) );
  XNOR U23872 ( .A(n23640), .B(n23543), .Z(n18618) );
  ANDN U23873 ( .B(n23641), .A(n22721), .Z(n23640) );
  IV U23874 ( .A(n23642), .Z(n22721) );
  XNOR U23875 ( .A(n23643), .B(n23548), .Z(n19308) );
  ANDN U23876 ( .B(n23644), .A(n22712), .Z(n23643) );
  XOR U23877 ( .A(n23645), .B(n23553), .Z(n19665) );
  ANDN U23878 ( .B(n23646), .A(n22708), .Z(n23645) );
  XOR U23879 ( .A(n23647), .B(n23648), .Z(n20251) );
  XOR U23880 ( .A(n19200), .B(n21347), .Z(n23648) );
  XOR U23881 ( .A(n23649), .B(n23539), .Z(n21347) );
  XNOR U23882 ( .A(n23651), .B(n23535), .Z(n19200) );
  XOR U23883 ( .A(n17295), .B(n23653), .Z(n23647) );
  XOR U23884 ( .A(n17550), .B(n15697), .Z(n23653) );
  XNOR U23885 ( .A(n23654), .B(n23528), .Z(n15697) );
  ANDN U23886 ( .B(n22732), .A(n23655), .Z(n23654) );
  XNOR U23887 ( .A(n23656), .B(n23537), .Z(n17550) );
  XOR U23888 ( .A(n23658), .B(n23531), .Z(n17295) );
  ANDN U23889 ( .B(n23659), .A(n23660), .Z(n23658) );
  ANDN U23890 ( .B(n15159), .A(n23661), .Z(n23632) );
  XOR U23891 ( .A(n23662), .B(n16700), .Z(n12523) );
  XOR U23892 ( .A(n18161), .B(n23663), .Z(n16700) );
  IV U23893 ( .A(n21532), .Z(n18161) );
  XOR U23894 ( .A(n23664), .B(n19167), .Z(n21532) );
  XNOR U23895 ( .A(n23665), .B(n23666), .Z(n19167) );
  XNOR U23896 ( .A(n19169), .B(n19028), .Z(n23666) );
  XNOR U23897 ( .A(n23667), .B(n23668), .Z(n19028) );
  ANDN U23898 ( .B(n23469), .A(n23669), .Z(n23667) );
  XOR U23899 ( .A(n23670), .B(n23671), .Z(n19169) );
  ANDN U23900 ( .B(n23461), .A(n23672), .Z(n23670) );
  XOR U23901 ( .A(n18786), .B(n23673), .Z(n23665) );
  XOR U23902 ( .A(n23674), .B(n20489), .Z(n23673) );
  XNOR U23903 ( .A(n23675), .B(n23676), .Z(n20489) );
  ANDN U23904 ( .B(n23677), .A(n23452), .Z(n23675) );
  XNOR U23905 ( .A(n23678), .B(n23679), .Z(n18786) );
  NOR U23906 ( .A(n23465), .B(n23680), .Z(n23678) );
  IV U23907 ( .A(n23681), .Z(n23465) );
  ANDN U23908 ( .B(n15145), .A(n19471), .Z(n23662) );
  IV U23909 ( .A(n16701), .Z(n19471) );
  XNOR U23910 ( .A(n18563), .B(n23127), .Z(n16701) );
  XNOR U23911 ( .A(n23682), .B(n22848), .Z(n23127) );
  ANDN U23912 ( .B(n21760), .A(n21762), .Z(n23682) );
  XOR U23913 ( .A(n23683), .B(n23684), .Z(n19877) );
  XNOR U23914 ( .A(n20359), .B(n17741), .Z(n23684) );
  XNOR U23915 ( .A(n23685), .B(n22269), .Z(n17741) );
  XOR U23916 ( .A(n23686), .B(n23687), .Z(n22269) );
  AND U23917 ( .A(n20118), .B(n22817), .Z(n23685) );
  XNOR U23918 ( .A(n23688), .B(n23689), .Z(n22817) );
  XOR U23919 ( .A(n23690), .B(n23691), .Z(n20118) );
  XNOR U23920 ( .A(n23692), .B(n22262), .Z(n20359) );
  XNOR U23921 ( .A(n23693), .B(n23013), .Z(n22262) );
  ANDN U23922 ( .B(n20110), .A(n22835), .Z(n23692) );
  XNOR U23923 ( .A(n23694), .B(n23695), .Z(n22835) );
  XOR U23924 ( .A(n22886), .B(n23696), .Z(n20110) );
  XOR U23925 ( .A(n18379), .B(n23697), .Z(n23683) );
  XNOR U23926 ( .A(n19282), .B(n17285), .Z(n23697) );
  XNOR U23927 ( .A(n23698), .B(n22826), .Z(n17285) );
  IV U23928 ( .A(n22274), .Z(n22826) );
  XOR U23929 ( .A(n23699), .B(n23700), .Z(n22274) );
  AND U23930 ( .A(n20114), .B(n22827), .Z(n23698) );
  XOR U23931 ( .A(n23701), .B(n23702), .Z(n22827) );
  XNOR U23932 ( .A(n23703), .B(n23704), .Z(n20114) );
  XOR U23933 ( .A(n23705), .B(n22265), .Z(n19282) );
  XNOR U23934 ( .A(n23706), .B(n23482), .Z(n22265) );
  ANDN U23935 ( .B(n22821), .A(n23148), .Z(n23705) );
  IV U23936 ( .A(n20101), .Z(n23148) );
  XNOR U23937 ( .A(n23707), .B(n23708), .Z(n20101) );
  XOR U23938 ( .A(n23709), .B(n23710), .Z(n22821) );
  XNOR U23939 ( .A(n23711), .B(n22271), .Z(n18379) );
  XNOR U23940 ( .A(n23712), .B(n23713), .Z(n22271) );
  AND U23941 ( .A(n22831), .B(n20105), .Z(n23711) );
  XNOR U23942 ( .A(n23714), .B(n23715), .Z(n20105) );
  XOR U23943 ( .A(n23716), .B(n22227), .Z(n22831) );
  XOR U23944 ( .A(n23717), .B(n23718), .Z(n19459) );
  XOR U23945 ( .A(n17963), .B(n17667), .Z(n23718) );
  NOR U23946 ( .A(n21766), .B(n22839), .Z(n23719) );
  XOR U23947 ( .A(n23720), .B(n23721), .Z(n22839) );
  XNOR U23948 ( .A(n23722), .B(n23710), .Z(n21766) );
  XNOR U23949 ( .A(n23723), .B(n22843), .Z(n17963) );
  ANDN U23950 ( .B(n23130), .A(n22844), .Z(n23723) );
  XNOR U23951 ( .A(n23724), .B(n23725), .Z(n22844) );
  XNOR U23952 ( .A(n23726), .B(n23727), .Z(n23130) );
  XNOR U23953 ( .A(n14998), .B(n23728), .Z(n23717) );
  XNOR U23954 ( .A(n22811), .B(n18331), .Z(n23728) );
  XNOR U23955 ( .A(n23729), .B(n22847), .Z(n18331) );
  NOR U23956 ( .A(n22848), .B(n21760), .Z(n23729) );
  XOR U23957 ( .A(n23730), .B(n23731), .Z(n21760) );
  XOR U23958 ( .A(n23732), .B(n23733), .Z(n22848) );
  XOR U23959 ( .A(n23734), .B(n23735), .Z(n22811) );
  NOR U23960 ( .A(n21770), .B(n22850), .Z(n23734) );
  XOR U23961 ( .A(n23736), .B(n23737), .Z(n22850) );
  XOR U23962 ( .A(n23738), .B(n23739), .Z(n21770) );
  XOR U23963 ( .A(n23740), .B(n22854), .Z(n14998) );
  IV U23964 ( .A(n23741), .Z(n22854) );
  NOR U23965 ( .A(n22853), .B(n21756), .Z(n23740) );
  XNOR U23966 ( .A(n23742), .B(n23743), .Z(n21756) );
  XNOR U23967 ( .A(n23744), .B(n23745), .Z(n22853) );
  XOR U23968 ( .A(n23746), .B(n16056), .Z(n15145) );
  IV U23969 ( .A(n17177), .Z(n16056) );
  XNOR U23970 ( .A(n23747), .B(n23748), .Z(n20252) );
  XOR U23971 ( .A(n19120), .B(n15643), .Z(n23748) );
  XNOR U23972 ( .A(n23749), .B(n20530), .Z(n15643) );
  XOR U23973 ( .A(n23750), .B(n23751), .Z(n20530) );
  ANDN U23974 ( .B(n21821), .A(n21362), .Z(n23749) );
  IV U23975 ( .A(n23752), .Z(n21362) );
  XNOR U23976 ( .A(n23753), .B(n20541), .Z(n19120) );
  XOR U23977 ( .A(n23754), .B(n23442), .Z(n20541) );
  ANDN U23978 ( .B(n21831), .A(n21360), .Z(n23753) );
  IV U23979 ( .A(n23755), .Z(n21360) );
  XOR U23980 ( .A(n16991), .B(n23756), .Z(n23747) );
  XOR U23981 ( .A(n19700), .B(n17018), .Z(n23756) );
  XOR U23982 ( .A(n23757), .B(n20537), .Z(n17018) );
  XOR U23983 ( .A(n23758), .B(n22017), .Z(n20537) );
  ANDN U23984 ( .B(n21827), .A(n23759), .Z(n23757) );
  XNOR U23985 ( .A(n23760), .B(n21345), .Z(n19700) );
  XOR U23986 ( .A(n23761), .B(n23708), .Z(n21345) );
  ANDN U23987 ( .B(n23762), .A(n21354), .Z(n23760) );
  XNOR U23988 ( .A(n23763), .B(n21358), .Z(n16991) );
  IV U23989 ( .A(n20527), .Z(n21358) );
  XOR U23990 ( .A(n23764), .B(n23765), .Z(n20527) );
  NOR U23991 ( .A(n23766), .B(n21357), .Z(n23763) );
  XOR U23992 ( .A(n23767), .B(n23768), .Z(n20013) );
  XNOR U23993 ( .A(n18376), .B(n17952), .Z(n23768) );
  XOR U23994 ( .A(n23769), .B(n23770), .Z(n17952) );
  ANDN U23995 ( .B(n23771), .A(n21452), .Z(n23769) );
  IV U23996 ( .A(n23772), .Z(n21452) );
  XNOR U23997 ( .A(n23773), .B(n20062), .Z(n18376) );
  IV U23998 ( .A(n23774), .Z(n20062) );
  ANDN U23999 ( .B(n21445), .A(n20061), .Z(n23773) );
  XOR U24000 ( .A(n20048), .B(n23775), .Z(n23767) );
  XNOR U24001 ( .A(n18895), .B(n15289), .Z(n23775) );
  XOR U24002 ( .A(n23776), .B(n22909), .Z(n15289) );
  NOR U24003 ( .A(n22908), .B(n21448), .Z(n23776) );
  XNOR U24004 ( .A(n23777), .B(n20065), .Z(n18895) );
  IV U24005 ( .A(n23778), .Z(n20065) );
  ANDN U24006 ( .B(n20066), .A(n21441), .Z(n23777) );
  XNOR U24007 ( .A(n23779), .B(n20055), .Z(n20048) );
  ANDN U24008 ( .B(n20056), .A(n23780), .Z(n23779) );
  XNOR U24009 ( .A(n14020), .B(n23781), .Z(n23630) );
  XNOR U24010 ( .A(n11300), .B(n16659), .Z(n23781) );
  XOR U24011 ( .A(n23782), .B(n16697), .Z(n16659) );
  XOR U24012 ( .A(n20619), .B(n16105), .Z(n16697) );
  IV U24013 ( .A(n16025), .Z(n16105) );
  XOR U24014 ( .A(n23783), .B(n21391), .Z(n16025) );
  XNOR U24015 ( .A(n23784), .B(n23785), .Z(n21391) );
  XNOR U24016 ( .A(n17749), .B(n18338), .Z(n23785) );
  XNOR U24017 ( .A(n23786), .B(n21803), .Z(n18338) );
  NOR U24018 ( .A(n23787), .B(n20611), .Z(n23786) );
  XOR U24019 ( .A(n23788), .B(n23789), .Z(n20611) );
  XNOR U24020 ( .A(n23790), .B(n21811), .Z(n17749) );
  ANDN U24021 ( .B(n20615), .A(n20616), .Z(n23790) );
  XOR U24022 ( .A(n23791), .B(n23792), .Z(n20615) );
  XNOR U24023 ( .A(n21774), .B(n23793), .Z(n23784) );
  XOR U24024 ( .A(n18971), .B(n19455), .Z(n23793) );
  XNOR U24025 ( .A(n23794), .B(n23795), .Z(n19455) );
  NOR U24026 ( .A(n20622), .B(n20621), .Z(n23794) );
  XNOR U24027 ( .A(n23796), .B(n21800), .Z(n18971) );
  NOR U24028 ( .A(n21799), .B(n23797), .Z(n23796) );
  XOR U24029 ( .A(n23798), .B(n23799), .Z(n21774) );
  ANDN U24030 ( .B(n20627), .A(n20625), .Z(n23798) );
  XOR U24031 ( .A(n23800), .B(n23139), .Z(n20625) );
  XNOR U24032 ( .A(n23801), .B(n21799), .Z(n20619) );
  XNOR U24033 ( .A(n23701), .B(n23802), .Z(n21799) );
  ANDN U24034 ( .B(n23797), .A(n23803), .Z(n23801) );
  ANDN U24035 ( .B(n19480), .A(n19478), .Z(n23782) );
  IV U24036 ( .A(n16698), .Z(n19478) );
  XOR U24037 ( .A(n23804), .B(n16086), .Z(n16698) );
  XNOR U24038 ( .A(n23805), .B(n20998), .Z(n16086) );
  XNOR U24039 ( .A(n23806), .B(n23807), .Z(n20998) );
  XNOR U24040 ( .A(n17904), .B(n18550), .Z(n23807) );
  XOR U24041 ( .A(n23808), .B(n19577), .Z(n18550) );
  XNOR U24042 ( .A(n23809), .B(n23810), .Z(n19577) );
  ANDN U24043 ( .B(n22094), .A(n22092), .Z(n23808) );
  IV U24044 ( .A(n19578), .Z(n22092) );
  XOR U24045 ( .A(n23811), .B(n23765), .Z(n19578) );
  IV U24046 ( .A(n23812), .Z(n23765) );
  XNOR U24047 ( .A(n23813), .B(n19585), .Z(n17904) );
  XOR U24048 ( .A(n23814), .B(n23815), .Z(n19585) );
  ANDN U24049 ( .B(n22087), .A(n22086), .Z(n23813) );
  IV U24050 ( .A(n19586), .Z(n22086) );
  XOR U24051 ( .A(n22217), .B(n23816), .Z(n19586) );
  XOR U24052 ( .A(n15197), .B(n23817), .Z(n23806) );
  XNOR U24053 ( .A(n17489), .B(n16610), .Z(n23817) );
  XNOR U24054 ( .A(n23818), .B(n20070), .Z(n16610) );
  XOR U24055 ( .A(n23819), .B(n23432), .Z(n20070) );
  ANDN U24056 ( .B(n22090), .A(n19581), .Z(n23818) );
  XOR U24057 ( .A(n23820), .B(n23821), .Z(n19581) );
  XOR U24058 ( .A(n23822), .B(n19569), .Z(n17489) );
  XOR U24059 ( .A(n23738), .B(n23823), .Z(n19569) );
  ANDN U24060 ( .B(n22096), .A(n19568), .Z(n23822) );
  XNOR U24061 ( .A(n23824), .B(n23825), .Z(n19568) );
  XNOR U24062 ( .A(n23826), .B(n19572), .Z(n15197) );
  XNOR U24063 ( .A(n23047), .B(n23827), .Z(n19572) );
  ANDN U24064 ( .B(n22084), .A(n19573), .Z(n23826) );
  XOR U24065 ( .A(n23828), .B(n23829), .Z(n19573) );
  XNOR U24066 ( .A(n17456), .B(n21293), .Z(n19480) );
  XNOR U24067 ( .A(n23830), .B(n23309), .Z(n21293) );
  XNOR U24068 ( .A(n23831), .B(n23832), .Z(n21852) );
  IV U24069 ( .A(n17268), .Z(n17456) );
  XNOR U24070 ( .A(n23004), .B(n18263), .Z(n17268) );
  XNOR U24071 ( .A(n23833), .B(n23834), .Z(n18263) );
  XOR U24072 ( .A(n16060), .B(n17923), .Z(n23834) );
  XOR U24073 ( .A(n23835), .B(n23308), .Z(n17923) );
  XNOR U24074 ( .A(n23836), .B(n23837), .Z(n23308) );
  ANDN U24075 ( .B(n23309), .A(n21850), .Z(n23835) );
  XOR U24076 ( .A(n23838), .B(n23839), .Z(n21850) );
  XOR U24077 ( .A(n23840), .B(n23841), .Z(n23309) );
  XOR U24078 ( .A(n23842), .B(n23444), .Z(n16060) );
  XOR U24079 ( .A(n23843), .B(n23844), .Z(n23444) );
  ANDN U24080 ( .B(n21295), .A(n21839), .Z(n23842) );
  IV U24081 ( .A(n21296), .Z(n21839) );
  XOR U24082 ( .A(n23845), .B(n21214), .Z(n21296) );
  XOR U24083 ( .A(n22654), .B(n23846), .Z(n21295) );
  XNOR U24084 ( .A(n22584), .B(n23847), .Z(n23833) );
  XOR U24085 ( .A(n16742), .B(n19739), .Z(n23847) );
  XNOR U24086 ( .A(n23848), .B(n23313), .Z(n19739) );
  XOR U24087 ( .A(n23849), .B(n23812), .Z(n23313) );
  ANDN U24088 ( .B(n21286), .A(n21285), .Z(n23848) );
  XOR U24089 ( .A(n23851), .B(n23852), .Z(n21286) );
  XNOR U24090 ( .A(n23853), .B(n23560), .Z(n16742) );
  XNOR U24091 ( .A(n23854), .B(n23855), .Z(n23560) );
  ANDN U24092 ( .B(n21299), .A(n21842), .Z(n23853) );
  IV U24093 ( .A(n21301), .Z(n21842) );
  XOR U24094 ( .A(n23856), .B(n23857), .Z(n21301) );
  XNOR U24095 ( .A(n23858), .B(n23136), .Z(n21299) );
  XNOR U24096 ( .A(n23859), .B(n23315), .Z(n22584) );
  XOR U24097 ( .A(n23860), .B(n21599), .Z(n23315) );
  NOR U24098 ( .A(n23316), .B(n21290), .Z(n23859) );
  XNOR U24099 ( .A(n23861), .B(n23862), .Z(n21290) );
  XOR U24100 ( .A(n23863), .B(n23864), .Z(n23316) );
  XOR U24101 ( .A(n23865), .B(n23866), .Z(n23004) );
  XNOR U24102 ( .A(n16607), .B(n17000), .Z(n23866) );
  XOR U24103 ( .A(n23867), .B(n22597), .Z(n17000) );
  NOR U24104 ( .A(n22598), .B(n23374), .Z(n23867) );
  XOR U24105 ( .A(n23868), .B(n23869), .Z(n22598) );
  XNOR U24106 ( .A(n23870), .B(n23871), .Z(n16607) );
  ANDN U24107 ( .B(n23368), .A(n23366), .Z(n23870) );
  XNOR U24108 ( .A(n17126), .B(n23872), .Z(n23865) );
  XNOR U24109 ( .A(n18970), .B(n19040), .Z(n23872) );
  XNOR U24110 ( .A(n23873), .B(n22602), .Z(n19040) );
  ANDN U24111 ( .B(n23371), .A(n22601), .Z(n23873) );
  XOR U24112 ( .A(n23856), .B(n23874), .Z(n22601) );
  XOR U24113 ( .A(n23875), .B(n22592), .Z(n18970) );
  ANDN U24114 ( .B(n23377), .A(n23876), .Z(n23875) );
  XNOR U24115 ( .A(n23877), .B(n23878), .Z(n23377) );
  XNOR U24116 ( .A(n23879), .B(n23880), .Z(n17126) );
  ANDN U24117 ( .B(n23381), .A(n23382), .Z(n23879) );
  XNOR U24118 ( .A(n23881), .B(n16694), .Z(n11300) );
  XNOR U24119 ( .A(n16770), .B(n23882), .Z(n16694) );
  ANDN U24120 ( .B(n16693), .A(n15149), .Z(n23881) );
  XNOR U24121 ( .A(n23883), .B(n16616), .Z(n15149) );
  XOR U24122 ( .A(n23884), .B(n23885), .Z(n23385) );
  XNOR U24123 ( .A(n18871), .B(n18978), .Z(n23885) );
  XOR U24124 ( .A(n23886), .B(n23887), .Z(n18978) );
  NOR U24125 ( .A(n23888), .B(n23889), .Z(n23886) );
  XOR U24126 ( .A(n23890), .B(n21262), .Z(n18871) );
  ANDN U24127 ( .B(n21263), .A(n23891), .Z(n23890) );
  XOR U24128 ( .A(n17234), .B(n23892), .Z(n23884) );
  XNOR U24129 ( .A(n21255), .B(n17636), .Z(n23892) );
  XOR U24130 ( .A(n23893), .B(n21527), .Z(n17636) );
  NOR U24131 ( .A(n23894), .B(n23895), .Z(n23893) );
  XNOR U24132 ( .A(n23896), .B(n23897), .Z(n21255) );
  NOR U24133 ( .A(n23898), .B(n23899), .Z(n23896) );
  XOR U24134 ( .A(n23900), .B(n21269), .Z(n17234) );
  AND U24135 ( .A(n21270), .B(n23901), .Z(n23900) );
  XOR U24136 ( .A(n23902), .B(n23903), .Z(n20141) );
  XNOR U24137 ( .A(n18217), .B(n17902), .Z(n23903) );
  XNOR U24138 ( .A(n23904), .B(n20356), .Z(n17902) );
  XNOR U24139 ( .A(n23905), .B(n23906), .Z(n20356) );
  ANDN U24140 ( .B(n20357), .A(n23907), .Z(n23904) );
  XNOR U24141 ( .A(n23908), .B(n21410), .Z(n18217) );
  IV U24142 ( .A(n20343), .Z(n21410) );
  XOR U24143 ( .A(n23909), .B(n23429), .Z(n20343) );
  NOR U24144 ( .A(n23910), .B(n20342), .Z(n23908) );
  XOR U24145 ( .A(n18904), .B(n23911), .Z(n23902) );
  XOR U24146 ( .A(n18055), .B(n19218), .Z(n23911) );
  XNOR U24147 ( .A(n23912), .B(n21406), .Z(n19218) );
  IV U24148 ( .A(n20347), .Z(n21406) );
  XOR U24149 ( .A(n23913), .B(n23914), .Z(n20347) );
  NOR U24150 ( .A(n23915), .B(n20346), .Z(n23912) );
  XOR U24151 ( .A(n23916), .B(n20352), .Z(n18055) );
  XOR U24152 ( .A(n23917), .B(n22012), .Z(n20352) );
  AND U24153 ( .A(n23918), .B(n20353), .Z(n23916) );
  XOR U24154 ( .A(n23919), .B(n20993), .Z(n18904) );
  XOR U24155 ( .A(n23047), .B(n23920), .Z(n20993) );
  ANDN U24156 ( .B(n20992), .A(n23921), .Z(n23919) );
  XOR U24157 ( .A(n21538), .B(n17514), .Z(n16693) );
  IV U24158 ( .A(n18422), .Z(n17514) );
  XNOR U24159 ( .A(n18551), .B(n20193), .Z(n18422) );
  XNOR U24160 ( .A(n23922), .B(n23923), .Z(n20193) );
  XNOR U24161 ( .A(n23924), .B(n15343), .Z(n23923) );
  XNOR U24162 ( .A(n23925), .B(n23926), .Z(n15343) );
  NOR U24163 ( .A(n21576), .B(n21577), .Z(n23925) );
  XOR U24164 ( .A(n18360), .B(n23927), .Z(n23922) );
  XOR U24165 ( .A(n17265), .B(n17791), .Z(n23927) );
  XOR U24166 ( .A(n23928), .B(n23929), .Z(n17791) );
  ANDN U24167 ( .B(n21563), .A(n21564), .Z(n23928) );
  XOR U24168 ( .A(n23930), .B(n23931), .Z(n17265) );
  NOR U24169 ( .A(n21568), .B(n21569), .Z(n23930) );
  XNOR U24170 ( .A(n23932), .B(n23933), .Z(n18360) );
  ANDN U24171 ( .B(n21574), .A(n21572), .Z(n23932) );
  IV U24172 ( .A(n23934), .Z(n21572) );
  XNOR U24173 ( .A(n23935), .B(n23936), .Z(n18551) );
  XNOR U24174 ( .A(n18214), .B(n19001), .Z(n23936) );
  XOR U24175 ( .A(n23937), .B(n21276), .Z(n19001) );
  ANDN U24176 ( .B(n21554), .A(n21553), .Z(n23937) );
  XOR U24177 ( .A(n23938), .B(n23812), .Z(n21553) );
  XNOR U24178 ( .A(n23939), .B(n20863), .Z(n18214) );
  IV U24179 ( .A(n20862), .Z(n21540) );
  XOR U24180 ( .A(n23940), .B(n23941), .Z(n20862) );
  XNOR U24181 ( .A(n20851), .B(n23942), .Z(n23935) );
  XNOR U24182 ( .A(n17941), .B(n16089), .Z(n23942) );
  XNOR U24183 ( .A(n23943), .B(n23944), .Z(n16089) );
  ANDN U24184 ( .B(n21545), .A(n21546), .Z(n23943) );
  XOR U24185 ( .A(n23945), .B(n22329), .Z(n17941) );
  NOR U24186 ( .A(n22330), .B(n21550), .Z(n23945) );
  XOR U24187 ( .A(n23946), .B(n23947), .Z(n22330) );
  XNOR U24188 ( .A(n23948), .B(n20937), .Z(n20851) );
  ANDN U24189 ( .B(n20936), .A(n23949), .Z(n23948) );
  XNOR U24190 ( .A(n23950), .B(n20936), .Z(n21538) );
  XOR U24191 ( .A(n23951), .B(n23952), .Z(n20936) );
  XOR U24192 ( .A(n23954), .B(n16687), .Z(n14020) );
  XOR U24193 ( .A(n22588), .B(n16830), .Z(n16687) );
  IV U24194 ( .A(n17031), .Z(n16830) );
  XOR U24195 ( .A(n23955), .B(n23956), .Z(n22588) );
  ANDN U24196 ( .B(n23366), .A(n23871), .Z(n23955) );
  XNOR U24197 ( .A(n23957), .B(n23958), .Z(n23366) );
  NOR U24198 ( .A(n15155), .B(n16686), .Z(n23954) );
  XOR U24199 ( .A(n23959), .B(n17574), .Z(n16686) );
  XNOR U24200 ( .A(n20044), .B(n19948), .Z(n17574) );
  XNOR U24201 ( .A(n23960), .B(n23961), .Z(n19948) );
  XNOR U24202 ( .A(n18661), .B(n18875), .Z(n23961) );
  XNOR U24203 ( .A(n23962), .B(n21743), .Z(n18875) );
  XOR U24204 ( .A(n23963), .B(n23964), .Z(n21743) );
  ANDN U24205 ( .B(n21654), .A(n21744), .Z(n23962) );
  XNOR U24206 ( .A(n23965), .B(n22663), .Z(n18661) );
  XNOR U24207 ( .A(n23966), .B(n23914), .Z(n22663) );
  NOR U24208 ( .A(n21662), .B(n22662), .Z(n23965) );
  XNOR U24209 ( .A(n21736), .B(n23967), .Z(n23960) );
  XNOR U24210 ( .A(n17473), .B(n17146), .Z(n23967) );
  XNOR U24211 ( .A(n23968), .B(n21752), .Z(n17146) );
  XOR U24212 ( .A(n23969), .B(n23970), .Z(n21752) );
  NOR U24213 ( .A(n23971), .B(n21751), .Z(n23968) );
  XNOR U24214 ( .A(n23972), .B(n21740), .Z(n17473) );
  XOR U24215 ( .A(n23973), .B(n23063), .Z(n21740) );
  IV U24216 ( .A(n23974), .Z(n23063) );
  ANDN U24217 ( .B(n21741), .A(n23975), .Z(n23972) );
  XOR U24218 ( .A(n23976), .B(n21749), .Z(n21736) );
  XOR U24219 ( .A(n23977), .B(n23978), .Z(n21749) );
  ANDN U24220 ( .B(n21645), .A(n21748), .Z(n23976) );
  XOR U24221 ( .A(n23979), .B(n23980), .Z(n20044) );
  XOR U24222 ( .A(n17315), .B(n16100), .Z(n23980) );
  XOR U24223 ( .A(n23981), .B(n21758), .Z(n16100) );
  XOR U24224 ( .A(n23982), .B(n23983), .Z(n21758) );
  NOR U24225 ( .A(n23741), .B(n21757), .Z(n23981) );
  XNOR U24226 ( .A(n23984), .B(n23985), .Z(n21757) );
  XOR U24227 ( .A(n23986), .B(n23987), .Z(n23741) );
  XNOR U24228 ( .A(n23988), .B(n21768), .Z(n17315) );
  XOR U24229 ( .A(n23699), .B(n23989), .Z(n21768) );
  ANDN U24230 ( .B(n22840), .A(n21767), .Z(n23988) );
  XNOR U24231 ( .A(n23831), .B(n23990), .Z(n21767) );
  XOR U24232 ( .A(n23991), .B(n23992), .Z(n22840) );
  XOR U24233 ( .A(n18779), .B(n23993), .Z(n23979) );
  XNOR U24234 ( .A(n19013), .B(n17010), .Z(n23993) );
  XOR U24235 ( .A(n23994), .B(n21762), .Z(n17010) );
  XOR U24236 ( .A(n23995), .B(n23996), .Z(n21762) );
  ANDN U24237 ( .B(n22847), .A(n21761), .Z(n23994) );
  XNOR U24238 ( .A(n23997), .B(n23969), .Z(n21761) );
  XNOR U24239 ( .A(n23998), .B(n23999), .Z(n22847) );
  XOR U24240 ( .A(n24000), .B(n23129), .Z(n19013) );
  XOR U24241 ( .A(n22624), .B(n24001), .Z(n23129) );
  AND U24242 ( .A(n22842), .B(n22843), .Z(n24000) );
  XNOR U24243 ( .A(n21603), .B(n24002), .Z(n22843) );
  XOR U24244 ( .A(n23843), .B(n24003), .Z(n22842) );
  XOR U24245 ( .A(n24004), .B(n21771), .Z(n18779) );
  XOR U24246 ( .A(n24005), .B(n24006), .Z(n21771) );
  ANDN U24247 ( .B(n22851), .A(n21773), .Z(n24004) );
  XOR U24248 ( .A(n24007), .B(n24008), .Z(n21773) );
  IV U24249 ( .A(n23735), .Z(n22851) );
  XOR U24250 ( .A(n24009), .B(n24010), .Z(n23735) );
  XOR U24251 ( .A(n20316), .B(n18834), .Z(n15155) );
  IV U24252 ( .A(n20039), .Z(n18834) );
  XNOR U24253 ( .A(n24011), .B(n24012), .Z(n20316) );
  NOR U24254 ( .A(n24013), .B(n19354), .Z(n24011) );
  XOR U24255 ( .A(n24014), .B(n24015), .Z(n16554) );
  XOR U24256 ( .A(n9546), .B(n12392), .Z(n24015) );
  XOR U24257 ( .A(n24016), .B(n13339), .Z(n12392) );
  XOR U24258 ( .A(n20057), .B(n18150), .Z(n13339) );
  XOR U24259 ( .A(n20521), .B(n24017), .Z(n18150) );
  XOR U24260 ( .A(n24018), .B(n24019), .Z(n20521) );
  XOR U24261 ( .A(n19506), .B(n16077), .Z(n24019) );
  XNOR U24262 ( .A(n24020), .B(n21446), .Z(n16077) );
  NOR U24263 ( .A(n23774), .B(n20060), .Z(n24020) );
  XNOR U24264 ( .A(n24021), .B(n23964), .Z(n20060) );
  XOR U24265 ( .A(n24022), .B(n22613), .Z(n23774) );
  XNOR U24266 ( .A(n24023), .B(n24024), .Z(n19506) );
  XNOR U24267 ( .A(n24025), .B(n24026), .Z(n20055) );
  XNOR U24268 ( .A(n18333), .B(n24027), .Z(n24018) );
  XNOR U24269 ( .A(n21419), .B(n18298), .Z(n24027) );
  XNOR U24270 ( .A(n24028), .B(n21442), .Z(n18298) );
  NOR U24271 ( .A(n23778), .B(n20064), .Z(n24028) );
  XOR U24272 ( .A(n24029), .B(n22406), .Z(n20064) );
  XOR U24273 ( .A(n24030), .B(n24031), .Z(n23778) );
  XNOR U24274 ( .A(n24032), .B(n21449), .Z(n21419) );
  ANDN U24275 ( .B(n21450), .A(n22909), .Z(n24032) );
  XOR U24276 ( .A(n24033), .B(n23985), .Z(n22909) );
  XNOR U24277 ( .A(n24036), .B(n21453), .Z(n18333) );
  NOR U24278 ( .A(n23770), .B(n21454), .Z(n24036) );
  XNOR U24279 ( .A(n24037), .B(n21454), .Z(n20057) );
  XOR U24280 ( .A(n24038), .B(n24039), .Z(n21454) );
  ANDN U24281 ( .B(n23770), .A(n23771), .Z(n24037) );
  XOR U24282 ( .A(n24040), .B(n24041), .Z(n23770) );
  NOR U24283 ( .A(n16665), .B(n15042), .Z(n24016) );
  XNOR U24284 ( .A(n24042), .B(n17140), .Z(n15042) );
  XNOR U24285 ( .A(n24043), .B(n24044), .Z(n20703) );
  XNOR U24286 ( .A(n18573), .B(n18280), .Z(n24044) );
  XNOR U24287 ( .A(n24045), .B(n22073), .Z(n18280) );
  NOR U24288 ( .A(n24046), .B(n24047), .Z(n24045) );
  XOR U24289 ( .A(n24048), .B(n22077), .Z(n18573) );
  NOR U24290 ( .A(n24049), .B(n24050), .Z(n24048) );
  XOR U24291 ( .A(n20599), .B(n24051), .Z(n24043) );
  XNOR U24292 ( .A(n17012), .B(n24052), .Z(n24051) );
  XNOR U24293 ( .A(n24053), .B(n23475), .Z(n17012) );
  ANDN U24294 ( .B(n24054), .A(n24055), .Z(n24053) );
  XNOR U24295 ( .A(n24056), .B(n22063), .Z(n20599) );
  IV U24296 ( .A(n24057), .Z(n22063) );
  NOR U24297 ( .A(n24058), .B(n24059), .Z(n24056) );
  XNOR U24298 ( .A(n24060), .B(n24061), .Z(n20153) );
  XOR U24299 ( .A(n19084), .B(n17950), .Z(n24061) );
  XNOR U24300 ( .A(n24062), .B(n22053), .Z(n17950) );
  ANDN U24301 ( .B(n22159), .A(n22158), .Z(n24062) );
  XNOR U24302 ( .A(n24063), .B(n24064), .Z(n22159) );
  XOR U24303 ( .A(n24065), .B(n22057), .Z(n19084) );
  NOR U24304 ( .A(n22151), .B(n22152), .Z(n24065) );
  XNOR U24305 ( .A(n22318), .B(n24066), .Z(n22152) );
  XNOR U24306 ( .A(n18040), .B(n24067), .Z(n24060) );
  XNOR U24307 ( .A(n18470), .B(n17915), .Z(n24067) );
  XOR U24308 ( .A(n24068), .B(n22044), .Z(n17915) );
  NOR U24309 ( .A(n22163), .B(n22162), .Z(n24068) );
  XOR U24310 ( .A(n24069), .B(n24070), .Z(n22163) );
  XNOR U24311 ( .A(n24071), .B(n22048), .Z(n18470) );
  NOR U24312 ( .A(n22149), .B(n22148), .Z(n24071) );
  XOR U24313 ( .A(n24072), .B(n24073), .Z(n22149) );
  XNOR U24314 ( .A(n24074), .B(n22039), .Z(n18040) );
  ANDN U24315 ( .B(n22155), .A(n22156), .Z(n24074) );
  XOR U24316 ( .A(n24075), .B(n24076), .Z(n22156) );
  XOR U24317 ( .A(n24077), .B(n16045), .Z(n16665) );
  XOR U24318 ( .A(n22362), .B(n24078), .Z(n16045) );
  XNOR U24319 ( .A(n24079), .B(n24080), .Z(n22362) );
  XNOR U24320 ( .A(n18612), .B(n19464), .Z(n24080) );
  XOR U24321 ( .A(n24081), .B(n23268), .Z(n19464) );
  XNOR U24322 ( .A(n24083), .B(n23273), .Z(n18612) );
  NOR U24323 ( .A(n23274), .B(n24084), .Z(n24083) );
  XOR U24324 ( .A(n19127), .B(n24085), .Z(n24079) );
  XOR U24325 ( .A(n18905), .B(n18516), .Z(n24085) );
  XNOR U24326 ( .A(n24086), .B(n24087), .Z(n18516) );
  NOR U24327 ( .A(n24088), .B(n23278), .Z(n24086) );
  XNOR U24328 ( .A(n24089), .B(n23282), .Z(n18905) );
  NOR U24329 ( .A(n23283), .B(n24090), .Z(n24089) );
  XNOR U24330 ( .A(n24091), .B(n24092), .Z(n19127) );
  NOR U24331 ( .A(n24093), .B(n23286), .Z(n24091) );
  XNOR U24332 ( .A(n24094), .B(n16670), .Z(n9546) );
  IV U24333 ( .A(n13345), .Z(n16670) );
  XOR U24334 ( .A(n21264), .B(n18234), .Z(n13345) );
  XOR U24335 ( .A(n24095), .B(n24096), .Z(n21264) );
  ANDN U24336 ( .B(n23898), .A(n24097), .Z(n24095) );
  NOR U24337 ( .A(n16669), .B(n15040), .Z(n24094) );
  XOR U24338 ( .A(n24098), .B(n16744), .Z(n15040) );
  XNOR U24339 ( .A(n20012), .B(n20570), .Z(n16744) );
  XNOR U24340 ( .A(n24099), .B(n24100), .Z(n20570) );
  XNOR U24341 ( .A(n17993), .B(n18067), .Z(n24100) );
  XOR U24342 ( .A(n24101), .B(n24102), .Z(n18067) );
  ANDN U24343 ( .B(n22304), .A(n24103), .Z(n24101) );
  XNOR U24344 ( .A(n24104), .B(n24105), .Z(n17993) );
  ANDN U24345 ( .B(n24106), .A(n22300), .Z(n24104) );
  XNOR U24346 ( .A(n18629), .B(n24107), .Z(n24099) );
  XOR U24347 ( .A(n15872), .B(n19134), .Z(n24107) );
  XNOR U24348 ( .A(n24108), .B(n24109), .Z(n19134) );
  NOR U24349 ( .A(n22287), .B(n24110), .Z(n24108) );
  XNOR U24350 ( .A(n24111), .B(n24112), .Z(n15872) );
  XNOR U24351 ( .A(n24114), .B(n24115), .Z(n18629) );
  AND U24352 ( .A(n24116), .B(n22296), .Z(n24114) );
  XOR U24353 ( .A(n24117), .B(n24118), .Z(n20012) );
  XNOR U24354 ( .A(n24119), .B(n19445), .Z(n24118) );
  XNOR U24355 ( .A(n24120), .B(n24121), .Z(n19445) );
  NOR U24356 ( .A(n22276), .B(n24122), .Z(n24120) );
  XNOR U24357 ( .A(n17860), .B(n24123), .Z(n24117) );
  XOR U24358 ( .A(n18549), .B(n20388), .Z(n24123) );
  XNOR U24359 ( .A(n24124), .B(n24125), .Z(n20388) );
  ANDN U24360 ( .B(n24126), .A(n21434), .Z(n24124) );
  IV U24361 ( .A(n24127), .Z(n21434) );
  XOR U24362 ( .A(n24128), .B(n24129), .Z(n18549) );
  NOR U24363 ( .A(n24130), .B(n21423), .Z(n24128) );
  XOR U24364 ( .A(n24131), .B(n24132), .Z(n17860) );
  ANDN U24365 ( .B(n24133), .A(n24134), .Z(n24131) );
  XOR U24366 ( .A(n18578), .B(n24135), .Z(n16669) );
  IV U24367 ( .A(n17246), .Z(n18578) );
  XOR U24368 ( .A(n22003), .B(n20704), .Z(n17246) );
  XOR U24369 ( .A(n24136), .B(n24137), .Z(n20704) );
  XNOR U24370 ( .A(n23180), .B(n18520), .Z(n24137) );
  XNOR U24371 ( .A(n24138), .B(n23894), .Z(n18520) );
  IV U24372 ( .A(n21528), .Z(n23894) );
  XOR U24373 ( .A(n22217), .B(n24139), .Z(n21528) );
  ANDN U24374 ( .B(n23895), .A(n24140), .Z(n24138) );
  XNOR U24375 ( .A(n24141), .B(n23889), .Z(n23180) );
  AND U24376 ( .A(n23888), .B(n24142), .Z(n24141) );
  XNOR U24377 ( .A(n23384), .B(n24143), .Z(n24136) );
  XOR U24378 ( .A(n18723), .B(n17545), .Z(n24143) );
  XNOR U24379 ( .A(n24144), .B(n21270), .Z(n17545) );
  XOR U24380 ( .A(n24145), .B(n24146), .Z(n21270) );
  NOR U24381 ( .A(n24147), .B(n23901), .Z(n24144) );
  XNOR U24382 ( .A(n24148), .B(n21263), .Z(n18723) );
  XNOR U24383 ( .A(n24149), .B(n24150), .Z(n21263) );
  ANDN U24384 ( .B(n23891), .A(n24151), .Z(n24148) );
  XNOR U24385 ( .A(n24152), .B(n23898), .Z(n23384) );
  XOR U24386 ( .A(n24153), .B(n24154), .Z(n23898) );
  XOR U24387 ( .A(n24156), .B(n24157), .Z(n22003) );
  XNOR U24388 ( .A(n17459), .B(n16615), .Z(n24157) );
  XOR U24389 ( .A(n24158), .B(n20346), .Z(n16615) );
  XOR U24390 ( .A(n24159), .B(n22021), .Z(n20346) );
  ANDN U24391 ( .B(n23915), .A(n21405), .Z(n24158) );
  XOR U24392 ( .A(n24160), .B(n20353), .Z(n17459) );
  XNOR U24393 ( .A(n24161), .B(n24162), .Z(n20353) );
  NOR U24394 ( .A(n21412), .B(n23918), .Z(n24160) );
  XNOR U24395 ( .A(n23883), .B(n24163), .Z(n24156) );
  XNOR U24396 ( .A(n19698), .B(n18251), .Z(n24163) );
  XNOR U24397 ( .A(n24164), .B(n20342), .Z(n18251) );
  XNOR U24398 ( .A(n24165), .B(n24166), .Z(n20342) );
  ANDN U24399 ( .B(n23910), .A(n24167), .Z(n24164) );
  XNOR U24400 ( .A(n24168), .B(n20992), .Z(n19698) );
  XOR U24401 ( .A(n22409), .B(n24169), .Z(n20992) );
  XOR U24402 ( .A(n24170), .B(n20357), .Z(n23883) );
  XOR U24403 ( .A(n24171), .B(n24172), .Z(n20357) );
  ANDN U24404 ( .B(n21414), .A(n24173), .Z(n24170) );
  XOR U24405 ( .A(n13441), .B(n24174), .Z(n24014) );
  XOR U24406 ( .A(n9567), .B(n12218), .Z(n24174) );
  XOR U24407 ( .A(n24175), .B(n14875), .Z(n12218) );
  XOR U24408 ( .A(n21077), .B(n19389), .Z(n14875) );
  XOR U24409 ( .A(n19792), .B(n18180), .Z(n19389) );
  XNOR U24410 ( .A(n24176), .B(n24177), .Z(n18180) );
  XOR U24411 ( .A(n20132), .B(n15898), .Z(n24177) );
  XNOR U24412 ( .A(n24178), .B(n21128), .Z(n15898) );
  XOR U24413 ( .A(n24179), .B(n24180), .Z(n21128) );
  ANDN U24414 ( .B(n21082), .A(n21080), .Z(n24178) );
  XOR U24415 ( .A(n24181), .B(n24182), .Z(n21080) );
  XNOR U24416 ( .A(n24183), .B(n21123), .Z(n20132) );
  IV U24417 ( .A(n22755), .Z(n21123) );
  XOR U24418 ( .A(n24184), .B(n24185), .Z(n22755) );
  NOR U24419 ( .A(n21070), .B(n21072), .Z(n24183) );
  XOR U24420 ( .A(n24186), .B(n23708), .Z(n21070) );
  XNOR U24421 ( .A(n19023), .B(n24187), .Z(n24176) );
  XNOR U24422 ( .A(n18346), .B(n16397), .Z(n24187) );
  ANDN U24423 ( .B(n21076), .A(n21074), .Z(n24188) );
  XOR U24424 ( .A(n24009), .B(n24189), .Z(n21074) );
  IV U24425 ( .A(n24190), .Z(n21076) );
  XNOR U24426 ( .A(n24191), .B(n21120), .Z(n18346) );
  XNOR U24427 ( .A(n24192), .B(n24193), .Z(n21120) );
  NOR U24428 ( .A(n21084), .B(n21086), .Z(n24191) );
  XOR U24429 ( .A(n24194), .B(n24172), .Z(n21084) );
  XNOR U24430 ( .A(n24195), .B(n21132), .Z(n19023) );
  XNOR U24431 ( .A(n24196), .B(n24197), .Z(n21132) );
  NOR U24432 ( .A(n21131), .B(n24198), .Z(n24195) );
  XOR U24433 ( .A(n24199), .B(n24200), .Z(n19792) );
  XNOR U24434 ( .A(n17517), .B(n21038), .Z(n24200) );
  XOR U24435 ( .A(n24201), .B(n22764), .Z(n21038) );
  XNOR U24436 ( .A(n24202), .B(n22770), .Z(n17517) );
  NOR U24437 ( .A(n21051), .B(n21052), .Z(n24202) );
  XOR U24438 ( .A(n20838), .B(n24203), .Z(n24199) );
  XOR U24439 ( .A(n16530), .B(n24204), .Z(n24203) );
  XNOR U24440 ( .A(n24205), .B(n22773), .Z(n16530) );
  NOR U24441 ( .A(n21057), .B(n21056), .Z(n24205) );
  XNOR U24442 ( .A(n24206), .B(n22762), .Z(n20838) );
  NOR U24443 ( .A(n24207), .B(n21060), .Z(n24206) );
  XNOR U24444 ( .A(n24208), .B(n21131), .Z(n21077) );
  XOR U24445 ( .A(n24209), .B(n24210), .Z(n21131) );
  AND U24446 ( .A(n22757), .B(n24198), .Z(n24208) );
  ANDN U24447 ( .B(n16675), .A(n15034), .Z(n24175) );
  XNOR U24448 ( .A(n24211), .B(n18275), .Z(n15034) );
  IV U24449 ( .A(n20849), .Z(n18275) );
  XNOR U24450 ( .A(n22578), .B(n24212), .Z(n20849) );
  XOR U24451 ( .A(n24213), .B(n24214), .Z(n22578) );
  XNOR U24452 ( .A(n20671), .B(n16867), .Z(n24214) );
  XOR U24453 ( .A(n24215), .B(n22481), .Z(n16867) );
  XNOR U24454 ( .A(n24216), .B(n22484), .Z(n20671) );
  ANDN U24455 ( .B(n22249), .A(n22483), .Z(n24216) );
  XOR U24456 ( .A(n17129), .B(n24217), .Z(n24213) );
  XOR U24457 ( .A(n19383), .B(n20298), .Z(n24217) );
  XOR U24458 ( .A(n24218), .B(n22472), .Z(n20298) );
  NOR U24459 ( .A(n24219), .B(n22245), .Z(n24218) );
  XNOR U24460 ( .A(n24220), .B(n22478), .Z(n19383) );
  ANDN U24461 ( .B(n24221), .A(n24222), .Z(n24220) );
  XNOR U24462 ( .A(n24223), .B(n22470), .Z(n17129) );
  ANDN U24463 ( .B(n22235), .A(n22469), .Z(n24223) );
  XOR U24464 ( .A(n22973), .B(n17640), .Z(n16675) );
  IV U24465 ( .A(n15879), .Z(n17640) );
  XNOR U24466 ( .A(n24224), .B(n24225), .Z(n18977) );
  XNOR U24467 ( .A(n18825), .B(n20305), .Z(n24225) );
  XNOR U24468 ( .A(n24226), .B(n19936), .Z(n20305) );
  XOR U24469 ( .A(n24227), .B(n24228), .Z(n19936) );
  ANDN U24470 ( .B(n19978), .A(n22351), .Z(n24226) );
  XOR U24471 ( .A(n24229), .B(n23015), .Z(n22351) );
  XNOR U24472 ( .A(n24230), .B(n24231), .Z(n19978) );
  XNOR U24473 ( .A(n24232), .B(n22356), .Z(n18825) );
  XOR U24474 ( .A(n24233), .B(n24234), .Z(n22356) );
  NOR U24475 ( .A(n22355), .B(n20835), .Z(n24232) );
  XNOR U24476 ( .A(n23503), .B(n24235), .Z(n20835) );
  XOR U24477 ( .A(n24236), .B(n24237), .Z(n22355) );
  XOR U24478 ( .A(n20772), .B(n24238), .Z(n24224) );
  XNOR U24479 ( .A(n19544), .B(n18501), .Z(n24238) );
  XNOR U24480 ( .A(n24239), .B(n19927), .Z(n18501) );
  XNOR U24481 ( .A(n24240), .B(n22621), .Z(n19927) );
  AND U24482 ( .A(n22343), .B(n19976), .Z(n24239) );
  XOR U24483 ( .A(n24241), .B(n24242), .Z(n19976) );
  XOR U24484 ( .A(n24243), .B(n23253), .Z(n22343) );
  XNOR U24485 ( .A(n24244), .B(n19933), .Z(n19544) );
  XNOR U24486 ( .A(n24025), .B(n24245), .Z(n19933) );
  ANDN U24487 ( .B(n22348), .A(n19972), .Z(n24244) );
  XOR U24488 ( .A(n24246), .B(n24247), .Z(n19972) );
  XNOR U24489 ( .A(n23695), .B(n24248), .Z(n22348) );
  XNOR U24490 ( .A(n24249), .B(n19923), .Z(n20772) );
  XOR U24491 ( .A(n24250), .B(n24251), .Z(n19923) );
  ANDN U24492 ( .B(n19980), .A(n22993), .Z(n24249) );
  IV U24493 ( .A(n22339), .Z(n22993) );
  XOR U24494 ( .A(n23856), .B(n24252), .Z(n22339) );
  XOR U24495 ( .A(n24253), .B(n21225), .Z(n19980) );
  XOR U24496 ( .A(n24254), .B(n24255), .Z(n23520) );
  XNOR U24497 ( .A(n16072), .B(n19873), .Z(n24255) );
  XNOR U24498 ( .A(n24256), .B(n23119), .Z(n19873) );
  NOR U24499 ( .A(n22969), .B(n22970), .Z(n24256) );
  XNOR U24500 ( .A(n24257), .B(n24258), .Z(n22970) );
  XOR U24501 ( .A(n23335), .B(n24259), .Z(n22969) );
  XNOR U24502 ( .A(n24260), .B(n23114), .Z(n16072) );
  NOR U24503 ( .A(n23115), .B(n22189), .Z(n24260) );
  XOR U24504 ( .A(n24261), .B(n24262), .Z(n22189) );
  XOR U24505 ( .A(n24263), .B(n24146), .Z(n23115) );
  XNOR U24506 ( .A(n17448), .B(n24264), .Z(n24254) );
  XNOR U24507 ( .A(n21279), .B(n22332), .Z(n24264) );
  XNOR U24508 ( .A(n24265), .B(n23109), .Z(n22332) );
  NOR U24509 ( .A(n24266), .B(n23110), .Z(n24265) );
  XOR U24510 ( .A(n24267), .B(n23117), .Z(n21279) );
  IV U24511 ( .A(n24268), .Z(n23117) );
  ANDN U24512 ( .B(n22967), .A(n22203), .Z(n24267) );
  XOR U24513 ( .A(n24269), .B(n24270), .Z(n22203) );
  XOR U24514 ( .A(n24271), .B(n24272), .Z(n22967) );
  XOR U24515 ( .A(n24273), .B(n23106), .Z(n17448) );
  ANDN U24516 ( .B(n22977), .A(n22199), .Z(n24273) );
  XOR U24517 ( .A(n24274), .B(n24275), .Z(n22199) );
  XNOR U24518 ( .A(n24276), .B(n23482), .Z(n22977) );
  XNOR U24519 ( .A(n24277), .B(n23110), .Z(n22973) );
  XOR U24520 ( .A(n24278), .B(n24279), .Z(n23110) );
  NOR U24521 ( .A(n22193), .B(n22194), .Z(n24277) );
  IV U24522 ( .A(n24266), .Z(n22193) );
  XOR U24523 ( .A(n24280), .B(n24281), .Z(n24266) );
  XOR U24524 ( .A(n24282), .B(n13350), .Z(n9567) );
  IV U24525 ( .A(n16678), .Z(n13350) );
  XOR U24526 ( .A(n22593), .B(n17031), .Z(n16678) );
  XOR U24527 ( .A(n20382), .B(n23561), .Z(n17031) );
  XNOR U24528 ( .A(n24283), .B(n24284), .Z(n23561) );
  XNOR U24529 ( .A(n16728), .B(n18770), .Z(n24284) );
  XOR U24530 ( .A(n24285), .B(n23383), .Z(n18770) );
  ANDN U24531 ( .B(n23880), .A(n24286), .Z(n24285) );
  XNOR U24532 ( .A(n24287), .B(n23375), .Z(n16728) );
  ANDN U24533 ( .B(n22596), .A(n22597), .Z(n24287) );
  XOR U24534 ( .A(n24288), .B(n24289), .Z(n22597) );
  XOR U24535 ( .A(n19603), .B(n24290), .Z(n24283) );
  XNOR U24536 ( .A(n19755), .B(n24291), .Z(n24290) );
  XNOR U24537 ( .A(n24292), .B(n23378), .Z(n19755) );
  ANDN U24538 ( .B(n22590), .A(n22592), .Z(n24292) );
  XOR U24539 ( .A(n24293), .B(n23978), .Z(n22592) );
  XNOR U24540 ( .A(n24294), .B(n23370), .Z(n19603) );
  AND U24541 ( .A(n22600), .B(n22602), .Z(n24294) );
  XOR U24542 ( .A(n24295), .B(n24296), .Z(n22602) );
  XOR U24543 ( .A(n24297), .B(n24298), .Z(n20382) );
  XOR U24544 ( .A(n24299), .B(n18336), .Z(n24298) );
  XOR U24545 ( .A(n24300), .B(n24301), .Z(n18336) );
  ANDN U24546 ( .B(n22567), .A(n22566), .Z(n24300) );
  XOR U24547 ( .A(n20903), .B(n24302), .Z(n24297) );
  XNOR U24548 ( .A(n17960), .B(n20033), .Z(n24302) );
  XNOR U24549 ( .A(n24303), .B(n23361), .Z(n20033) );
  ANDN U24550 ( .B(n24304), .A(n24305), .Z(n24303) );
  XNOR U24551 ( .A(n24306), .B(n24307), .Z(n17960) );
  ANDN U24552 ( .B(n22570), .A(n24308), .Z(n24306) );
  XNOR U24553 ( .A(n24309), .B(n24310), .Z(n20903) );
  AND U24554 ( .A(n22575), .B(n22574), .Z(n24309) );
  XOR U24555 ( .A(n24311), .B(n24286), .Z(n22593) );
  NOR U24556 ( .A(n23381), .B(n23880), .Z(n24311) );
  XOR U24557 ( .A(n23738), .B(n24313), .Z(n23381) );
  IV U24558 ( .A(n22886), .Z(n23738) );
  XOR U24559 ( .A(n24314), .B(n24315), .Z(n22886) );
  NOR U24560 ( .A(n16677), .B(n17725), .Z(n24282) );
  XOR U24561 ( .A(n19783), .B(n20696), .Z(n17725) );
  XOR U24562 ( .A(n24316), .B(n20281), .Z(n19783) );
  ANDN U24563 ( .B(n19537), .A(n24317), .Z(n24316) );
  XNOR U24564 ( .A(n24318), .B(n23436), .Z(n19537) );
  XOR U24565 ( .A(n21865), .B(n18456), .Z(n16677) );
  IV U24566 ( .A(n19263), .Z(n18456) );
  XNOR U24567 ( .A(n19522), .B(n19764), .Z(n19263) );
  XNOR U24568 ( .A(n24319), .B(n24320), .Z(n19764) );
  XNOR U24569 ( .A(n18066), .B(n18956), .Z(n24320) );
  XNOR U24570 ( .A(n24321), .B(n24322), .Z(n18956) );
  NOR U24571 ( .A(n21861), .B(n21862), .Z(n24321) );
  XNOR U24572 ( .A(n24323), .B(n24324), .Z(n18066) );
  ANDN U24573 ( .B(n24325), .A(n24326), .Z(n24323) );
  XOR U24574 ( .A(n19827), .B(n24327), .Z(n24319) );
  XOR U24575 ( .A(n17917), .B(n18727), .Z(n24327) );
  XNOR U24576 ( .A(n24328), .B(n24329), .Z(n18727) );
  NOR U24577 ( .A(n21868), .B(n21867), .Z(n24328) );
  XNOR U24578 ( .A(n24330), .B(n24331), .Z(n17917) );
  ANDN U24579 ( .B(n21872), .A(n21871), .Z(n24330) );
  XOR U24580 ( .A(n24332), .B(n24333), .Z(n19827) );
  ANDN U24581 ( .B(n22874), .A(n22875), .Z(n24332) );
  XOR U24582 ( .A(n24334), .B(n24335), .Z(n19522) );
  XNOR U24583 ( .A(n19768), .B(n20812), .Z(n24335) );
  XNOR U24584 ( .A(n24336), .B(n21498), .Z(n20812) );
  AND U24585 ( .A(n21499), .B(n21892), .Z(n24336) );
  XOR U24586 ( .A(n24337), .B(n24338), .Z(n21499) );
  XOR U24587 ( .A(n24339), .B(n24340), .Z(n19768) );
  NOR U24588 ( .A(n21481), .B(n21888), .Z(n24339) );
  XNOR U24589 ( .A(n24341), .B(n24275), .Z(n21481) );
  XNOR U24590 ( .A(n15192), .B(n24342), .Z(n24334) );
  XNOR U24591 ( .A(n20094), .B(n21475), .Z(n24342) );
  XNOR U24592 ( .A(n24343), .B(n21494), .Z(n21475) );
  AND U24593 ( .A(n21495), .B(n21886), .Z(n24343) );
  XOR U24594 ( .A(n24344), .B(n24345), .Z(n21495) );
  XOR U24595 ( .A(n24346), .B(n24347), .Z(n20094) );
  AND U24596 ( .A(n21486), .B(n21878), .Z(n24346) );
  XOR U24597 ( .A(n24348), .B(n24349), .Z(n21486) );
  XNOR U24598 ( .A(n24350), .B(n21491), .Z(n15192) );
  ANDN U24599 ( .B(n21882), .A(n21880), .Z(n24350) );
  NOR U24600 ( .A(n24325), .B(n24353), .Z(n24352) );
  XNOR U24601 ( .A(n24354), .B(n14486), .Z(n13441) );
  IV U24602 ( .A(n16682), .Z(n14486) );
  XOR U24603 ( .A(n20559), .B(n18289), .Z(n16682) );
  IV U24604 ( .A(n16103), .Z(n18289) );
  XNOR U24605 ( .A(n21457), .B(n20666), .Z(n16103) );
  XOR U24606 ( .A(n24355), .B(n24356), .Z(n20666) );
  XOR U24607 ( .A(n18413), .B(n20707), .Z(n24356) );
  NOR U24608 ( .A(n20563), .B(n20562), .Z(n24357) );
  XOR U24609 ( .A(n24358), .B(n24162), .Z(n20562) );
  XNOR U24610 ( .A(n24359), .B(n20746), .Z(n18413) );
  ANDN U24611 ( .B(n20556), .A(n20557), .Z(n24359) );
  XOR U24612 ( .A(n24360), .B(n24349), .Z(n20556) );
  XOR U24613 ( .A(n20603), .B(n24361), .Z(n24355) );
  XNOR U24614 ( .A(n19230), .B(n19244), .Z(n24361) );
  XNOR U24615 ( .A(n24362), .B(n20736), .Z(n19244) );
  AND U24616 ( .A(n20737), .B(n24363), .Z(n24362) );
  XOR U24617 ( .A(n24364), .B(n20743), .Z(n19230) );
  ANDN U24618 ( .B(n20567), .A(n20566), .Z(n24364) );
  IV U24619 ( .A(n20742), .Z(n20566) );
  XOR U24620 ( .A(n24365), .B(n24366), .Z(n20742) );
  XOR U24621 ( .A(n24367), .B(n23258), .Z(n20603) );
  NOR U24622 ( .A(n20553), .B(n20552), .Z(n24367) );
  XNOR U24623 ( .A(n22495), .B(n24368), .Z(n20552) );
  XOR U24624 ( .A(n24369), .B(n24370), .Z(n21457) );
  XOR U24625 ( .A(n18943), .B(n18211), .Z(n24370) );
  XOR U24626 ( .A(n24371), .B(n20729), .Z(n18211) );
  XOR U24627 ( .A(n24372), .B(n24193), .Z(n20729) );
  NOR U24628 ( .A(n20730), .B(n22115), .Z(n24371) );
  XNOR U24629 ( .A(n24373), .B(n24374), .Z(n22115) );
  XOR U24630 ( .A(n24375), .B(n24376), .Z(n20730) );
  XNOR U24631 ( .A(n24377), .B(n20717), .Z(n18943) );
  XOR U24632 ( .A(n24378), .B(n24379), .Z(n20717) );
  ANDN U24633 ( .B(n22127), .A(n20716), .Z(n24377) );
  XNOR U24634 ( .A(n24380), .B(n24381), .Z(n20716) );
  XNOR U24635 ( .A(n23745), .B(n24382), .Z(n22127) );
  XOR U24636 ( .A(n19039), .B(n24383), .Z(n24369) );
  XOR U24637 ( .A(n18794), .B(n19053), .Z(n24383) );
  XOR U24638 ( .A(n24384), .B(n20713), .Z(n19053) );
  XOR U24639 ( .A(n24385), .B(n22949), .Z(n20713) );
  ANDN U24640 ( .B(n23420), .A(n20712), .Z(n24384) );
  XOR U24641 ( .A(n24386), .B(n22825), .Z(n20712) );
  XOR U24642 ( .A(n23505), .B(n24387), .Z(n23420) );
  XNOR U24643 ( .A(n24388), .B(n20726), .Z(n18794) );
  XOR U24644 ( .A(n24389), .B(n21601), .Z(n20726) );
  ANDN U24645 ( .B(n22118), .A(n20725), .Z(n24388) );
  XNOR U24646 ( .A(n24390), .B(n24391), .Z(n20725) );
  XOR U24647 ( .A(n24392), .B(n23964), .Z(n22118) );
  XNOR U24648 ( .A(n24393), .B(n20722), .Z(n19039) );
  XNOR U24649 ( .A(n24394), .B(n24395), .Z(n20722) );
  NOR U24650 ( .A(n20721), .B(n22123), .Z(n24393) );
  XOR U24651 ( .A(n24396), .B(n24397), .Z(n22123) );
  XOR U24652 ( .A(n24398), .B(n24399), .Z(n20721) );
  XOR U24653 ( .A(n24400), .B(n20737), .Z(n20559) );
  XOR U24654 ( .A(n24401), .B(n24402), .Z(n20737) );
  NOR U24655 ( .A(n24403), .B(n24363), .Z(n24400) );
  ANDN U24656 ( .B(n15036), .A(n16681), .Z(n24354) );
  XOR U24657 ( .A(n21628), .B(n19664), .Z(n16681) );
  XNOR U24658 ( .A(n19310), .B(n20123), .Z(n19664) );
  XOR U24659 ( .A(n24404), .B(n24405), .Z(n20123) );
  XOR U24660 ( .A(n18947), .B(n18315), .Z(n24405) );
  XNOR U24661 ( .A(n24406), .B(n22253), .Z(n18315) );
  IV U24662 ( .A(n20246), .Z(n22253) );
  XOR U24663 ( .A(n24407), .B(n24408), .Z(n20246) );
  NOR U24664 ( .A(n24409), .B(n20245), .Z(n24406) );
  XNOR U24665 ( .A(n24410), .B(n24411), .Z(n20245) );
  XOR U24666 ( .A(n24412), .B(n20471), .Z(n18947) );
  XOR U24667 ( .A(n24413), .B(n24414), .Z(n20471) );
  NOR U24668 ( .A(n24415), .B(n20478), .Z(n24412) );
  XNOR U24669 ( .A(n18722), .B(n24416), .Z(n24404) );
  XOR U24670 ( .A(n19946), .B(n17023), .Z(n24416) );
  XOR U24671 ( .A(n24417), .B(n20236), .Z(n17023) );
  XOR U24672 ( .A(n24418), .B(n24399), .Z(n20236) );
  NOR U24673 ( .A(n20235), .B(n21630), .Z(n24417) );
  XNOR U24674 ( .A(n24419), .B(n24420), .Z(n20235) );
  XNOR U24675 ( .A(n24421), .B(n20241), .Z(n19946) );
  XNOR U24676 ( .A(n23840), .B(n24422), .Z(n20241) );
  ANDN U24677 ( .B(n20242), .A(n21637), .Z(n24421) );
  XOR U24678 ( .A(n24423), .B(n24424), .Z(n20242) );
  XOR U24679 ( .A(n24425), .B(n20232), .Z(n18722) );
  XNOR U24680 ( .A(n24426), .B(n23597), .Z(n20232) );
  XOR U24681 ( .A(n24427), .B(n24428), .Z(n20231) );
  XOR U24682 ( .A(n24429), .B(n24430), .Z(n19310) );
  XNOR U24683 ( .A(n23959), .B(n21926), .Z(n24430) );
  XOR U24684 ( .A(n24431), .B(n21751), .Z(n21926) );
  XNOR U24685 ( .A(n24432), .B(n24433), .Z(n21751) );
  ANDN U24686 ( .B(n23971), .A(n23501), .Z(n24431) );
  IV U24687 ( .A(n21660), .Z(n23501) );
  XOR U24688 ( .A(n23422), .B(n24434), .Z(n21660) );
  IV U24689 ( .A(n21658), .Z(n23971) );
  XOR U24690 ( .A(n24435), .B(n23821), .Z(n21658) );
  XNOR U24691 ( .A(n24436), .B(n21748), .Z(n23959) );
  XOR U24692 ( .A(n24437), .B(n24438), .Z(n21748) );
  ANDN U24693 ( .B(n21647), .A(n21645), .Z(n24436) );
  XNOR U24694 ( .A(n24439), .B(n24440), .Z(n21645) );
  XOR U24695 ( .A(n24441), .B(n24427), .Z(n21647) );
  IV U24696 ( .A(n24442), .Z(n24427) );
  XOR U24697 ( .A(n17573), .B(n24443), .Z(n24429) );
  XNOR U24698 ( .A(n18730), .B(n22806), .Z(n24443) );
  XOR U24699 ( .A(n24444), .B(n21741), .Z(n22806) );
  ANDN U24700 ( .B(n21650), .A(n21649), .Z(n24444) );
  IV U24701 ( .A(n23975), .Z(n21649) );
  XOR U24702 ( .A(n24446), .B(n24447), .Z(n23975) );
  XOR U24703 ( .A(n24448), .B(n24449), .Z(n21650) );
  XOR U24704 ( .A(n24450), .B(n22662), .Z(n18730) );
  XOR U24705 ( .A(n23831), .B(n24451), .Z(n22662) );
  ANDN U24706 ( .B(n21662), .A(n21663), .Z(n24450) );
  XOR U24707 ( .A(n24452), .B(n24453), .Z(n21663) );
  XNOR U24708 ( .A(n24454), .B(n24455), .Z(n21662) );
  XNOR U24709 ( .A(n24456), .B(n21744), .Z(n17573) );
  XOR U24710 ( .A(n21713), .B(n24457), .Z(n21744) );
  XOR U24711 ( .A(n24458), .B(n24459), .Z(n21654) );
  XOR U24712 ( .A(n24460), .B(n24461), .Z(n21655) );
  XNOR U24713 ( .A(n24462), .B(n20478), .Z(n21628) );
  XOR U24714 ( .A(n24463), .B(n22892), .Z(n20478) );
  ANDN U24715 ( .B(n24415), .A(n24464), .Z(n24462) );
  XNOR U24716 ( .A(n20868), .B(n15256), .Z(n15036) );
  XOR U24717 ( .A(n24465), .B(n24466), .Z(n20868) );
  ANDN U24718 ( .B(n21674), .A(n24467), .Z(n24465) );
  XNOR U24719 ( .A(n24468), .B(n16689), .Z(n19474) );
  IV U24720 ( .A(n23661), .Z(n16689) );
  XNOR U24721 ( .A(n15342), .B(n23924), .Z(n23661) );
  XOR U24722 ( .A(n24469), .B(n24470), .Z(n23924) );
  ANDN U24723 ( .B(n21561), .A(n24471), .Z(n24469) );
  XOR U24724 ( .A(n21184), .B(n20852), .Z(n15342) );
  XNOR U24725 ( .A(n24472), .B(n24473), .Z(n20852) );
  XNOR U24726 ( .A(n16667), .B(n17002), .Z(n24473) );
  XNOR U24727 ( .A(n24474), .B(n24475), .Z(n17002) );
  ANDN U24728 ( .B(n21576), .A(n23926), .Z(n24474) );
  XOR U24729 ( .A(n24476), .B(n23974), .Z(n21576) );
  XNOR U24730 ( .A(n24477), .B(n24478), .Z(n16667) );
  ANDN U24731 ( .B(n24470), .A(n21559), .Z(n24477) );
  IV U24732 ( .A(n24471), .Z(n21559) );
  XOR U24733 ( .A(n22829), .B(n24479), .Z(n24471) );
  XOR U24734 ( .A(n16406), .B(n24480), .Z(n24472) );
  XOR U24735 ( .A(n18916), .B(n18532), .Z(n24480) );
  XNOR U24736 ( .A(n24481), .B(n24482), .Z(n18532) );
  ANDN U24737 ( .B(n24483), .A(n23934), .Z(n24481) );
  XOR U24738 ( .A(n24484), .B(n24485), .Z(n23934) );
  XNOR U24739 ( .A(n24486), .B(n24487), .Z(n18916) );
  XOR U24740 ( .A(n24488), .B(n23077), .Z(n21568) );
  XNOR U24741 ( .A(n24489), .B(n24490), .Z(n16406) );
  ANDN U24742 ( .B(n23929), .A(n21563), .Z(n24489) );
  XNOR U24743 ( .A(n24491), .B(n24492), .Z(n21563) );
  XOR U24744 ( .A(n24493), .B(n24494), .Z(n21184) );
  XNOR U24745 ( .A(n16148), .B(n18620), .Z(n24494) );
  XNOR U24746 ( .A(n24495), .B(n20616), .Z(n18620) );
  XNOR U24747 ( .A(n21229), .B(n24496), .Z(n20616) );
  XNOR U24748 ( .A(n24497), .B(n20627), .Z(n16148) );
  XOR U24749 ( .A(n24498), .B(n24499), .Z(n20627) );
  ANDN U24750 ( .B(n20626), .A(n21807), .Z(n24497) );
  IV U24751 ( .A(n24500), .Z(n21807) );
  XOR U24752 ( .A(n19504), .B(n24501), .Z(n24493) );
  XOR U24753 ( .A(n18790), .B(n20606), .Z(n24501) );
  XOR U24754 ( .A(n24502), .B(n23797), .Z(n20606) );
  XNOR U24755 ( .A(n24503), .B(n24438), .Z(n23797) );
  XOR U24756 ( .A(n24504), .B(n20622), .Z(n18790) );
  XNOR U24757 ( .A(n24505), .B(n23057), .Z(n20622) );
  IV U24758 ( .A(n24506), .Z(n23057) );
  ANDN U24759 ( .B(n20623), .A(n24507), .Z(n24504) );
  XNOR U24760 ( .A(n24508), .B(n23787), .Z(n19504) );
  IV U24761 ( .A(n20612), .Z(n23787) );
  XOR U24762 ( .A(n24509), .B(n23721), .Z(n20612) );
  ANDN U24763 ( .B(n15160), .A(n15159), .Z(n24468) );
  XOR U24764 ( .A(n15885), .B(n24510), .Z(n15159) );
  XNOR U24765 ( .A(n20597), .B(n19712), .Z(n15885) );
  XOR U24766 ( .A(n24511), .B(n24512), .Z(n19712) );
  XNOR U24767 ( .A(n18153), .B(n18253), .Z(n24512) );
  XOR U24768 ( .A(n24513), .B(n20563), .Z(n18253) );
  XOR U24769 ( .A(n24514), .B(n24515), .Z(n20563) );
  XNOR U24770 ( .A(n24516), .B(n20557), .Z(n18153) );
  XOR U24771 ( .A(n24517), .B(n24518), .Z(n20557) );
  ANDN U24772 ( .B(n20745), .A(n20558), .Z(n24516) );
  XOR U24773 ( .A(n20256), .B(n24519), .Z(n24511) );
  XOR U24774 ( .A(n17943), .B(n20378), .Z(n24519) );
  XOR U24775 ( .A(n24520), .B(n24363), .Z(n20378) );
  XNOR U24776 ( .A(n24521), .B(n23436), .Z(n24363) );
  ANDN U24777 ( .B(n20735), .A(n24522), .Z(n24520) );
  XNOR U24778 ( .A(n24523), .B(n20567), .Z(n17943) );
  XNOR U24779 ( .A(n24524), .B(n24525), .Z(n20567) );
  ANDN U24780 ( .B(n20568), .A(n20741), .Z(n24523) );
  XNOR U24781 ( .A(n24526), .B(n20553), .Z(n20256) );
  XNOR U24782 ( .A(n22346), .B(n24527), .Z(n20553) );
  IV U24783 ( .A(n24528), .Z(n22346) );
  ANDN U24784 ( .B(n20554), .A(n23257), .Z(n24526) );
  XOR U24785 ( .A(n24529), .B(n24530), .Z(n20597) );
  XNOR U24786 ( .A(n19518), .B(n20547), .Z(n24530) );
  XOR U24787 ( .A(n24531), .B(n24532), .Z(n20547) );
  NOR U24788 ( .A(n24533), .B(n24534), .Z(n24531) );
  XNOR U24789 ( .A(n24535), .B(n22865), .Z(n19518) );
  NOR U24790 ( .A(n24536), .B(n22370), .Z(n24535) );
  XOR U24791 ( .A(n19441), .B(n24537), .Z(n24529) );
  XNOR U24792 ( .A(n19401), .B(n18622), .Z(n24537) );
  XOR U24793 ( .A(n24538), .B(n22872), .Z(n18622) );
  NOR U24794 ( .A(n22376), .B(n24539), .Z(n24538) );
  IV U24795 ( .A(n24540), .Z(n22376) );
  XOR U24796 ( .A(n24541), .B(n22862), .Z(n19401) );
  NOR U24797 ( .A(n22380), .B(n24542), .Z(n24541) );
  IV U24798 ( .A(n24543), .Z(n22380) );
  XNOR U24799 ( .A(n24544), .B(n22860), .Z(n19441) );
  ANDN U24800 ( .B(n24545), .A(n22366), .Z(n24544) );
  IV U24801 ( .A(n24546), .Z(n22366) );
  XNOR U24802 ( .A(n19864), .B(n18830), .Z(n15160) );
  XOR U24803 ( .A(n23497), .B(n24547), .Z(n18830) );
  XOR U24804 ( .A(n24548), .B(n24549), .Z(n23497) );
  XOR U24805 ( .A(n18776), .B(n20040), .Z(n24549) );
  XNOR U24806 ( .A(n24550), .B(n21637), .Z(n20040) );
  XOR U24807 ( .A(n23326), .B(n24551), .Z(n21637) );
  ANDN U24808 ( .B(n20240), .A(n20475), .Z(n24550) );
  IV U24809 ( .A(n21638), .Z(n20475) );
  XOR U24810 ( .A(n24552), .B(n24150), .Z(n21638) );
  XNOR U24811 ( .A(n24553), .B(n24554), .Z(n20240) );
  XNOR U24812 ( .A(n24555), .B(n24415), .Z(n18776) );
  XNOR U24813 ( .A(n24556), .B(n23429), .Z(n24415) );
  NOR U24814 ( .A(n20469), .B(n20470), .Z(n24555) );
  XNOR U24815 ( .A(n24557), .B(n24558), .Z(n20470) );
  IV U24816 ( .A(n24464), .Z(n20469) );
  XOR U24817 ( .A(n22223), .B(n24559), .Z(n24464) );
  XNOR U24818 ( .A(n20633), .B(n24560), .Z(n24548) );
  XNOR U24819 ( .A(n19633), .B(n21625), .Z(n24560) );
  XNOR U24820 ( .A(n24561), .B(n21630), .Z(n21625) );
  XOR U24821 ( .A(n24562), .B(n24563), .Z(n21630) );
  ANDN U24822 ( .B(n20234), .A(n20473), .Z(n24561) );
  IV U24823 ( .A(n21631), .Z(n20473) );
  XOR U24824 ( .A(n24564), .B(n24381), .Z(n21631) );
  XOR U24825 ( .A(n24565), .B(n24566), .Z(n20234) );
  XOR U24826 ( .A(n24567), .B(n24409), .Z(n19633) );
  IV U24827 ( .A(n21634), .Z(n24409) );
  XOR U24828 ( .A(n24458), .B(n24568), .Z(n21634) );
  ANDN U24829 ( .B(n21635), .A(n20244), .Z(n24567) );
  XOR U24830 ( .A(n24569), .B(n24570), .Z(n20244) );
  XOR U24831 ( .A(n24571), .B(n24572), .Z(n21635) );
  XOR U24832 ( .A(n24573), .B(n21641), .Z(n20633) );
  XOR U24833 ( .A(n24574), .B(n24575), .Z(n21641) );
  NOR U24834 ( .A(n20230), .B(n21640), .Z(n24573) );
  XOR U24835 ( .A(n24576), .B(n24577), .Z(n21640) );
  XOR U24836 ( .A(n22495), .B(n24578), .Z(n20230) );
  XNOR U24837 ( .A(n24579), .B(n24580), .Z(n19864) );
  AND U24838 ( .A(n21588), .B(n20401), .Z(n24579) );
  XOR U24839 ( .A(n24581), .B(n24582), .Z(n20401) );
  ANDN U24840 ( .B(n7132), .A(n9323), .Z(n23629) );
  XOR U24841 ( .A(n15175), .B(n11842), .Z(n9323) );
  IV U24842 ( .A(n11714), .Z(n11842) );
  XOR U24843 ( .A(n14475), .B(n12625), .Z(n11714) );
  XOR U24844 ( .A(n24583), .B(n24584), .Z(n12625) );
  XNOR U24845 ( .A(n12760), .B(n12974), .Z(n24584) );
  XNOR U24846 ( .A(n24585), .B(n15310), .Z(n12974) );
  XOR U24847 ( .A(n18277), .B(n23636), .Z(n15310) );
  XNOR U24848 ( .A(n24586), .B(n23545), .Z(n23636) );
  NOR U24849 ( .A(n22725), .B(n24587), .Z(n24586) );
  XNOR U24850 ( .A(n20016), .B(n21348), .Z(n18277) );
  XOR U24851 ( .A(n24588), .B(n24589), .Z(n21348) );
  XNOR U24852 ( .A(n20027), .B(n18928), .Z(n24589) );
  XNOR U24853 ( .A(n24590), .B(n22739), .Z(n18928) );
  XOR U24854 ( .A(n24591), .B(n24420), .Z(n22739) );
  NOR U24855 ( .A(n23650), .B(n23539), .Z(n24590) );
  XNOR U24856 ( .A(n24592), .B(n22990), .Z(n23539) );
  XOR U24857 ( .A(n24593), .B(n22742), .Z(n20027) );
  XNOR U24858 ( .A(n24594), .B(n24595), .Z(n22742) );
  NOR U24859 ( .A(n23535), .B(n23652), .Z(n24593) );
  XOR U24860 ( .A(n24596), .B(n24597), .Z(n23535) );
  XOR U24861 ( .A(n20486), .B(n24598), .Z(n24588) );
  XNOR U24862 ( .A(n19486), .B(n16612), .Z(n24598) );
  XNOR U24863 ( .A(n24599), .B(n22734), .Z(n16612) );
  NOR U24864 ( .A(n24601), .B(n23528), .Z(n24599) );
  XNOR U24865 ( .A(n24602), .B(n23584), .Z(n23528) );
  XOR U24866 ( .A(n24603), .B(n22747), .Z(n19486) );
  XOR U24867 ( .A(n24604), .B(n24278), .Z(n22747) );
  NOR U24868 ( .A(n23657), .B(n23537), .Z(n24603) );
  XOR U24869 ( .A(n24605), .B(n24606), .Z(n23537) );
  XNOR U24870 ( .A(n24607), .B(n23532), .Z(n20486) );
  ANDN U24871 ( .B(n23660), .A(n23531), .Z(n24607) );
  XOR U24872 ( .A(n24446), .B(n24608), .Z(n23531) );
  XOR U24873 ( .A(n24609), .B(n24610), .Z(n20016) );
  XNOR U24874 ( .A(n16508), .B(n23524), .Z(n24610) );
  XNOR U24875 ( .A(n24611), .B(n22713), .Z(n23524) );
  XOR U24876 ( .A(n24072), .B(n24612), .Z(n22713) );
  IV U24877 ( .A(n24613), .Z(n24072) );
  XOR U24878 ( .A(n24614), .B(n22337), .Z(n23548) );
  XOR U24879 ( .A(n24615), .B(n22727), .Z(n16508) );
  XNOR U24880 ( .A(n24241), .B(n24616), .Z(n22727) );
  ANDN U24881 ( .B(n24587), .A(n23545), .Z(n24615) );
  XOR U24882 ( .A(n24617), .B(n24618), .Z(n23545) );
  XNOR U24883 ( .A(n19258), .B(n24619), .Z(n24609) );
  XOR U24884 ( .A(n19554), .B(n19226), .Z(n24619) );
  XNOR U24885 ( .A(n24620), .B(n22722), .Z(n19226) );
  XOR U24886 ( .A(n24621), .B(n24622), .Z(n22722) );
  NOR U24887 ( .A(n23641), .B(n23543), .Z(n24620) );
  XOR U24888 ( .A(n24623), .B(n24624), .Z(n23543) );
  XOR U24889 ( .A(n24625), .B(n22719), .Z(n19554) );
  XOR U24890 ( .A(n24626), .B(n24627), .Z(n22719) );
  NOR U24891 ( .A(n23638), .B(n23550), .Z(n24625) );
  XOR U24892 ( .A(n24628), .B(n24629), .Z(n23550) );
  XNOR U24893 ( .A(n24630), .B(n22710), .Z(n19258) );
  XOR U24894 ( .A(n24631), .B(n24632), .Z(n22710) );
  ANDN U24895 ( .B(n23553), .A(n23646), .Z(n24630) );
  XOR U24896 ( .A(n24633), .B(n24634), .Z(n23553) );
  NOR U24897 ( .A(n15311), .B(n16587), .Z(n24585) );
  XNOR U24898 ( .A(n21259), .B(n18234), .Z(n16587) );
  XNOR U24899 ( .A(n24635), .B(n24636), .Z(n20988) );
  XNOR U24900 ( .A(n18173), .B(n17296), .Z(n24636) );
  XNOR U24901 ( .A(n24637), .B(n24155), .Z(n17296) );
  NOR U24902 ( .A(n23897), .B(n24096), .Z(n24637) );
  IV U24903 ( .A(n24097), .Z(n23897) );
  XOR U24904 ( .A(n24528), .B(n24638), .Z(n24097) );
  XNOR U24905 ( .A(n24639), .B(n24640), .Z(n18173) );
  NOR U24906 ( .A(n21268), .B(n21269), .Z(n24639) );
  XNOR U24907 ( .A(n24571), .B(n24641), .Z(n21269) );
  XOR U24908 ( .A(n24642), .B(n24643), .Z(n24635) );
  XNOR U24909 ( .A(n19251), .B(n19096), .Z(n24643) );
  XOR U24910 ( .A(n24644), .B(n24140), .Z(n19096) );
  ANDN U24911 ( .B(n21526), .A(n21527), .Z(n24644) );
  XNOR U24912 ( .A(n23335), .B(n24645), .Z(n21527) );
  XNOR U24913 ( .A(n24646), .B(n24142), .Z(n19251) );
  ANDN U24914 ( .B(n24647), .A(n23887), .Z(n24646) );
  IV U24915 ( .A(n24648), .Z(n23887) );
  XNOR U24916 ( .A(n24649), .B(n24650), .Z(n23477) );
  XNOR U24917 ( .A(n18647), .B(n17981), .Z(n24650) );
  XOR U24918 ( .A(n24651), .B(n24054), .Z(n17981) );
  AND U24919 ( .A(n23476), .B(n23474), .Z(n24651) );
  XOR U24920 ( .A(n24652), .B(n24653), .Z(n18647) );
  NOR U24921 ( .A(n24654), .B(n22065), .Z(n24652) );
  XOR U24922 ( .A(n19723), .B(n24655), .Z(n24649) );
  XNOR U24923 ( .A(n16857), .B(n18960), .Z(n24655) );
  XNOR U24924 ( .A(n24656), .B(n24050), .Z(n18960) );
  ANDN U24925 ( .B(n22075), .A(n22076), .Z(n24656) );
  XNOR U24926 ( .A(n24657), .B(n24059), .Z(n16857) );
  ANDN U24927 ( .B(n22061), .A(n22062), .Z(n24657) );
  XOR U24928 ( .A(n24658), .B(n24047), .Z(n19723) );
  NOR U24929 ( .A(n22072), .B(n22071), .Z(n24658) );
  XOR U24930 ( .A(n24659), .B(n24647), .Z(n21259) );
  ANDN U24931 ( .B(n23889), .A(n24648), .Z(n24659) );
  XOR U24932 ( .A(n24660), .B(n24661), .Z(n24648) );
  XNOR U24933 ( .A(n24662), .B(n24663), .Z(n23889) );
  XOR U24934 ( .A(n21825), .B(n17744), .Z(n15311) );
  XNOR U24935 ( .A(n24666), .B(n23762), .Z(n21825) );
  ANDN U24936 ( .B(n21343), .A(n21344), .Z(n24666) );
  XOR U24937 ( .A(n24667), .B(n23710), .Z(n21344) );
  XNOR U24938 ( .A(n24668), .B(n15328), .Z(n12760) );
  XOR U24939 ( .A(n24119), .B(n17861), .Z(n15328) );
  XNOR U24940 ( .A(n19135), .B(n20049), .Z(n17861) );
  XNOR U24941 ( .A(n24669), .B(n24670), .Z(n20049) );
  XNOR U24942 ( .A(n22657), .B(n18381), .Z(n24670) );
  XNOR U24943 ( .A(n24671), .B(n24672), .Z(n18381) );
  NOR U24944 ( .A(n24673), .B(n24133), .Z(n24671) );
  XOR U24945 ( .A(n24674), .B(n21429), .Z(n22657) );
  ANDN U24946 ( .B(n24675), .A(n24676), .Z(n24674) );
  XOR U24947 ( .A(n18104), .B(n24677), .Z(n24669) );
  XOR U24948 ( .A(n19789), .B(n24678), .Z(n24677) );
  XNOR U24949 ( .A(n24679), .B(n21424), .Z(n19789) );
  XNOR U24950 ( .A(n24680), .B(n22277), .Z(n18104) );
  ANDN U24951 ( .B(n24122), .A(n24121), .Z(n24680) );
  XOR U24952 ( .A(n24681), .B(n24682), .Z(n19135) );
  XOR U24953 ( .A(n16393), .B(n24683), .Z(n24682) );
  XNOR U24954 ( .A(n24684), .B(n22302), .Z(n16393) );
  ANDN U24955 ( .B(n24105), .A(n24106), .Z(n24684) );
  XOR U24956 ( .A(n16031), .B(n24685), .Z(n24681) );
  XNOR U24957 ( .A(n18870), .B(n17651), .Z(n24685) );
  XNOR U24958 ( .A(n24686), .B(n22292), .Z(n17651) );
  ANDN U24959 ( .B(n24113), .A(n24687), .Z(n24686) );
  XNOR U24960 ( .A(n24688), .B(n22306), .Z(n18870) );
  AND U24961 ( .A(n24103), .B(n24102), .Z(n24688) );
  XOR U24962 ( .A(n24689), .B(n22298), .Z(n16031) );
  NOR U24963 ( .A(n24116), .B(n24115), .Z(n24689) );
  XOR U24964 ( .A(n24690), .B(n24675), .Z(n24119) );
  ANDN U24965 ( .B(n24676), .A(n24691), .Z(n24690) );
  NOR U24966 ( .A(n16573), .B(n15327), .Z(n24668) );
  XOR U24967 ( .A(n21272), .B(n20857), .Z(n15327) );
  XNOR U24968 ( .A(n24692), .B(n24693), .Z(n20857) );
  NOR U24969 ( .A(n23944), .B(n21545), .Z(n24692) );
  XOR U24970 ( .A(n24694), .B(n24695), .Z(n21545) );
  XNOR U24971 ( .A(n18917), .B(n23154), .Z(n21272) );
  XNOR U24972 ( .A(n24696), .B(n24697), .Z(n23154) );
  XOR U24973 ( .A(n14167), .B(n17731), .Z(n24697) );
  XOR U24974 ( .A(n24698), .B(n23953), .Z(n17731) );
  AND U24975 ( .A(n20937), .B(n20935), .Z(n24698) );
  XOR U24976 ( .A(n24699), .B(n24700), .Z(n20937) );
  XNOR U24977 ( .A(n24701), .B(n21555), .Z(n14167) );
  AND U24978 ( .A(n21274), .B(n21276), .Z(n24701) );
  XNOR U24979 ( .A(n24702), .B(n24703), .Z(n21276) );
  XOR U24980 ( .A(n18913), .B(n24704), .Z(n24696) );
  XOR U24981 ( .A(n17971), .B(n24705), .Z(n24704) );
  XOR U24982 ( .A(n24706), .B(n21547), .Z(n17971) );
  IV U24983 ( .A(n24707), .Z(n21547) );
  AND U24984 ( .A(n23944), .B(n24693), .Z(n24706) );
  XOR U24985 ( .A(n24708), .B(n24709), .Z(n23944) );
  XNOR U24986 ( .A(n24710), .B(n21551), .Z(n18913) );
  ANDN U24987 ( .B(n22328), .A(n22329), .Z(n24710) );
  XOR U24988 ( .A(n24711), .B(n24712), .Z(n22329) );
  XOR U24989 ( .A(n24713), .B(n24714), .Z(n18917) );
  XNOR U24990 ( .A(n18196), .B(n18795), .Z(n24714) );
  XNOR U24991 ( .A(n24715), .B(n21570), .Z(n18795) );
  ANDN U24992 ( .B(n24487), .A(n23931), .Z(n24715) );
  XOR U24993 ( .A(n24716), .B(n24709), .Z(n23931) );
  XNOR U24994 ( .A(n24717), .B(n21578), .Z(n18196) );
  XNOR U24995 ( .A(n24718), .B(n22396), .Z(n23926) );
  XNOR U24996 ( .A(n21389), .B(n24719), .Z(n24713) );
  XNOR U24997 ( .A(n19429), .B(n16510), .Z(n24719) );
  XOR U24998 ( .A(n24720), .B(n21573), .Z(n16510) );
  ANDN U24999 ( .B(n24482), .A(n24483), .Z(n24720) );
  IV U25000 ( .A(n23933), .Z(n24483) );
  XOR U25001 ( .A(n24721), .B(n24182), .Z(n23933) );
  XOR U25002 ( .A(n24722), .B(n21565), .Z(n19429) );
  ANDN U25003 ( .B(n24490), .A(n23929), .Z(n24722) );
  XNOR U25004 ( .A(n23998), .B(n24723), .Z(n23929) );
  XOR U25005 ( .A(n24724), .B(n21560), .Z(n21389) );
  ANDN U25006 ( .B(n24478), .A(n24470), .Z(n24724) );
  XOR U25007 ( .A(n24725), .B(n22012), .Z(n24470) );
  XNOR U25008 ( .A(n24299), .B(n18337), .Z(n16573) );
  IV U25009 ( .A(n17961), .Z(n18337) );
  XOR U25010 ( .A(n24726), .B(n22880), .Z(n17961) );
  XNOR U25011 ( .A(n24727), .B(n24728), .Z(n22880) );
  XNOR U25012 ( .A(n16734), .B(n14993), .Z(n24728) );
  XNOR U25013 ( .A(n24729), .B(n21204), .Z(n14993) );
  ANDN U25014 ( .B(n21205), .A(n22541), .Z(n24729) );
  XOR U25015 ( .A(n24730), .B(n20945), .Z(n16734) );
  ANDN U25016 ( .B(n20946), .A(n24731), .Z(n24730) );
  XOR U25017 ( .A(n19043), .B(n24732), .Z(n24727) );
  XOR U25018 ( .A(n19821), .B(n17783), .Z(n24732) );
  XNOR U25019 ( .A(n24733), .B(n20955), .Z(n17783) );
  ANDN U25020 ( .B(n20956), .A(n22552), .Z(n24733) );
  XNOR U25021 ( .A(n24734), .B(n20950), .Z(n19821) );
  NOR U25022 ( .A(n22544), .B(n20949), .Z(n24734) );
  XOR U25023 ( .A(n24735), .B(n20959), .Z(n19043) );
  ANDN U25024 ( .B(n24736), .A(n20960), .Z(n24735) );
  XOR U25025 ( .A(n24737), .B(n24738), .Z(n24299) );
  ANDN U25026 ( .B(n22559), .A(n22557), .Z(n24737) );
  XOR U25027 ( .A(n15282), .B(n24739), .Z(n24583) );
  XOR U25028 ( .A(n9621), .B(n11179), .Z(n24739) );
  XNOR U25029 ( .A(n24740), .B(n15324), .Z(n11179) );
  XNOR U25030 ( .A(n24052), .B(n17013), .Z(n15324) );
  XNOR U25031 ( .A(n19085), .B(n23386), .Z(n17013) );
  XNOR U25032 ( .A(n24741), .B(n24742), .Z(n23386) );
  XNOR U25033 ( .A(n18453), .B(n19984), .Z(n24742) );
  XNOR U25034 ( .A(n24743), .B(n22076), .Z(n19984) );
  XNOR U25035 ( .A(n24744), .B(n24745), .Z(n22076) );
  XOR U25036 ( .A(n24746), .B(n24747), .Z(n22077) );
  XOR U25037 ( .A(n24748), .B(n23476), .Z(n18453) );
  XOR U25038 ( .A(n24749), .B(n24750), .Z(n23476) );
  NOR U25039 ( .A(n24751), .B(n23475), .Z(n24748) );
  XOR U25040 ( .A(n24076), .B(n24752), .Z(n23475) );
  IV U25041 ( .A(n22829), .Z(n24076) );
  XNOR U25042 ( .A(n22034), .B(n24753), .Z(n24741) );
  XNOR U25043 ( .A(n15695), .B(n19396), .Z(n24753) );
  XOR U25044 ( .A(n24754), .B(n22072), .Z(n19396) );
  XOR U25045 ( .A(n24755), .B(n24756), .Z(n22072) );
  XOR U25046 ( .A(n24605), .B(n24757), .Z(n22073) );
  XNOR U25047 ( .A(n24758), .B(n22062), .Z(n15695) );
  XNOR U25048 ( .A(n24759), .B(n22394), .Z(n22062) );
  ANDN U25049 ( .B(n24058), .A(n24057), .Z(n24758) );
  XOR U25050 ( .A(n24760), .B(n24761), .Z(n24057) );
  XOR U25051 ( .A(n24762), .B(n22067), .Z(n22034) );
  IV U25052 ( .A(n24654), .Z(n22067) );
  XOR U25053 ( .A(n23951), .B(n24763), .Z(n24654) );
  NOR U25054 ( .A(n24764), .B(n22066), .Z(n24762) );
  XOR U25055 ( .A(n24765), .B(n24766), .Z(n19085) );
  XOR U25056 ( .A(n20883), .B(n18176), .Z(n24766) );
  XNOR U25057 ( .A(n24767), .B(n22052), .Z(n18176) );
  XOR U25058 ( .A(n24768), .B(n24769), .Z(n22052) );
  ANDN U25059 ( .B(n22158), .A(n22053), .Z(n24767) );
  XOR U25060 ( .A(n24770), .B(n23788), .Z(n22053) );
  XNOR U25061 ( .A(n24771), .B(n24772), .Z(n22158) );
  XNOR U25062 ( .A(n24773), .B(n22056), .Z(n20883) );
  XOR U25063 ( .A(n24774), .B(n23566), .Z(n22056) );
  XOR U25064 ( .A(n24775), .B(n24776), .Z(n22151) );
  XOR U25065 ( .A(n24777), .B(n24778), .Z(n22057) );
  XOR U25066 ( .A(n18632), .B(n24779), .Z(n24765) );
  XOR U25067 ( .A(n18866), .B(n18585), .Z(n24779) );
  XOR U25068 ( .A(n24780), .B(n22043), .Z(n18585) );
  XOR U25069 ( .A(n22223), .B(n24781), .Z(n22043) );
  XOR U25070 ( .A(n24782), .B(n24783), .Z(n22044) );
  XNOR U25071 ( .A(n24784), .B(n24247), .Z(n22162) );
  XNOR U25072 ( .A(n24785), .B(n22049), .Z(n18866) );
  XOR U25073 ( .A(n24786), .B(n24595), .Z(n22049) );
  IV U25074 ( .A(n21721), .Z(n24595) );
  ANDN U25075 ( .B(n22148), .A(n22048), .Z(n24785) );
  XNOR U25076 ( .A(n24787), .B(n24788), .Z(n22048) );
  XOR U25077 ( .A(n23946), .B(n24789), .Z(n22148) );
  NOR U25078 ( .A(n22039), .B(n22155), .Z(n24790) );
  XOR U25079 ( .A(n24792), .B(n24793), .Z(n22155) );
  XNOR U25080 ( .A(n24794), .B(n24795), .Z(n22039) );
  XNOR U25081 ( .A(n24796), .B(n22066), .Z(n24052) );
  XNOR U25082 ( .A(n24797), .B(n24798), .Z(n22066) );
  NOR U25083 ( .A(n15323), .B(n16577), .Z(n24740) );
  XOR U25084 ( .A(n24799), .B(n18419), .Z(n16577) );
  XOR U25085 ( .A(n20582), .B(n18508), .Z(n15323) );
  IV U25086 ( .A(n18219), .Z(n18508) );
  XOR U25087 ( .A(n24547), .B(n19136), .Z(n18219) );
  XOR U25088 ( .A(n24800), .B(n24801), .Z(n19136) );
  XOR U25089 ( .A(n17865), .B(n17581), .Z(n24801) );
  XNOR U25090 ( .A(n24802), .B(n22326), .Z(n17581) );
  XOR U25091 ( .A(n23035), .B(n24803), .Z(n20576) );
  IV U25092 ( .A(n24439), .Z(n23035) );
  XNOR U25093 ( .A(n24804), .B(n22311), .Z(n17865) );
  XNOR U25094 ( .A(n14175), .B(n24806), .Z(n24800) );
  XNOR U25095 ( .A(n16891), .B(n18924), .Z(n24806) );
  XNOR U25096 ( .A(n24807), .B(n22322), .Z(n18924) );
  ANDN U25097 ( .B(n24808), .A(n21615), .Z(n24807) );
  XNOR U25098 ( .A(n24809), .B(n22320), .Z(n16891) );
  XOR U25099 ( .A(n24810), .B(n23864), .Z(n20585) );
  XOR U25100 ( .A(n24811), .B(n24812), .Z(n14175) );
  NOR U25101 ( .A(n20588), .B(n20589), .Z(n24811) );
  XOR U25102 ( .A(n24040), .B(n24813), .Z(n20589) );
  XOR U25103 ( .A(n24814), .B(n24815), .Z(n24547) );
  XOR U25104 ( .A(n18158), .B(n17029), .Z(n24815) );
  XNOR U25105 ( .A(n24816), .B(n20127), .Z(n17029) );
  XOR U25106 ( .A(n24817), .B(n24172), .Z(n20127) );
  ANDN U25107 ( .B(n19870), .A(n19871), .Z(n24816) );
  XOR U25108 ( .A(n22223), .B(n24818), .Z(n19871) );
  XOR U25109 ( .A(n24819), .B(n24820), .Z(n19870) );
  XNOR U25110 ( .A(n24821), .B(n20004), .Z(n18158) );
  XOR U25111 ( .A(n24822), .B(n24823), .Z(n20004) );
  NOR U25112 ( .A(n24580), .B(n21588), .Z(n24821) );
  XNOR U25113 ( .A(n24824), .B(n24825), .Z(n21588) );
  IV U25114 ( .A(n20005), .Z(n24580) );
  XOR U25115 ( .A(n24826), .B(n24827), .Z(n20005) );
  XOR U25116 ( .A(n19988), .B(n24828), .Z(n24814) );
  XOR U25117 ( .A(n19259), .B(n18284), .Z(n24828) );
  XNOR U25118 ( .A(n24829), .B(n20001), .Z(n18284) );
  XOR U25119 ( .A(n24830), .B(n23582), .Z(n20001) );
  ANDN U25120 ( .B(n19862), .A(n19860), .Z(n24829) );
  XOR U25121 ( .A(n24831), .B(n22025), .Z(n19860) );
  XNOR U25122 ( .A(n24832), .B(n24570), .Z(n19862) );
  XNOR U25123 ( .A(n24833), .B(n19996), .Z(n19259) );
  XOR U25124 ( .A(n24834), .B(n24835), .Z(n19996) );
  ANDN U25125 ( .B(n19856), .A(n19858), .Z(n24833) );
  XOR U25126 ( .A(n24836), .B(n24837), .Z(n19858) );
  XNOR U25127 ( .A(n24838), .B(n24839), .Z(n19856) );
  XNOR U25128 ( .A(n24840), .B(n19993), .Z(n19988) );
  XOR U25129 ( .A(n24841), .B(n24842), .Z(n19993) );
  ANDN U25130 ( .B(n19868), .A(n19866), .Z(n24840) );
  XOR U25131 ( .A(n24843), .B(n24844), .Z(n19866) );
  XOR U25132 ( .A(n24845), .B(n24846), .Z(n19868) );
  XNOR U25133 ( .A(n24847), .B(n24808), .Z(n20582) );
  ANDN U25134 ( .B(n21615), .A(n21616), .Z(n24847) );
  XOR U25135 ( .A(n24848), .B(n24849), .Z(n21616) );
  XOR U25136 ( .A(n24851), .B(n15314), .Z(n9621) );
  XOR U25137 ( .A(n23290), .B(n18033), .Z(n15314) );
  IV U25138 ( .A(n18949), .Z(n18033) );
  XNOR U25139 ( .A(n20248), .B(n20596), .Z(n18949) );
  XNOR U25140 ( .A(n24852), .B(n24853), .Z(n20596) );
  XNOR U25141 ( .A(n17927), .B(n19560), .Z(n24853) );
  XOR U25142 ( .A(n24854), .B(n24855), .Z(n19560) );
  NOR U25143 ( .A(n24087), .B(n23277), .Z(n24854) );
  IV U25144 ( .A(n23279), .Z(n24087) );
  XOR U25145 ( .A(n24856), .B(n24857), .Z(n23279) );
  XOR U25146 ( .A(n24858), .B(n24859), .Z(n17927) );
  ANDN U25147 ( .B(n23268), .A(n23266), .Z(n24858) );
  XOR U25148 ( .A(n24860), .B(n24861), .Z(n23268) );
  XOR U25149 ( .A(n24862), .B(n24863), .Z(n24852) );
  XNOR U25150 ( .A(n19290), .B(n17620), .Z(n24863) );
  XOR U25151 ( .A(n24864), .B(n24865), .Z(n17620) );
  ANDN U25152 ( .B(n23285), .A(n24092), .Z(n24864) );
  IV U25153 ( .A(n23287), .Z(n24092) );
  XOR U25154 ( .A(n24866), .B(n23059), .Z(n23287) );
  XOR U25155 ( .A(n24867), .B(n24868), .Z(n19290) );
  ANDN U25156 ( .B(n23281), .A(n23282), .Z(n24867) );
  XOR U25157 ( .A(n24869), .B(n22536), .Z(n23282) );
  XOR U25158 ( .A(n24870), .B(n24871), .Z(n20248) );
  XOR U25159 ( .A(n19007), .B(n20701), .Z(n24871) );
  XOR U25160 ( .A(n24872), .B(n23166), .Z(n20701) );
  XOR U25161 ( .A(n24873), .B(n24874), .Z(n23167) );
  XNOR U25162 ( .A(n24875), .B(n24876), .Z(n19007) );
  ANDN U25163 ( .B(n24877), .A(n24878), .Z(n24875) );
  XNOR U25164 ( .A(n19660), .B(n24879), .Z(n24870) );
  XOR U25165 ( .A(n23157), .B(n18556), .Z(n24879) );
  XNOR U25166 ( .A(n24880), .B(n23177), .Z(n18556) );
  NOR U25167 ( .A(n23178), .B(n23299), .Z(n24880) );
  XOR U25168 ( .A(n21713), .B(n24881), .Z(n23178) );
  XNOR U25169 ( .A(n24882), .B(n23173), .Z(n23157) );
  XOR U25170 ( .A(n24883), .B(n24884), .Z(n23172) );
  XOR U25171 ( .A(n24885), .B(n23163), .Z(n19660) );
  NOR U25172 ( .A(n23303), .B(n23162), .Z(n24885) );
  XOR U25173 ( .A(n22643), .B(n24886), .Z(n23162) );
  XNOR U25174 ( .A(n24887), .B(n24888), .Z(n23290) );
  ANDN U25175 ( .B(n24889), .A(n24877), .Z(n24887) );
  ANDN U25176 ( .B(n18205), .A(n18250), .Z(n24851) );
  XOR U25177 ( .A(n20271), .B(n16954), .Z(n18250) );
  XOR U25178 ( .A(n24890), .B(n23006), .Z(n16954) );
  XOR U25179 ( .A(n24891), .B(n24892), .Z(n23006) );
  XNOR U25180 ( .A(n24893), .B(n17631), .Z(n24892) );
  XOR U25181 ( .A(n24894), .B(n23624), .Z(n17631) );
  ANDN U25182 ( .B(n24895), .A(n21939), .Z(n24894) );
  IV U25183 ( .A(n24896), .Z(n21939) );
  XOR U25184 ( .A(n19500), .B(n24897), .Z(n24891) );
  XOR U25185 ( .A(n19433), .B(n20142), .Z(n24897) );
  XNOR U25186 ( .A(n24898), .B(n23622), .Z(n20142) );
  ANDN U25187 ( .B(n20264), .A(n20262), .Z(n24898) );
  XOR U25188 ( .A(n24899), .B(n24900), .Z(n20264) );
  XNOR U25189 ( .A(n24901), .B(n23618), .Z(n19433) );
  NOR U25190 ( .A(n21946), .B(n22701), .Z(n24901) );
  IV U25191 ( .A(n22702), .Z(n21946) );
  XOR U25192 ( .A(n24903), .B(n23628), .Z(n19500) );
  ANDN U25193 ( .B(n20275), .A(n20273), .Z(n24903) );
  XNOR U25194 ( .A(n24904), .B(n24905), .Z(n20275) );
  XNOR U25195 ( .A(n24906), .B(n24895), .Z(n20271) );
  ANDN U25196 ( .B(n21940), .A(n24896), .Z(n24906) );
  XOR U25197 ( .A(n24907), .B(n24700), .Z(n24896) );
  IV U25198 ( .A(n24908), .Z(n24700) );
  XOR U25199 ( .A(n24909), .B(n21819), .Z(n21940) );
  XOR U25200 ( .A(n24910), .B(n17853), .Z(n18205) );
  XNOR U25201 ( .A(n24911), .B(n15320), .Z(n15282) );
  XNOR U25202 ( .A(n20448), .B(n17093), .Z(n15320) );
  XNOR U25203 ( .A(n21092), .B(n21835), .Z(n17093) );
  XNOR U25204 ( .A(n24912), .B(n24913), .Z(n21835) );
  XOR U25205 ( .A(n15649), .B(n17997), .Z(n24913) );
  XOR U25206 ( .A(n24914), .B(n19417), .Z(n17997) );
  XOR U25207 ( .A(n24915), .B(n24916), .Z(n19417) );
  XOR U25208 ( .A(n24917), .B(n23582), .Z(n21854) );
  XOR U25209 ( .A(n24918), .B(n23244), .Z(n21855) );
  XOR U25210 ( .A(n24919), .B(n22673), .Z(n15649) );
  XOR U25211 ( .A(n24626), .B(n24920), .Z(n22673) );
  AND U25212 ( .A(n20512), .B(n20511), .Z(n24919) );
  XNOR U25213 ( .A(n24921), .B(n23494), .Z(n20511) );
  IV U25214 ( .A(n23024), .Z(n23494) );
  XNOR U25215 ( .A(n23145), .B(n24922), .Z(n20512) );
  XOR U25216 ( .A(n17396), .B(n24923), .Z(n24912) );
  XOR U25217 ( .A(n16495), .B(n21280), .Z(n24923) );
  XOR U25218 ( .A(n24924), .B(n22680), .Z(n21280) );
  XOR U25219 ( .A(n24925), .B(n24926), .Z(n22680) );
  AND U25220 ( .A(n20503), .B(n20501), .Z(n24924) );
  XNOR U25221 ( .A(n24927), .B(n24399), .Z(n20501) );
  XOR U25222 ( .A(n24928), .B(n23568), .Z(n20503) );
  XNOR U25223 ( .A(n24929), .B(n21042), .Z(n16495) );
  IV U25224 ( .A(n22677), .Z(n21042) );
  XOR U25225 ( .A(n24930), .B(n24931), .Z(n22677) );
  ANDN U25226 ( .B(n20505), .A(n20506), .Z(n24929) );
  XOR U25227 ( .A(n24932), .B(n22342), .Z(n20506) );
  XOR U25228 ( .A(n22939), .B(n24933), .Z(n20505) );
  XNOR U25229 ( .A(n24934), .B(n19410), .Z(n17396) );
  XNOR U25230 ( .A(n24904), .B(n24935), .Z(n19410) );
  AND U25231 ( .A(n20516), .B(n20515), .Z(n24934) );
  XOR U25232 ( .A(n24936), .B(n24937), .Z(n20515) );
  XOR U25233 ( .A(n24938), .B(n24374), .Z(n20516) );
  XOR U25234 ( .A(n24939), .B(n24940), .Z(n21092) );
  XNOR U25235 ( .A(n18748), .B(n17478), .Z(n24940) );
  XOR U25236 ( .A(n24941), .B(n22699), .Z(n17478) );
  XNOR U25237 ( .A(n24942), .B(n24943), .Z(n22699) );
  ANDN U25238 ( .B(n24944), .A(n20450), .Z(n24941) );
  XOR U25239 ( .A(n24945), .B(n24946), .Z(n20450) );
  XOR U25240 ( .A(n24947), .B(n22693), .Z(n18748) );
  XOR U25241 ( .A(n24948), .B(n24949), .Z(n22693) );
  ANDN U25242 ( .B(n24950), .A(n22692), .Z(n24947) );
  XOR U25243 ( .A(n19033), .B(n24951), .Z(n24939) );
  XOR U25244 ( .A(n22667), .B(n17608), .Z(n24951) );
  XOR U25245 ( .A(n24953), .B(n23015), .Z(n22696) );
  NOR U25246 ( .A(n20457), .B(n20456), .Z(n24952) );
  XNOR U25247 ( .A(n24954), .B(n22500), .Z(n20456) );
  XNOR U25248 ( .A(n24955), .B(n22685), .Z(n22667) );
  XOR U25249 ( .A(n24956), .B(n24379), .Z(n22685) );
  ANDN U25250 ( .B(n22358), .A(n22359), .Z(n24955) );
  XOR U25251 ( .A(n21593), .B(n24957), .Z(n22358) );
  XNOR U25252 ( .A(n24958), .B(n22688), .Z(n19033) );
  XNOR U25253 ( .A(n24959), .B(n24960), .Z(n22688) );
  ANDN U25254 ( .B(n20460), .A(n20461), .Z(n24958) );
  XNOR U25255 ( .A(n24961), .B(n24761), .Z(n20460) );
  XOR U25256 ( .A(n24963), .B(n24964), .Z(n22692) );
  NOR U25257 ( .A(n24950), .B(n23400), .Z(n24962) );
  ANDN U25258 ( .B(n16583), .A(n18241), .Z(n24911) );
  XOR U25259 ( .A(n22547), .B(n17578), .Z(n18241) );
  XOR U25260 ( .A(n20383), .B(n21336), .Z(n17578) );
  XNOR U25261 ( .A(n24965), .B(n24966), .Z(n21336) );
  XNOR U25262 ( .A(n18892), .B(n15691), .Z(n24966) );
  XNOR U25263 ( .A(n24967), .B(n20437), .Z(n15691) );
  XOR U25264 ( .A(n24968), .B(n22988), .Z(n20437) );
  ANDN U25265 ( .B(n21194), .A(n22896), .Z(n24967) );
  XNOR U25266 ( .A(n24969), .B(n20423), .Z(n18892) );
  XOR U25267 ( .A(n24618), .B(n24970), .Z(n20423) );
  IV U25268 ( .A(n24971), .Z(n24618) );
  ANDN U25269 ( .B(n21197), .A(n24972), .Z(n24969) );
  XNOR U25270 ( .A(n19093), .B(n24973), .Z(n24965) );
  XOR U25271 ( .A(n17450), .B(n17669), .Z(n24973) );
  XNOR U25272 ( .A(n24974), .B(n20433), .Z(n17669) );
  XNOR U25273 ( .A(n24975), .B(n21599), .Z(n20433) );
  ANDN U25274 ( .B(n24976), .A(n22884), .Z(n24974) );
  XNOR U25275 ( .A(n24977), .B(n20427), .Z(n17450) );
  XNOR U25276 ( .A(n23991), .B(n24978), .Z(n20427) );
  NOR U25277 ( .A(n21200), .B(n22888), .Z(n24977) );
  XOR U25278 ( .A(n24979), .B(n20441), .Z(n19093) );
  XOR U25279 ( .A(n24980), .B(n23558), .Z(n20441) );
  ANDN U25280 ( .B(n22900), .A(n21190), .Z(n24979) );
  XNOR U25281 ( .A(n24981), .B(n24982), .Z(n20383) );
  XNOR U25282 ( .A(n18001), .B(n16116), .Z(n24982) );
  XOR U25283 ( .A(n24983), .B(n20949), .Z(n16116) );
  XOR U25284 ( .A(n24040), .B(n24984), .Z(n20949) );
  AND U25285 ( .A(n22544), .B(n22545), .Z(n24983) );
  XNOR U25286 ( .A(n24985), .B(n24986), .Z(n22544) );
  XNOR U25287 ( .A(n24987), .B(n20956), .Z(n18001) );
  XOR U25288 ( .A(n24988), .B(n24989), .Z(n20956) );
  ANDN U25289 ( .B(n22552), .A(n24990), .Z(n24987) );
  XOR U25290 ( .A(n23831), .B(n24991), .Z(n22552) );
  XOR U25291 ( .A(n18494), .B(n24992), .Z(n24981) );
  XOR U25292 ( .A(n22879), .B(n16073), .Z(n24992) );
  XNOR U25293 ( .A(n24993), .B(n20946), .Z(n16073) );
  XOR U25294 ( .A(n24994), .B(n24995), .Z(n20946) );
  ANDN U25295 ( .B(n24996), .A(n22549), .Z(n24993) );
  IV U25296 ( .A(n24731), .Z(n22549) );
  XNOR U25297 ( .A(n24997), .B(n24998), .Z(n24731) );
  XNOR U25298 ( .A(n24999), .B(n20960), .Z(n22879) );
  XOR U25299 ( .A(n23503), .B(n25000), .Z(n20960) );
  IV U25300 ( .A(n25001), .Z(n23503) );
  ANDN U25301 ( .B(n25002), .A(n24736), .Z(n24999) );
  XNOR U25302 ( .A(n25003), .B(n21205), .Z(n18494) );
  XOR U25303 ( .A(n25004), .B(n24908), .Z(n21205) );
  AND U25304 ( .A(n22541), .B(n22542), .Z(n25003) );
  XNOR U25305 ( .A(n25005), .B(n21586), .Z(n22541) );
  XOR U25306 ( .A(n25006), .B(n24736), .Z(n22547) );
  XOR U25307 ( .A(n25007), .B(n25008), .Z(n24736) );
  ANDN U25308 ( .B(n20958), .A(n25002), .Z(n25006) );
  XOR U25309 ( .A(n21900), .B(n21029), .Z(n16583) );
  XNOR U25310 ( .A(n25009), .B(n21167), .Z(n21029) );
  ANDN U25311 ( .B(n25010), .A(n25011), .Z(n25009) );
  IV U25312 ( .A(n17338), .Z(n21900) );
  XNOR U25313 ( .A(n25012), .B(n25013), .Z(n23341) );
  XNOR U25314 ( .A(n18402), .B(n16098), .Z(n25013) );
  XOR U25315 ( .A(n25014), .B(n21170), .Z(n16098) );
  XOR U25316 ( .A(n25015), .B(n22536), .Z(n21170) );
  NOR U25317 ( .A(n21031), .B(n21032), .Z(n25014) );
  XOR U25318 ( .A(n25016), .B(n25017), .Z(n21031) );
  XOR U25319 ( .A(n25018), .B(n21174), .Z(n18402) );
  NOR U25320 ( .A(n21175), .B(n21027), .Z(n25018) );
  XOR U25321 ( .A(n25019), .B(n24162), .Z(n21175) );
  XOR U25322 ( .A(n20820), .B(n25020), .Z(n25012) );
  XOR U25323 ( .A(n21150), .B(n17004), .Z(n25020) );
  XNOR U25324 ( .A(n25021), .B(n21178), .Z(n17004) );
  XNOR U25325 ( .A(n25022), .B(n25023), .Z(n21178) );
  ANDN U25326 ( .B(n21035), .A(n25024), .Z(n25021) );
  XNOR U25327 ( .A(n25025), .B(n25026), .Z(n21035) );
  XOR U25328 ( .A(n25027), .B(n21166), .Z(n21150) );
  XNOR U25329 ( .A(n25028), .B(n21368), .Z(n21166) );
  NOR U25330 ( .A(n25010), .B(n21167), .Z(n25027) );
  XNOR U25331 ( .A(n25029), .B(n22982), .Z(n21167) );
  XNOR U25332 ( .A(n25030), .B(n21181), .Z(n20820) );
  XNOR U25333 ( .A(n25031), .B(n23432), .Z(n21181) );
  IV U25334 ( .A(n25032), .Z(n23432) );
  ANDN U25335 ( .B(n21182), .A(n21902), .Z(n25030) );
  XOR U25336 ( .A(n25033), .B(n23983), .Z(n21182) );
  XOR U25337 ( .A(n25035), .B(n25036), .Z(n14475) );
  XNOR U25338 ( .A(n12199), .B(n10191), .Z(n25036) );
  XOR U25339 ( .A(n25037), .B(n14628), .Z(n10191) );
  XOR U25340 ( .A(n22374), .B(n16878), .Z(n14628) );
  XOR U25341 ( .A(n23239), .B(n19465), .Z(n16878) );
  XNOR U25342 ( .A(n25038), .B(n25039), .Z(n19465) );
  XOR U25343 ( .A(n17792), .B(n17036), .Z(n25039) );
  XNOR U25344 ( .A(n25040), .B(n24534), .Z(n17036) );
  ANDN U25345 ( .B(n24533), .A(n22867), .Z(n25040) );
  XOR U25346 ( .A(n25041), .B(n24545), .Z(n17792) );
  NOR U25347 ( .A(n24546), .B(n22367), .Z(n25041) );
  XOR U25348 ( .A(n25042), .B(n25043), .Z(n22367) );
  XOR U25349 ( .A(n25044), .B(n25045), .Z(n24546) );
  XOR U25350 ( .A(n15886), .B(n25046), .Z(n25038) );
  XOR U25351 ( .A(n16467), .B(n24510), .Z(n25046) );
  XNOR U25352 ( .A(n25047), .B(n24542), .Z(n24510) );
  NOR U25353 ( .A(n24543), .B(n22382), .Z(n25047) );
  XOR U25354 ( .A(n23592), .B(n25048), .Z(n22382) );
  XNOR U25355 ( .A(n25049), .B(n25050), .Z(n24543) );
  XNOR U25356 ( .A(n25051), .B(n24536), .Z(n16467) );
  ANDN U25357 ( .B(n22370), .A(n22371), .Z(n25051) );
  XOR U25358 ( .A(n24772), .B(n25052), .Z(n22371) );
  IV U25359 ( .A(n25053), .Z(n24772) );
  XOR U25360 ( .A(n25054), .B(n24908), .Z(n22370) );
  XNOR U25361 ( .A(n25055), .B(n24539), .Z(n15886) );
  NOR U25362 ( .A(n24540), .B(n22377), .Z(n25055) );
  XOR U25363 ( .A(n23969), .B(n25056), .Z(n22377) );
  IV U25364 ( .A(n25057), .Z(n23969) );
  XOR U25365 ( .A(n25058), .B(n23482), .Z(n24540) );
  XNOR U25366 ( .A(n25059), .B(n25060), .Z(n23239) );
  XNOR U25367 ( .A(n16838), .B(n19710), .Z(n25060) );
  XOR U25368 ( .A(n25061), .B(n20568), .Z(n19710) );
  XOR U25369 ( .A(n25062), .B(n21725), .Z(n20568) );
  AND U25370 ( .A(n20743), .B(n20741), .Z(n25061) );
  XOR U25371 ( .A(n25063), .B(n22892), .Z(n20741) );
  XNOR U25372 ( .A(n25064), .B(n24825), .Z(n20743) );
  XOR U25373 ( .A(n25065), .B(n20558), .Z(n16838) );
  XOR U25374 ( .A(n21593), .B(n25066), .Z(n20558) );
  NOR U25375 ( .A(n20746), .B(n20745), .Z(n25065) );
  XNOR U25376 ( .A(n25057), .B(n25067), .Z(n20745) );
  XOR U25377 ( .A(n25068), .B(n25069), .Z(n20746) );
  XNOR U25378 ( .A(n17442), .B(n25070), .Z(n25059) );
  XOR U25379 ( .A(n16067), .B(n18224), .Z(n25070) );
  XNOR U25380 ( .A(n25071), .B(n20564), .Z(n18224) );
  XOR U25381 ( .A(n25072), .B(n22396), .Z(n20564) );
  ANDN U25382 ( .B(n21972), .A(n21969), .Z(n25071) );
  XOR U25383 ( .A(n25073), .B(n21216), .Z(n21969) );
  XNOR U25384 ( .A(n25074), .B(n25050), .Z(n21972) );
  XNOR U25385 ( .A(n25075), .B(n20554), .Z(n16067) );
  XOR U25386 ( .A(n23745), .B(n25076), .Z(n20554) );
  IV U25387 ( .A(n23690), .Z(n23745) );
  AND U25388 ( .A(n23258), .B(n23257), .Z(n25075) );
  XNOR U25389 ( .A(n25077), .B(n24399), .Z(n23257) );
  XOR U25390 ( .A(n25078), .B(n25079), .Z(n23258) );
  XOR U25391 ( .A(n25080), .B(n24522), .Z(n17442) );
  IV U25392 ( .A(n24403), .Z(n24522) );
  XOR U25393 ( .A(n25081), .B(n24835), .Z(n24403) );
  NOR U25394 ( .A(n20736), .B(n20735), .Z(n25080) );
  XOR U25395 ( .A(n25082), .B(n22021), .Z(n20735) );
  IV U25396 ( .A(n25083), .Z(n22021) );
  XOR U25397 ( .A(n25084), .B(n24695), .Z(n20736) );
  IV U25398 ( .A(n25085), .Z(n24695) );
  XNOR U25399 ( .A(n25086), .B(n24533), .Z(n22374) );
  XOR U25400 ( .A(n25087), .B(n24499), .Z(n24533) );
  ANDN U25401 ( .B(n22867), .A(n22868), .Z(n25086) );
  XOR U25402 ( .A(n25088), .B(n24237), .Z(n22867) );
  IV U25403 ( .A(n24661), .Z(n24237) );
  ANDN U25404 ( .B(n16599), .A(n19647), .Z(n25037) );
  XOR U25405 ( .A(n17474), .B(n20794), .Z(n19647) );
  XNOR U25406 ( .A(n25089), .B(n25090), .Z(n20794) );
  NOR U25407 ( .A(n23227), .B(n23228), .Z(n25089) );
  XOR U25408 ( .A(n23664), .B(n23155), .Z(n17474) );
  XOR U25409 ( .A(n25091), .B(n25092), .Z(n23155) );
  XOR U25410 ( .A(n19540), .B(n18185), .Z(n25092) );
  XOR U25411 ( .A(n25093), .B(n22094), .Z(n18185) );
  XNOR U25412 ( .A(n25094), .B(n23573), .Z(n22094) );
  ANDN U25413 ( .B(n19576), .A(n19692), .Z(n25093) );
  IV U25414 ( .A(n22093), .Z(n19692) );
  XOR U25415 ( .A(n25095), .B(n23150), .Z(n22093) );
  XOR U25416 ( .A(n25097), .B(n22084), .Z(n19540) );
  XNOR U25417 ( .A(n25098), .B(n25099), .Z(n22084) );
  XOR U25418 ( .A(n25100), .B(n22511), .Z(n19571) );
  XOR U25419 ( .A(n25101), .B(n24399), .Z(n22083) );
  XNOR U25420 ( .A(n19248), .B(n25104), .Z(n25091) );
  XOR U25421 ( .A(n20148), .B(n21732), .Z(n25104) );
  XOR U25422 ( .A(n22096), .B(n25105), .Z(n21732) );
  XOR U25423 ( .A(n25106), .B(n4407), .Z(n25105) );
  ANDN U25424 ( .B(n19687), .A(n19567), .Z(n25106) );
  XNOR U25425 ( .A(n25107), .B(n23914), .Z(n19567) );
  XOR U25426 ( .A(n25108), .B(n25109), .Z(n19687) );
  XOR U25427 ( .A(n25110), .B(n25111), .Z(n22096) );
  XOR U25428 ( .A(n25112), .B(n22090), .Z(n20148) );
  XNOR U25429 ( .A(n25113), .B(n25114), .Z(n22090) );
  AND U25430 ( .A(n20069), .B(n19580), .Z(n25112) );
  XOR U25431 ( .A(n23690), .B(n25115), .Z(n19580) );
  XNOR U25432 ( .A(n25118), .B(n23072), .Z(n20069) );
  XNOR U25433 ( .A(n25119), .B(n22087), .Z(n19248) );
  XNOR U25434 ( .A(n25120), .B(n24499), .Z(n22087) );
  ANDN U25435 ( .B(n20029), .A(n19584), .Z(n25119) );
  XOR U25436 ( .A(n24819), .B(n25121), .Z(n19584) );
  IV U25437 ( .A(n22641), .Z(n24819) );
  XOR U25438 ( .A(n25122), .B(n23878), .Z(n20029) );
  XOR U25439 ( .A(n25123), .B(n25124), .Z(n23664) );
  XOR U25440 ( .A(n16888), .B(n19767), .Z(n25124) );
  XNOR U25441 ( .A(n25125), .B(n25126), .Z(n19767) );
  NOR U25442 ( .A(n23232), .B(n20805), .Z(n25125) );
  XOR U25443 ( .A(n25127), .B(n24860), .Z(n23232) );
  IV U25444 ( .A(n23033), .Z(n24860) );
  XNOR U25445 ( .A(n25128), .B(n25129), .Z(n16888) );
  ANDN U25446 ( .B(n20810), .A(n20809), .Z(n25128) );
  XNOR U25447 ( .A(n22217), .B(n25130), .Z(n20810) );
  XNOR U25448 ( .A(n25131), .B(n25132), .Z(n22217) );
  XOR U25449 ( .A(n22078), .B(n25133), .Z(n25123) );
  XNOR U25450 ( .A(n20839), .B(n19386), .Z(n25133) );
  XNOR U25451 ( .A(n25134), .B(n25135), .Z(n19386) );
  NOR U25452 ( .A(n23224), .B(n20801), .Z(n25134) );
  XOR U25453 ( .A(n25136), .B(n24554), .Z(n23224) );
  XOR U25454 ( .A(n25137), .B(n25138), .Z(n20839) );
  NOR U25455 ( .A(n23237), .B(n20796), .Z(n25137) );
  XOR U25456 ( .A(n24632), .B(n25139), .Z(n23237) );
  XNOR U25457 ( .A(n25140), .B(n25141), .Z(n22078) );
  ANDN U25458 ( .B(n23227), .A(n25090), .Z(n25140) );
  IV U25459 ( .A(n25142), .Z(n25090) );
  XOR U25460 ( .A(n25143), .B(n25144), .Z(n23227) );
  XNOR U25461 ( .A(n24642), .B(n17297), .Z(n16599) );
  XNOR U25462 ( .A(n19724), .B(n19192), .Z(n17297) );
  XOR U25463 ( .A(n25145), .B(n25146), .Z(n19192) );
  XOR U25464 ( .A(n17645), .B(n20081), .Z(n25146) );
  XOR U25465 ( .A(n25147), .B(n23901), .Z(n20081) );
  XNOR U25466 ( .A(n25148), .B(n21829), .Z(n23901) );
  ANDN U25467 ( .B(n21268), .A(n24640), .Z(n25147) );
  IV U25468 ( .A(n24147), .Z(n24640) );
  XOR U25469 ( .A(n25149), .B(n25150), .Z(n24147) );
  XNOR U25470 ( .A(n25151), .B(n25152), .Z(n21268) );
  XNOR U25471 ( .A(n25153), .B(n23888), .Z(n17645) );
  XOR U25472 ( .A(n25154), .B(n24798), .Z(n23888) );
  NOR U25473 ( .A(n24647), .B(n24142), .Z(n25153) );
  XOR U25474 ( .A(n23737), .B(n25155), .Z(n24142) );
  XOR U25475 ( .A(n25156), .B(n24281), .Z(n24647) );
  XOR U25476 ( .A(n17850), .B(n25157), .Z(n25145) );
  XNOR U25477 ( .A(n15701), .B(n20702), .Z(n25157) );
  XNOR U25478 ( .A(n25158), .B(n23891), .Z(n20702) );
  XNOR U25479 ( .A(n25159), .B(n25111), .Z(n23891) );
  AND U25480 ( .A(n21261), .B(n24151), .Z(n25158) );
  XNOR U25481 ( .A(n25160), .B(n23895), .Z(n15701) );
  XOR U25482 ( .A(n24233), .B(n25161), .Z(n23895) );
  XOR U25483 ( .A(n25162), .B(n25163), .Z(n21526) );
  XOR U25484 ( .A(n25164), .B(n25165), .Z(n24140) );
  XNOR U25485 ( .A(n25166), .B(n23899), .Z(n17850) );
  XNOR U25486 ( .A(n25167), .B(n23914), .Z(n23899) );
  ANDN U25487 ( .B(n24096), .A(n24155), .Z(n25166) );
  XNOR U25488 ( .A(n25169), .B(n25170), .Z(n24096) );
  XOR U25489 ( .A(n25171), .B(n25172), .Z(n19724) );
  XOR U25490 ( .A(n17139), .B(n17205), .Z(n25172) );
  XNOR U25491 ( .A(n25173), .B(n24751), .Z(n17205) );
  IV U25492 ( .A(n24055), .Z(n24751) );
  XOR U25493 ( .A(n25174), .B(n25175), .Z(n24055) );
  NOR U25494 ( .A(n24054), .B(n23474), .Z(n25173) );
  XOR U25495 ( .A(n25176), .B(n25177), .Z(n23474) );
  XNOR U25496 ( .A(n25178), .B(n22396), .Z(n24054) );
  XOR U25497 ( .A(n25179), .B(n24764), .Z(n17139) );
  XOR U25498 ( .A(n25180), .B(n23839), .Z(n24764) );
  ANDN U25499 ( .B(n22065), .A(n24653), .Z(n25179) );
  XOR U25500 ( .A(n25181), .B(n25182), .Z(n24653) );
  XOR U25501 ( .A(n25183), .B(n25184), .Z(n22065) );
  XNOR U25502 ( .A(n18869), .B(n25185), .Z(n25171) );
  XOR U25503 ( .A(n24042), .B(n18189), .Z(n25185) );
  XNOR U25504 ( .A(n25186), .B(n24049), .Z(n18189) );
  XNOR U25505 ( .A(n25187), .B(n24154), .Z(n24049) );
  ANDN U25506 ( .B(n24050), .A(n22075), .Z(n25186) );
  XOR U25507 ( .A(n25188), .B(n25189), .Z(n22075) );
  XNOR U25508 ( .A(n23742), .B(n25190), .Z(n24050) );
  XNOR U25509 ( .A(n24702), .B(n25192), .Z(n24058) );
  ANDN U25510 ( .B(n24059), .A(n22061), .Z(n25191) );
  XOR U25511 ( .A(n25193), .B(n23573), .Z(n22061) );
  XNOR U25512 ( .A(n25194), .B(n23571), .Z(n24059) );
  IV U25513 ( .A(n22342), .Z(n23571) );
  XNOR U25514 ( .A(n25195), .B(n24046), .Z(n18869) );
  XNOR U25515 ( .A(n25196), .B(n23513), .Z(n24046) );
  AND U25516 ( .A(n24047), .B(n22071), .Z(n25195) );
  XNOR U25517 ( .A(n22223), .B(n25197), .Z(n22071) );
  XOR U25518 ( .A(n25200), .B(n25201), .Z(n24047) );
  XNOR U25519 ( .A(n25202), .B(n24151), .Z(n24642) );
  XOR U25520 ( .A(n25203), .B(n25204), .Z(n24151) );
  NOR U25521 ( .A(n21261), .B(n21262), .Z(n25202) );
  XOR U25522 ( .A(n25207), .B(n23244), .Z(n21261) );
  IV U25523 ( .A(n24943), .Z(n23244) );
  XOR U25524 ( .A(n25208), .B(n14623), .Z(n12199) );
  XNOR U25525 ( .A(n19779), .B(n17870), .Z(n14623) );
  IV U25526 ( .A(n20696), .Z(n17870) );
  XOR U25527 ( .A(n21399), .B(n22905), .Z(n20696) );
  XNOR U25528 ( .A(n25209), .B(n25210), .Z(n22905) );
  XNOR U25529 ( .A(n17008), .B(n20276), .Z(n25210) );
  XOR U25530 ( .A(n25211), .B(n19534), .Z(n20276) );
  XOR U25531 ( .A(n25212), .B(n22227), .Z(n19534) );
  ANDN U25532 ( .B(n20285), .A(n21723), .Z(n25211) );
  XNOR U25533 ( .A(n25213), .B(n19528), .Z(n17008) );
  ANDN U25534 ( .B(n19785), .A(n19786), .Z(n25213) );
  XOR U25535 ( .A(n25216), .B(n22025), .Z(n19785) );
  XOR U25536 ( .A(n14988), .B(n25217), .Z(n25209) );
  XOR U25537 ( .A(n17491), .B(n18642), .Z(n25217) );
  XOR U25538 ( .A(n25218), .B(n20288), .Z(n18642) );
  XOR U25539 ( .A(n25219), .B(n25220), .Z(n20288) );
  NOR U25540 ( .A(n20289), .B(n21339), .Z(n25218) );
  XOR U25541 ( .A(n25221), .B(n25222), .Z(n21339) );
  XOR U25542 ( .A(n25223), .B(n25224), .Z(n20289) );
  XOR U25543 ( .A(n25225), .B(n19538), .Z(n17491) );
  XOR U25544 ( .A(n25226), .B(n25227), .Z(n19538) );
  ANDN U25545 ( .B(n20281), .A(n21708), .Z(n25225) );
  IV U25546 ( .A(n24317), .Z(n21708) );
  XOR U25547 ( .A(n25228), .B(n24270), .Z(n24317) );
  IV U25548 ( .A(n21372), .Z(n24270) );
  XOR U25549 ( .A(n25229), .B(n25230), .Z(n20281) );
  XNOR U25550 ( .A(n25231), .B(n20292), .Z(n14988) );
  XOR U25551 ( .A(n25232), .B(n24849), .Z(n20292) );
  ANDN U25552 ( .B(n20293), .A(n20698), .Z(n25231) );
  XOR U25553 ( .A(n24936), .B(n25233), .Z(n20698) );
  XNOR U25554 ( .A(n25234), .B(n25206), .Z(n20293) );
  XOR U25555 ( .A(n25235), .B(n25236), .Z(n21399) );
  XOR U25556 ( .A(n18827), .B(n19761), .Z(n25236) );
  XNOR U25557 ( .A(n25237), .B(n25238), .Z(n19761) );
  ANDN U25558 ( .B(n20327), .A(n20325), .Z(n25237) );
  XOR U25559 ( .A(n25239), .B(n25240), .Z(n20327) );
  XNOR U25560 ( .A(n25241), .B(n22018), .Z(n18827) );
  NOR U25561 ( .A(n21416), .B(n21417), .Z(n25241) );
  XOR U25562 ( .A(n25242), .B(n24180), .Z(n21417) );
  XOR U25563 ( .A(n21731), .B(n25243), .Z(n25235) );
  XOR U25564 ( .A(n16408), .B(n25244), .Z(n25243) );
  XNOR U25565 ( .A(n25245), .B(n22022), .Z(n16408) );
  NOR U25566 ( .A(n20335), .B(n20336), .Z(n25245) );
  XNOR U25567 ( .A(n25246), .B(n25247), .Z(n20336) );
  XNOR U25568 ( .A(n25248), .B(n25249), .Z(n21731) );
  ANDN U25569 ( .B(n21701), .A(n25250), .Z(n25248) );
  XOR U25570 ( .A(n25251), .B(n25252), .Z(n21701) );
  XNOR U25571 ( .A(n25253), .B(n20285), .Z(n19779) );
  XNOR U25572 ( .A(n25254), .B(n25255), .Z(n20285) );
  AND U25573 ( .A(n19533), .B(n21723), .Z(n25253) );
  XOR U25574 ( .A(n24025), .B(n25256), .Z(n21723) );
  XNOR U25575 ( .A(n25257), .B(n25045), .Z(n19533) );
  XOR U25576 ( .A(n21439), .B(n17874), .Z(n15178) );
  IV U25577 ( .A(n20130), .Z(n17874) );
  XNOR U25578 ( .A(n25258), .B(n25259), .Z(n24664) );
  XOR U25579 ( .A(n20011), .B(n18721), .Z(n25259) );
  XOR U25580 ( .A(n25260), .B(n20061), .Z(n18721) );
  XOR U25581 ( .A(n25261), .B(n23812), .Z(n20061) );
  NOR U25582 ( .A(n21446), .B(n21445), .Z(n25260) );
  XNOR U25583 ( .A(n25264), .B(n24989), .Z(n21445) );
  XOR U25584 ( .A(n25265), .B(n22231), .Z(n21446) );
  XNOR U25585 ( .A(n25266), .B(n20066), .Z(n20011) );
  XOR U25586 ( .A(n22654), .B(n25267), .Z(n20066) );
  IV U25587 ( .A(n25268), .Z(n22654) );
  ANDN U25588 ( .B(n21441), .A(n21442), .Z(n25266) );
  XNOR U25589 ( .A(n25269), .B(n22899), .Z(n21442) );
  XNOR U25590 ( .A(n25270), .B(n24745), .Z(n21441) );
  XOR U25591 ( .A(n19749), .B(n25271), .Z(n25258) );
  XOR U25592 ( .A(n18044), .B(n17400), .Z(n25271) );
  XNOR U25593 ( .A(n25272), .B(n20056), .Z(n17400) );
  XOR U25594 ( .A(n23695), .B(n25273), .Z(n20056) );
  ANDN U25595 ( .B(n23780), .A(n24024), .Z(n25272) );
  XOR U25596 ( .A(n25274), .B(n23771), .Z(n18044) );
  XOR U25597 ( .A(n25275), .B(n25276), .Z(n23771) );
  NOR U25598 ( .A(n23772), .B(n21453), .Z(n25274) );
  XNOR U25599 ( .A(n25277), .B(n25278), .Z(n21453) );
  XOR U25600 ( .A(n25053), .B(n25279), .Z(n23772) );
  XNOR U25601 ( .A(n25280), .B(n22908), .Z(n19749) );
  XOR U25602 ( .A(n25281), .B(n24916), .Z(n22908) );
  ANDN U25603 ( .B(n21448), .A(n21449), .Z(n25280) );
  XNOR U25604 ( .A(n25282), .B(n25283), .Z(n21449) );
  XOR U25605 ( .A(n25284), .B(n23013), .Z(n21448) );
  XNOR U25606 ( .A(n25286), .B(n23780), .Z(n21439) );
  XOR U25607 ( .A(n25287), .B(n23568), .Z(n23780) );
  AND U25608 ( .A(n20054), .B(n24024), .Z(n25286) );
  XOR U25609 ( .A(n24930), .B(n25288), .Z(n24024) );
  XNOR U25610 ( .A(n25289), .B(n25290), .Z(n20054) );
  XOR U25611 ( .A(n18103), .B(n24678), .Z(n14622) );
  XNOR U25612 ( .A(n25291), .B(n21436), .Z(n24678) );
  NOR U25613 ( .A(n24126), .B(n24125), .Z(n25291) );
  IV U25614 ( .A(n18380), .Z(n18103) );
  XNOR U25615 ( .A(n25292), .B(n24017), .Z(n18380) );
  XNOR U25616 ( .A(n25293), .B(n25294), .Z(n24017) );
  XNOR U25617 ( .A(n16022), .B(n18802), .Z(n25294) );
  XOR U25618 ( .A(n25295), .B(n21435), .Z(n18802) );
  AND U25619 ( .A(n21436), .B(n24125), .Z(n25295) );
  XOR U25620 ( .A(n21593), .B(n25296), .Z(n24125) );
  XOR U25621 ( .A(n25297), .B(n23731), .Z(n21436) );
  XNOR U25622 ( .A(n25298), .B(n25299), .Z(n16022) );
  ANDN U25623 ( .B(n24672), .A(n24132), .Z(n25298) );
  IV U25624 ( .A(n24673), .Z(n24132) );
  XOR U25625 ( .A(n25300), .B(n25301), .Z(n24673) );
  XOR U25626 ( .A(n19178), .B(n25302), .Z(n25293) );
  XNOR U25627 ( .A(n18610), .B(n17175), .Z(n25302) );
  XNOR U25628 ( .A(n25303), .B(n21425), .Z(n17175) );
  ANDN U25629 ( .B(n21424), .A(n24129), .Z(n25303) );
  XOR U25630 ( .A(n25304), .B(n25305), .Z(n24129) );
  XOR U25631 ( .A(n25306), .B(n25307), .Z(n21424) );
  XNOR U25632 ( .A(n25308), .B(n25309), .Z(n18610) );
  ANDN U25633 ( .B(n24121), .A(n22277), .Z(n25308) );
  XOR U25634 ( .A(n25310), .B(n24035), .Z(n22277) );
  XOR U25635 ( .A(n24337), .B(n25311), .Z(n24121) );
  XOR U25636 ( .A(n25312), .B(n21428), .Z(n19178) );
  ANDN U25637 ( .B(n21429), .A(n24675), .Z(n25312) );
  XOR U25638 ( .A(n25313), .B(n23852), .Z(n24675) );
  XNOR U25639 ( .A(n25314), .B(n22958), .Z(n21429) );
  XOR U25640 ( .A(n11410), .B(n25315), .Z(n25035) );
  XNOR U25641 ( .A(n12848), .B(n9816), .Z(n25315) );
  XOR U25642 ( .A(n25316), .B(n14631), .Z(n9816) );
  XOR U25643 ( .A(n17619), .B(n24862), .Z(n14631) );
  XNOR U25644 ( .A(n25317), .B(n25318), .Z(n24862) );
  NOR U25645 ( .A(n25319), .B(n23273), .Z(n25317) );
  XNOR U25646 ( .A(n24063), .B(n25320), .Z(n23273) );
  XOR U25647 ( .A(n20548), .B(n23179), .Z(n17619) );
  XNOR U25648 ( .A(n25321), .B(n25322), .Z(n23179) );
  XNOR U25649 ( .A(n18236), .B(n18964), .Z(n25322) );
  XNOR U25650 ( .A(n25323), .B(n24088), .Z(n18964) );
  IV U25651 ( .A(n25324), .Z(n24088) );
  ANDN U25652 ( .B(n23277), .A(n24855), .Z(n25323) );
  XNOR U25653 ( .A(n22313), .B(n25325), .Z(n23277) );
  XNOR U25654 ( .A(n25326), .B(n24093), .Z(n18236) );
  ANDN U25655 ( .B(n24865), .A(n23285), .Z(n25326) );
  XOR U25656 ( .A(n25327), .B(n24844), .Z(n23285) );
  XOR U25657 ( .A(n18504), .B(n25328), .Z(n25321) );
  XOR U25658 ( .A(n22855), .B(n19790), .Z(n25328) );
  XNOR U25659 ( .A(n25329), .B(n24084), .Z(n19790) );
  ANDN U25660 ( .B(n25318), .A(n23269), .Z(n25329) );
  IV U25661 ( .A(n25319), .Z(n23269) );
  XOR U25662 ( .A(n25330), .B(n23721), .Z(n25319) );
  IV U25663 ( .A(n22526), .Z(n23721) );
  XNOR U25664 ( .A(n25331), .B(n24090), .Z(n22855) );
  ANDN U25665 ( .B(n24868), .A(n23281), .Z(n25331) );
  XOR U25666 ( .A(n23592), .B(n25332), .Z(n23281) );
  XNOR U25667 ( .A(n25333), .B(n24082), .Z(n18504) );
  ANDN U25668 ( .B(n23266), .A(n24859), .Z(n25333) );
  XNOR U25669 ( .A(n25334), .B(n23253), .Z(n23266) );
  XOR U25670 ( .A(n25335), .B(n25336), .Z(n20548) );
  XOR U25671 ( .A(n20665), .B(n19327), .Z(n25336) );
  XNOR U25672 ( .A(n25337), .B(n22381), .Z(n19327) );
  XNOR U25673 ( .A(n25338), .B(n25227), .Z(n22381) );
  ANDN U25674 ( .B(n24542), .A(n22862), .Z(n25337) );
  XOR U25675 ( .A(n24241), .B(n25339), .Z(n22862) );
  XOR U25676 ( .A(n25340), .B(n23050), .Z(n24542) );
  XOR U25677 ( .A(n22868), .B(n25341), .Z(n20665) );
  XOR U25678 ( .A(n25342), .B(n4407), .Z(n25341) );
  ANDN U25679 ( .B(n24534), .A(n24532), .Z(n25342) );
  IV U25680 ( .A(n22869), .Z(n24532) );
  XOR U25681 ( .A(n22635), .B(n25343), .Z(n22869) );
  XOR U25682 ( .A(n25344), .B(n23040), .Z(n24534) );
  XOR U25683 ( .A(n25345), .B(n22834), .Z(n22868) );
  XOR U25684 ( .A(n18630), .B(n25346), .Z(n25335) );
  XOR U25685 ( .A(n17612), .B(n18305), .Z(n25346) );
  XNOR U25686 ( .A(n25347), .B(n22368), .Z(n18305) );
  XOR U25687 ( .A(n25348), .B(n24986), .Z(n22368) );
  NOR U25688 ( .A(n24545), .B(n22860), .Z(n25347) );
  XNOR U25689 ( .A(n25349), .B(n25350), .Z(n22860) );
  XOR U25690 ( .A(n25351), .B(n25352), .Z(n24545) );
  XNOR U25691 ( .A(n25353), .B(n22378), .Z(n17612) );
  IV U25692 ( .A(n22871), .Z(n22378) );
  XOR U25693 ( .A(n25354), .B(n24835), .Z(n22871) );
  AND U25694 ( .A(n24539), .B(n22872), .Z(n25353) );
  XNOR U25695 ( .A(n25355), .B(n25356), .Z(n22872) );
  XOR U25696 ( .A(n25357), .B(n21606), .Z(n24539) );
  XOR U25697 ( .A(n25358), .B(n22372), .Z(n18630) );
  XOR U25698 ( .A(n24442), .B(n25359), .Z(n22372) );
  ANDN U25699 ( .B(n24536), .A(n22865), .Z(n25358) );
  XOR U25700 ( .A(n25360), .B(n25361), .Z(n22865) );
  XNOR U25701 ( .A(n25362), .B(n25363), .Z(n24536) );
  ANDN U25702 ( .B(n14632), .A(n16594), .Z(n25316) );
  XNOR U25703 ( .A(n25364), .B(n16614), .Z(n12848) );
  IV U25704 ( .A(n15471), .Z(n16614) );
  XNOR U25705 ( .A(n25365), .B(n18419), .Z(n15471) );
  XNOR U25706 ( .A(n18637), .B(n19241), .Z(n18419) );
  XNOR U25707 ( .A(n25366), .B(n25367), .Z(n19241) );
  XNOR U25708 ( .A(n17969), .B(n18362), .Z(n25367) );
  XNOR U25709 ( .A(n25368), .B(n21885), .Z(n18362) );
  ANDN U25710 ( .B(n21494), .A(n21493), .Z(n25368) );
  XNOR U25711 ( .A(n23145), .B(n25369), .Z(n21494) );
  XNOR U25712 ( .A(n25370), .B(n21877), .Z(n17969) );
  IV U25713 ( .A(n25371), .Z(n21877) );
  ANDN U25714 ( .B(n21484), .A(n24347), .Z(n25370) );
  IV U25715 ( .A(n21485), .Z(n24347) );
  XOR U25716 ( .A(n25372), .B(n25373), .Z(n21485) );
  XNOR U25717 ( .A(n18764), .B(n25374), .Z(n25366) );
  XOR U25718 ( .A(n20389), .B(n22903), .Z(n25374) );
  XNOR U25719 ( .A(n25375), .B(n21889), .Z(n22903) );
  ANDN U25720 ( .B(n21480), .A(n24340), .Z(n25375) );
  IV U25721 ( .A(n21482), .Z(n24340) );
  XOR U25722 ( .A(n25376), .B(n24857), .Z(n21482) );
  XOR U25723 ( .A(n25377), .B(n21881), .Z(n20389) );
  AND U25724 ( .A(n21491), .B(n21489), .Z(n25377) );
  XNOR U25725 ( .A(n23066), .B(n25378), .Z(n21491) );
  XNOR U25726 ( .A(n25379), .B(n21891), .Z(n18764) );
  ANDN U25727 ( .B(n21498), .A(n25380), .Z(n25379) );
  XOR U25728 ( .A(n25381), .B(n25382), .Z(n21498) );
  XOR U25729 ( .A(n25383), .B(n25384), .Z(n18637) );
  XNOR U25730 ( .A(n17634), .B(n21114), .Z(n25384) );
  XOR U25731 ( .A(n25385), .B(n21863), .Z(n21114) );
  XOR U25732 ( .A(n25387), .B(n24353), .Z(n17634) );
  ANDN U25733 ( .B(n25388), .A(n25389), .Z(n25387) );
  XOR U25734 ( .A(n19509), .B(n25390), .Z(n25383) );
  XOR U25735 ( .A(n15961), .B(n25391), .Z(n25390) );
  XNOR U25736 ( .A(n25392), .B(n22876), .Z(n15961) );
  XOR U25737 ( .A(n25394), .B(n21873), .Z(n19509) );
  ANDN U25738 ( .B(n25395), .A(n25396), .Z(n25394) );
  ANDN U25739 ( .B(n15167), .A(n15169), .Z(n25364) );
  XOR U25740 ( .A(n16374), .B(n25397), .Z(n15169) );
  IV U25741 ( .A(n17063), .Z(n16374) );
  XOR U25742 ( .A(n24212), .B(n22282), .Z(n17063) );
  XNOR U25743 ( .A(n25398), .B(n25399), .Z(n22282) );
  XOR U25744 ( .A(n19198), .B(n18599), .Z(n25399) );
  XNOR U25745 ( .A(n25400), .B(n23646), .Z(n18599) );
  XOR U25746 ( .A(n25401), .B(n23568), .Z(n23646) );
  IV U25747 ( .A(n24839), .Z(n23568) );
  XOR U25748 ( .A(n25402), .B(n25403), .Z(n24839) );
  ANDN U25749 ( .B(n22708), .A(n23552), .Z(n25400) );
  IV U25750 ( .A(n22709), .Z(n23552) );
  XOR U25751 ( .A(n25404), .B(n25405), .Z(n22709) );
  XNOR U25752 ( .A(n25406), .B(n21221), .Z(n22708) );
  XNOR U25753 ( .A(n25407), .B(n23644), .Z(n19198) );
  XNOR U25754 ( .A(n25408), .B(n24702), .Z(n23644) );
  XOR U25755 ( .A(n25409), .B(n25410), .Z(n22712) );
  XNOR U25756 ( .A(n25411), .B(n23573), .Z(n22714) );
  XOR U25757 ( .A(n18071), .B(n25412), .Z(n25398) );
  XNOR U25758 ( .A(n19760), .B(n23633), .Z(n25412) );
  XNOR U25759 ( .A(n25413), .B(n23641), .Z(n23633) );
  XOR U25760 ( .A(n25414), .B(n25415), .Z(n23641) );
  ANDN U25761 ( .B(n22723), .A(n23642), .Z(n25413) );
  XOR U25762 ( .A(n25416), .B(n23602), .Z(n23642) );
  XNOR U25763 ( .A(n25417), .B(n22008), .Z(n22723) );
  XNOR U25764 ( .A(n25418), .B(n23638), .Z(n19760) );
  XNOR U25765 ( .A(n25419), .B(n21606), .Z(n23638) );
  AND U25766 ( .A(n22718), .B(n22717), .Z(n25418) );
  XOR U25767 ( .A(n25420), .B(n22391), .Z(n22717) );
  XOR U25768 ( .A(n24458), .B(n25421), .Z(n22718) );
  XNOR U25769 ( .A(n25422), .B(n24587), .Z(n18071) );
  XOR U25770 ( .A(n25423), .B(n25424), .Z(n24587) );
  AND U25771 ( .A(n22726), .B(n22725), .Z(n25422) );
  XOR U25772 ( .A(n24432), .B(n25425), .Z(n22725) );
  XOR U25773 ( .A(n25426), .B(n25427), .Z(n22726) );
  XNOR U25774 ( .A(n25428), .B(n25429), .Z(n24212) );
  XOR U25775 ( .A(n19428), .B(n19438), .Z(n25429) );
  XNOR U25776 ( .A(n25430), .B(n20678), .Z(n19438) );
  XOR U25777 ( .A(n25431), .B(n25307), .Z(n20678) );
  ANDN U25778 ( .B(n22225), .A(n25432), .Z(n25430) );
  XNOR U25779 ( .A(n25433), .B(n20695), .Z(n19428) );
  XOR U25780 ( .A(n25434), .B(n21382), .Z(n20695) );
  NOR U25781 ( .A(n25435), .B(n20694), .Z(n25433) );
  XNOR U25782 ( .A(n16087), .B(n25436), .Z(n25428) );
  XOR U25783 ( .A(n19593), .B(n19512), .Z(n25436) );
  XNOR U25784 ( .A(n25437), .B(n20690), .Z(n19512) );
  XOR U25785 ( .A(n25438), .B(n24558), .Z(n20690) );
  ANDN U25786 ( .B(n22221), .A(n20691), .Z(n25437) );
  XNOR U25787 ( .A(n25439), .B(n20686), .Z(n19593) );
  XNOR U25788 ( .A(n25440), .B(n24769), .Z(n20686) );
  IV U25789 ( .A(n22394), .Z(n24769) );
  ANDN U25790 ( .B(n20687), .A(n22216), .Z(n25439) );
  XOR U25791 ( .A(n25441), .B(n22029), .Z(n16087) );
  IV U25792 ( .A(n20682), .Z(n22029) );
  XOR U25793 ( .A(n23033), .B(n25442), .Z(n20682) );
  ANDN U25794 ( .B(n22229), .A(n20681), .Z(n25441) );
  IV U25795 ( .A(n25443), .Z(n20681) );
  XOR U25796 ( .A(n25444), .B(n19757), .Z(n15167) );
  XOR U25797 ( .A(n19671), .B(n20198), .Z(n19757) );
  XOR U25798 ( .A(n25445), .B(n25446), .Z(n20198) );
  XNOR U25799 ( .A(n20079), .B(n20909), .Z(n25446) );
  XNOR U25800 ( .A(n25447), .B(n20916), .Z(n20909) );
  XOR U25801 ( .A(n25448), .B(n25449), .Z(n20916) );
  ANDN U25802 ( .B(n20915), .A(n22440), .Z(n25447) );
  XNOR U25803 ( .A(n25450), .B(n20928), .Z(n20079) );
  XOR U25804 ( .A(n25451), .B(n25224), .Z(n20928) );
  XOR U25805 ( .A(n17484), .B(n25452), .Z(n25445) );
  XOR U25806 ( .A(n19274), .B(n19252), .Z(n25452) );
  XOR U25807 ( .A(n25453), .B(n20932), .Z(n19252) );
  XOR U25808 ( .A(n24971), .B(n25454), .Z(n20932) );
  ANDN U25809 ( .B(n20933), .A(n22443), .Z(n25453) );
  XOR U25810 ( .A(n25455), .B(n20919), .Z(n19274) );
  XNOR U25811 ( .A(n25456), .B(n25457), .Z(n20919) );
  AND U25812 ( .A(n25458), .B(n20920), .Z(n25455) );
  XNOR U25813 ( .A(n25459), .B(n20924), .Z(n17484) );
  IV U25814 ( .A(n22519), .Z(n20924) );
  XOR U25815 ( .A(n25460), .B(n25361), .Z(n22519) );
  XOR U25816 ( .A(n25461), .B(n25462), .Z(n19671) );
  XNOR U25817 ( .A(n18490), .B(n21975), .Z(n25462) );
  XOR U25818 ( .A(n25463), .B(n21979), .Z(n21975) );
  XNOR U25819 ( .A(n25464), .B(n25465), .Z(n21979) );
  XOR U25820 ( .A(n25466), .B(n21989), .Z(n18490) );
  XNOR U25821 ( .A(n25467), .B(n21590), .Z(n21989) );
  NOR U25822 ( .A(n23344), .B(n21988), .Z(n25466) );
  XNOR U25823 ( .A(n19117), .B(n25468), .Z(n25461) );
  XOR U25824 ( .A(n19221), .B(n18091), .Z(n25468) );
  XOR U25825 ( .A(n25469), .B(n21991), .Z(n18091) );
  XNOR U25826 ( .A(n23840), .B(n25470), .Z(n21991) );
  ANDN U25827 ( .B(n21992), .A(n25471), .Z(n25469) );
  XOR U25828 ( .A(n25472), .B(n22800), .Z(n19221) );
  XOR U25829 ( .A(n25473), .B(n25144), .Z(n22800) );
  ANDN U25830 ( .B(n23038), .A(n22805), .Z(n25472) );
  XNOR U25831 ( .A(n25474), .B(n21983), .Z(n19117) );
  ANDN U25832 ( .B(n21011), .A(n21982), .Z(n25474) );
  XOR U25833 ( .A(n25477), .B(n14635), .Z(n11410) );
  XOR U25834 ( .A(n25244), .B(n18828), .Z(n14635) );
  XNOR U25835 ( .A(n25478), .B(n25479), .Z(n20277) );
  XOR U25836 ( .A(n18247), .B(n22002), .Z(n25479) );
  XOR U25837 ( .A(n25480), .B(n21702), .Z(n22002) );
  XOR U25838 ( .A(n25481), .B(n25182), .Z(n21702) );
  ANDN U25839 ( .B(n25250), .A(n25249), .Z(n25480) );
  IV U25840 ( .A(n22026), .Z(n25249) );
  XOR U25841 ( .A(n25482), .B(n23864), .Z(n22026) );
  IV U25842 ( .A(n20841), .Z(n25250) );
  XOR U25843 ( .A(n25483), .B(n23727), .Z(n20841) );
  XOR U25844 ( .A(n25484), .B(n21697), .Z(n18247) );
  XNOR U25845 ( .A(n25485), .B(n24825), .Z(n21697) );
  ANDN U25846 ( .B(n22009), .A(n20331), .Z(n25484) );
  XOR U25847 ( .A(n19750), .B(n25486), .Z(n25478) );
  XOR U25848 ( .A(n19453), .B(n18880), .Z(n25486) );
  XNOR U25849 ( .A(n25487), .B(n21692), .Z(n18880) );
  XOR U25850 ( .A(n25488), .B(n25489), .Z(n21692) );
  ANDN U25851 ( .B(n20335), .A(n22022), .Z(n25487) );
  XNOR U25852 ( .A(n25490), .B(n25491), .Z(n22022) );
  XNOR U25853 ( .A(n25492), .B(n24395), .Z(n20335) );
  XNOR U25854 ( .A(n25493), .B(n21694), .Z(n19453) );
  XNOR U25855 ( .A(n24423), .B(n25494), .Z(n21694) );
  ANDN U25856 ( .B(n20325), .A(n22013), .Z(n25493) );
  IV U25857 ( .A(n25238), .Z(n22013) );
  XOR U25858 ( .A(n25495), .B(n22401), .Z(n25238) );
  XNOR U25859 ( .A(n25496), .B(n23577), .Z(n20325) );
  XNOR U25860 ( .A(n25497), .B(n21699), .Z(n19750) );
  XNOR U25861 ( .A(n25498), .B(n23815), .Z(n21699) );
  XOR U25862 ( .A(n25499), .B(n23040), .Z(n22018) );
  XOR U25863 ( .A(n25500), .B(n25501), .Z(n21416) );
  XOR U25864 ( .A(n25502), .B(n25503), .Z(n19193) );
  XNOR U25865 ( .A(n24135), .B(n17247), .Z(n25503) );
  XNOR U25866 ( .A(n25504), .B(n23915), .Z(n17247) );
  XOR U25867 ( .A(n25505), .B(n23878), .Z(n23915) );
  XOR U25868 ( .A(n25506), .B(n23792), .Z(n20345) );
  XOR U25869 ( .A(n25507), .B(n22613), .Z(n21405) );
  IV U25870 ( .A(n25405), .Z(n22613) );
  XOR U25871 ( .A(n25508), .B(n23918), .Z(n24135) );
  XNOR U25872 ( .A(n25509), .B(n25382), .Z(n23918) );
  XOR U25873 ( .A(n25510), .B(n21584), .Z(n21412) );
  XNOR U25874 ( .A(n25511), .B(n24554), .Z(n20351) );
  IV U25875 ( .A(n22899), .Z(n24554) );
  XOR U25876 ( .A(n25512), .B(n25513), .Z(n22899) );
  XOR U25877 ( .A(n18579), .B(n25514), .Z(n25502) );
  XOR U25878 ( .A(n21145), .B(n18299), .Z(n25514) );
  XNOR U25879 ( .A(n25515), .B(n23921), .Z(n18299) );
  XOR U25880 ( .A(n25516), .B(n24949), .Z(n23921) );
  ANDN U25881 ( .B(n20991), .A(n21403), .Z(n25515) );
  XOR U25882 ( .A(n24963), .B(n25517), .Z(n21403) );
  XOR U25883 ( .A(n25518), .B(n24397), .Z(n20991) );
  XNOR U25884 ( .A(n25519), .B(n23907), .Z(n21145) );
  IV U25885 ( .A(n24173), .Z(n23907) );
  XOR U25886 ( .A(n25520), .B(n23482), .Z(n24173) );
  XNOR U25887 ( .A(n25403), .B(n25521), .Z(n23482) );
  XOR U25888 ( .A(n25522), .B(n25523), .Z(n25403) );
  XNOR U25889 ( .A(n25524), .B(n25525), .Z(n25523) );
  XNOR U25890 ( .A(n25526), .B(n25527), .Z(n25522) );
  XNOR U25891 ( .A(n24434), .B(n23423), .Z(n25527) );
  XOR U25892 ( .A(n25528), .B(n25529), .Z(n23423) );
  AND U25893 ( .A(n25530), .B(n25531), .Z(n25528) );
  XNOR U25894 ( .A(n25532), .B(n25533), .Z(n24434) );
  ANDN U25895 ( .B(n25534), .A(n25535), .Z(n25532) );
  ANDN U25896 ( .B(n20355), .A(n21414), .Z(n25519) );
  XOR U25897 ( .A(n25536), .B(n25152), .Z(n21414) );
  XNOR U25898 ( .A(n24423), .B(n25537), .Z(n20355) );
  XNOR U25899 ( .A(n25538), .B(n23910), .Z(n18579) );
  XOR U25900 ( .A(n25539), .B(n21601), .Z(n23910) );
  NOR U25901 ( .A(n21409), .B(n20341), .Z(n25538) );
  XOR U25902 ( .A(n23025), .B(n25540), .Z(n20341) );
  IV U25903 ( .A(n24167), .Z(n21409) );
  XOR U25904 ( .A(n24209), .B(n25541), .Z(n24167) );
  XNOR U25905 ( .A(n25542), .B(n22009), .Z(n25244) );
  XOR U25906 ( .A(n25543), .B(n21716), .Z(n22009) );
  ANDN U25907 ( .B(n20331), .A(n20332), .Z(n25542) );
  XOR U25908 ( .A(n24390), .B(n25544), .Z(n20332) );
  XOR U25909 ( .A(n25545), .B(n24525), .Z(n20331) );
  NOR U25910 ( .A(n15171), .B(n15172), .Z(n25477) );
  XNOR U25911 ( .A(n25546), .B(n15948), .Z(n15172) );
  IV U25912 ( .A(n22666), .Z(n15948) );
  XNOR U25913 ( .A(n23783), .B(n24078), .Z(n22666) );
  XNOR U25914 ( .A(n25547), .B(n25548), .Z(n24078) );
  XOR U25915 ( .A(n18005), .B(n19505), .Z(n25548) );
  XOR U25916 ( .A(n25549), .B(n23292), .Z(n19505) );
  XOR U25917 ( .A(n25550), .B(n25551), .Z(n23292) );
  AND U25918 ( .A(n23293), .B(n23171), .Z(n25549) );
  XNOR U25919 ( .A(n25552), .B(n23303), .Z(n18005) );
  XOR U25920 ( .A(n25553), .B(n23021), .Z(n23303) );
  NOR U25921 ( .A(n23161), .B(n23302), .Z(n25552) );
  XOR U25922 ( .A(n19758), .B(n25554), .Z(n25547) );
  XOR U25923 ( .A(n23262), .B(n18303), .Z(n25554) );
  XNOR U25924 ( .A(n25555), .B(n24877), .Z(n18303) );
  XOR U25925 ( .A(n24662), .B(n25556), .Z(n24877) );
  NOR U25926 ( .A(n25557), .B(n24889), .Z(n25555) );
  XOR U25927 ( .A(n25558), .B(n23299), .Z(n23262) );
  XNOR U25928 ( .A(n25559), .B(n24844), .Z(n23299) );
  IV U25929 ( .A(n24566), .Z(n24844) );
  ANDN U25930 ( .B(n23175), .A(n25560), .Z(n25558) );
  XNOR U25931 ( .A(n25561), .B(n23297), .Z(n19758) );
  XNOR U25932 ( .A(n25562), .B(n23577), .Z(n23297) );
  NOR U25933 ( .A(n23296), .B(n23165), .Z(n25561) );
  XOR U25934 ( .A(n25563), .B(n25564), .Z(n23783) );
  XNOR U25935 ( .A(n18522), .B(n20600), .Z(n25564) );
  XOR U25936 ( .A(n25565), .B(n21790), .Z(n20600) );
  ANDN U25937 ( .B(n21522), .A(n21789), .Z(n25565) );
  XOR U25938 ( .A(n25566), .B(n21786), .Z(n18522) );
  NOR U25939 ( .A(n25567), .B(n21518), .Z(n25566) );
  XOR U25940 ( .A(n16411), .B(n25568), .Z(n25563) );
  XOR U25941 ( .A(n17583), .B(n16901), .Z(n25568) );
  XOR U25942 ( .A(n25569), .B(n21782), .Z(n16901) );
  ANDN U25943 ( .B(n21783), .A(n23082), .Z(n25569) );
  XNOR U25944 ( .A(n25570), .B(n21794), .Z(n17583) );
  NOR U25945 ( .A(n21793), .B(n25571), .Z(n25570) );
  XOR U25946 ( .A(n25572), .B(n21778), .Z(n16411) );
  ANDN U25947 ( .B(n21512), .A(n21779), .Z(n25572) );
  XNOR U25948 ( .A(n20893), .B(n18692), .Z(n15171) );
  XNOR U25949 ( .A(n19774), .B(n18668), .Z(n18692) );
  XNOR U25950 ( .A(n25573), .B(n25574), .Z(n18668) );
  XNOR U25951 ( .A(n21393), .B(n18576), .Z(n25574) );
  XNOR U25952 ( .A(n25575), .B(n22142), .Z(n18576) );
  XOR U25953 ( .A(n24613), .B(n25576), .Z(n22142) );
  XNOR U25954 ( .A(n25577), .B(n25578), .Z(n20888) );
  XOR U25955 ( .A(n21593), .B(n25579), .Z(n19805) );
  XOR U25956 ( .A(n25582), .B(n22144), .Z(n21393) );
  XOR U25957 ( .A(n25583), .B(n24257), .Z(n22144) );
  NOR U25958 ( .A(n19814), .B(n20890), .Z(n25582) );
  XOR U25959 ( .A(n25584), .B(n23602), .Z(n20890) );
  IV U25960 ( .A(n20891), .Z(n19814) );
  XNOR U25961 ( .A(n25585), .B(n22227), .Z(n20891) );
  XNOR U25962 ( .A(n19082), .B(n25586), .Z(n25573) );
  XOR U25963 ( .A(n18908), .B(n17243), .Z(n25586) );
  XNOR U25964 ( .A(n25587), .B(n22137), .Z(n17243) );
  XOR U25965 ( .A(n25588), .B(n24792), .Z(n22137) );
  IV U25966 ( .A(n24458), .Z(n24792) );
  XNOR U25967 ( .A(n25589), .B(n25590), .Z(n24458) );
  ANDN U25968 ( .B(n19810), .A(n20898), .Z(n25587) );
  XNOR U25969 ( .A(n23695), .B(n25591), .Z(n20898) );
  XNOR U25970 ( .A(n25592), .B(n25382), .Z(n19810) );
  XOR U25971 ( .A(n25593), .B(n22140), .Z(n18908) );
  XOR U25972 ( .A(n25594), .B(n22213), .Z(n22140) );
  NOR U25973 ( .A(n19801), .B(n20895), .Z(n25593) );
  XNOR U25974 ( .A(n25595), .B(n25596), .Z(n20895) );
  IV U25975 ( .A(n20896), .Z(n19801) );
  XOR U25976 ( .A(n25597), .B(n21823), .Z(n20896) );
  XOR U25977 ( .A(n25598), .B(n22656), .Z(n19082) );
  IV U25978 ( .A(n22651), .Z(n22656) );
  XNOR U25979 ( .A(n25599), .B(n23145), .Z(n22651) );
  NOR U25980 ( .A(n19818), .B(n22655), .Z(n25598) );
  XNOR U25981 ( .A(n25600), .B(n25601), .Z(n19774) );
  XOR U25982 ( .A(n16057), .B(n17511), .Z(n25601) );
  XNOR U25983 ( .A(n25602), .B(n22614), .Z(n17511) );
  ANDN U25984 ( .B(n22176), .A(n22177), .Z(n25602) );
  XOR U25985 ( .A(n25603), .B(n25604), .Z(n22177) );
  XOR U25986 ( .A(n25605), .B(n22610), .Z(n16057) );
  NOR U25987 ( .A(n22174), .B(n21316), .Z(n25605) );
  XOR U25988 ( .A(n25606), .B(n23065), .Z(n21316) );
  XNOR U25989 ( .A(n18388), .B(n25607), .Z(n25600) );
  XNOR U25990 ( .A(n18537), .B(n25608), .Z(n25607) );
  XNOR U25991 ( .A(n25609), .B(n22622), .Z(n18537) );
  ANDN U25992 ( .B(n21320), .A(n22180), .Z(n25609) );
  XNOR U25993 ( .A(n22635), .B(n25610), .Z(n21320) );
  XOR U25994 ( .A(n25611), .B(n25612), .Z(n18388) );
  ANDN U25995 ( .B(n22168), .A(n21310), .Z(n25611) );
  XOR U25996 ( .A(n25613), .B(n22949), .Z(n21310) );
  XNOR U25997 ( .A(n25614), .B(n22655), .Z(n20893) );
  XOR U25998 ( .A(n24899), .B(n25615), .Z(n22655) );
  ANDN U25999 ( .B(n19818), .A(n22650), .Z(n25614) );
  XOR U26000 ( .A(n25616), .B(n21229), .Z(n22650) );
  XOR U26001 ( .A(n22624), .B(n25617), .Z(n19818) );
  XOR U26002 ( .A(n25618), .B(n14632), .Z(n15175) );
  XNOR U26003 ( .A(n22914), .B(n17392), .Z(n14632) );
  IV U26004 ( .A(n15663), .Z(n17392) );
  XNOR U26005 ( .A(n21504), .B(n18394), .Z(n15663) );
  XNOR U26006 ( .A(n25619), .B(n25620), .Z(n18394) );
  XNOR U26007 ( .A(n23882), .B(n18671), .Z(n25620) );
  XNOR U26008 ( .A(n25621), .B(n25622), .Z(n18671) );
  ANDN U26009 ( .B(n22921), .A(n25623), .Z(n25621) );
  XNOR U26010 ( .A(n25624), .B(n23186), .Z(n23882) );
  ANDN U26011 ( .B(n22925), .A(n25625), .Z(n25624) );
  XOR U26012 ( .A(n25626), .B(n25627), .Z(n25619) );
  XOR U26013 ( .A(n21238), .B(n16771), .Z(n25627) );
  XOR U26014 ( .A(n25628), .B(n23195), .Z(n16771) );
  ANDN U26015 ( .B(n22916), .A(n22917), .Z(n25628) );
  XNOR U26016 ( .A(n25629), .B(n23190), .Z(n21238) );
  ANDN U26017 ( .B(n22929), .A(n22930), .Z(n25629) );
  XNOR U26018 ( .A(n25630), .B(n25631), .Z(n21504) );
  XNOR U26019 ( .A(n16810), .B(n22997), .Z(n25631) );
  XNOR U26020 ( .A(n25632), .B(n23215), .Z(n22997) );
  ANDN U26021 ( .B(n22453), .A(n25633), .Z(n25632) );
  XNOR U26022 ( .A(n25634), .B(n23210), .Z(n16810) );
  ANDN U26023 ( .B(n25635), .A(n22463), .Z(n25634) );
  XNOR U26024 ( .A(n18497), .B(n25636), .Z(n25630) );
  XNOR U26025 ( .A(n19378), .B(n17463), .Z(n25636) );
  XNOR U26026 ( .A(n25637), .B(n23207), .Z(n17463) );
  ANDN U26027 ( .B(n25638), .A(n25639), .Z(n25637) );
  XNOR U26028 ( .A(n25640), .B(n23213), .Z(n19378) );
  ANDN U26029 ( .B(n25641), .A(n25642), .Z(n25640) );
  XOR U26030 ( .A(n25643), .B(n23218), .Z(n18497) );
  NOR U26031 ( .A(n22459), .B(n25644), .Z(n25643) );
  IV U26032 ( .A(n25645), .Z(n22459) );
  XOR U26033 ( .A(n25646), .B(n25647), .Z(n22914) );
  ANDN U26034 ( .B(n25648), .A(n23200), .Z(n25646) );
  ANDN U26035 ( .B(n16594), .A(n15476), .Z(n25618) );
  XNOR U26036 ( .A(n23359), .B(n17432), .Z(n15476) );
  XNOR U26037 ( .A(n25649), .B(n22572), .Z(n23359) );
  ANDN U26038 ( .B(n24307), .A(n25650), .Z(n25649) );
  XOR U26039 ( .A(n23405), .B(n17898), .Z(n16594) );
  XOR U26040 ( .A(n24890), .B(n19677), .Z(n17898) );
  XNOR U26041 ( .A(n25651), .B(n25652), .Z(n19677) );
  XNOR U26042 ( .A(n15646), .B(n18940), .Z(n25652) );
  XOR U26043 ( .A(n25653), .B(n20461), .Z(n18940) );
  XOR U26044 ( .A(n25654), .B(n23869), .Z(n20461) );
  ANDN U26045 ( .B(n22687), .A(n23402), .Z(n25653) );
  XOR U26046 ( .A(n25655), .B(n22504), .Z(n23402) );
  XOR U26047 ( .A(n25656), .B(n24162), .Z(n22687) );
  XOR U26048 ( .A(n25657), .B(n20451), .Z(n15646) );
  IV U26049 ( .A(n24944), .Z(n20451) );
  XNOR U26050 ( .A(n25658), .B(n23442), .Z(n24944) );
  XOR U26051 ( .A(n25659), .B(n25660), .Z(n22698) );
  XOR U26052 ( .A(n25001), .B(n25661), .Z(n20452) );
  XOR U26053 ( .A(n18265), .B(n25662), .Z(n25651) );
  XNOR U26054 ( .A(n19297), .B(n15683), .Z(n25662) );
  XOR U26055 ( .A(n25663), .B(n22359), .Z(n15683) );
  XOR U26056 ( .A(n24632), .B(n25664), .Z(n22359) );
  ANDN U26057 ( .B(n22360), .A(n23394), .Z(n25663) );
  IV U26058 ( .A(n22684), .Z(n23394) );
  XNOR U26059 ( .A(n25665), .B(n21833), .Z(n22684) );
  XOR U26060 ( .A(n25666), .B(n24835), .Z(n22360) );
  XOR U26061 ( .A(n25668), .B(n24558), .Z(n20457) );
  ANDN U26062 ( .B(n20458), .A(n22695), .Z(n25667) );
  XOR U26063 ( .A(n23991), .B(n25669), .Z(n22695) );
  IV U26064 ( .A(n23398), .Z(n20458) );
  XOR U26065 ( .A(n24605), .B(n25670), .Z(n23398) );
  XNOR U26066 ( .A(n25671), .B(n24950), .Z(n18265) );
  XNOR U26067 ( .A(n25672), .B(n25673), .Z(n24950) );
  AND U26068 ( .A(n22691), .B(n23400), .Z(n25671) );
  XOR U26069 ( .A(n24069), .B(n25674), .Z(n23400) );
  XNOR U26070 ( .A(n25675), .B(n21216), .Z(n22691) );
  XOR U26071 ( .A(n25676), .B(n25677), .Z(n24890) );
  XNOR U26072 ( .A(n17979), .B(n19334), .Z(n25677) );
  XNOR U26073 ( .A(n25678), .B(n25679), .Z(n19334) );
  ANDN U26074 ( .B(n21966), .A(n23407), .Z(n25678) );
  XOR U26075 ( .A(n25680), .B(n25085), .Z(n21966) );
  XNOR U26076 ( .A(n25681), .B(n23606), .Z(n17979) );
  ANDN U26077 ( .B(n25682), .A(n21952), .Z(n25681) );
  XOR U26078 ( .A(n20444), .B(n25683), .Z(n25676) );
  XNOR U26079 ( .A(n19944), .B(n17101), .Z(n25683) );
  XNOR U26080 ( .A(n25684), .B(n23603), .Z(n17101) );
  ANDN U26081 ( .B(n23410), .A(n23388), .Z(n25684) );
  XOR U26082 ( .A(n25685), .B(n21590), .Z(n23388) );
  IV U26083 ( .A(n25686), .Z(n21590) );
  XOR U26084 ( .A(n25687), .B(n23594), .Z(n19944) );
  ANDN U26085 ( .B(n23412), .A(n21956), .Z(n25687) );
  IV U26086 ( .A(n23413), .Z(n21956) );
  XOR U26087 ( .A(n25688), .B(n21382), .Z(n23413) );
  XOR U26088 ( .A(n25689), .B(n23609), .Z(n20444) );
  NOR U26089 ( .A(n21962), .B(n23415), .Z(n25689) );
  IV U26090 ( .A(n23416), .Z(n21962) );
  XNOR U26091 ( .A(n25690), .B(n23584), .Z(n23416) );
  XNOR U26092 ( .A(n25691), .B(n25682), .Z(n23405) );
  AND U26093 ( .A(n21952), .B(n21953), .Z(n25691) );
  XOR U26094 ( .A(n25692), .B(n24745), .Z(n21953) );
  XOR U26095 ( .A(n25693), .B(n24035), .Z(n21952) );
  XOR U26096 ( .A(n9107), .B(n13490), .Z(n7132) );
  XOR U26097 ( .A(n25694), .B(n14727), .Z(n13490) );
  ANDN U26098 ( .B(n16726), .A(n16213), .Z(n25694) );
  XNOR U26099 ( .A(n25695), .B(n18074), .Z(n16213) );
  XOR U26100 ( .A(n25696), .B(n25697), .Z(n12768) );
  XNOR U26101 ( .A(n9887), .B(n11443), .Z(n25697) );
  XNOR U26102 ( .A(n25698), .B(n18129), .Z(n11443) );
  XOR U26103 ( .A(n16822), .B(n23095), .Z(n18129) );
  XOR U26104 ( .A(n25699), .B(n25700), .Z(n23095) );
  ANDN U26105 ( .B(n25701), .A(n21909), .Z(n25699) );
  IV U26106 ( .A(n22901), .Z(n16822) );
  XOR U26107 ( .A(n20865), .B(n19558), .Z(n22901) );
  XOR U26108 ( .A(n25702), .B(n25703), .Z(n19558) );
  XOR U26109 ( .A(n18771), .B(n17248), .Z(n25703) );
  XOR U26110 ( .A(n25704), .B(n22971), .Z(n17248) );
  XOR U26111 ( .A(n25705), .B(n24349), .Z(n22971) );
  IV U26112 ( .A(n25706), .Z(n24349) );
  ANDN U26113 ( .B(n22996), .A(n23119), .Z(n25704) );
  XNOR U26114 ( .A(n25707), .B(n22790), .Z(n23119) );
  XNOR U26115 ( .A(n23033), .B(n25708), .Z(n22996) );
  XOR U26116 ( .A(n25709), .B(n25710), .Z(n23033) );
  XNOR U26117 ( .A(n25711), .B(n22194), .Z(n18771) );
  XNOR U26118 ( .A(n25712), .B(n23878), .Z(n22194) );
  NOR U26119 ( .A(n23108), .B(n23109), .Z(n25711) );
  XOR U26120 ( .A(n25713), .B(n24506), .Z(n23109) );
  IV U26121 ( .A(n22195), .Z(n23108) );
  XOR U26122 ( .A(n25714), .B(n23597), .Z(n22195) );
  XNOR U26123 ( .A(n18719), .B(n25715), .Z(n25702) );
  XOR U26124 ( .A(n19275), .B(n19966), .Z(n25715) );
  XNOR U26125 ( .A(n25716), .B(n22190), .Z(n19966) );
  XOR U26126 ( .A(n25476), .B(n25717), .Z(n22190) );
  ANDN U26127 ( .B(n23114), .A(n23113), .Z(n25716) );
  IV U26128 ( .A(n22191), .Z(n23113) );
  XOR U26129 ( .A(n25718), .B(n22521), .Z(n22191) );
  XOR U26130 ( .A(n25719), .B(n21225), .Z(n23114) );
  XOR U26131 ( .A(n25720), .B(n22200), .Z(n19275) );
  XOR U26132 ( .A(n23699), .B(n25721), .Z(n22200) );
  IV U26133 ( .A(n24783), .Z(n23699) );
  NOR U26134 ( .A(n23106), .B(n22201), .Z(n25720) );
  XOR U26135 ( .A(n25722), .B(n21728), .Z(n22201) );
  XNOR U26136 ( .A(n25723), .B(n21221), .Z(n23106) );
  XOR U26137 ( .A(n25724), .B(n22205), .Z(n18719) );
  XOR U26138 ( .A(n25725), .B(n22342), .Z(n22205) );
  NOR U26139 ( .A(n24268), .B(n22204), .Z(n25724) );
  XOR U26140 ( .A(n25728), .B(n23139), .Z(n22204) );
  XOR U26141 ( .A(n24613), .B(n25729), .Z(n24268) );
  XOR U26142 ( .A(n25730), .B(n25731), .Z(n20865) );
  XOR U26143 ( .A(n17305), .B(n18327), .Z(n25731) );
  XOR U26144 ( .A(n25732), .B(n23523), .Z(n18327) );
  AND U26145 ( .A(n23097), .B(n23099), .Z(n25732) );
  XNOR U26146 ( .A(n25733), .B(n21925), .Z(n17305) );
  ANDN U26147 ( .B(n23102), .A(n23101), .Z(n25733) );
  XNOR U26148 ( .A(n21501), .B(n25734), .Z(n25730) );
  XNOR U26149 ( .A(n22184), .B(n18313), .Z(n25734) );
  XOR U26150 ( .A(n25735), .B(n21911), .Z(n18313) );
  NOR U26151 ( .A(n25700), .B(n25701), .Z(n25735) );
  IV U26152 ( .A(n25736), .Z(n25700) );
  NOR U26153 ( .A(n25738), .B(n23089), .Z(n25737) );
  IV U26154 ( .A(n23088), .Z(n25738) );
  XNOR U26155 ( .A(n25739), .B(n21914), .Z(n21501) );
  ANDN U26156 ( .B(n23092), .A(n25740), .Z(n25739) );
  ANDN U26157 ( .B(n15927), .A(n15928), .Z(n25698) );
  XOR U26158 ( .A(n21432), .B(n18865), .Z(n15928) );
  IV U26159 ( .A(n18058), .Z(n18865) );
  XOR U26160 ( .A(n20085), .B(n25285), .Z(n18058) );
  XOR U26161 ( .A(n25741), .B(n25742), .Z(n25285) );
  XOR U26162 ( .A(n18410), .B(n16743), .Z(n25742) );
  XOR U26163 ( .A(n25743), .B(n24133), .Z(n16743) );
  XNOR U26164 ( .A(n25426), .B(n25744), .Z(n24133) );
  IV U26165 ( .A(n25745), .Z(n25426) );
  AND U26166 ( .A(n25299), .B(n24134), .Z(n25743) );
  XNOR U26167 ( .A(n25746), .B(n24676), .Z(n18410) );
  XOR U26168 ( .A(n25747), .B(n23855), .Z(n24676) );
  ANDN U26169 ( .B(n21428), .A(n21427), .Z(n25746) );
  IV U26170 ( .A(n24691), .Z(n21427) );
  XOR U26171 ( .A(n25748), .B(n25749), .Z(n24691) );
  XNOR U26172 ( .A(n25750), .B(n21716), .Z(n21428) );
  IV U26173 ( .A(n22406), .Z(n21716) );
  XOR U26174 ( .A(n25751), .B(n25752), .Z(n22406) );
  XOR U26175 ( .A(n17664), .B(n25753), .Z(n25741) );
  XNOR U26176 ( .A(n24098), .B(n18335), .Z(n25753) );
  XOR U26177 ( .A(n25754), .B(n24122), .Z(n18335) );
  XOR U26178 ( .A(n25755), .B(n25111), .Z(n24122) );
  ANDN U26179 ( .B(n22276), .A(n25309), .Z(n25754) );
  IV U26180 ( .A(n22278), .Z(n25309) );
  XNOR U26181 ( .A(n25756), .B(n25757), .Z(n22278) );
  XOR U26182 ( .A(n25758), .B(n24166), .Z(n22276) );
  XOR U26183 ( .A(n25759), .B(n24130), .Z(n24098) );
  XOR U26184 ( .A(n25760), .B(n24998), .Z(n24130) );
  AND U26185 ( .A(n21423), .B(n21425), .Z(n25759) );
  XOR U26186 ( .A(n25761), .B(n25762), .Z(n21425) );
  XOR U26187 ( .A(n25763), .B(n25673), .Z(n21423) );
  XNOR U26188 ( .A(n25764), .B(n24126), .Z(n17664) );
  XNOR U26189 ( .A(n25765), .B(n25766), .Z(n24126) );
  NOR U26190 ( .A(n24127), .B(n21435), .Z(n25764) );
  XOR U26191 ( .A(n24822), .B(n25767), .Z(n21435) );
  XOR U26192 ( .A(n25768), .B(n24031), .Z(n24127) );
  XOR U26193 ( .A(n25769), .B(n25770), .Z(n20085) );
  XNOR U26194 ( .A(n20136), .B(n17439), .Z(n25770) );
  XOR U26195 ( .A(n25771), .B(n24116), .Z(n17439) );
  XOR U26196 ( .A(n25772), .B(n21227), .Z(n24116) );
  NOR U26197 ( .A(n22297), .B(n22296), .Z(n25771) );
  XOR U26198 ( .A(n23686), .B(n25773), .Z(n22296) );
  XNOR U26199 ( .A(n25774), .B(n24110), .Z(n20136) );
  AND U26200 ( .A(n22287), .B(n22288), .Z(n25774) );
  XOR U26201 ( .A(n25775), .B(n25776), .Z(n22287) );
  XOR U26202 ( .A(n18703), .B(n25777), .Z(n25769) );
  XOR U26203 ( .A(n20569), .B(n18148), .Z(n25777) );
  XOR U26204 ( .A(n25778), .B(n24103), .Z(n18148) );
  XOR U26205 ( .A(n25779), .B(n21730), .Z(n24103) );
  ANDN U26206 ( .B(n22305), .A(n22304), .Z(n25778) );
  XOR U26207 ( .A(n24621), .B(n25780), .Z(n22304) );
  XNOR U26208 ( .A(n25781), .B(n24113), .Z(n20569) );
  XNOR U26209 ( .A(n25782), .B(n25045), .Z(n24113) );
  ANDN U26210 ( .B(n22293), .A(n22291), .Z(n25781) );
  XNOR U26211 ( .A(n25783), .B(n25673), .Z(n22291) );
  XNOR U26212 ( .A(n25784), .B(n24106), .Z(n18703) );
  XOR U26213 ( .A(n25785), .B(n24166), .Z(n24106) );
  ANDN U26214 ( .B(n22300), .A(n22301), .Z(n25784) );
  XOR U26215 ( .A(n25786), .B(n22534), .Z(n22300) );
  XNOR U26216 ( .A(n25787), .B(n24134), .Z(n21432) );
  XNOR U26217 ( .A(n23725), .B(n25788), .Z(n24134) );
  NOR U26218 ( .A(n24672), .B(n25299), .Z(n25787) );
  XOR U26219 ( .A(n24662), .B(n25789), .Z(n25299) );
  XOR U26220 ( .A(n25790), .B(n25278), .Z(n24672) );
  XOR U26221 ( .A(n24893), .B(n20143), .Z(n15927) );
  IV U26222 ( .A(n17632), .Z(n20143) );
  XOR U26223 ( .A(n20638), .B(n20445), .Z(n17632) );
  XNOR U26224 ( .A(n25791), .B(n25792), .Z(n20445) );
  XNOR U26225 ( .A(n19610), .B(n16049), .Z(n25792) );
  XOR U26226 ( .A(n25793), .B(n21963), .Z(n16049) );
  XOR U26227 ( .A(n25794), .B(n23040), .Z(n21963) );
  AND U26228 ( .A(n23609), .B(n23415), .Z(n25793) );
  XOR U26229 ( .A(n25448), .B(n25795), .Z(n23415) );
  XOR U26230 ( .A(n25796), .B(n21599), .Z(n23609) );
  XNOR U26231 ( .A(n25797), .B(n21954), .Z(n19610) );
  XOR U26232 ( .A(n25798), .B(n22834), .Z(n21954) );
  NOR U26233 ( .A(n23606), .B(n25682), .Z(n25797) );
  XNOR U26234 ( .A(n25799), .B(n25247), .Z(n25682) );
  XOR U26235 ( .A(n25800), .B(n25801), .Z(n23606) );
  XOR U26236 ( .A(n19439), .B(n25802), .Z(n25791) );
  XOR U26237 ( .A(n21091), .B(n15300), .Z(n25802) );
  XOR U26238 ( .A(n25803), .B(n21958), .Z(n15300) );
  XOR U26239 ( .A(n25804), .B(n25805), .Z(n21958) );
  ANDN U26240 ( .B(n23594), .A(n23412), .Z(n25803) );
  XOR U26241 ( .A(n25053), .B(n25806), .Z(n23412) );
  XOR U26242 ( .A(n25807), .B(n24518), .Z(n23594) );
  XOR U26243 ( .A(n25808), .B(n21968), .Z(n21091) );
  XOR U26244 ( .A(n25809), .B(n25810), .Z(n21968) );
  ANDN U26245 ( .B(n23407), .A(n25679), .Z(n25808) );
  IV U26246 ( .A(n23598), .Z(n25679) );
  XNOR U26247 ( .A(n25811), .B(n24162), .Z(n23598) );
  XOR U26248 ( .A(n25812), .B(n25813), .Z(n24162) );
  XOR U26249 ( .A(n25814), .B(n25745), .Z(n23407) );
  XNOR U26250 ( .A(n25815), .B(n23390), .Z(n19439) );
  IV U26251 ( .A(n23604), .Z(n23390) );
  XOR U26252 ( .A(n25816), .B(n23513), .Z(n23604) );
  NOR U26253 ( .A(n23603), .B(n23410), .Z(n25815) );
  XNOR U26254 ( .A(n25817), .B(n25305), .Z(n23410) );
  XOR U26255 ( .A(n25476), .B(n25818), .Z(n23603) );
  XOR U26256 ( .A(n25819), .B(n25820), .Z(n20638) );
  XNOR U26257 ( .A(n20995), .B(n22256), .Z(n25820) );
  XNOR U26258 ( .A(n25821), .B(n21947), .Z(n22256) );
  XNOR U26259 ( .A(n25268), .B(n25822), .Z(n21947) );
  AND U26260 ( .A(n23618), .B(n22701), .Z(n25821) );
  XNOR U26261 ( .A(n25823), .B(n22526), .Z(n22701) );
  XOR U26262 ( .A(n25824), .B(n25825), .Z(n22526) );
  XNOR U26263 ( .A(n25826), .B(n21829), .Z(n23618) );
  XNOR U26264 ( .A(n25827), .B(n21941), .Z(n20995) );
  XOR U26265 ( .A(n25828), .B(n25829), .Z(n21941) );
  ANDN U26266 ( .B(n23624), .A(n24895), .Z(n25827) );
  XOR U26267 ( .A(n25745), .B(n25830), .Z(n24895) );
  XOR U26268 ( .A(n25831), .B(n25832), .Z(n23624) );
  XOR U26269 ( .A(n23588), .B(n25833), .Z(n25819) );
  XOR U26270 ( .A(n23518), .B(n18188), .Z(n25833) );
  XOR U26271 ( .A(n25834), .B(n21936), .Z(n18188) );
  XOR U26272 ( .A(n25835), .B(n25836), .Z(n21936) );
  AND U26273 ( .A(n20273), .B(n23628), .Z(n25834) );
  XOR U26274 ( .A(n25837), .B(n22951), .Z(n23628) );
  XOR U26275 ( .A(n25838), .B(n25222), .Z(n20273) );
  IV U26276 ( .A(n25839), .Z(n25222) );
  XNOR U26277 ( .A(n25840), .B(n21943), .Z(n23518) );
  IV U26278 ( .A(n23614), .Z(n21943) );
  XOR U26279 ( .A(n24241), .B(n25841), .Z(n23614) );
  IV U26280 ( .A(n25113), .Z(n24241) );
  XOR U26281 ( .A(n25842), .B(n25199), .Z(n25113) );
  XOR U26282 ( .A(n25843), .B(n25844), .Z(n25199) );
  XOR U26283 ( .A(n24803), .B(n23578), .Z(n25844) );
  XOR U26284 ( .A(n25845), .B(n25846), .Z(n23578) );
  ANDN U26285 ( .B(n25847), .A(n25848), .Z(n25845) );
  XNOR U26286 ( .A(n25849), .B(n25850), .Z(n24803) );
  ANDN U26287 ( .B(n25851), .A(n25852), .Z(n25849) );
  XNOR U26288 ( .A(n25853), .B(n25854), .Z(n25843) );
  XNOR U26289 ( .A(n24440), .B(n23036), .Z(n25854) );
  XNOR U26290 ( .A(n25855), .B(n25856), .Z(n23036) );
  ANDN U26291 ( .B(n25857), .A(n25858), .Z(n25855) );
  XNOR U26292 ( .A(n25859), .B(n25860), .Z(n24440) );
  ANDN U26293 ( .B(n25861), .A(n25862), .Z(n25859) );
  AND U26294 ( .A(n20266), .B(n23615), .Z(n25840) );
  XOR U26295 ( .A(n25863), .B(n21934), .Z(n23588) );
  XNOR U26296 ( .A(n25864), .B(n25865), .Z(n21934) );
  XOR U26297 ( .A(n25866), .B(n25170), .Z(n20262) );
  XOR U26298 ( .A(n24778), .B(n25867), .Z(n23622) );
  XNOR U26299 ( .A(n25868), .B(n23615), .Z(n24893) );
  XOR U26300 ( .A(n25869), .B(n23996), .Z(n23615) );
  NOR U26301 ( .A(n20267), .B(n20266), .Z(n25868) );
  XOR U26302 ( .A(n25870), .B(n25801), .Z(n20266) );
  XNOR U26303 ( .A(n25871), .B(n23040), .Z(n20267) );
  XNOR U26304 ( .A(n25872), .B(n25873), .Z(n23040) );
  XOR U26305 ( .A(n25874), .B(n19110), .Z(n9887) );
  XOR U26306 ( .A(n20314), .B(n20039), .Z(n19110) );
  XOR U26307 ( .A(n25875), .B(n25034), .Z(n20039) );
  XNOR U26308 ( .A(n25876), .B(n25877), .Z(n25034) );
  XNOR U26309 ( .A(n20194), .B(n17293), .Z(n25877) );
  XNOR U26310 ( .A(n25878), .B(n21135), .Z(n17293) );
  XOR U26311 ( .A(n25879), .B(n21730), .Z(n21135) );
  IV U26312 ( .A(n24262), .Z(n21730) );
  ANDN U26313 ( .B(n20985), .A(n20983), .Z(n25878) );
  XNOR U26314 ( .A(n24971), .B(n25880), .Z(n20983) );
  XNOR U26315 ( .A(n25881), .B(n19341), .Z(n20194) );
  XOR U26316 ( .A(n24009), .B(n25882), .Z(n19341) );
  IV U26317 ( .A(n24994), .Z(n24009) );
  NOR U26318 ( .A(n20313), .B(n20312), .Z(n25881) );
  XOR U26319 ( .A(n24196), .B(n25883), .Z(n20312) );
  XNOR U26320 ( .A(n20483), .B(n25884), .Z(n25876) );
  XNOR U26321 ( .A(n17504), .B(n18416), .Z(n25884) );
  XNOR U26322 ( .A(n25885), .B(n19346), .Z(n18416) );
  XNOR U26323 ( .A(n25886), .B(n22391), .Z(n19346) );
  IV U26324 ( .A(n25836), .Z(n22391) );
  XNOR U26325 ( .A(n25887), .B(n25888), .Z(n25836) );
  NOR U26326 ( .A(n21158), .B(n20319), .Z(n25885) );
  XOR U26327 ( .A(n25889), .B(n23510), .Z(n21158) );
  XNOR U26328 ( .A(n25890), .B(n19352), .Z(n17504) );
  XOR U26329 ( .A(n25891), .B(n24515), .Z(n19352) );
  NOR U26330 ( .A(n25892), .B(n21160), .Z(n25890) );
  XNOR U26331 ( .A(n25893), .B(n19356), .Z(n20483) );
  XNOR U26332 ( .A(n24461), .B(n25894), .Z(n19356) );
  IV U26333 ( .A(n24626), .Z(n24461) );
  ANDN U26334 ( .B(n21154), .A(n25895), .Z(n25893) );
  IV U26335 ( .A(n24012), .Z(n21154) );
  XOR U26336 ( .A(n25896), .B(n25897), .Z(n24012) );
  XNOR U26337 ( .A(n25898), .B(n21160), .Z(n20314) );
  XNOR U26338 ( .A(n25899), .B(n23864), .Z(n21160) );
  NOR U26339 ( .A(n25900), .B(n19350), .Z(n25898) );
  NOR U26340 ( .A(n15915), .B(n15914), .Z(n25874) );
  XNOR U26341 ( .A(n23674), .B(n19170), .Z(n15914) );
  IV U26342 ( .A(n18787), .Z(n19170) );
  XOR U26343 ( .A(n22079), .B(n19747), .Z(n18787) );
  XOR U26344 ( .A(n25901), .B(n25902), .Z(n19747) );
  XOR U26345 ( .A(n19555), .B(n17852), .Z(n25902) );
  XOR U26346 ( .A(n25903), .B(n23471), .Z(n17852) );
  ANDN U26347 ( .B(n23669), .A(n23668), .Z(n25903) );
  XNOR U26348 ( .A(n25904), .B(n23463), .Z(n19555) );
  XNOR U26349 ( .A(n25905), .B(n25906), .Z(n25901) );
  XOR U26350 ( .A(n24910), .B(n18367), .Z(n25906) );
  XNOR U26351 ( .A(n25907), .B(n23454), .Z(n18367) );
  NOR U26352 ( .A(n23676), .B(n23677), .Z(n25907) );
  XOR U26353 ( .A(n25908), .B(n23458), .Z(n24910) );
  ANDN U26354 ( .B(n25909), .A(n25910), .Z(n25908) );
  XOR U26355 ( .A(n25911), .B(n25912), .Z(n22079) );
  XOR U26356 ( .A(n19183), .B(n23804), .Z(n25912) );
  XNOR U26357 ( .A(n25913), .B(n23225), .Z(n23804) );
  ANDN U26358 ( .B(n20801), .A(n25135), .Z(n25913) );
  XOR U26359 ( .A(n25603), .B(n25914), .Z(n20801) );
  XOR U26360 ( .A(n25915), .B(n23238), .Z(n19183) );
  ANDN U26361 ( .B(n20796), .A(n25138), .Z(n25915) );
  XOR U26362 ( .A(n25916), .B(n25917), .Z(n20796) );
  XOR U26363 ( .A(n16085), .B(n25918), .Z(n25911) );
  XNOR U26364 ( .A(n18930), .B(n19493), .Z(n25918) );
  XOR U26365 ( .A(n25919), .B(n23235), .Z(n19493) );
  IV U26366 ( .A(n25920), .Z(n23235) );
  ANDN U26367 ( .B(n20809), .A(n25921), .Z(n25919) );
  XNOR U26368 ( .A(n25922), .B(n25099), .Z(n20809) );
  XOR U26369 ( .A(n25923), .B(n23233), .Z(n18930) );
  XOR U26370 ( .A(n25924), .B(n24577), .Z(n20805) );
  XNOR U26371 ( .A(n25925), .B(n25926), .Z(n16085) );
  NOR U26372 ( .A(n25142), .B(n25141), .Z(n25925) );
  XOR U26373 ( .A(n25927), .B(n25928), .Z(n25142) );
  XNOR U26374 ( .A(n25929), .B(n25910), .Z(n23674) );
  NOR U26375 ( .A(n23456), .B(n25909), .Z(n25929) );
  XOR U26376 ( .A(n23358), .B(n17432), .Z(n15915) );
  XNOR U26377 ( .A(n23005), .B(n21201), .Z(n17432) );
  XOR U26378 ( .A(n25930), .B(n25931), .Z(n21201) );
  XOR U26379 ( .A(n17739), .B(n15670), .Z(n25931) );
  XNOR U26380 ( .A(n25932), .B(n25002), .Z(n15670) );
  XNOR U26381 ( .A(n25933), .B(n21225), .Z(n25002) );
  ANDN U26382 ( .B(n20959), .A(n20958), .Z(n25932) );
  XOR U26383 ( .A(n22815), .B(n25934), .Z(n20958) );
  XNOR U26384 ( .A(n25935), .B(n22396), .Z(n20959) );
  XOR U26385 ( .A(n25936), .B(n25937), .Z(n22396) );
  XNOR U26386 ( .A(n25938), .B(n22545), .Z(n17739) );
  XNOR U26387 ( .A(n25939), .B(n25940), .Z(n22545) );
  NOR U26388 ( .A(n20950), .B(n20948), .Z(n25938) );
  XNOR U26389 ( .A(n25941), .B(n25942), .Z(n20948) );
  XNOR U26390 ( .A(n25943), .B(n22809), .Z(n20950) );
  XOR U26391 ( .A(n18641), .B(n25944), .Z(n25930) );
  XNOR U26392 ( .A(n18817), .B(n18320), .Z(n25944) );
  XOR U26393 ( .A(n25945), .B(n22550), .Z(n18320) );
  IV U26394 ( .A(n24996), .Z(n22550) );
  XNOR U26395 ( .A(n24904), .B(n25946), .Z(n24996) );
  XOR U26396 ( .A(n25164), .B(n25947), .Z(n20944) );
  XOR U26397 ( .A(n25948), .B(n25307), .Z(n20945) );
  IV U26398 ( .A(n23837), .Z(n25307) );
  XNOR U26399 ( .A(n25949), .B(n24990), .Z(n18817) );
  IV U26400 ( .A(n22553), .Z(n24990) );
  XNOR U26401 ( .A(n25950), .B(n23513), .Z(n22553) );
  NOR U26402 ( .A(n20954), .B(n20955), .Z(n25949) );
  XOR U26403 ( .A(n25951), .B(n25952), .Z(n20955) );
  XNOR U26404 ( .A(n25953), .B(n22982), .Z(n20954) );
  XNOR U26405 ( .A(n25954), .B(n22542), .Z(n18641) );
  XOR U26406 ( .A(n25955), .B(n23143), .Z(n22542) );
  NOR U26407 ( .A(n21204), .B(n21203), .Z(n25954) );
  XOR U26408 ( .A(n25956), .B(n22621), .Z(n21203) );
  XOR U26409 ( .A(n25957), .B(n25958), .Z(n21204) );
  XNOR U26410 ( .A(n25959), .B(n25960), .Z(n23005) );
  XNOR U26411 ( .A(n22537), .B(n18929), .Z(n25960) );
  XNOR U26412 ( .A(n25961), .B(n22562), .Z(n18929) );
  IV U26413 ( .A(n24305), .Z(n22562) );
  XOR U26414 ( .A(n25962), .B(n25963), .Z(n24305) );
  XOR U26415 ( .A(n23326), .B(n25964), .Z(n22563) );
  XNOR U26416 ( .A(n25965), .B(n24308), .Z(n22537) );
  IV U26417 ( .A(n22571), .Z(n24308) );
  XOR U26418 ( .A(n25966), .B(n23597), .Z(n22571) );
  IV U26419 ( .A(n23689), .Z(n23597) );
  XNOR U26420 ( .A(n25967), .B(n25968), .Z(n23689) );
  ANDN U26421 ( .B(n22572), .A(n25969), .Z(n25965) );
  XOR U26422 ( .A(n25970), .B(n25776), .Z(n22572) );
  XOR U26423 ( .A(n15640), .B(n25971), .Z(n25959) );
  XNOR U26424 ( .A(n19294), .B(n19604), .Z(n25971) );
  XOR U26425 ( .A(n25972), .B(n22575), .Z(n19604) );
  XOR U26426 ( .A(n25973), .B(n25974), .Z(n22575) );
  ANDN U26427 ( .B(n22576), .A(n23352), .Z(n25972) );
  XNOR U26428 ( .A(n25219), .B(n25975), .Z(n22576) );
  XNOR U26429 ( .A(n25976), .B(n22559), .Z(n19294) );
  XNOR U26430 ( .A(n25977), .B(n23978), .Z(n22559) );
  ANDN U26431 ( .B(n22558), .A(n25978), .Z(n25976) );
  XOR U26432 ( .A(n22313), .B(n25979), .Z(n22558) );
  IV U26433 ( .A(n22337), .Z(n22313) );
  XOR U26434 ( .A(n25980), .B(n25981), .Z(n22337) );
  XNOR U26435 ( .A(n25982), .B(n22567), .Z(n15640) );
  XOR U26436 ( .A(n25983), .B(n23510), .Z(n22567) );
  ANDN U26437 ( .B(n22568), .A(n25984), .Z(n25982) );
  XOR U26438 ( .A(n25985), .B(n22568), .Z(n23358) );
  XOR U26439 ( .A(n25986), .B(n25987), .Z(n22568) );
  ANDN U26440 ( .B(n24301), .A(n25988), .Z(n25985) );
  XOR U26441 ( .A(n18119), .B(n25989), .Z(n25696) );
  XNOR U26442 ( .A(n10831), .B(n10610), .Z(n25989) );
  XOR U26443 ( .A(n25990), .B(n18123), .Z(n10610) );
  XOR U26444 ( .A(n22243), .B(n17108), .Z(n18123) );
  XOR U26445 ( .A(n22999), .B(n19734), .Z(n17108) );
  XNOR U26446 ( .A(n25991), .B(n25992), .Z(n19734) );
  XNOR U26447 ( .A(n16375), .B(n25397), .Z(n25992) );
  XNOR U26448 ( .A(n25993), .B(n25443), .Z(n25397) );
  XOR U26449 ( .A(n25994), .B(n25940), .Z(n25443) );
  NOR U26450 ( .A(n22028), .B(n22229), .Z(n25993) );
  XOR U26451 ( .A(n25995), .B(n25996), .Z(n22229) );
  XNOR U26452 ( .A(n25997), .B(n24575), .Z(n22028) );
  IV U26453 ( .A(n21601), .Z(n24575) );
  XOR U26454 ( .A(n25998), .B(n25999), .Z(n21601) );
  XNOR U26455 ( .A(n26000), .B(n20694), .Z(n16375) );
  XOR U26456 ( .A(n26001), .B(n25032), .Z(n20694) );
  NOR U26457 ( .A(n22212), .B(n21243), .Z(n26000) );
  XNOR U26458 ( .A(n26002), .B(n22820), .Z(n21243) );
  IV U26459 ( .A(n25435), .Z(n22212) );
  XNOR U26460 ( .A(n26003), .B(n21833), .Z(n25435) );
  XOR U26461 ( .A(n26004), .B(n26005), .Z(n21833) );
  XOR U26462 ( .A(n23495), .B(n26006), .Z(n25991) );
  XOR U26463 ( .A(n17062), .B(n18901), .Z(n26006) );
  XNOR U26464 ( .A(n26007), .B(n20677), .Z(n18901) );
  IV U26465 ( .A(n25432), .Z(n20677) );
  XOR U26466 ( .A(n26008), .B(n25424), .Z(n25432) );
  NOR U26467 ( .A(n22225), .B(n21250), .Z(n26007) );
  XNOR U26468 ( .A(n23905), .B(n26009), .Z(n21250) );
  XOR U26469 ( .A(n26010), .B(n26011), .Z(n22225) );
  XOR U26470 ( .A(n26012), .B(n20691), .Z(n17062) );
  XOR U26471 ( .A(n26013), .B(n23602), .Z(n20691) );
  XOR U26472 ( .A(n26014), .B(n26015), .Z(n23602) );
  ANDN U26473 ( .B(n21252), .A(n22221), .Z(n26012) );
  XOR U26474 ( .A(n26016), .B(n26017), .Z(n22221) );
  XNOR U26475 ( .A(n26019), .B(n20687), .Z(n23495) );
  XOR U26476 ( .A(n26020), .B(n24272), .Z(n20687) );
  ANDN U26477 ( .B(n22216), .A(n21246), .Z(n26019) );
  XNOR U26478 ( .A(n26021), .B(n26022), .Z(n21246) );
  XOR U26479 ( .A(n26023), .B(n25163), .Z(n22216) );
  XOR U26480 ( .A(n26024), .B(n26025), .Z(n22999) );
  XNOR U26481 ( .A(n24211), .B(n20848), .Z(n26025) );
  XOR U26482 ( .A(n26026), .B(n22483), .Z(n20848) );
  XNOR U26483 ( .A(n26027), .B(n26028), .Z(n22483) );
  NOR U26484 ( .A(n22249), .B(n22250), .Z(n26026) );
  XNOR U26485 ( .A(n26029), .B(n26030), .Z(n22249) );
  XOR U26486 ( .A(n26031), .B(n22477), .Z(n24211) );
  IV U26487 ( .A(n24222), .Z(n22477) );
  XOR U26488 ( .A(n26032), .B(n24582), .Z(n24222) );
  NOR U26489 ( .A(n24221), .B(n26033), .Z(n26031) );
  XOR U26490 ( .A(n19205), .B(n26034), .Z(n26024) );
  XOR U26491 ( .A(n18274), .B(n20019), .Z(n26034) );
  XNOR U26492 ( .A(n26035), .B(n22480), .Z(n20019) );
  XNOR U26493 ( .A(n24776), .B(n26036), .Z(n22480) );
  IV U26494 ( .A(n24005), .Z(n24776) );
  NOR U26495 ( .A(n22239), .B(n22240), .Z(n26035) );
  XOR U26496 ( .A(n26037), .B(n24916), .Z(n22239) );
  XNOR U26497 ( .A(n26038), .B(n22469), .Z(n18274) );
  XOR U26498 ( .A(n26039), .B(n21721), .Z(n22469) );
  NOR U26499 ( .A(n26040), .B(n22235), .Z(n26038) );
  XOR U26500 ( .A(n26041), .B(n25829), .Z(n22235) );
  XNOR U26501 ( .A(n26042), .B(n22473), .Z(n19205) );
  IV U26502 ( .A(n24219), .Z(n22473) );
  XOR U26503 ( .A(n24963), .B(n26043), .Z(n24219) );
  ANDN U26504 ( .B(n22245), .A(n22246), .Z(n26042) );
  XOR U26505 ( .A(n24233), .B(n26044), .Z(n22245) );
  XNOR U26506 ( .A(n26045), .B(n24221), .Z(n22243) );
  XOR U26507 ( .A(n26046), .B(n25686), .Z(n24221) );
  ANDN U26508 ( .B(n26033), .A(n26047), .Z(n26045) );
  NOR U26509 ( .A(n15918), .B(n15919), .Z(n25990) );
  XOR U26510 ( .A(n21188), .B(n16112), .Z(n15919) );
  XOR U26511 ( .A(n23448), .B(n18818), .Z(n16112) );
  XNOR U26512 ( .A(n26048), .B(n26049), .Z(n18818) );
  XNOR U26513 ( .A(n18471), .B(n18172), .Z(n26049) );
  XOR U26514 ( .A(n26050), .B(n22893), .Z(n18172) );
  IV U26515 ( .A(n24972), .Z(n22893) );
  XOR U26516 ( .A(n26051), .B(n25829), .Z(n24972) );
  IV U26517 ( .A(n26022), .Z(n25829) );
  NOR U26518 ( .A(n20422), .B(n21197), .Z(n26050) );
  XNOR U26519 ( .A(n26052), .B(n26053), .Z(n21197) );
  XOR U26520 ( .A(n22815), .B(n26054), .Z(n20422) );
  IV U26521 ( .A(n24822), .Z(n22815) );
  XOR U26522 ( .A(n26055), .B(n26056), .Z(n24822) );
  XOR U26523 ( .A(n26057), .B(n22884), .Z(n18471) );
  XNOR U26524 ( .A(n26058), .B(n26059), .Z(n22884) );
  NOR U26525 ( .A(n24976), .B(n20431), .Z(n26057) );
  XOR U26526 ( .A(n18782), .B(n26060), .Z(n26048) );
  XOR U26527 ( .A(n21334), .B(n18718), .Z(n26060) );
  XOR U26528 ( .A(n26061), .B(n22888), .Z(n18718) );
  XNOR U26529 ( .A(n24344), .B(n26062), .Z(n22888) );
  XOR U26530 ( .A(n26063), .B(n25301), .Z(n20426) );
  XNOR U26531 ( .A(n26064), .B(n23019), .Z(n21200) );
  XNOR U26532 ( .A(n26065), .B(n22900), .Z(n21334) );
  XOR U26533 ( .A(n26066), .B(n22809), .Z(n22900) );
  ANDN U26534 ( .B(n21190), .A(n20439), .Z(n26065) );
  IV U26535 ( .A(n21191), .Z(n20439) );
  XNOR U26536 ( .A(n26067), .B(n24518), .Z(n21191) );
  XOR U26537 ( .A(n26068), .B(n22943), .Z(n21190) );
  XNOR U26538 ( .A(n26069), .B(n22896), .Z(n18782) );
  XOR U26539 ( .A(n26070), .B(n24414), .Z(n22896) );
  NOR U26540 ( .A(n20435), .B(n21194), .Z(n26069) );
  XOR U26541 ( .A(n24375), .B(n26071), .Z(n21194) );
  IV U26542 ( .A(n21195), .Z(n20435) );
  XOR U26543 ( .A(n22939), .B(n26072), .Z(n21195) );
  XNOR U26544 ( .A(n26073), .B(n26074), .Z(n23448) );
  XNOR U26545 ( .A(n18805), .B(n25695), .Z(n26074) );
  XNOR U26546 ( .A(n26075), .B(n19162), .Z(n25695) );
  IV U26547 ( .A(n26076), .Z(n19162) );
  NOR U26548 ( .A(n20410), .B(n21380), .Z(n26075) );
  XOR U26549 ( .A(n26077), .B(n26078), .Z(n20410) );
  XNOR U26550 ( .A(n26079), .B(n19156), .Z(n18805) );
  ANDN U26551 ( .B(n20415), .A(n21370), .Z(n26079) );
  XOR U26552 ( .A(n23145), .B(n26080), .Z(n20415) );
  XOR U26553 ( .A(n26081), .B(n26082), .Z(n23145) );
  XNOR U26554 ( .A(n20404), .B(n26083), .Z(n26073) );
  XNOR U26555 ( .A(n18073), .B(n26084), .Z(n26083) );
  XNOR U26556 ( .A(n26085), .B(n19152), .Z(n18073) );
  ANDN U26557 ( .B(n21378), .A(n21376), .Z(n26085) );
  IV U26558 ( .A(n26086), .Z(n21376) );
  XOR U26559 ( .A(n26087), .B(n23059), .Z(n21378) );
  XOR U26560 ( .A(n26088), .B(n19745), .Z(n20404) );
  ANDN U26561 ( .B(n20418), .A(n23446), .Z(n26088) );
  XNOR U26562 ( .A(n26089), .B(n26090), .Z(n20418) );
  XNOR U26563 ( .A(n26091), .B(n24976), .Z(n21188) );
  XOR U26564 ( .A(n26092), .B(n26093), .Z(n24976) );
  ANDN U26565 ( .B(n20431), .A(n20432), .Z(n26091) );
  XNOR U26566 ( .A(n26094), .B(n23053), .Z(n20432) );
  XNOR U26567 ( .A(n26095), .B(n23143), .Z(n20431) );
  IV U26568 ( .A(n24185), .Z(n23143) );
  XOR U26569 ( .A(n20874), .B(n15256), .Z(n15918) );
  XNOR U26570 ( .A(n26096), .B(n26097), .Z(n19956) );
  XOR U26571 ( .A(n17998), .B(n18198), .Z(n26097) );
  XNOR U26572 ( .A(n26098), .B(n22109), .Z(n18198) );
  NOR U26573 ( .A(n20876), .B(n20877), .Z(n26098) );
  XOR U26574 ( .A(n26099), .B(n23862), .Z(n20877) );
  IV U26575 ( .A(n23050), .Z(n23862) );
  XOR U26576 ( .A(n25577), .B(n26100), .Z(n20876) );
  XNOR U26577 ( .A(n26101), .B(n22105), .Z(n17998) );
  NOR U26578 ( .A(n20870), .B(n20871), .Z(n26101) );
  XNOR U26579 ( .A(n26102), .B(n22825), .Z(n20871) );
  XNOR U26580 ( .A(n24439), .B(n25853), .Z(n20870) );
  XOR U26581 ( .A(n26103), .B(n26104), .Z(n25853) );
  ANDN U26582 ( .B(n26105), .A(n26106), .Z(n26103) );
  XNOR U26583 ( .A(n26107), .B(n26108), .Z(n24439) );
  XOR U26584 ( .A(n18982), .B(n26109), .Z(n26096) );
  XNOR U26585 ( .A(n17587), .B(n17563), .Z(n26109) );
  XNOR U26586 ( .A(n26110), .B(n22103), .Z(n17563) );
  ANDN U26587 ( .B(n21679), .A(n22102), .Z(n26110) );
  XNOR U26588 ( .A(n26111), .B(n26112), .Z(n17587) );
  NOR U26589 ( .A(n21672), .B(n24466), .Z(n26111) );
  IV U26590 ( .A(n24467), .Z(n21672) );
  XNOR U26591 ( .A(n23725), .B(n26113), .Z(n24467) );
  XNOR U26592 ( .A(n26114), .B(n22111), .Z(n18982) );
  IV U26593 ( .A(n26115), .Z(n22111) );
  NOR U26594 ( .A(n20881), .B(n20880), .Z(n26114) );
  XOR U26595 ( .A(n23505), .B(n26116), .Z(n20880) );
  XNOR U26596 ( .A(n26117), .B(n25174), .Z(n20881) );
  IV U26597 ( .A(n24233), .Z(n25174) );
  XOR U26598 ( .A(n26118), .B(n26119), .Z(n24233) );
  XOR U26599 ( .A(n26120), .B(n26121), .Z(n22185) );
  XNOR U26600 ( .A(n15894), .B(n21392), .Z(n26121) );
  XNOR U26601 ( .A(n26122), .B(n23522), .Z(n21392) );
  ANDN U26602 ( .B(n23523), .A(n23097), .Z(n26122) );
  XOR U26603 ( .A(n24344), .B(n26123), .Z(n23097) );
  XNOR U26604 ( .A(n26124), .B(n23855), .Z(n23523) );
  XNOR U26605 ( .A(n26125), .B(n21924), .Z(n15894) );
  ANDN U26606 ( .B(n23101), .A(n21925), .Z(n26125) );
  XOR U26607 ( .A(n26126), .B(n24949), .Z(n21925) );
  XNOR U26608 ( .A(n26127), .B(n23566), .Z(n23101) );
  XOR U26609 ( .A(n21904), .B(n26128), .Z(n26120) );
  XNOR U26610 ( .A(n15637), .B(n18812), .Z(n26128) );
  XNOR U26611 ( .A(n26129), .B(n21910), .Z(n18812) );
  ANDN U26612 ( .B(n21911), .A(n25736), .Z(n26129) );
  XNOR U26613 ( .A(n24623), .B(n26130), .Z(n25736) );
  XOR U26614 ( .A(n26131), .B(n23727), .Z(n21911) );
  XNOR U26615 ( .A(n26132), .B(n21921), .Z(n15637) );
  ANDN U26616 ( .B(n21920), .A(n23088), .Z(n26132) );
  XOR U26617 ( .A(n23703), .B(n26133), .Z(n23088) );
  XOR U26618 ( .A(n24209), .B(n26134), .Z(n21920) );
  IV U26619 ( .A(n26135), .Z(n24209) );
  XNOR U26620 ( .A(n26136), .B(n26137), .Z(n21904) );
  NOR U26621 ( .A(n23092), .B(n21914), .Z(n26136) );
  XNOR U26622 ( .A(n25414), .B(n26138), .Z(n21914) );
  XOR U26623 ( .A(n26139), .B(n25083), .Z(n23092) );
  XNOR U26624 ( .A(n26140), .B(n22102), .Z(n20874) );
  XOR U26625 ( .A(n26141), .B(n21235), .Z(n22102) );
  ANDN U26626 ( .B(n21680), .A(n21679), .Z(n26140) );
  XNOR U26627 ( .A(n23998), .B(n26142), .Z(n21679) );
  XNOR U26628 ( .A(n26143), .B(n18125), .Z(n10831) );
  XOR U26629 ( .A(n21516), .B(n23080), .Z(n18125) );
  IV U26630 ( .A(n17498), .Z(n23080) );
  XNOR U26631 ( .A(n20607), .B(n26144), .Z(n17498) );
  XOR U26632 ( .A(n26145), .B(n26146), .Z(n20607) );
  XNOR U26633 ( .A(n25546), .B(n18157), .Z(n26146) );
  XNOR U26634 ( .A(n26147), .B(n21793), .Z(n18157) );
  XOR U26635 ( .A(n26148), .B(n24039), .Z(n21793) );
  ANDN U26636 ( .B(n25571), .A(n26149), .Z(n26147) );
  XOR U26637 ( .A(n26150), .B(n21787), .Z(n25546) );
  IV U26638 ( .A(n25567), .Z(n21787) );
  XOR U26639 ( .A(n23586), .B(n26151), .Z(n25567) );
  ANDN U26640 ( .B(n21518), .A(n21519), .Z(n26150) );
  XOR U26641 ( .A(n26152), .B(n25405), .Z(n21518) );
  XOR U26642 ( .A(n26154), .B(n26155), .Z(n24315) );
  XOR U26643 ( .A(n25178), .B(n22395), .Z(n26155) );
  XOR U26644 ( .A(n26156), .B(n26157), .Z(n22395) );
  ANDN U26645 ( .B(n26158), .A(n26159), .Z(n26156) );
  XNOR U26646 ( .A(n26160), .B(n26161), .Z(n25178) );
  ANDN U26647 ( .B(n26162), .A(n26163), .Z(n26160) );
  XNOR U26648 ( .A(n24718), .B(n26164), .Z(n26154) );
  XOR U26649 ( .A(n25072), .B(n25935), .Z(n26164) );
  XNOR U26650 ( .A(n26165), .B(n26166), .Z(n25935) );
  ANDN U26651 ( .B(n26167), .A(n26168), .Z(n26165) );
  XNOR U26652 ( .A(n26169), .B(n26170), .Z(n25072) );
  XNOR U26653 ( .A(n26173), .B(n26174), .Z(n24718) );
  NOR U26654 ( .A(n26175), .B(n26176), .Z(n26173) );
  XOR U26655 ( .A(n22665), .B(n26177), .Z(n26145) );
  XOR U26656 ( .A(n19949), .B(n15947), .Z(n26177) );
  XNOR U26657 ( .A(n26178), .B(n21789), .Z(n15947) );
  XOR U26658 ( .A(n26179), .B(n26180), .Z(n21789) );
  NOR U26659 ( .A(n21522), .B(n21523), .Z(n26178) );
  XOR U26660 ( .A(n21718), .B(n26181), .Z(n21522) );
  XOR U26661 ( .A(n26182), .B(n21783), .Z(n19949) );
  XNOR U26662 ( .A(n26183), .B(n23429), .Z(n21783) );
  ANDN U26663 ( .B(n23082), .A(n23083), .Z(n26182) );
  XOR U26664 ( .A(n26184), .B(n22325), .Z(n23082) );
  XNOR U26665 ( .A(n26185), .B(n21779), .Z(n22665) );
  XNOR U26666 ( .A(n23489), .B(n26186), .Z(n21779) );
  ANDN U26667 ( .B(n21513), .A(n21512), .Z(n26185) );
  XOR U26668 ( .A(n26187), .B(n26188), .Z(n21512) );
  XNOR U26669 ( .A(n26189), .B(n25571), .Z(n21516) );
  XOR U26670 ( .A(n26190), .B(n22960), .Z(n25571) );
  ANDN U26671 ( .B(n26149), .A(n21792), .Z(n26189) );
  NOR U26672 ( .A(n15925), .B(n15923), .Z(n26143) );
  XOR U26673 ( .A(n18286), .B(n20824), .Z(n15923) );
  XNOR U26674 ( .A(n26191), .B(n20782), .Z(n20824) );
  IV U26675 ( .A(n26192), .Z(n20782) );
  NOR U26676 ( .A(n19905), .B(n22388), .Z(n26191) );
  IV U26677 ( .A(n22389), .Z(n19905) );
  XOR U26678 ( .A(n26193), .B(n21584), .Z(n22389) );
  IV U26679 ( .A(n18048), .Z(n18286) );
  XNOR U26680 ( .A(n19707), .B(n18976), .Z(n18048) );
  XNOR U26681 ( .A(n26194), .B(n26195), .Z(n18976) );
  XOR U26682 ( .A(n15185), .B(n20544), .Z(n26195) );
  XOR U26683 ( .A(n26196), .B(n19918), .Z(n20544) );
  XOR U26684 ( .A(n26197), .B(n25382), .Z(n19918) );
  AND U26685 ( .A(n20784), .B(n21002), .Z(n26196) );
  XOR U26686 ( .A(n26198), .B(n25201), .Z(n21002) );
  IV U26687 ( .A(n22949), .Z(n25201) );
  XOR U26688 ( .A(n25813), .B(n26199), .Z(n22949) );
  XOR U26689 ( .A(n26200), .B(n26201), .Z(n25813) );
  XOR U26690 ( .A(n25343), .B(n26202), .Z(n26201) );
  XNOR U26691 ( .A(n26203), .B(n26204), .Z(n25343) );
  ANDN U26692 ( .B(n26205), .A(n26206), .Z(n26203) );
  XOR U26693 ( .A(n25610), .B(n26207), .Z(n26200) );
  XNOR U26694 ( .A(n22634), .B(n26208), .Z(n26207) );
  XNOR U26695 ( .A(n26209), .B(n26210), .Z(n22634) );
  ANDN U26696 ( .B(n26211), .A(n26212), .Z(n26209) );
  XNOR U26697 ( .A(n26213), .B(n26214), .Z(n25610) );
  ANDN U26698 ( .B(n26215), .A(n26216), .Z(n26213) );
  XOR U26699 ( .A(n26217), .B(n24563), .Z(n20784) );
  XOR U26700 ( .A(n26218), .B(n19911), .Z(n15185) );
  XOR U26701 ( .A(n22939), .B(n26219), .Z(n19911) );
  IV U26702 ( .A(n23987), .Z(n22939) );
  XNOR U26703 ( .A(n26220), .B(n26221), .Z(n23987) );
  ANDN U26704 ( .B(n20779), .A(n20832), .Z(n26218) );
  XNOR U26705 ( .A(n26222), .B(n24031), .Z(n20832) );
  XOR U26706 ( .A(n26223), .B(n26224), .Z(n20779) );
  XOR U26707 ( .A(n16526), .B(n26225), .Z(n26194) );
  XOR U26708 ( .A(n17257), .B(n18760), .Z(n26225) );
  XNOR U26709 ( .A(n26226), .B(n20493), .Z(n18760) );
  XNOR U26710 ( .A(n26227), .B(n25085), .Z(n20493) );
  AND U26711 ( .A(n22399), .B(n20777), .Z(n26226) );
  XOR U26712 ( .A(n24344), .B(n26228), .Z(n20777) );
  XOR U26713 ( .A(n23856), .B(n26229), .Z(n22399) );
  IV U26714 ( .A(n24788), .Z(n23856) );
  XNOR U26715 ( .A(n26230), .B(n26231), .Z(n24788) );
  XNOR U26716 ( .A(n26232), .B(n19907), .Z(n17257) );
  XNOR U26717 ( .A(n26233), .B(n23346), .Z(n19907) );
  ANDN U26718 ( .B(n22388), .A(n26192), .Z(n26232) );
  XOR U26719 ( .A(n26234), .B(n23059), .Z(n26192) );
  XNOR U26720 ( .A(n26235), .B(n24247), .Z(n22388) );
  XNOR U26721 ( .A(n26236), .B(n20787), .Z(n16526) );
  XNOR U26722 ( .A(n26237), .B(n26238), .Z(n20787) );
  AND U26723 ( .A(n20788), .B(n20830), .Z(n26236) );
  XOR U26724 ( .A(n26239), .B(n24827), .Z(n20830) );
  XOR U26725 ( .A(n26240), .B(n26028), .Z(n20788) );
  XOR U26726 ( .A(n26241), .B(n26242), .Z(n19707) );
  XNOR U26727 ( .A(n19091), .B(n19644), .Z(n26242) );
  XNOR U26728 ( .A(n26243), .B(n25625), .Z(n19644) );
  IV U26729 ( .A(n22926), .Z(n25625) );
  XNOR U26730 ( .A(n26247), .B(n24150), .Z(n22927) );
  XNOR U26731 ( .A(n26248), .B(n22930), .Z(n19091) );
  XOR U26732 ( .A(n26249), .B(n25757), .Z(n22930) );
  ANDN U26733 ( .B(n23191), .A(n23189), .Z(n26248) );
  IV U26734 ( .A(n22931), .Z(n23189) );
  XOR U26735 ( .A(n24613), .B(n26250), .Z(n22931) );
  XOR U26736 ( .A(n26251), .B(n26252), .Z(n24613) );
  XNOR U26737 ( .A(n19320), .B(n26253), .Z(n26241) );
  XOR U26738 ( .A(n18835), .B(n22910), .Z(n26253) );
  XNOR U26739 ( .A(n26254), .B(n22917), .Z(n22910) );
  XOR U26740 ( .A(n26255), .B(n25596), .Z(n22917) );
  AND U26741 ( .A(n22918), .B(n23194), .Z(n26254) );
  XNOR U26742 ( .A(n26256), .B(n21710), .Z(n22918) );
  IV U26743 ( .A(n26053), .Z(n21710) );
  XNOR U26744 ( .A(n26259), .B(n25623), .Z(n18835) );
  IV U26745 ( .A(n22922), .Z(n25623) );
  XOR U26746 ( .A(n26260), .B(n24795), .Z(n22922) );
  IV U26747 ( .A(n23079), .Z(n24795) );
  ANDN U26748 ( .B(n22923), .A(n23197), .Z(n26259) );
  IV U26749 ( .A(n26261), .Z(n23197) );
  XOR U26750 ( .A(n26262), .B(n24166), .Z(n22923) );
  IV U26751 ( .A(n25252), .Z(n24166) );
  XNOR U26752 ( .A(n26265), .B(n25648), .Z(n19320) );
  ANDN U26753 ( .B(n23200), .A(n23201), .Z(n26265) );
  XNOR U26754 ( .A(n26266), .B(n23829), .Z(n23200) );
  IV U26755 ( .A(n25163), .Z(n23829) );
  XOR U26756 ( .A(n26084), .B(n18806), .Z(n15925) );
  IV U26757 ( .A(n18074), .Z(n18806) );
  XNOR U26758 ( .A(n21335), .B(n20791), .Z(n18074) );
  XNOR U26759 ( .A(n26267), .B(n26268), .Z(n20791) );
  XNOR U26760 ( .A(n18162), .B(n20072), .Z(n26268) );
  XOR U26761 ( .A(n26269), .B(n23680), .Z(n20072) );
  NOR U26762 ( .A(n23681), .B(n23466), .Z(n26269) );
  XOR U26763 ( .A(n26270), .B(n21214), .Z(n23681) );
  IV U26764 ( .A(n25230), .Z(n21214) );
  XNOR U26765 ( .A(n26271), .B(n26272), .Z(n25230) );
  XNOR U26766 ( .A(n26273), .B(n23677), .Z(n18162) );
  XOR U26767 ( .A(n24442), .B(n26274), .Z(n23677) );
  XOR U26768 ( .A(n26275), .B(n25361), .Z(n23452) );
  XOR U26769 ( .A(n21533), .B(n26276), .Z(n26267) );
  XOR U26770 ( .A(n19303), .B(n23663), .Z(n26276) );
  XOR U26771 ( .A(n26277), .B(n25909), .Z(n23663) );
  XOR U26772 ( .A(n23725), .B(n26278), .Z(n25909) );
  XOR U26773 ( .A(n26279), .B(n26280), .Z(n23456) );
  XOR U26774 ( .A(n26281), .B(n23669), .Z(n19303) );
  XOR U26775 ( .A(n24007), .B(n26282), .Z(n23669) );
  IV U26776 ( .A(n23951), .Z(n24007) );
  NOR U26777 ( .A(n23470), .B(n23469), .Z(n26281) );
  XOR U26778 ( .A(n26283), .B(n26284), .Z(n23469) );
  XOR U26779 ( .A(n26285), .B(n23672), .Z(n21533) );
  XNOR U26780 ( .A(n26286), .B(n26287), .Z(n23672) );
  NOR U26781 ( .A(n26288), .B(n23461), .Z(n26285) );
  XNOR U26782 ( .A(n23326), .B(n26289), .Z(n23461) );
  IV U26783 ( .A(n24449), .Z(n23326) );
  XNOR U26784 ( .A(n26290), .B(n26291), .Z(n24449) );
  XOR U26785 ( .A(n26292), .B(n26293), .Z(n21335) );
  XNOR U26786 ( .A(n19146), .B(n18526), .Z(n26293) );
  XOR U26787 ( .A(n26294), .B(n19744), .Z(n18526) );
  XNOR U26788 ( .A(n26179), .B(n26295), .Z(n19744) );
  IV U26789 ( .A(n22511), .Z(n26179) );
  XOR U26790 ( .A(n25580), .B(n25752), .Z(n22511) );
  XNOR U26791 ( .A(n26296), .B(n26297), .Z(n25752) );
  XNOR U26792 ( .A(n25425), .B(n24641), .Z(n26297) );
  XNOR U26793 ( .A(n26298), .B(n26299), .Z(n24641) );
  ANDN U26794 ( .B(n26300), .A(n26301), .Z(n26298) );
  XNOR U26795 ( .A(n26302), .B(n26303), .Z(n25425) );
  NOR U26796 ( .A(n26304), .B(n26305), .Z(n26302) );
  XOR U26797 ( .A(n26306), .B(n26307), .Z(n26296) );
  XNOR U26798 ( .A(n24433), .B(n24572), .Z(n26307) );
  XNOR U26799 ( .A(n26308), .B(n26309), .Z(n24572) );
  NOR U26800 ( .A(n26310), .B(n26311), .Z(n26308) );
  XNOR U26801 ( .A(n26312), .B(n26313), .Z(n24433) );
  NOR U26802 ( .A(n26314), .B(n26315), .Z(n26312) );
  XOR U26803 ( .A(n26316), .B(n26317), .Z(n25580) );
  XNOR U26804 ( .A(n23034), .B(n25442), .Z(n26317) );
  XNOR U26805 ( .A(n26318), .B(n26319), .Z(n25442) );
  ANDN U26806 ( .B(n26320), .A(n26321), .Z(n26318) );
  XNOR U26807 ( .A(n26322), .B(n26323), .Z(n23034) );
  NOR U26808 ( .A(n26324), .B(n26325), .Z(n26322) );
  XOR U26809 ( .A(n24861), .B(n26326), .Z(n26316) );
  XOR U26810 ( .A(n25127), .B(n25708), .Z(n26326) );
  XOR U26811 ( .A(n26327), .B(n26328), .Z(n25708) );
  XOR U26812 ( .A(n26331), .B(n26332), .Z(n25127) );
  NOR U26813 ( .A(n26333), .B(n26334), .Z(n26331) );
  XOR U26814 ( .A(n26335), .B(n26336), .Z(n24861) );
  NOR U26815 ( .A(n26337), .B(n26338), .Z(n26335) );
  ANDN U26816 ( .B(n23446), .A(n19745), .Z(n26294) );
  XOR U26817 ( .A(n26339), .B(n24379), .Z(n19745) );
  XOR U26818 ( .A(n26340), .B(n24453), .Z(n23446) );
  IV U26819 ( .A(n25111), .Z(n24453) );
  XOR U26820 ( .A(n26341), .B(n26342), .Z(n25111) );
  XOR U26821 ( .A(n26343), .B(n19166), .Z(n19146) );
  XNOR U26822 ( .A(n25219), .B(n26344), .Z(n19166) );
  XOR U26823 ( .A(n16528), .B(n26346), .Z(n26292) );
  XOR U26824 ( .A(n16605), .B(n18734), .Z(n26346) );
  XNOR U26825 ( .A(n26347), .B(n19151), .Z(n18734) );
  XNOR U26826 ( .A(n25577), .B(n26348), .Z(n19151) );
  ANDN U26827 ( .B(n19152), .A(n26086), .Z(n26347) );
  XOR U26828 ( .A(n26349), .B(n24566), .Z(n26086) );
  XOR U26829 ( .A(n26272), .B(n26350), .Z(n24566) );
  XNOR U26830 ( .A(n26351), .B(n26352), .Z(n26272) );
  XNOR U26831 ( .A(n25345), .B(n26353), .Z(n26352) );
  XNOR U26832 ( .A(n26354), .B(n26355), .Z(n25345) );
  ANDN U26833 ( .B(n26356), .A(n26357), .Z(n26354) );
  XOR U26834 ( .A(n26358), .B(n26359), .Z(n26351) );
  XOR U26835 ( .A(n25798), .B(n22833), .Z(n26359) );
  XOR U26836 ( .A(n26360), .B(n26361), .Z(n22833) );
  ANDN U26837 ( .B(n26362), .A(n26363), .Z(n26360) );
  XNOR U26838 ( .A(n26364), .B(n26365), .Z(n25798) );
  ANDN U26839 ( .B(n26366), .A(n26367), .Z(n26364) );
  XNOR U26840 ( .A(n26368), .B(n22494), .Z(n19152) );
  IV U26841 ( .A(n23136), .Z(n22494) );
  XNOR U26842 ( .A(n26369), .B(n19161), .Z(n16605) );
  XOR U26843 ( .A(n26370), .B(n25247), .Z(n19161) );
  ANDN U26844 ( .B(n21380), .A(n26076), .Z(n26369) );
  XOR U26845 ( .A(n26371), .B(n24414), .Z(n26076) );
  IV U26846 ( .A(n21227), .Z(n24414) );
  XOR U26847 ( .A(n26372), .B(n26373), .Z(n21227) );
  XOR U26848 ( .A(n26374), .B(n23964), .Z(n21380) );
  XNOR U26849 ( .A(n26375), .B(n19155), .Z(n16528) );
  XOR U26850 ( .A(n26376), .B(n26022), .Z(n19155) );
  XOR U26851 ( .A(n26377), .B(n26378), .Z(n26022) );
  XOR U26852 ( .A(n23712), .B(n26379), .Z(n21370) );
  XOR U26853 ( .A(n25831), .B(n26380), .Z(n19156) );
  IV U26854 ( .A(n26381), .Z(n25831) );
  XNOR U26855 ( .A(n26382), .B(n19165), .Z(n26084) );
  XOR U26856 ( .A(n26383), .B(n23558), .Z(n19165) );
  ANDN U26857 ( .B(n20413), .A(n26345), .Z(n26382) );
  IV U26858 ( .A(n21366), .Z(n26345) );
  XOR U26859 ( .A(n26384), .B(n25373), .Z(n21366) );
  IV U26860 ( .A(n24849), .Z(n25373) );
  XOR U26861 ( .A(n26385), .B(n24960), .Z(n20413) );
  XNOR U26862 ( .A(n26386), .B(n18131), .Z(n18119) );
  XNOR U26863 ( .A(n15962), .B(n25391), .Z(n18131) );
  XNOR U26864 ( .A(n26387), .B(n21869), .Z(n25391) );
  ANDN U26865 ( .B(n24329), .A(n26388), .Z(n26387) );
  XOR U26866 ( .A(n26389), .B(n26390), .Z(n22904) );
  XOR U26867 ( .A(n19651), .B(n17214), .Z(n26390) );
  XNOR U26868 ( .A(n26391), .B(n21878), .Z(n17214) );
  XNOR U26869 ( .A(n26392), .B(n24379), .Z(n21878) );
  NOR U26870 ( .A(n25371), .B(n21484), .Z(n26391) );
  XNOR U26871 ( .A(n26393), .B(n25109), .Z(n21484) );
  XNOR U26872 ( .A(n24702), .B(n26394), .Z(n25371) );
  XNOR U26873 ( .A(n26395), .B(n21882), .Z(n19651) );
  XOR U26874 ( .A(n26396), .B(n24146), .Z(n21882) );
  ANDN U26875 ( .B(n21881), .A(n21489), .Z(n26395) );
  XOR U26876 ( .A(n24621), .B(n26397), .Z(n21489) );
  IV U26877 ( .A(n26092), .Z(n24621) );
  XOR U26878 ( .A(n23703), .B(n26398), .Z(n21881) );
  XOR U26879 ( .A(n19367), .B(n26399), .Z(n26389) );
  XOR U26880 ( .A(n19227), .B(n18244), .Z(n26399) );
  XNOR U26881 ( .A(n26400), .B(n21888), .Z(n18244) );
  XOR U26882 ( .A(n26401), .B(n25757), .Z(n21888) );
  ANDN U26883 ( .B(n21889), .A(n21480), .Z(n26400) );
  XOR U26884 ( .A(n24005), .B(n26402), .Z(n21480) );
  XOR U26885 ( .A(n26403), .B(n25043), .Z(n21889) );
  XNOR U26886 ( .A(n26404), .B(n21886), .Z(n19227) );
  XNOR U26887 ( .A(n26405), .B(n25050), .Z(n21886) );
  AND U26888 ( .A(n21493), .B(n21885), .Z(n26404) );
  XNOR U26889 ( .A(n26406), .B(n22809), .Z(n21885) );
  XOR U26890 ( .A(n26407), .B(n23253), .Z(n21493) );
  XNOR U26891 ( .A(n26410), .B(n21892), .Z(n19367) );
  XNOR U26892 ( .A(n26411), .B(n23429), .Z(n21892) );
  XNOR U26893 ( .A(n26412), .B(n26413), .Z(n23429) );
  ANDN U26894 ( .B(n21891), .A(n21497), .Z(n26410) );
  IV U26895 ( .A(n25380), .Z(n21497) );
  XOR U26896 ( .A(n26414), .B(n23053), .Z(n25380) );
  XOR U26897 ( .A(n24025), .B(n26415), .Z(n21891) );
  XNOR U26898 ( .A(n26416), .B(n26417), .Z(n21461) );
  XNOR U26899 ( .A(n20155), .B(n19089), .Z(n26417) );
  XNOR U26900 ( .A(n26418), .B(n21872), .Z(n19089) );
  XNOR U26901 ( .A(n26419), .B(n24247), .Z(n21872) );
  IV U26902 ( .A(n25501), .Z(n24247) );
  XNOR U26903 ( .A(n26420), .B(n25824), .Z(n25501) );
  XOR U26904 ( .A(n26421), .B(n26422), .Z(n25824) );
  XOR U26905 ( .A(n21213), .B(n22617), .Z(n26422) );
  XOR U26906 ( .A(n26423), .B(n26424), .Z(n22617) );
  NOR U26907 ( .A(n26425), .B(n26426), .Z(n26423) );
  XOR U26908 ( .A(n26427), .B(n26428), .Z(n21213) );
  ANDN U26909 ( .B(n26429), .A(n26430), .Z(n26427) );
  XOR U26910 ( .A(n23845), .B(n26431), .Z(n26421) );
  XNOR U26911 ( .A(n25229), .B(n26270), .Z(n26431) );
  XNOR U26912 ( .A(n26432), .B(n26433), .Z(n26270) );
  NOR U26913 ( .A(n26434), .B(n26435), .Z(n26432) );
  XNOR U26914 ( .A(n26436), .B(n26437), .Z(n25229) );
  ANDN U26915 ( .B(n26438), .A(n26439), .Z(n26436) );
  XNOR U26916 ( .A(n26440), .B(n26441), .Z(n23845) );
  ANDN U26917 ( .B(n26442), .A(n26443), .Z(n26440) );
  ANDN U26918 ( .B(n21873), .A(n25395), .Z(n26418) );
  IV U26919 ( .A(n26444), .Z(n25395) );
  XNOR U26920 ( .A(n26445), .B(n24745), .Z(n21873) );
  XNOR U26921 ( .A(n26446), .B(n21862), .Z(n20155) );
  XNOR U26922 ( .A(n26447), .B(n23053), .Z(n21862) );
  IV U26923 ( .A(n26448), .Z(n23053) );
  AND U26924 ( .A(n21863), .B(n25386), .Z(n26446) );
  XOR U26925 ( .A(n25362), .B(n26449), .Z(n21863) );
  XNOR U26926 ( .A(n21856), .B(n26450), .Z(n26416) );
  XOR U26927 ( .A(n18017), .B(n20904), .Z(n26450) );
  XNOR U26928 ( .A(n26451), .B(n24325), .Z(n20904) );
  XOR U26929 ( .A(n26089), .B(n26452), .Z(n24325) );
  ANDN U26930 ( .B(n24353), .A(n25388), .Z(n26451) );
  IV U26931 ( .A(n26453), .Z(n25388) );
  XOR U26932 ( .A(n26454), .B(n26455), .Z(n24353) );
  XNOR U26933 ( .A(n26456), .B(n22875), .Z(n18017) );
  XOR U26934 ( .A(n26457), .B(n25749), .Z(n22875) );
  IV U26935 ( .A(n23810), .Z(n25749) );
  ANDN U26936 ( .B(n22876), .A(n25393), .Z(n26456) );
  XNOR U26937 ( .A(n24623), .B(n26458), .Z(n22876) );
  XOR U26938 ( .A(n23991), .B(n26460), .Z(n21868) );
  XNOR U26939 ( .A(n26461), .B(n26462), .Z(n23991) );
  ANDN U26940 ( .B(n26388), .A(n21869), .Z(n26459) );
  XNOR U26941 ( .A(n26463), .B(n22982), .Z(n21869) );
  ANDN U26942 ( .B(n15931), .A(n15932), .Z(n26386) );
  XOR U26943 ( .A(n24683), .B(n16032), .Z(n15932) );
  XOR U26944 ( .A(n25292), .B(n18925), .Z(n16032) );
  XNOR U26945 ( .A(n26464), .B(n26465), .Z(n18925) );
  XOR U26946 ( .A(n17973), .B(n20390), .Z(n26465) );
  XNOR U26947 ( .A(n26466), .B(n21617), .Z(n20390) );
  XNOR U26948 ( .A(n26467), .B(n21599), .Z(n21617) );
  XNOR U26949 ( .A(n26468), .B(n26469), .Z(n21599) );
  ANDN U26950 ( .B(n22322), .A(n24808), .Z(n26466) );
  XOR U26951 ( .A(n26470), .B(n26471), .Z(n24808) );
  XOR U26952 ( .A(n26472), .B(n24180), .Z(n22322) );
  IV U26953 ( .A(n24228), .Z(n24180) );
  XOR U26954 ( .A(n26473), .B(n21612), .Z(n17973) );
  XOR U26955 ( .A(n26474), .B(n25350), .Z(n21612) );
  XOR U26956 ( .A(n26475), .B(n22506), .Z(n20588) );
  IV U26957 ( .A(n24812), .Z(n22315) );
  XOR U26958 ( .A(n26476), .B(n25152), .Z(n24812) );
  XOR U26959 ( .A(n19546), .B(n26477), .Z(n26464) );
  XOR U26960 ( .A(n17322), .B(n19080), .Z(n26477) );
  XNOR U26961 ( .A(n26478), .B(n21621), .Z(n19080) );
  XNOR U26962 ( .A(n26479), .B(n25045), .Z(n21621) );
  XOR U26963 ( .A(n21385), .B(n26480), .Z(n22326) );
  XOR U26964 ( .A(n26481), .B(n26017), .Z(n20574) );
  XNOR U26965 ( .A(n26482), .B(n21610), .Z(n17322) );
  XOR U26966 ( .A(n26483), .B(n24582), .Z(n21610) );
  IV U26967 ( .A(n24154), .Z(n24582) );
  XOR U26968 ( .A(n26485), .B(n26486), .Z(n25710) );
  XOR U26969 ( .A(n24564), .B(n23320), .Z(n26486) );
  XNOR U26970 ( .A(n26487), .B(n26488), .Z(n23320) );
  ANDN U26971 ( .B(n26489), .A(n26490), .Z(n26487) );
  XNOR U26972 ( .A(n26491), .B(n26492), .Z(n24564) );
  NOR U26973 ( .A(n26493), .B(n26494), .Z(n26491) );
  XOR U26974 ( .A(n26495), .B(n26496), .Z(n26485) );
  XOR U26975 ( .A(n24380), .B(n26497), .Z(n26496) );
  XNOR U26976 ( .A(n26498), .B(n26499), .Z(n24380) );
  NOR U26977 ( .A(n26500), .B(n26501), .Z(n26498) );
  ANDN U26978 ( .B(n22320), .A(n20584), .Z(n26482) );
  XOR U26979 ( .A(n24904), .B(n26502), .Z(n20584) );
  XNOR U26980 ( .A(n26503), .B(n24846), .Z(n22320) );
  XNOR U26981 ( .A(n26504), .B(n21619), .Z(n19546) );
  XOR U26982 ( .A(n26505), .B(n21221), .Z(n21619) );
  ANDN U26983 ( .B(n22311), .A(n20578), .Z(n26504) );
  XOR U26984 ( .A(n25053), .B(n26509), .Z(n22311) );
  XNOR U26985 ( .A(n26510), .B(n26511), .Z(n25053) );
  XOR U26986 ( .A(n26512), .B(n26513), .Z(n25292) );
  XOR U26987 ( .A(n18220), .B(n19231), .Z(n26513) );
  XNOR U26988 ( .A(n26514), .B(n22293), .Z(n19231) );
  XOR U26989 ( .A(n24936), .B(n26515), .Z(n22293) );
  XOR U26990 ( .A(n23951), .B(n26516), .Z(n22292) );
  XOR U26991 ( .A(n26517), .B(n26518), .Z(n23951) );
  IV U26992 ( .A(n24112), .Z(n24687) );
  XOR U26993 ( .A(n26519), .B(n25152), .Z(n24112) );
  XOR U26994 ( .A(n26520), .B(n22301), .Z(n18220) );
  ANDN U26995 ( .B(n22302), .A(n24105), .Z(n26520) );
  XNOR U26996 ( .A(n26522), .B(n24857), .Z(n24105) );
  XOR U26997 ( .A(n26523), .B(n24272), .Z(n22302) );
  XOR U26998 ( .A(n19045), .B(n26524), .Z(n26512) );
  XOR U26999 ( .A(n22283), .B(n19460), .Z(n26524) );
  XNOR U27000 ( .A(n26525), .B(n22288), .Z(n19460) );
  XNOR U27001 ( .A(n26381), .B(n26526), .Z(n22288) );
  ANDN U27002 ( .B(n22289), .A(n24109), .Z(n26525) );
  IV U27003 ( .A(n26527), .Z(n24109) );
  XNOR U27004 ( .A(n26528), .B(n22305), .Z(n22283) );
  XOR U27005 ( .A(n26529), .B(n22954), .Z(n22305) );
  IV U27006 ( .A(n22500), .Z(n22954) );
  XOR U27007 ( .A(n25980), .B(n26530), .Z(n22500) );
  XOR U27008 ( .A(n26531), .B(n26532), .Z(n25980) );
  XNOR U27009 ( .A(n26533), .B(n26534), .Z(n26532) );
  XNOR U27010 ( .A(n26535), .B(n26536), .Z(n26531) );
  XOR U27011 ( .A(n26537), .B(n26538), .Z(n26536) );
  ANDN U27012 ( .B(n22306), .A(n24102), .Z(n26528) );
  XOR U27013 ( .A(n24904), .B(n26539), .Z(n24102) );
  XOR U27014 ( .A(n26542), .B(n26448), .Z(n22306) );
  XOR U27015 ( .A(n26543), .B(n26544), .Z(n26448) );
  XOR U27016 ( .A(n26545), .B(n22297), .Z(n19045) );
  XOR U27017 ( .A(n26495), .B(n24381), .Z(n22297) );
  IV U27018 ( .A(n23321), .Z(n24381) );
  XNOR U27019 ( .A(n26546), .B(n26547), .Z(n26495) );
  AND U27020 ( .A(n26548), .B(n26549), .Z(n26546) );
  ANDN U27021 ( .B(n24115), .A(n22298), .Z(n26545) );
  XOR U27022 ( .A(n26550), .B(n25008), .Z(n22298) );
  XNOR U27023 ( .A(n26551), .B(n25757), .Z(n24115) );
  XOR U27024 ( .A(n26552), .B(n22289), .Z(n24683) );
  XOR U27025 ( .A(n26553), .B(n25805), .Z(n22289) );
  ANDN U27026 ( .B(n24110), .A(n26527), .Z(n26552) );
  XNOR U27027 ( .A(n26554), .B(n22820), .Z(n26527) );
  XOR U27028 ( .A(n26555), .B(n25177), .Z(n24110) );
  XOR U27029 ( .A(n16727), .B(n24291), .Z(n15931) );
  XOR U27030 ( .A(n26556), .B(n23367), .Z(n24291) );
  ANDN U27031 ( .B(n23871), .A(n23956), .Z(n26556) );
  XNOR U27032 ( .A(n26557), .B(n22412), .Z(n23871) );
  XNOR U27033 ( .A(n26558), .B(n26559), .Z(n24726) );
  XNOR U27034 ( .A(n19491), .B(n20939), .Z(n26559) );
  XNOR U27035 ( .A(n26560), .B(n25650), .Z(n20939) );
  IV U27036 ( .A(n25969), .Z(n25650) );
  XNOR U27037 ( .A(n26561), .B(n23139), .Z(n25969) );
  NOR U27038 ( .A(n24307), .B(n22570), .Z(n26560) );
  XNOR U27039 ( .A(n26562), .B(n24661), .Z(n22570) );
  XOR U27040 ( .A(n24040), .B(n26563), .Z(n24307) );
  IV U27041 ( .A(n23733), .Z(n24040) );
  XOR U27042 ( .A(n26564), .B(n26565), .Z(n23733) );
  XNOR U27043 ( .A(n26566), .B(n23356), .Z(n19491) );
  IV U27044 ( .A(n25978), .Z(n23356) );
  XNOR U27045 ( .A(n26567), .B(n26568), .Z(n25978) );
  ANDN U27046 ( .B(n22557), .A(n23355), .Z(n26566) );
  IV U27047 ( .A(n24738), .Z(n23355) );
  XOR U27048 ( .A(n26569), .B(n26570), .Z(n24738) );
  XOR U27049 ( .A(n26571), .B(n22621), .Z(n22557) );
  XOR U27050 ( .A(n18879), .B(n26572), .Z(n26558) );
  XOR U27051 ( .A(n16840), .B(n16986), .Z(n26572) );
  XNOR U27052 ( .A(n26573), .B(n25988), .Z(n16986) );
  IV U27053 ( .A(n25984), .Z(n25988) );
  XOR U27054 ( .A(n26574), .B(n25673), .Z(n25984) );
  ANDN U27055 ( .B(n22566), .A(n24301), .Z(n26573) );
  XOR U27056 ( .A(n23047), .B(n26575), .Z(n24301) );
  IV U27057 ( .A(n23626), .Z(n23047) );
  XOR U27058 ( .A(n26576), .B(n26577), .Z(n23626) );
  XOR U27059 ( .A(n26578), .B(n24916), .Z(n22566) );
  IV U27060 ( .A(n26579), .Z(n24916) );
  XNOR U27061 ( .A(n26580), .B(n23362), .Z(n16840) );
  XOR U27062 ( .A(n26581), .B(n24408), .Z(n23362) );
  NOR U27063 ( .A(n24304), .B(n23361), .Z(n26580) );
  XOR U27064 ( .A(n26582), .B(n22790), .Z(n23361) );
  IV U27065 ( .A(n22561), .Z(n24304) );
  XOR U27066 ( .A(n26583), .B(n22412), .Z(n22561) );
  IV U27067 ( .A(n25596), .Z(n22412) );
  XOR U27068 ( .A(n26584), .B(n26585), .Z(n25596) );
  XNOR U27069 ( .A(n26586), .B(n23352), .Z(n18879) );
  XOR U27070 ( .A(n24994), .B(n26587), .Z(n23352) );
  XOR U27071 ( .A(n26251), .B(n26588), .Z(n24994) );
  XOR U27072 ( .A(n26589), .B(n26590), .Z(n26251) );
  XOR U27073 ( .A(n26384), .B(n25232), .Z(n26590) );
  XNOR U27074 ( .A(n26591), .B(n26592), .Z(n25232) );
  ANDN U27075 ( .B(n26593), .A(n26594), .Z(n26591) );
  XOR U27076 ( .A(n26595), .B(n26596), .Z(n26384) );
  NOR U27077 ( .A(n26597), .B(n26598), .Z(n26595) );
  XOR U27078 ( .A(n26599), .B(n26600), .Z(n26589) );
  XNOR U27079 ( .A(n24848), .B(n25372), .Z(n26600) );
  XNOR U27080 ( .A(n26601), .B(n26602), .Z(n25372) );
  ANDN U27081 ( .B(n26603), .A(n26604), .Z(n26601) );
  XOR U27082 ( .A(n26605), .B(n26606), .Z(n24848) );
  ANDN U27083 ( .B(n26607), .A(n26608), .Z(n26605) );
  NOR U27084 ( .A(n24310), .B(n22574), .Z(n26586) );
  XOR U27085 ( .A(n26609), .B(n26610), .Z(n22574) );
  IV U27086 ( .A(n23353), .Z(n24310) );
  XOR U27087 ( .A(n23957), .B(n26611), .Z(n23353) );
  XNOR U27088 ( .A(n26612), .B(n26613), .Z(n19983) );
  XNOR U27089 ( .A(n18597), .B(n23348), .Z(n26613) );
  XNOR U27090 ( .A(n26614), .B(n23368), .Z(n23348) );
  XNOR U27091 ( .A(n26615), .B(n23852), .Z(n23368) );
  IV U27092 ( .A(n24420), .Z(n23852) );
  XNOR U27093 ( .A(n26616), .B(n26617), .Z(n24420) );
  ANDN U27094 ( .B(n23956), .A(n23367), .Z(n26614) );
  XOR U27095 ( .A(n26618), .B(n26619), .Z(n23367) );
  XNOR U27096 ( .A(n26535), .B(n26620), .Z(n23956) );
  XNOR U27097 ( .A(n26621), .B(n26622), .Z(n26535) );
  ANDN U27098 ( .B(n26623), .A(n26624), .Z(n26621) );
  XNOR U27099 ( .A(n26625), .B(n23371), .Z(n18597) );
  XOR U27100 ( .A(n23946), .B(n26626), .Z(n23371) );
  NOR U27101 ( .A(n22600), .B(n23370), .Z(n26625) );
  XOR U27102 ( .A(n26627), .B(n24960), .Z(n23370) );
  IV U27103 ( .A(n24570), .Z(n24960) );
  XNOR U27104 ( .A(n26628), .B(n26629), .Z(n24570) );
  XOR U27105 ( .A(n26630), .B(n26631), .Z(n22600) );
  XOR U27106 ( .A(n22582), .B(n26632), .Z(n26612) );
  XNOR U27107 ( .A(n19304), .B(n19952), .Z(n26632) );
  XNOR U27108 ( .A(n26633), .B(n23379), .Z(n19952) );
  IV U27109 ( .A(n23876), .Z(n23379) );
  XOR U27110 ( .A(n26634), .B(n24842), .Z(n23876) );
  NOR U27111 ( .A(n23378), .B(n22590), .Z(n26633) );
  XNOR U27112 ( .A(n23998), .B(n26635), .Z(n22590) );
  XOR U27113 ( .A(n26636), .B(n25278), .Z(n23378) );
  XNOR U27114 ( .A(n26637), .B(n23374), .Z(n19304) );
  XOR U27115 ( .A(n26638), .B(n26639), .Z(n23374) );
  XOR U27116 ( .A(n26640), .B(n24035), .Z(n22596) );
  XNOR U27117 ( .A(n26641), .B(n23708), .Z(n23375) );
  XNOR U27118 ( .A(n26642), .B(n23382), .Z(n22582) );
  XOR U27119 ( .A(n25603), .B(n26643), .Z(n23382) );
  ANDN U27120 ( .B(n24286), .A(n23383), .Z(n26642) );
  XOR U27121 ( .A(n26092), .B(n26644), .Z(n23383) );
  XOR U27122 ( .A(n25132), .B(n26645), .Z(n26092) );
  XNOR U27123 ( .A(n26646), .B(n26647), .Z(n25132) );
  XOR U27124 ( .A(n23018), .B(n25941), .Z(n26647) );
  XNOR U27125 ( .A(n26648), .B(n26649), .Z(n25941) );
  NOR U27126 ( .A(n26650), .B(n26651), .Z(n26648) );
  XNOR U27127 ( .A(n26652), .B(n26653), .Z(n23018) );
  ANDN U27128 ( .B(n26654), .A(n26655), .Z(n26652) );
  XOR U27129 ( .A(n26656), .B(n26657), .Z(n26646) );
  XOR U27130 ( .A(n26658), .B(n26064), .Z(n26657) );
  XNOR U27131 ( .A(n26659), .B(n26660), .Z(n26064) );
  ANDN U27132 ( .B(n26661), .A(n26662), .Z(n26659) );
  XNOR U27133 ( .A(n26663), .B(n23510), .Z(n24286) );
  XOR U27134 ( .A(n26664), .B(n26665), .Z(n15046) );
  XOR U27135 ( .A(n13269), .B(n14043), .Z(n26665) );
  XNOR U27136 ( .A(n26666), .B(n14728), .Z(n14043) );
  XOR U27137 ( .A(n25608), .B(n16058), .Z(n14728) );
  XOR U27138 ( .A(n21395), .B(n18936), .Z(n16058) );
  XNOR U27139 ( .A(n26667), .B(n26668), .Z(n18936) );
  XOR U27140 ( .A(n20961), .B(n20092), .Z(n26668) );
  XNOR U27141 ( .A(n26669), .B(n20980), .Z(n20092) );
  XOR U27142 ( .A(n26670), .B(n24172), .Z(n20980) );
  IV U27143 ( .A(n26631), .Z(n24172) );
  XOR U27144 ( .A(n26671), .B(n25263), .Z(n26631) );
  XNOR U27145 ( .A(n26672), .B(n26673), .Z(n25263) );
  XOR U27146 ( .A(n26674), .B(n23715), .Z(n26673) );
  XNOR U27147 ( .A(n26675), .B(n26676), .Z(n23715) );
  XNOR U27148 ( .A(n22319), .B(n26679), .Z(n26672) );
  XNOR U27149 ( .A(n24066), .B(n26680), .Z(n26679) );
  XNOR U27150 ( .A(n26681), .B(n26682), .Z(n24066) );
  ANDN U27151 ( .B(n26683), .A(n26684), .Z(n26681) );
  XOR U27152 ( .A(n26685), .B(n26686), .Z(n22319) );
  AND U27153 ( .A(n26687), .B(n26688), .Z(n26685) );
  ANDN U27154 ( .B(n20647), .A(n20981), .Z(n26669) );
  XOR U27155 ( .A(n26689), .B(n23079), .Z(n20981) );
  XNOR U27156 ( .A(n26690), .B(n23710), .Z(n20647) );
  XNOR U27157 ( .A(n26691), .B(n20970), .Z(n20961) );
  XOR U27158 ( .A(n26692), .B(n23436), .Z(n20970) );
  NOR U27159 ( .A(n20655), .B(n20656), .Z(n26691) );
  XNOR U27160 ( .A(n26695), .B(n23751), .Z(n20656) );
  IV U27161 ( .A(n26028), .Z(n23751) );
  XOR U27162 ( .A(n26696), .B(n25839), .Z(n20655) );
  XOR U27163 ( .A(n17410), .B(n26697), .Z(n26667) );
  XOR U27164 ( .A(n16604), .B(n18322), .Z(n26697) );
  XNOR U27165 ( .A(n26698), .B(n20974), .Z(n18322) );
  XOR U27166 ( .A(n26699), .B(n23065), .Z(n20974) );
  NOR U27167 ( .A(n20642), .B(n20643), .Z(n26698) );
  XNOR U27168 ( .A(n25488), .B(n26700), .Z(n20643) );
  XNOR U27169 ( .A(n26701), .B(n25673), .Z(n20642) );
  XNOR U27170 ( .A(n26702), .B(n26703), .Z(n25673) );
  XNOR U27171 ( .A(n26704), .B(n20967), .Z(n16604) );
  XNOR U27172 ( .A(n26705), .B(n22231), .Z(n20967) );
  AND U27173 ( .A(n20651), .B(n20653), .Z(n26704) );
  XOR U27174 ( .A(n24662), .B(n26706), .Z(n20653) );
  XOR U27175 ( .A(n26707), .B(n23825), .Z(n20651) );
  XNOR U27176 ( .A(n26708), .B(n20977), .Z(n17410) );
  XOR U27177 ( .A(n26709), .B(n23974), .Z(n20977) );
  ANDN U27178 ( .B(n20659), .A(n20660), .Z(n26708) );
  XNOR U27179 ( .A(n26710), .B(n22809), .Z(n20660) );
  XOR U27180 ( .A(n26713), .B(n25050), .Z(n20659) );
  XOR U27181 ( .A(n26714), .B(n26715), .Z(n21395) );
  XNOR U27182 ( .A(n20662), .B(n17081), .Z(n26715) );
  XOR U27183 ( .A(n26716), .B(n21317), .Z(n17081) );
  XOR U27184 ( .A(n26717), .B(n26718), .Z(n21317) );
  ANDN U27185 ( .B(n22174), .A(n22610), .Z(n26716) );
  XOR U27186 ( .A(n26497), .B(n23321), .Z(n22610) );
  XNOR U27187 ( .A(n26719), .B(n26720), .Z(n23321) );
  XNOR U27188 ( .A(n26721), .B(n26722), .Z(n26497) );
  ANDN U27189 ( .B(n26723), .A(n26724), .Z(n26721) );
  XOR U27190 ( .A(n26725), .B(n25050), .Z(n22174) );
  XNOR U27191 ( .A(n26726), .B(n26727), .Z(n25050) );
  XNOR U27192 ( .A(n26728), .B(n21322), .Z(n20662) );
  XOR U27193 ( .A(n24629), .B(n26729), .Z(n21322) );
  IV U27194 ( .A(n24605), .Z(n24629) );
  XOR U27195 ( .A(n25116), .B(n26730), .Z(n24605) );
  XOR U27196 ( .A(n26731), .B(n26732), .Z(n25116) );
  XNOR U27197 ( .A(n26733), .B(n26237), .Z(n26732) );
  XOR U27198 ( .A(n26734), .B(n26735), .Z(n26237) );
  XNOR U27199 ( .A(n26738), .B(n26739), .Z(n26731) );
  XOR U27200 ( .A(n24968), .B(n22987), .Z(n26739) );
  XOR U27201 ( .A(n26740), .B(n26741), .Z(n22987) );
  ANDN U27202 ( .B(n26742), .A(n26743), .Z(n26740) );
  XNOR U27203 ( .A(n26744), .B(n26745), .Z(n24968) );
  AND U27204 ( .A(n22622), .B(n22180), .Z(n26728) );
  XOR U27205 ( .A(n26748), .B(n26749), .Z(n22180) );
  XOR U27206 ( .A(n26750), .B(n22008), .Z(n22622) );
  XNOR U27207 ( .A(n16758), .B(n26751), .Z(n26714) );
  XNOR U27208 ( .A(n18206), .B(n17460), .Z(n26751) );
  XOR U27209 ( .A(n26752), .B(n22183), .Z(n17460) );
  XOR U27210 ( .A(n26753), .B(n25952), .Z(n22183) );
  ANDN U27211 ( .B(n22614), .A(n22176), .Z(n26752) );
  XOR U27212 ( .A(n26754), .B(n26028), .Z(n22176) );
  XOR U27213 ( .A(n26755), .B(n26756), .Z(n26028) );
  XOR U27214 ( .A(n26757), .B(n24989), .Z(n22614) );
  XNOR U27215 ( .A(n26758), .B(n21308), .Z(n18206) );
  XOR U27216 ( .A(n25476), .B(n26759), .Z(n21308) );
  ANDN U27217 ( .B(n22618), .A(n22170), .Z(n26758) );
  XNOR U27218 ( .A(n26760), .B(n21312), .Z(n16758) );
  XOR U27219 ( .A(n26761), .B(n22404), .Z(n21312) );
  NOR U27220 ( .A(n25612), .B(n22168), .Z(n26760) );
  XNOR U27221 ( .A(n26762), .B(n23864), .Z(n22168) );
  IV U27222 ( .A(n22626), .Z(n25612) );
  XOR U27223 ( .A(n26765), .B(n25206), .Z(n22626) );
  XNOR U27224 ( .A(n26766), .B(n22618), .Z(n25608) );
  XOR U27225 ( .A(n26767), .B(n23710), .Z(n22618) );
  XNOR U27226 ( .A(n26768), .B(n26769), .Z(n23710) );
  AND U27227 ( .A(n22170), .B(n21306), .Z(n26766) );
  XOR U27228 ( .A(n26770), .B(n24035), .Z(n21306) );
  XOR U27229 ( .A(n26771), .B(n26772), .Z(n24035) );
  XNOR U27230 ( .A(n26454), .B(n26773), .Z(n22170) );
  ANDN U27231 ( .B(n14727), .A(n16726), .Z(n26666) );
  XOR U27232 ( .A(n21998), .B(n16852), .Z(n16726) );
  IV U27233 ( .A(n17470), .Z(n16852) );
  XNOR U27234 ( .A(n21115), .B(n22785), .Z(n17470) );
  XNOR U27235 ( .A(n26774), .B(n26775), .Z(n22785) );
  XNOR U27236 ( .A(n15527), .B(n17044), .Z(n26775) );
  XNOR U27237 ( .A(n26776), .B(n21902), .Z(n17044) );
  XOR U27238 ( .A(n23703), .B(n26777), .Z(n21902) );
  IV U27239 ( .A(n25761), .Z(n23703) );
  XOR U27240 ( .A(n26778), .B(n26779), .Z(n25761) );
  ANDN U27241 ( .B(n21180), .A(n21903), .Z(n26776) );
  XOR U27242 ( .A(n26780), .B(n23072), .Z(n21903) );
  IV U27243 ( .A(n25940), .Z(n23072) );
  XOR U27244 ( .A(n26781), .B(n26782), .Z(n25940) );
  XNOR U27245 ( .A(n26783), .B(n26784), .Z(n21180) );
  XNOR U27246 ( .A(n26785), .B(n21027), .Z(n15527) );
  XNOR U27247 ( .A(n26786), .B(n24499), .Z(n21027) );
  IV U27248 ( .A(n26787), .Z(n24499) );
  ANDN U27249 ( .B(n21173), .A(n21026), .Z(n26785) );
  XNOR U27250 ( .A(n20306), .B(n26788), .Z(n26774) );
  XNOR U27251 ( .A(n18375), .B(n19502), .Z(n26788) );
  XNOR U27252 ( .A(n26789), .B(n21032), .Z(n19502) );
  XNOR U27253 ( .A(n26790), .B(n23015), .Z(n21032) );
  ANDN U27254 ( .B(n21033), .A(n21169), .Z(n26789) );
  XNOR U27255 ( .A(n26793), .B(n24423), .Z(n21169) );
  XNOR U27256 ( .A(n23840), .B(n26794), .Z(n21033) );
  IV U27257 ( .A(n26638), .Z(n23840) );
  XNOR U27258 ( .A(n26118), .B(n26795), .Z(n26638) );
  XOR U27259 ( .A(n26796), .B(n26797), .Z(n26118) );
  XNOR U27260 ( .A(n24997), .B(n26798), .Z(n26797) );
  XNOR U27261 ( .A(n26799), .B(n26800), .Z(n24997) );
  ANDN U27262 ( .B(n26801), .A(n26802), .Z(n26799) );
  XOR U27263 ( .A(n26803), .B(n26804), .Z(n26796) );
  XOR U27264 ( .A(n25760), .B(n26805), .Z(n26804) );
  XOR U27265 ( .A(n26806), .B(n26807), .Z(n25760) );
  NOR U27266 ( .A(n26808), .B(n26809), .Z(n26806) );
  XNOR U27267 ( .A(n26810), .B(n25010), .Z(n18375) );
  XOR U27268 ( .A(n26811), .B(n23510), .Z(n25010) );
  XOR U27269 ( .A(n26812), .B(n26813), .Z(n23510) );
  ANDN U27270 ( .B(n21165), .A(n22000), .Z(n26810) );
  IV U27271 ( .A(n25011), .Z(n22000) );
  XOR U27272 ( .A(n24626), .B(n26814), .Z(n25011) );
  XNOR U27273 ( .A(n26815), .B(n26816), .Z(n24626) );
  XOR U27274 ( .A(n26817), .B(n25144), .Z(n21165) );
  XOR U27275 ( .A(n26818), .B(n21036), .Z(n20306) );
  IV U27276 ( .A(n25024), .Z(n21036) );
  XNOR U27277 ( .A(n26819), .B(n24558), .Z(n25024) );
  XOR U27278 ( .A(n24005), .B(n26820), .Z(n21177) );
  XOR U27279 ( .A(n26821), .B(n25727), .Z(n24005) );
  XOR U27280 ( .A(n26822), .B(n26823), .Z(n25727) );
  XNOR U27281 ( .A(n25654), .B(n26824), .Z(n26823) );
  XOR U27282 ( .A(n26825), .B(n26826), .Z(n25654) );
  ANDN U27283 ( .B(n26827), .A(n26828), .Z(n26825) );
  XOR U27284 ( .A(n26829), .B(n26830), .Z(n26822) );
  XOR U27285 ( .A(n26831), .B(n23868), .Z(n26830) );
  XNOR U27286 ( .A(n26832), .B(n26833), .Z(n23868) );
  ANDN U27287 ( .B(n26834), .A(n26835), .Z(n26832) );
  XOR U27288 ( .A(n26836), .B(n23439), .Z(n21037) );
  IV U27289 ( .A(n21725), .Z(n23439) );
  XOR U27290 ( .A(n26837), .B(n26838), .Z(n21115) );
  XOR U27291 ( .A(n19420), .B(n19330), .Z(n26838) );
  XNOR U27292 ( .A(n26839), .B(n20313), .Z(n19330) );
  XOR U27293 ( .A(n26840), .B(n26787), .Z(n20313) );
  XOR U27294 ( .A(n26841), .B(n26484), .Z(n26787) );
  XNOR U27295 ( .A(n26842), .B(n26843), .Z(n26484) );
  XNOR U27296 ( .A(n25591), .B(n26844), .Z(n26843) );
  XNOR U27297 ( .A(n26845), .B(n25851), .Z(n25591) );
  XOR U27298 ( .A(n25273), .B(n26848), .Z(n26842) );
  XNOR U27299 ( .A(n23694), .B(n24248), .Z(n26848) );
  XNOR U27300 ( .A(n26849), .B(n25858), .Z(n24248) );
  IV U27301 ( .A(n26850), .Z(n25858) );
  AND U27302 ( .A(n26851), .B(n26852), .Z(n26849) );
  XNOR U27303 ( .A(n26853), .B(n25861), .Z(n23694) );
  ANDN U27304 ( .B(n26854), .A(n26855), .Z(n26853) );
  XNOR U27305 ( .A(n26856), .B(n26857), .Z(n25273) );
  ANDN U27306 ( .B(n26858), .A(n26859), .Z(n26856) );
  ANDN U27307 ( .B(n19342), .A(n19340), .Z(n26839) );
  XOR U27308 ( .A(n22648), .B(n26860), .Z(n19340) );
  IV U27309 ( .A(n23586), .Z(n22648) );
  XNOR U27310 ( .A(n24344), .B(n26861), .Z(n19342) );
  XNOR U27311 ( .A(n26862), .B(n26863), .Z(n24344) );
  XOR U27312 ( .A(n26864), .B(n20319), .Z(n19420) );
  XNOR U27313 ( .A(n26865), .B(n23914), .Z(n20319) );
  AND U27314 ( .A(n19345), .B(n19344), .Z(n26864) );
  XNOR U27315 ( .A(n26868), .B(n25356), .Z(n19344) );
  XOR U27316 ( .A(n26869), .B(n26017), .Z(n19345) );
  XOR U27317 ( .A(n16093), .B(n26870), .Z(n26837) );
  XNOR U27318 ( .A(n17784), .B(n17480), .Z(n26870) );
  XOR U27319 ( .A(n26871), .B(n20985), .Z(n17480) );
  XOR U27320 ( .A(n26872), .B(n25352), .Z(n20985) );
  ANDN U27321 ( .B(n21134), .A(n20984), .Z(n26871) );
  XOR U27322 ( .A(n26010), .B(n26873), .Z(n20984) );
  XOR U27323 ( .A(n23074), .B(n26874), .Z(n21134) );
  XNOR U27324 ( .A(n26875), .B(n25900), .Z(n17784) );
  IV U27325 ( .A(n25892), .Z(n25900) );
  XOR U27326 ( .A(n26876), .B(n24374), .Z(n25892) );
  AND U27327 ( .A(n19351), .B(n19350), .Z(n26875) );
  XNOR U27328 ( .A(n26877), .B(n23792), .Z(n19350) );
  IV U27329 ( .A(n25204), .Z(n23792) );
  XNOR U27330 ( .A(n26878), .B(n24943), .Z(n19351) );
  XNOR U27331 ( .A(n26881), .B(n25895), .Z(n16093) );
  IV U27332 ( .A(n24013), .Z(n25895) );
  XNOR U27333 ( .A(n26882), .B(n22227), .Z(n24013) );
  XNOR U27334 ( .A(n26230), .B(n26883), .Z(n22227) );
  XOR U27335 ( .A(n26884), .B(n26885), .Z(n26230) );
  XOR U27336 ( .A(n24915), .B(n26886), .Z(n26885) );
  XNOR U27337 ( .A(n26887), .B(n26888), .Z(n24915) );
  AND U27338 ( .A(n26889), .B(n26890), .Z(n26887) );
  XOR U27339 ( .A(n25281), .B(n26891), .Z(n26884) );
  XOR U27340 ( .A(n26037), .B(n26578), .Z(n26891) );
  XNOR U27341 ( .A(n26892), .B(n26893), .Z(n26578) );
  ANDN U27342 ( .B(n26894), .A(n26895), .Z(n26892) );
  XNOR U27343 ( .A(n26896), .B(n26897), .Z(n26037) );
  ANDN U27344 ( .B(n26898), .A(n26899), .Z(n26896) );
  XNOR U27345 ( .A(n26900), .B(n26901), .Z(n25281) );
  AND U27346 ( .A(n19355), .B(n19354), .Z(n26881) );
  XNOR U27347 ( .A(n26904), .B(n26905), .Z(n19354) );
  XNOR U27348 ( .A(n26906), .B(n26907), .Z(n19355) );
  XOR U27349 ( .A(n26908), .B(n21026), .Z(n21998) );
  XOR U27350 ( .A(n24936), .B(n26909), .Z(n21026) );
  IV U27351 ( .A(n22631), .Z(n24936) );
  XOR U27352 ( .A(n26910), .B(n26911), .Z(n22631) );
  NOR U27353 ( .A(n21173), .B(n21174), .Z(n26908) );
  XNOR U27354 ( .A(n26912), .B(n22012), .Z(n21174) );
  IV U27355 ( .A(n26913), .Z(n22012) );
  XOR U27356 ( .A(n26914), .B(n21216), .Z(n21173) );
  XNOR U27357 ( .A(n22438), .B(n19451), .Z(n14727) );
  XOR U27358 ( .A(n23042), .B(n23342), .Z(n19451) );
  XNOR U27359 ( .A(n26915), .B(n26916), .Z(n23342) );
  XNOR U27360 ( .A(n19322), .B(n19669), .Z(n26916) );
  XOR U27361 ( .A(n26917), .B(n21988), .Z(n19669) );
  XNOR U27362 ( .A(n26918), .B(n25043), .Z(n21988) );
  XOR U27363 ( .A(n25183), .B(n26919), .Z(n23344) );
  XNOR U27364 ( .A(n26920), .B(n26078), .Z(n22802) );
  XNOR U27365 ( .A(n26921), .B(n21980), .Z(n19322) );
  XNOR U27366 ( .A(n26568), .B(n26922), .Z(n21980) );
  ANDN U27367 ( .B(n21020), .A(n21018), .Z(n26921) );
  XOR U27368 ( .A(n26923), .B(n24231), .Z(n21018) );
  XOR U27369 ( .A(n26924), .B(n26925), .Z(n21020) );
  XOR U27370 ( .A(n16832), .B(n26926), .Z(n26915) );
  XOR U27371 ( .A(n19058), .B(n16501), .Z(n26926) );
  XOR U27372 ( .A(n26927), .B(n22805), .Z(n16501) );
  XOR U27373 ( .A(n24337), .B(n26928), .Z(n22805) );
  IV U27374 ( .A(n24069), .Z(n24337) );
  XNOR U27375 ( .A(n25131), .B(n26929), .Z(n24069) );
  XOR U27376 ( .A(n26930), .B(n26931), .Z(n25131) );
  XNOR U27377 ( .A(n26932), .B(n26933), .Z(n26931) );
  XNOR U27378 ( .A(n25355), .B(n26934), .Z(n26930) );
  XNOR U27379 ( .A(n26868), .B(n26935), .Z(n26934) );
  XNOR U27380 ( .A(n26936), .B(n26937), .Z(n26868) );
  ANDN U27381 ( .B(n26938), .A(n26939), .Z(n26936) );
  XOR U27382 ( .A(n26940), .B(n26941), .Z(n25355) );
  ANDN U27383 ( .B(n26942), .A(n26943), .Z(n26940) );
  NOR U27384 ( .A(n22798), .B(n23038), .Z(n26927) );
  XNOR U27385 ( .A(n26353), .B(n22834), .Z(n23038) );
  IV U27386 ( .A(n26944), .Z(n22834) );
  XNOR U27387 ( .A(n26945), .B(n26946), .Z(n26353) );
  NOR U27388 ( .A(n26947), .B(n26948), .Z(n26945) );
  XOR U27389 ( .A(n26949), .B(n23815), .Z(n22798) );
  XNOR U27390 ( .A(n26951), .B(n24558), .Z(n21992) );
  XNOR U27391 ( .A(n26221), .B(n26952), .Z(n24558) );
  XOR U27392 ( .A(n26953), .B(n26954), .Z(n26221) );
  XOR U27393 ( .A(n25304), .B(n26955), .Z(n26954) );
  XNOR U27394 ( .A(n26956), .B(n26957), .Z(n25304) );
  NOR U27395 ( .A(n26958), .B(n26959), .Z(n26956) );
  XNOR U27396 ( .A(n22950), .B(n26960), .Z(n26953) );
  XNOR U27397 ( .A(n25837), .B(n25817), .Z(n26960) );
  XOR U27398 ( .A(n26961), .B(n26962), .Z(n25817) );
  NOR U27399 ( .A(n26963), .B(n26964), .Z(n26961) );
  XNOR U27400 ( .A(n26965), .B(n26966), .Z(n25837) );
  ANDN U27401 ( .B(n26967), .A(n26968), .Z(n26965) );
  XOR U27402 ( .A(n26969), .B(n26970), .Z(n22950) );
  ANDN U27403 ( .B(n26971), .A(n26972), .Z(n26969) );
  ANDN U27404 ( .B(n25471), .A(n21008), .Z(n26950) );
  XOR U27405 ( .A(n26973), .B(n26059), .Z(n21008) );
  IV U27406 ( .A(n21007), .Z(n25471) );
  XOR U27407 ( .A(n26974), .B(n26975), .Z(n21007) );
  XNOR U27408 ( .A(n26976), .B(n21982), .Z(n16832) );
  XNOR U27409 ( .A(n26977), .B(n23582), .Z(n21982) );
  ANDN U27410 ( .B(n21013), .A(n21011), .Z(n26976) );
  XOR U27411 ( .A(n26978), .B(n26287), .Z(n21011) );
  IV U27412 ( .A(n22025), .Z(n26287) );
  XOR U27413 ( .A(n26979), .B(n26980), .Z(n22025) );
  XNOR U27414 ( .A(n26981), .B(n22960), .Z(n21013) );
  XNOR U27415 ( .A(n26982), .B(n26983), .Z(n23042) );
  XOR U27416 ( .A(n22207), .B(n20628), .Z(n26983) );
  XOR U27417 ( .A(n26984), .B(n20925), .Z(n20628) );
  XOR U27418 ( .A(n26985), .B(n23150), .Z(n20925) );
  IV U27419 ( .A(n24577), .Z(n23150) );
  XNOR U27420 ( .A(n26986), .B(n26987), .Z(n24577) );
  ANDN U27421 ( .B(n22433), .A(n22431), .Z(n26984) );
  XOR U27422 ( .A(n23422), .B(n25525), .Z(n22431) );
  XOR U27423 ( .A(n26988), .B(n26989), .Z(n25525) );
  ANDN U27424 ( .B(n26990), .A(n26991), .Z(n26988) );
  XNOR U27425 ( .A(n26534), .B(n26620), .Z(n22433) );
  XOR U27426 ( .A(n26992), .B(n26993), .Z(n26534) );
  NOR U27427 ( .A(n26994), .B(n26995), .Z(n26992) );
  XNOR U27428 ( .A(n26996), .B(n20920), .Z(n22207) );
  XNOR U27429 ( .A(n26997), .B(n24438), .Z(n20920) );
  NOR U27430 ( .A(n26998), .B(n25458), .Z(n26996) );
  XOR U27431 ( .A(n19756), .B(n26999), .Z(n26982) );
  XOR U27432 ( .A(n22583), .B(n25444), .Z(n26999) );
  XNOR U27433 ( .A(n27000), .B(n20933), .Z(n25444) );
  XOR U27434 ( .A(n27001), .B(n24231), .Z(n20933) );
  ANDN U27435 ( .B(n22443), .A(n22444), .Z(n27000) );
  XOR U27436 ( .A(n26935), .B(n27002), .Z(n22444) );
  XNOR U27437 ( .A(n27003), .B(n27004), .Z(n26935) );
  ANDN U27438 ( .B(n27005), .A(n27006), .Z(n27003) );
  XOR U27439 ( .A(n27007), .B(n22506), .Z(n22443) );
  XNOR U27440 ( .A(n27008), .B(n20929), .Z(n22583) );
  XOR U27441 ( .A(n27009), .B(n25839), .Z(n20929) );
  ANDN U27442 ( .B(n22436), .A(n22435), .Z(n27008) );
  XOR U27443 ( .A(n27010), .B(n26975), .Z(n22435) );
  IV U27444 ( .A(n22524), .Z(n22436) );
  XNOR U27445 ( .A(n27011), .B(n24745), .Z(n22524) );
  XNOR U27446 ( .A(n27012), .B(n27013), .Z(n26377) );
  XNOR U27447 ( .A(n27014), .B(n21585), .Z(n27013) );
  XNOR U27448 ( .A(n27015), .B(n26942), .Z(n21585) );
  ANDN U27449 ( .B(n27016), .A(n27017), .Z(n27015) );
  XOR U27450 ( .A(n25005), .B(n27018), .Z(n27012) );
  XNOR U27451 ( .A(n22016), .B(n23758), .Z(n27018) );
  XNOR U27452 ( .A(n27019), .B(n27020), .Z(n23758) );
  ANDN U27453 ( .B(n27021), .A(n27022), .Z(n27019) );
  XNOR U27454 ( .A(n27023), .B(n27024), .Z(n22016) );
  AND U27455 ( .A(n27025), .B(n27026), .Z(n27023) );
  XNOR U27456 ( .A(n27027), .B(n27028), .Z(n25005) );
  ANDN U27457 ( .B(n27029), .A(n27030), .Z(n27027) );
  XNOR U27458 ( .A(n27032), .B(n20915), .Z(n19756) );
  XNOR U27459 ( .A(n27033), .B(n24296), .Z(n20915) );
  ANDN U27460 ( .B(n22440), .A(n22528), .Z(n27032) );
  IV U27461 ( .A(n22441), .Z(n22528) );
  XOR U27462 ( .A(n27034), .B(n25686), .Z(n22441) );
  XOR U27463 ( .A(n27035), .B(n25981), .Z(n25686) );
  XNOR U27464 ( .A(n27036), .B(n27037), .Z(n25981) );
  XNOR U27465 ( .A(n24360), .B(n27038), .Z(n27037) );
  XOR U27466 ( .A(n27039), .B(n26958), .Z(n24360) );
  NOR U27467 ( .A(n27040), .B(n27041), .Z(n27039) );
  XOR U27468 ( .A(n27042), .B(n27043), .Z(n27036) );
  XOR U27469 ( .A(n25705), .B(n24348), .Z(n27043) );
  XOR U27470 ( .A(n27044), .B(n26963), .Z(n24348) );
  NOR U27471 ( .A(n27045), .B(n27046), .Z(n27044) );
  XNOR U27472 ( .A(n27047), .B(n26967), .Z(n25705) );
  ANDN U27473 ( .B(n27048), .A(n27049), .Z(n27047) );
  XNOR U27474 ( .A(n27050), .B(n23582), .Z(n22440) );
  XNOR U27475 ( .A(n27051), .B(n27052), .Z(n23582) );
  XOR U27476 ( .A(n27053), .B(n25458), .Z(n22438) );
  XNOR U27477 ( .A(n27054), .B(n27055), .Z(n25458) );
  ANDN U27478 ( .B(n20918), .A(n22531), .Z(n27053) );
  IV U27479 ( .A(n26998), .Z(n22531) );
  XOR U27480 ( .A(n27056), .B(n22504), .Z(n26998) );
  XNOR U27481 ( .A(n27057), .B(n27058), .Z(n22504) );
  XOR U27482 ( .A(n26599), .B(n24849), .Z(n20918) );
  XNOR U27483 ( .A(n27061), .B(n27062), .Z(n26599) );
  ANDN U27484 ( .B(n27063), .A(n27064), .Z(n27061) );
  XOR U27485 ( .A(n27065), .B(n14731), .Z(n13269) );
  XNOR U27486 ( .A(n24705), .B(n17732), .Z(n14731) );
  IV U27487 ( .A(n14168), .Z(n17732) );
  XOR U27488 ( .A(n21390), .B(n21734), .Z(n14168) );
  XNOR U27489 ( .A(n27066), .B(n27067), .Z(n21734) );
  XOR U27490 ( .A(n21535), .B(n18707), .Z(n27067) );
  XNOR U27491 ( .A(n27068), .B(n21542), .Z(n18707) );
  XOR U27492 ( .A(n27069), .B(n24661), .Z(n21542) );
  NOR U27493 ( .A(n20861), .B(n21541), .Z(n27068) );
  XNOR U27494 ( .A(n27072), .B(n23949), .Z(n21535) );
  XOR U27495 ( .A(n27073), .B(n23815), .Z(n23949) );
  XNOR U27496 ( .A(n26005), .B(n27074), .Z(n23815) );
  XNOR U27497 ( .A(n27075), .B(n27076), .Z(n26005) );
  XNOR U27498 ( .A(n27077), .B(n24496), .Z(n27076) );
  XNOR U27499 ( .A(n27078), .B(n27079), .Z(n24496) );
  NOR U27500 ( .A(n27080), .B(n27081), .Z(n27078) );
  XNOR U27501 ( .A(n21230), .B(n27082), .Z(n27075) );
  XNOR U27502 ( .A(n25616), .B(n23485), .Z(n27082) );
  XNOR U27503 ( .A(n27083), .B(n27084), .Z(n23485) );
  NOR U27504 ( .A(n27085), .B(n27086), .Z(n27083) );
  XOR U27505 ( .A(n27087), .B(n27088), .Z(n25616) );
  XOR U27506 ( .A(n27091), .B(n27092), .Z(n21230) );
  ANDN U27507 ( .B(n27093), .A(n27094), .Z(n27091) );
  NOR U27508 ( .A(n23953), .B(n20935), .Z(n27072) );
  XOR U27509 ( .A(n26610), .B(n27095), .Z(n20935) );
  IV U27510 ( .A(n23712), .Z(n26610) );
  XOR U27511 ( .A(n23737), .B(n27096), .Z(n23953) );
  XOR U27512 ( .A(n18741), .B(n27097), .Z(n27066) );
  XOR U27513 ( .A(n19278), .B(n19674), .Z(n27097) );
  XOR U27514 ( .A(n27098), .B(n21550), .Z(n19674) );
  XOR U27515 ( .A(n27099), .B(n21219), .Z(n21550) );
  IV U27516 ( .A(n23821), .Z(n21219) );
  XOR U27517 ( .A(n27100), .B(n27101), .Z(n23821) );
  NOR U27518 ( .A(n21551), .B(n22328), .Z(n27098) );
  XNOR U27519 ( .A(n27102), .B(n24857), .Z(n22328) );
  XNOR U27520 ( .A(n22990), .B(n27103), .Z(n21551) );
  IV U27521 ( .A(n24836), .Z(n22990) );
  XNOR U27522 ( .A(n27104), .B(n21554), .Z(n19278) );
  XNOR U27523 ( .A(n23505), .B(n27105), .Z(n21554) );
  XNOR U27524 ( .A(n27106), .B(n27107), .Z(n26577) );
  XOR U27525 ( .A(n25181), .B(n25481), .Z(n27107) );
  XNOR U27526 ( .A(n27108), .B(n27109), .Z(n25481) );
  NOR U27527 ( .A(n27110), .B(n27111), .Z(n27108) );
  XNOR U27528 ( .A(n27112), .B(n27113), .Z(n25181) );
  ANDN U27529 ( .B(n27114), .A(n27115), .Z(n27112) );
  XOR U27530 ( .A(n27116), .B(n27117), .Z(n27106) );
  XOR U27531 ( .A(n23028), .B(n27118), .Z(n27117) );
  XOR U27532 ( .A(n27119), .B(n27120), .Z(n23028) );
  ANDN U27533 ( .B(n27121), .A(n27122), .Z(n27119) );
  XOR U27534 ( .A(n27123), .B(n27124), .Z(n25825) );
  XOR U27535 ( .A(n24565), .B(n25327), .Z(n27124) );
  XOR U27536 ( .A(n27125), .B(n26356), .Z(n25327) );
  ANDN U27537 ( .B(n26357), .A(n27126), .Z(n27125) );
  XNOR U27538 ( .A(n27127), .B(n26947), .Z(n24565) );
  IV U27539 ( .A(n27128), .Z(n26947) );
  ANDN U27540 ( .B(n26948), .A(n27129), .Z(n27127) );
  XOR U27541 ( .A(n26349), .B(n27130), .Z(n27123) );
  XNOR U27542 ( .A(n25559), .B(n24843), .Z(n27130) );
  XNOR U27543 ( .A(n27131), .B(n26362), .Z(n24843) );
  XOR U27544 ( .A(n27133), .B(n26367), .Z(n25559) );
  IV U27545 ( .A(n27134), .Z(n26367) );
  NOR U27546 ( .A(n27135), .B(n26366), .Z(n27133) );
  XOR U27547 ( .A(n27136), .B(n27137), .Z(n26349) );
  ANDN U27548 ( .B(n27138), .A(n27139), .Z(n27136) );
  NOR U27549 ( .A(n21555), .B(n21274), .Z(n27104) );
  XOR U27550 ( .A(n25164), .B(n27140), .Z(n21274) );
  IV U27551 ( .A(n25448), .Z(n25164) );
  XOR U27552 ( .A(n27141), .B(n25117), .Z(n25448) );
  XNOR U27553 ( .A(n27142), .B(n27143), .Z(n25117) );
  XOR U27554 ( .A(n23861), .B(n27144), .Z(n27143) );
  XNOR U27555 ( .A(n27145), .B(n27146), .Z(n23861) );
  NOR U27556 ( .A(n27147), .B(n27148), .Z(n27145) );
  XOR U27557 ( .A(n23049), .B(n27149), .Z(n27142) );
  XOR U27558 ( .A(n25340), .B(n26099), .Z(n27149) );
  XNOR U27559 ( .A(n27150), .B(n27151), .Z(n26099) );
  ANDN U27560 ( .B(n27152), .A(n27153), .Z(n27150) );
  XNOR U27561 ( .A(n27154), .B(n27155), .Z(n25340) );
  NOR U27562 ( .A(n27156), .B(n27157), .Z(n27154) );
  XOR U27563 ( .A(n27158), .B(n27159), .Z(n23049) );
  AND U27564 ( .A(n27160), .B(n27161), .Z(n27158) );
  XOR U27565 ( .A(n27162), .B(n26975), .Z(n21555) );
  XNOR U27566 ( .A(n27163), .B(n21546), .Z(n18741) );
  XNOR U27567 ( .A(n24971), .B(n27164), .Z(n21546) );
  XOR U27568 ( .A(n27165), .B(n27166), .Z(n24971) );
  NOR U27569 ( .A(n24707), .B(n24693), .Z(n27163) );
  XOR U27570 ( .A(n24633), .B(n27167), .Z(n24693) );
  XOR U27571 ( .A(n27168), .B(n22825), .Z(n24707) );
  XOR U27572 ( .A(n27169), .B(n27170), .Z(n21390) );
  XOR U27573 ( .A(n19795), .B(n15295), .Z(n27170) );
  XOR U27574 ( .A(n27171), .B(n21574), .Z(n15295) );
  XNOR U27575 ( .A(n27172), .B(n27173), .Z(n21574) );
  NOR U27576 ( .A(n24482), .B(n21573), .Z(n27171) );
  XOR U27577 ( .A(n23074), .B(n27174), .Z(n21573) );
  IV U27578 ( .A(n23701), .Z(n23074) );
  XOR U27579 ( .A(n25726), .B(n27175), .Z(n23701) );
  XOR U27580 ( .A(n27176), .B(n27177), .Z(n25726) );
  XOR U27581 ( .A(n23447), .B(n23617), .Z(n27177) );
  XOR U27582 ( .A(n27178), .B(n26902), .Z(n23617) );
  ANDN U27583 ( .B(n27179), .A(n27180), .Z(n27178) );
  XNOR U27584 ( .A(n27181), .B(n27182), .Z(n23447) );
  NOR U27585 ( .A(n27183), .B(n27184), .Z(n27181) );
  XNOR U27586 ( .A(n26256), .B(n27185), .Z(n27176) );
  XOR U27587 ( .A(n26052), .B(n21709), .Z(n27185) );
  XNOR U27588 ( .A(n27186), .B(n26899), .Z(n21709) );
  ANDN U27589 ( .B(n27187), .A(n27188), .Z(n27186) );
  XOR U27590 ( .A(n27189), .B(n26894), .Z(n26052) );
  NOR U27591 ( .A(n27190), .B(n27191), .Z(n27189) );
  XOR U27592 ( .A(n27192), .B(n26890), .Z(n26256) );
  ANDN U27593 ( .B(n27193), .A(n27194), .Z(n27192) );
  XOR U27594 ( .A(n27195), .B(n23442), .Z(n24482) );
  XNOR U27595 ( .A(n27196), .B(n21564), .Z(n19795) );
  XOR U27596 ( .A(n27197), .B(n24761), .Z(n21564) );
  IV U27597 ( .A(n26059), .Z(n24761) );
  XOR U27598 ( .A(n27198), .B(n27199), .Z(n26059) );
  NOR U27599 ( .A(n21565), .B(n24490), .Z(n27196) );
  XOR U27600 ( .A(n27200), .B(n24712), .Z(n24490) );
  IV U27601 ( .A(n25278), .Z(n24712) );
  XOR U27602 ( .A(n27201), .B(n27202), .Z(n25278) );
  XOR U27603 ( .A(n27203), .B(n21721), .Z(n21565) );
  XOR U27604 ( .A(n26291), .B(n27204), .Z(n21721) );
  XOR U27605 ( .A(n27205), .B(n27206), .Z(n26291) );
  XOR U27606 ( .A(n25505), .B(n25712), .Z(n27206) );
  XOR U27607 ( .A(n27207), .B(n27208), .Z(n25712) );
  ANDN U27608 ( .B(n27209), .A(n27210), .Z(n27207) );
  XNOR U27609 ( .A(n27211), .B(n27212), .Z(n25505) );
  ANDN U27610 ( .B(n27213), .A(n27214), .Z(n27211) );
  XOR U27611 ( .A(n25122), .B(n27215), .Z(n27205) );
  XNOR U27612 ( .A(n27216), .B(n23877), .Z(n27215) );
  XNOR U27613 ( .A(n27217), .B(n27218), .Z(n23877) );
  NOR U27614 ( .A(n27219), .B(n27220), .Z(n27217) );
  XNOR U27615 ( .A(n27221), .B(n27222), .Z(n25122) );
  ANDN U27616 ( .B(n27223), .A(n27224), .Z(n27221) );
  XOR U27617 ( .A(n18270), .B(n27225), .Z(n27169) );
  XNOR U27618 ( .A(n15882), .B(n20900), .Z(n27225) );
  XOR U27619 ( .A(n27226), .B(n21561), .Z(n20900) );
  XOR U27620 ( .A(n27227), .B(n27228), .Z(n21561) );
  NOR U27621 ( .A(n21560), .B(n24478), .Z(n27226) );
  XNOR U27622 ( .A(n22318), .B(n26674), .Z(n24478) );
  XNOR U27623 ( .A(n27229), .B(n27230), .Z(n26674) );
  IV U27624 ( .A(n23714), .Z(n22318) );
  XOR U27625 ( .A(n27233), .B(n24518), .Z(n21560) );
  XOR U27626 ( .A(n27234), .B(n21569), .Z(n15882) );
  XNOR U27627 ( .A(n27235), .B(n25255), .Z(n21569) );
  NOR U27628 ( .A(n21570), .B(n24487), .Z(n27234) );
  XOR U27629 ( .A(n27236), .B(n25963), .Z(n24487) );
  XOR U27630 ( .A(n27237), .B(n25766), .Z(n21570) );
  XNOR U27631 ( .A(n27238), .B(n21577), .Z(n18270) );
  XOR U27632 ( .A(n27239), .B(n25204), .Z(n21577) );
  XOR U27633 ( .A(n27240), .B(n26617), .Z(n25204) );
  XNOR U27634 ( .A(n27241), .B(n27242), .Z(n26617) );
  XNOR U27635 ( .A(n27243), .B(n26699), .Z(n27242) );
  XOR U27636 ( .A(n27244), .B(n27245), .Z(n26699) );
  NOR U27637 ( .A(n27246), .B(n26989), .Z(n27244) );
  XOR U27638 ( .A(n24351), .B(n27247), .Z(n27241) );
  XOR U27639 ( .A(n23064), .B(n25606), .Z(n27247) );
  XNOR U27640 ( .A(n27248), .B(n27249), .Z(n25606) );
  ANDN U27641 ( .B(n27250), .A(n27251), .Z(n27248) );
  XNOR U27642 ( .A(n27252), .B(n27253), .Z(n23064) );
  NOR U27643 ( .A(n27254), .B(n27255), .Z(n27252) );
  XOR U27644 ( .A(n27256), .B(n27257), .Z(n24351) );
  ANDN U27645 ( .B(n25533), .A(n27258), .Z(n27256) );
  ANDN U27646 ( .B(n21578), .A(n24475), .Z(n27238) );
  XNOR U27647 ( .A(n27259), .B(n24193), .Z(n24475) );
  XNOR U27648 ( .A(n23946), .B(n27260), .Z(n21578) );
  XNOR U27649 ( .A(n27261), .B(n21541), .Z(n24705) );
  XOR U27650 ( .A(n27262), .B(n26749), .Z(n21541) );
  XOR U27651 ( .A(n27263), .B(n26913), .Z(n20861) );
  XOR U27652 ( .A(n25402), .B(n27264), .Z(n26913) );
  XOR U27653 ( .A(n27265), .B(n27266), .Z(n25402) );
  XNOR U27654 ( .A(n27267), .B(n26773), .Z(n27266) );
  XOR U27655 ( .A(n27268), .B(n27269), .Z(n26773) );
  AND U27656 ( .A(n27270), .B(n27271), .Z(n27268) );
  XOR U27657 ( .A(n26455), .B(n27272), .Z(n27265) );
  XOR U27658 ( .A(n22637), .B(n27273), .Z(n27272) );
  XNOR U27659 ( .A(n27274), .B(n27275), .Z(n22637) );
  NOR U27660 ( .A(n27276), .B(n27277), .Z(n27274) );
  XNOR U27661 ( .A(n27278), .B(n27279), .Z(n26455) );
  NOR U27662 ( .A(n27280), .B(n27281), .Z(n27278) );
  XOR U27663 ( .A(n27282), .B(n23573), .Z(n20863) );
  XNOR U27664 ( .A(n27284), .B(n27285), .Z(n26911) );
  XNOR U27665 ( .A(n25042), .B(n26403), .Z(n27285) );
  XNOR U27666 ( .A(n27286), .B(n27287), .Z(n26403) );
  ANDN U27667 ( .B(n27288), .A(n27289), .Z(n27286) );
  XNOR U27668 ( .A(n27290), .B(n27291), .Z(n25042) );
  AND U27669 ( .A(n27292), .B(n27293), .Z(n27290) );
  XOR U27670 ( .A(n25078), .B(n27294), .Z(n27284) );
  XOR U27671 ( .A(n27295), .B(n26918), .Z(n27294) );
  XNOR U27672 ( .A(n27296), .B(n27297), .Z(n26918) );
  ANDN U27673 ( .B(n27298), .A(n27299), .Z(n27296) );
  XNOR U27674 ( .A(n27300), .B(n27301), .Z(n25078) );
  ANDN U27675 ( .B(n27302), .A(n27303), .Z(n27300) );
  ANDN U27676 ( .B(n13499), .A(n13497), .Z(n27065) );
  XNOR U27677 ( .A(n16390), .B(n22730), .Z(n13497) );
  XNOR U27678 ( .A(n27304), .B(n23659), .Z(n22730) );
  XNOR U27679 ( .A(n24623), .B(n27305), .Z(n23532) );
  XNOR U27680 ( .A(n22281), .B(n24665), .Z(n16390) );
  XNOR U27681 ( .A(n27306), .B(n27307), .Z(n24665) );
  XOR U27682 ( .A(n17176), .B(n22781), .Z(n27307) );
  XOR U27683 ( .A(n27308), .B(n21354), .Z(n22781) );
  XOR U27684 ( .A(n25268), .B(n27309), .Z(n21354) );
  XNOR U27685 ( .A(n26862), .B(n27310), .Z(n25268) );
  XOR U27686 ( .A(n27311), .B(n27312), .Z(n26862) );
  XOR U27687 ( .A(n27313), .B(n27314), .Z(n27312) );
  XOR U27688 ( .A(n25973), .B(n27315), .Z(n27311) );
  XNOR U27689 ( .A(n23824), .B(n26707), .Z(n27315) );
  XNOR U27690 ( .A(n27316), .B(n27317), .Z(n26707) );
  ANDN U27691 ( .B(n27318), .A(n27319), .Z(n27316) );
  XNOR U27692 ( .A(n27320), .B(n27321), .Z(n23824) );
  ANDN U27693 ( .B(n27322), .A(n27323), .Z(n27320) );
  XNOR U27694 ( .A(n27324), .B(n27325), .Z(n25973) );
  NOR U27695 ( .A(n27326), .B(n27327), .Z(n27324) );
  NOR U27696 ( .A(n21343), .B(n23762), .Z(n27308) );
  XOR U27697 ( .A(n23422), .B(n25526), .Z(n23762) );
  XNOR U27698 ( .A(n27328), .B(n27250), .Z(n25526) );
  XOR U27699 ( .A(n26829), .B(n23869), .Z(n21343) );
  XNOR U27700 ( .A(n27331), .B(n27332), .Z(n26829) );
  ANDN U27701 ( .B(n27333), .A(n27334), .Z(n27331) );
  XOR U27702 ( .A(n27335), .B(n23755), .Z(n17176) );
  XOR U27703 ( .A(n27336), .B(n26280), .Z(n23755) );
  NOR U27704 ( .A(n20539), .B(n21831), .Z(n27335) );
  XOR U27705 ( .A(n27337), .B(n27338), .Z(n21831) );
  XOR U27706 ( .A(n24783), .B(n27339), .Z(n20539) );
  XOR U27707 ( .A(n27340), .B(n27341), .Z(n25581) );
  XOR U27708 ( .A(n24581), .B(n25187), .Z(n27341) );
  XOR U27709 ( .A(n27342), .B(n26490), .Z(n25187) );
  NOR U27710 ( .A(n27343), .B(n26489), .Z(n27342) );
  XOR U27711 ( .A(n27344), .B(n26494), .Z(n24581) );
  AND U27712 ( .A(n26493), .B(n27345), .Z(n27344) );
  XNOR U27713 ( .A(n26032), .B(n27346), .Z(n27340) );
  XOR U27714 ( .A(n26483), .B(n24153), .Z(n27346) );
  XOR U27715 ( .A(n27347), .B(n26723), .Z(n24153) );
  ANDN U27716 ( .B(n26724), .A(n27348), .Z(n27347) );
  XNOR U27717 ( .A(n27349), .B(n27350), .Z(n26483) );
  ANDN U27718 ( .B(n26501), .A(n27351), .Z(n27349) );
  XNOR U27719 ( .A(n27352), .B(n26548), .Z(n26032) );
  XNOR U27720 ( .A(n23746), .B(n27355), .Z(n27306) );
  XOR U27721 ( .A(n17219), .B(n16055), .Z(n27355) );
  XNOR U27722 ( .A(n27356), .B(n23752), .Z(n16055) );
  XOR U27723 ( .A(n27357), .B(n22892), .Z(n23752) );
  ANDN U27724 ( .B(n20529), .A(n21821), .Z(n27356) );
  XOR U27725 ( .A(n25239), .B(n27358), .Z(n21821) );
  IV U27726 ( .A(n22213), .Z(n25239) );
  XOR U27727 ( .A(n27359), .B(n25099), .Z(n20529) );
  IV U27728 ( .A(n24926), .Z(n25099) );
  XNOR U27729 ( .A(n27360), .B(n21352), .Z(n17219) );
  IV U27730 ( .A(n23759), .Z(n21352) );
  XNOR U27731 ( .A(n24025), .B(n27361), .Z(n23759) );
  XNOR U27732 ( .A(n25936), .B(n27362), .Z(n24025) );
  XOR U27733 ( .A(n27363), .B(n27364), .Z(n25936) );
  XOR U27734 ( .A(n25789), .B(n26706), .Z(n27364) );
  XNOR U27735 ( .A(n27365), .B(n27366), .Z(n26706) );
  ANDN U27736 ( .B(n27367), .A(n27368), .Z(n27365) );
  XNOR U27737 ( .A(n27369), .B(n27370), .Z(n25789) );
  ANDN U27738 ( .B(n27371), .A(n27372), .Z(n27369) );
  XOR U27739 ( .A(n24663), .B(n27373), .Z(n27363) );
  XNOR U27740 ( .A(n27374), .B(n25556), .Z(n27373) );
  XNOR U27741 ( .A(n27375), .B(n27376), .Z(n25556) );
  ANDN U27742 ( .B(n27377), .A(n27378), .Z(n27375) );
  XNOR U27743 ( .A(n27379), .B(n27380), .Z(n24663) );
  ANDN U27744 ( .B(n27381), .A(n27382), .Z(n27379) );
  ANDN U27745 ( .B(n20535), .A(n21827), .Z(n27360) );
  XOR U27746 ( .A(n27383), .B(n24039), .Z(n21827) );
  IV U27747 ( .A(n22354), .Z(n24039) );
  XNOR U27748 ( .A(n27384), .B(n23024), .Z(n20535) );
  XNOR U27749 ( .A(n27385), .B(n21357), .Z(n23746) );
  XOR U27750 ( .A(n24278), .B(n27386), .Z(n21357) );
  NOR U27751 ( .A(n21817), .B(n20525), .Z(n27385) );
  XNOR U27752 ( .A(n27387), .B(n23077), .Z(n20525) );
  IV U27753 ( .A(n24563), .Z(n23077) );
  XOR U27754 ( .A(n27388), .B(n27059), .Z(n24563) );
  XNOR U27755 ( .A(n27389), .B(n27390), .Z(n27059) );
  XNOR U27756 ( .A(n22609), .B(n27391), .Z(n27390) );
  XNOR U27757 ( .A(n27392), .B(n27393), .Z(n22609) );
  ANDN U27758 ( .B(n27394), .A(n27395), .Z(n27392) );
  XOR U27759 ( .A(n27396), .B(n27397), .Z(n27389) );
  XOR U27760 ( .A(n22646), .B(n22994), .Z(n27397) );
  ANDN U27761 ( .B(n27400), .A(n27401), .Z(n27398) );
  IV U27762 ( .A(n27402), .Z(n27401) );
  XOR U27763 ( .A(n27403), .B(n27404), .Z(n22646) );
  ANDN U27764 ( .B(n27405), .A(n27406), .Z(n27403) );
  IV U27765 ( .A(n23766), .Z(n21817) );
  XOR U27766 ( .A(n27407), .B(n23978), .Z(n23766) );
  XNOR U27767 ( .A(n27409), .B(n27410), .Z(n26199) );
  XNOR U27768 ( .A(n26777), .B(n25762), .Z(n27410) );
  XNOR U27769 ( .A(n27411), .B(n27412), .Z(n25762) );
  NOR U27770 ( .A(n27413), .B(n27414), .Z(n27411) );
  XNOR U27771 ( .A(n27415), .B(n27416), .Z(n26777) );
  ANDN U27772 ( .B(n27417), .A(n27418), .Z(n27415) );
  XNOR U27773 ( .A(n23704), .B(n27419), .Z(n27409) );
  XOR U27774 ( .A(n26133), .B(n26398), .Z(n27419) );
  XOR U27775 ( .A(n27420), .B(n27421), .Z(n26398) );
  NOR U27776 ( .A(n27422), .B(n27423), .Z(n27420) );
  XOR U27777 ( .A(n27424), .B(n27425), .Z(n26133) );
  AND U27778 ( .A(n27426), .B(n27427), .Z(n27424) );
  XNOR U27779 ( .A(n27428), .B(n27429), .Z(n23704) );
  ANDN U27780 ( .B(n27430), .A(n27431), .Z(n27428) );
  XOR U27781 ( .A(n27432), .B(n27433), .Z(n22281) );
  XNOR U27782 ( .A(n19720), .B(n20250), .Z(n27433) );
  XNOR U27783 ( .A(n27434), .B(n23657), .Z(n20250) );
  XOR U27784 ( .A(n23025), .B(n27435), .Z(n23657) );
  IV U27785 ( .A(n22944), .Z(n23025) );
  NOR U27786 ( .A(n22745), .B(n22746), .Z(n27434) );
  XNOR U27787 ( .A(n27436), .B(n27338), .Z(n22746) );
  IV U27788 ( .A(n24275), .Z(n27338) );
  XOR U27789 ( .A(n25219), .B(n27437), .Z(n22745) );
  IV U27790 ( .A(n26470), .Z(n25219) );
  XOR U27791 ( .A(n27283), .B(n27438), .Z(n26470) );
  XNOR U27792 ( .A(n27439), .B(n27440), .Z(n27283) );
  XNOR U27793 ( .A(n26376), .B(n26021), .Z(n27440) );
  XOR U27794 ( .A(n27441), .B(n27016), .Z(n26021) );
  ANDN U27795 ( .B(n27017), .A(n26941), .Z(n27441) );
  XNOR U27796 ( .A(n27442), .B(n27443), .Z(n26376) );
  XOR U27797 ( .A(n25828), .B(n27445), .Z(n27439) );
  XOR U27798 ( .A(n26051), .B(n26041), .Z(n27445) );
  XNOR U27799 ( .A(n27446), .B(n27021), .Z(n26041) );
  XNOR U27800 ( .A(n27448), .B(n27026), .Z(n26051) );
  NOR U27801 ( .A(n27449), .B(n27025), .Z(n27448) );
  XNOR U27802 ( .A(n27450), .B(n27029), .Z(n25828) );
  XOR U27803 ( .A(n27452), .B(n24946), .Z(n23660) );
  NOR U27804 ( .A(n23530), .B(n23659), .Z(n27451) );
  XOR U27805 ( .A(n27453), .B(n25085), .Z(n23659) );
  XOR U27806 ( .A(n25589), .B(n27354), .Z(n25085) );
  XNOR U27807 ( .A(n27454), .B(n27455), .Z(n27354) );
  XOR U27808 ( .A(n24498), .B(n25120), .Z(n27455) );
  XNOR U27809 ( .A(n27456), .B(n26855), .Z(n25120) );
  IV U27810 ( .A(n27457), .Z(n26855) );
  ANDN U27811 ( .B(n25860), .A(n26854), .Z(n27456) );
  XNOR U27812 ( .A(n27458), .B(n26847), .Z(n24498) );
  ANDN U27813 ( .B(n26846), .A(n25850), .Z(n27458) );
  XOR U27814 ( .A(n26840), .B(n27459), .Z(n27454) );
  XNOR U27815 ( .A(n25087), .B(n26786), .Z(n27459) );
  XNOR U27816 ( .A(n27460), .B(n27461), .Z(n26786) );
  ANDN U27817 ( .B(n27462), .A(n26104), .Z(n27460) );
  XOR U27818 ( .A(n27463), .B(n26852), .Z(n25087) );
  ANDN U27819 ( .B(n25856), .A(n26851), .Z(n27463) );
  XOR U27820 ( .A(n27464), .B(n26859), .Z(n26840) );
  NOR U27821 ( .A(n25846), .B(n26858), .Z(n27464) );
  XOR U27822 ( .A(n27465), .B(n27466), .Z(n25589) );
  XOR U27823 ( .A(n27467), .B(n23995), .Z(n27466) );
  XOR U27824 ( .A(n27468), .B(n27469), .Z(n23995) );
  ANDN U27825 ( .B(n27470), .A(n27471), .Z(n27468) );
  XOR U27826 ( .A(n25869), .B(n27472), .Z(n27465) );
  XNOR U27827 ( .A(n24841), .B(n26634), .Z(n27472) );
  XOR U27828 ( .A(n27473), .B(n27474), .Z(n26634) );
  ANDN U27829 ( .B(n27475), .A(n27476), .Z(n27473) );
  XNOR U27830 ( .A(n27477), .B(n27478), .Z(n24841) );
  ANDN U27831 ( .B(n27479), .A(n27480), .Z(n27477) );
  XNOR U27832 ( .A(n27481), .B(n27482), .Z(n25869) );
  NOR U27833 ( .A(n27483), .B(n27484), .Z(n27481) );
  XOR U27834 ( .A(n27485), .B(n24182), .Z(n23530) );
  IV U27835 ( .A(n26078), .Z(n24182) );
  XOR U27836 ( .A(n27486), .B(n26544), .Z(n26078) );
  XNOR U27837 ( .A(n27487), .B(n27488), .Z(n26544) );
  XNOR U27838 ( .A(n24189), .B(n25882), .Z(n27488) );
  XNOR U27839 ( .A(n27489), .B(n27490), .Z(n25882) );
  ANDN U27840 ( .B(n27491), .A(n27492), .Z(n27489) );
  XNOR U27841 ( .A(n27493), .B(n27494), .Z(n24189) );
  ANDN U27842 ( .B(n27495), .A(n27496), .Z(n27493) );
  XOR U27843 ( .A(n24995), .B(n27497), .Z(n27487) );
  XNOR U27844 ( .A(n24010), .B(n26587), .Z(n27497) );
  XNOR U27845 ( .A(n27498), .B(n27499), .Z(n26587) );
  NOR U27846 ( .A(n27500), .B(n27501), .Z(n27498) );
  XNOR U27847 ( .A(n27502), .B(n27503), .Z(n24010) );
  ANDN U27848 ( .B(n27504), .A(n27505), .Z(n27502) );
  XOR U27849 ( .A(n27506), .B(n27507), .Z(n24995) );
  NOR U27850 ( .A(n27508), .B(n27509), .Z(n27506) );
  XOR U27851 ( .A(n19629), .B(n27510), .Z(n27432) );
  XOR U27852 ( .A(n19090), .B(n18399), .Z(n27510) );
  XNOR U27853 ( .A(n27511), .B(n23652), .Z(n18399) );
  XNOR U27854 ( .A(n23946), .B(n27512), .Z(n23652) );
  XOR U27855 ( .A(n27513), .B(n26764), .Z(n23946) );
  XOR U27856 ( .A(n27514), .B(n27515), .Z(n26764) );
  XOR U27857 ( .A(n25062), .B(n21724), .Z(n27515) );
  XNOR U27858 ( .A(n27516), .B(n27517), .Z(n21724) );
  ANDN U27859 ( .B(n27518), .A(n27519), .Z(n27516) );
  XOR U27860 ( .A(n27520), .B(n27521), .Z(n25062) );
  XOR U27861 ( .A(n23438), .B(n27524), .Z(n27514) );
  XOR U27862 ( .A(n27525), .B(n26836), .Z(n27524) );
  XOR U27863 ( .A(n27526), .B(n27527), .Z(n26836) );
  NOR U27864 ( .A(n27528), .B(n27529), .Z(n27526) );
  XNOR U27865 ( .A(n27530), .B(n27531), .Z(n23438) );
  ANDN U27866 ( .B(n27532), .A(n27533), .Z(n27530) );
  ANDN U27867 ( .B(n22743), .A(n22741), .Z(n27511) );
  XOR U27868 ( .A(n22608), .B(n27396), .Z(n22741) );
  XNOR U27869 ( .A(n27534), .B(n27535), .Z(n27396) );
  XOR U27870 ( .A(n27538), .B(n24986), .Z(n22743) );
  IV U27871 ( .A(n24827), .Z(n24986) );
  XOR U27872 ( .A(n27058), .B(n26952), .Z(n24827) );
  XNOR U27873 ( .A(n27539), .B(n27540), .Z(n26952) );
  XOR U27874 ( .A(n23252), .B(n25334), .Z(n27540) );
  XOR U27875 ( .A(n27541), .B(n27542), .Z(n25334) );
  NOR U27876 ( .A(n26993), .B(n27543), .Z(n27541) );
  XNOR U27877 ( .A(n27544), .B(n27545), .Z(n23252) );
  XOR U27878 ( .A(n26407), .B(n27548), .Z(n27539) );
  XOR U27879 ( .A(n24243), .B(n25215), .Z(n27548) );
  XNOR U27880 ( .A(n27549), .B(n27550), .Z(n25215) );
  XOR U27881 ( .A(n27553), .B(n27554), .Z(n24243) );
  ANDN U27882 ( .B(n26622), .A(n27555), .Z(n27553) );
  XOR U27883 ( .A(n27556), .B(n27557), .Z(n26407) );
  ANDN U27884 ( .B(n27558), .A(n27559), .Z(n27556) );
  XNOR U27885 ( .A(n27560), .B(n27561), .Z(n27058) );
  XOR U27886 ( .A(n26922), .B(n27562), .Z(n27561) );
  XNOR U27887 ( .A(n27563), .B(n27564), .Z(n26922) );
  ANDN U27888 ( .B(n27565), .A(n27566), .Z(n27563) );
  XOR U27889 ( .A(n27567), .B(n27568), .Z(n27560) );
  XOR U27890 ( .A(n26567), .B(n27569), .Z(n27568) );
  XNOR U27891 ( .A(n27570), .B(n27571), .Z(n26567) );
  ANDN U27892 ( .B(n27572), .A(n27573), .Z(n27570) );
  XNOR U27893 ( .A(n27574), .B(n24601), .Z(n19090) );
  IV U27894 ( .A(n23655), .Z(n24601) );
  XOR U27895 ( .A(n22624), .B(n27575), .Z(n23655) );
  XOR U27896 ( .A(n27576), .B(n27577), .Z(n22624) );
  NOR U27897 ( .A(n22732), .B(n22733), .Z(n27574) );
  XOR U27898 ( .A(n27578), .B(n23024), .Z(n22733) );
  XOR U27899 ( .A(n24196), .B(n27581), .Z(n22732) );
  IV U27900 ( .A(n23843), .Z(n24196) );
  XOR U27901 ( .A(n27582), .B(n27583), .Z(n23843) );
  XNOR U27902 ( .A(n27584), .B(n23650), .Z(n19629) );
  XNOR U27903 ( .A(n27374), .B(n24662), .Z(n23650) );
  XNOR U27904 ( .A(n25998), .B(n27585), .Z(n24662) );
  XOR U27905 ( .A(n27586), .B(n27587), .Z(n25998) );
  XNOR U27906 ( .A(n25750), .B(n25543), .Z(n27587) );
  XOR U27907 ( .A(n27588), .B(n27589), .Z(n25543) );
  ANDN U27908 ( .B(n27590), .A(n27591), .Z(n27588) );
  XOR U27909 ( .A(n27592), .B(n27593), .Z(n25750) );
  NOR U27910 ( .A(n27594), .B(n27595), .Z(n27592) );
  XNOR U27911 ( .A(n22405), .B(n27596), .Z(n27586) );
  XOR U27912 ( .A(n24029), .B(n21715), .Z(n27596) );
  XOR U27913 ( .A(n27597), .B(n27598), .Z(n21715) );
  XNOR U27914 ( .A(n27601), .B(n27602), .Z(n24029) );
  ANDN U27915 ( .B(n27603), .A(n27604), .Z(n27601) );
  XOR U27916 ( .A(n27605), .B(n27606), .Z(n22405) );
  ANDN U27917 ( .B(n27607), .A(n27608), .Z(n27605) );
  XNOR U27918 ( .A(n27609), .B(n27610), .Z(n27374) );
  ANDN U27919 ( .B(n27611), .A(n27612), .Z(n27609) );
  ANDN U27920 ( .B(n22738), .A(n22737), .Z(n27584) );
  XOR U27921 ( .A(n27613), .B(n24926), .Z(n22737) );
  XNOR U27922 ( .A(n27614), .B(n27615), .Z(n26763) );
  XNOR U27923 ( .A(n26516), .B(n23952), .Z(n27615) );
  XOR U27924 ( .A(n27616), .B(n27617), .Z(n23952) );
  ANDN U27925 ( .B(n27618), .A(n27619), .Z(n27616) );
  XNOR U27926 ( .A(n27620), .B(n27621), .Z(n26516) );
  ANDN U27927 ( .B(n27622), .A(n27623), .Z(n27620) );
  XNOR U27928 ( .A(n24763), .B(n27624), .Z(n27614) );
  XOR U27929 ( .A(n24008), .B(n26282), .Z(n27624) );
  XNOR U27930 ( .A(n27625), .B(n27626), .Z(n26282) );
  NOR U27931 ( .A(n27627), .B(n27628), .Z(n27625) );
  XNOR U27932 ( .A(n27629), .B(n27630), .Z(n24008) );
  XNOR U27933 ( .A(n27633), .B(n27634), .Z(n24763) );
  ANDN U27934 ( .B(n27635), .A(n27636), .Z(n27633) );
  XOR U27935 ( .A(n27172), .B(n27638), .Z(n22738) );
  IV U27936 ( .A(n25414), .Z(n27172) );
  XNOR U27937 ( .A(n15956), .B(n21804), .Z(n13499) );
  XOR U27938 ( .A(n27639), .B(n24507), .Z(n21804) );
  IV U27939 ( .A(n27640), .Z(n24507) );
  AND U27940 ( .A(n20621), .B(n23795), .Z(n27639) );
  XOR U27941 ( .A(n27641), .B(n25023), .Z(n20621) );
  IV U27942 ( .A(n26280), .Z(n25023) );
  XNOR U27943 ( .A(n20192), .B(n20249), .Z(n15956) );
  XNOR U27944 ( .A(n27642), .B(n27643), .Z(n20249) );
  XNOR U27945 ( .A(n18902), .B(n17653), .Z(n27643) );
  XNOR U27946 ( .A(n27644), .B(n21513), .Z(n17653) );
  XNOR U27947 ( .A(n25362), .B(n27645), .Z(n21513) );
  ANDN U27948 ( .B(n21514), .A(n21778), .Z(n27644) );
  XOR U27949 ( .A(n26358), .B(n26944), .Z(n21778) );
  XNOR U27950 ( .A(n27646), .B(n27647), .Z(n26245) );
  XNOR U27951 ( .A(n27648), .B(n26700), .Z(n27647) );
  XNOR U27952 ( .A(n27649), .B(n27650), .Z(n26700) );
  XOR U27953 ( .A(n27651), .B(n27652), .Z(n27128) );
  XOR U27954 ( .A(n25489), .B(n27653), .Z(n27646) );
  XOR U27955 ( .A(n27654), .B(n24289), .Z(n27653) );
  XOR U27956 ( .A(n27655), .B(n27656), .Z(n24289) );
  NOR U27957 ( .A(n27134), .B(n26365), .Z(n27655) );
  XOR U27958 ( .A(n27657), .B(n27658), .Z(n27134) );
  XOR U27959 ( .A(n27659), .B(n27660), .Z(n25489) );
  NOR U27960 ( .A(n26355), .B(n26356), .Z(n27659) );
  XNOR U27961 ( .A(n27661), .B(n27662), .Z(n26356) );
  XNOR U27962 ( .A(n27664), .B(n27665), .Z(n26358) );
  ANDN U27963 ( .B(n27139), .A(n27137), .Z(n27664) );
  XNOR U27964 ( .A(n25577), .B(n27666), .Z(n21514) );
  XNOR U27965 ( .A(n21523), .B(n27667), .Z(n18902) );
  XOR U27966 ( .A(n27668), .B(n4694), .Z(n27667) );
  NANDN U27967 ( .A(rc_i[1]), .B(n11417), .Z(n4694) );
  ANDN U27968 ( .B(n21790), .A(n21524), .Z(n27668) );
  XOR U27969 ( .A(n26454), .B(n27267), .Z(n21790) );
  XNOR U27970 ( .A(n27670), .B(n27671), .Z(n27267) );
  NOR U27971 ( .A(n27672), .B(n27673), .Z(n27670) );
  XOR U27972 ( .A(n27674), .B(n24411), .Z(n21523) );
  XOR U27973 ( .A(n21506), .B(n27675), .Z(n27642) );
  XNOR U27974 ( .A(n17959), .B(n19216), .Z(n27675) );
  XNOR U27975 ( .A(n27676), .B(n26149), .Z(n19216) );
  XOR U27976 ( .A(n27677), .B(n27678), .Z(n26149) );
  ANDN U27977 ( .B(n21792), .A(n21794), .Z(n27676) );
  XOR U27978 ( .A(n27679), .B(n22521), .Z(n21794) );
  XOR U27979 ( .A(n27680), .B(n27681), .Z(n26702) );
  XNOR U27980 ( .A(n25031), .B(n26001), .Z(n27681) );
  XNOR U27981 ( .A(n27682), .B(n27683), .Z(n26001) );
  NOR U27982 ( .A(n27684), .B(n27685), .Z(n27682) );
  XOR U27983 ( .A(n27686), .B(n27687), .Z(n25031) );
  ANDN U27984 ( .B(n27688), .A(n27689), .Z(n27686) );
  XOR U27985 ( .A(n23431), .B(n27690), .Z(n27680) );
  XNOR U27986 ( .A(n23819), .B(n27691), .Z(n27690) );
  XOR U27987 ( .A(n27692), .B(n27693), .Z(n23819) );
  ANDN U27988 ( .B(n27694), .A(n27695), .Z(n27692) );
  XNOR U27989 ( .A(n27696), .B(n27697), .Z(n23431) );
  ANDN U27990 ( .B(n27698), .A(n27699), .Z(n27696) );
  XNOR U27991 ( .A(n26904), .B(n27701), .Z(n21792) );
  XNOR U27992 ( .A(n27702), .B(n23083), .Z(n17959) );
  XOR U27993 ( .A(n27703), .B(n23021), .Z(n23083) );
  IV U27994 ( .A(n25301), .Z(n23021) );
  XOR U27995 ( .A(n26517), .B(n27704), .Z(n25301) );
  XOR U27996 ( .A(n27705), .B(n27706), .Z(n26517) );
  XOR U27997 ( .A(n23938), .B(n25261), .Z(n27706) );
  XNOR U27998 ( .A(n27707), .B(n26677), .Z(n25261) );
  ANDN U27999 ( .B(n27708), .A(n26678), .Z(n27707) );
  XOR U28000 ( .A(n27709), .B(n27232), .Z(n23938) );
  NOR U28001 ( .A(n27231), .B(n27710), .Z(n27709) );
  XOR U28002 ( .A(n23849), .B(n27711), .Z(n27705) );
  XOR U28003 ( .A(n23811), .B(n23764), .Z(n27711) );
  XNOR U28004 ( .A(n27712), .B(n26688), .Z(n23764) );
  NOR U28005 ( .A(n27713), .B(n26687), .Z(n27712) );
  XNOR U28006 ( .A(n27714), .B(n27715), .Z(n23811) );
  ANDN U28007 ( .B(n27716), .A(n26683), .Z(n27714) );
  XNOR U28008 ( .A(n27717), .B(n27718), .Z(n23849) );
  ANDN U28009 ( .B(n27719), .A(n27720), .Z(n27717) );
  ANDN U28010 ( .B(n21781), .A(n21782), .Z(n27702) );
  XNOR U28011 ( .A(n27721), .B(n22793), .Z(n21782) );
  XOR U28012 ( .A(n27722), .B(n25457), .Z(n21781) );
  IV U28013 ( .A(n27723), .Z(n25457) );
  XNOR U28014 ( .A(n27724), .B(n21519), .Z(n21506) );
  XNOR U28015 ( .A(n27725), .B(n25008), .Z(n21519) );
  ANDN U28016 ( .B(n21520), .A(n21786), .Z(n27724) );
  XOR U28017 ( .A(n27726), .B(n24515), .Z(n21786) );
  XOR U28018 ( .A(n27727), .B(n21225), .Z(n21520) );
  XNOR U28019 ( .A(n27728), .B(n27729), .Z(n21225) );
  XOR U28020 ( .A(n27730), .B(n27731), .Z(n20192) );
  XNOR U28021 ( .A(n17319), .B(n17196), .Z(n27731) );
  XNOR U28022 ( .A(n27732), .B(n20623), .Z(n17196) );
  XNOR U28023 ( .A(n24278), .B(n27733), .Z(n20623) );
  NOR U28024 ( .A(n27640), .B(n23795), .Z(n27732) );
  XOR U28025 ( .A(n24930), .B(n27734), .Z(n23795) );
  XOR U28026 ( .A(n27735), .B(n27723), .Z(n27640) );
  XNOR U28027 ( .A(n27736), .B(n23803), .Z(n17319) );
  XNOR U28028 ( .A(n27737), .B(n24825), .Z(n23803) );
  NOR U28029 ( .A(n21800), .B(n21798), .Z(n27736) );
  XOR U28030 ( .A(n27738), .B(n25008), .Z(n21798) );
  XOR U28031 ( .A(n26462), .B(n26246), .Z(n25008) );
  XNOR U28032 ( .A(n27739), .B(n27740), .Z(n26246) );
  XNOR U28033 ( .A(n24418), .B(n25077), .Z(n27740) );
  XNOR U28034 ( .A(n27741), .B(n27742), .Z(n25077) );
  XNOR U28035 ( .A(n27744), .B(n27745), .Z(n24418) );
  NOR U28036 ( .A(n27746), .B(n26428), .Z(n27744) );
  XOR U28037 ( .A(n25101), .B(n27747), .Z(n27739) );
  XNOR U28038 ( .A(n24398), .B(n24927), .Z(n27747) );
  XNOR U28039 ( .A(n27748), .B(n27749), .Z(n24927) );
  NOR U28040 ( .A(n27750), .B(n26433), .Z(n27748) );
  XNOR U28041 ( .A(n27751), .B(n27752), .Z(n24398) );
  NOR U28042 ( .A(n27753), .B(n26441), .Z(n27751) );
  XOR U28043 ( .A(n27754), .B(n27755), .Z(n25101) );
  ANDN U28044 ( .B(n27756), .A(n26424), .Z(n27754) );
  XOR U28045 ( .A(n27757), .B(n27758), .Z(n26462) );
  XOR U28046 ( .A(n27759), .B(n23062), .Z(n27758) );
  XOR U28047 ( .A(n27760), .B(n27761), .Z(n23062) );
  NOR U28048 ( .A(n27762), .B(n27763), .Z(n27760) );
  XOR U28049 ( .A(n24476), .B(n27764), .Z(n27757) );
  XOR U28050 ( .A(n26709), .B(n23973), .Z(n27764) );
  XNOR U28051 ( .A(n27765), .B(n27766), .Z(n23973) );
  ANDN U28052 ( .B(n27767), .A(n27768), .Z(n27765) );
  XNOR U28053 ( .A(n27769), .B(n27770), .Z(n26709) );
  ANDN U28054 ( .B(n27771), .A(n27772), .Z(n27769) );
  XNOR U28055 ( .A(n27773), .B(n27774), .Z(n24476) );
  ANDN U28056 ( .B(n27775), .A(n27776), .Z(n27773) );
  XOR U28057 ( .A(n27777), .B(n26188), .Z(n21800) );
  IV U28058 ( .A(n24989), .Z(n26188) );
  XOR U28059 ( .A(n26341), .B(n27778), .Z(n24989) );
  XOR U28060 ( .A(n27779), .B(n27780), .Z(n26341) );
  XNOR U28061 ( .A(n24925), .B(n25098), .Z(n27780) );
  XOR U28062 ( .A(n27781), .B(n27618), .Z(n25098) );
  ANDN U28063 ( .B(n27619), .A(n27782), .Z(n27781) );
  XNOR U28064 ( .A(n27783), .B(n27627), .Z(n24925) );
  ANDN U28065 ( .B(n27628), .A(n27784), .Z(n27783) );
  XOR U28066 ( .A(n27613), .B(n27785), .Z(n27779) );
  XOR U28067 ( .A(n27359), .B(n25922), .Z(n27785) );
  XNOR U28068 ( .A(n27786), .B(n27636), .Z(n25922) );
  NOR U28069 ( .A(n27787), .B(n27635), .Z(n27786) );
  XNOR U28070 ( .A(n27788), .B(n27632), .Z(n27359) );
  NOR U28071 ( .A(n27631), .B(n27789), .Z(n27788) );
  XNOR U28072 ( .A(n27790), .B(n27623), .Z(n27613) );
  ANDN U28073 ( .B(n27791), .A(n27622), .Z(n27790) );
  XNOR U28074 ( .A(n21183), .B(n27792), .Z(n27730) );
  XOR U28075 ( .A(n18041), .B(n19962), .Z(n27792) );
  XNOR U28076 ( .A(n27793), .B(n20613), .Z(n19962) );
  XNOR U28077 ( .A(n27794), .B(n24798), .Z(n20613) );
  NOR U28078 ( .A(n21802), .B(n21803), .Z(n27793) );
  XOR U28079 ( .A(n27797), .B(n21823), .Z(n21802) );
  IV U28080 ( .A(n25963), .Z(n21823) );
  XNOR U28081 ( .A(n25512), .B(n26671), .Z(n25963) );
  XNOR U28082 ( .A(n27798), .B(n27799), .Z(n26671) );
  XOR U28083 ( .A(n27800), .B(n25544), .Z(n27799) );
  XNOR U28084 ( .A(n27801), .B(n27791), .Z(n25544) );
  ANDN U28085 ( .B(n27802), .A(n27621), .Z(n27801) );
  XNOR U28086 ( .A(n25897), .B(n27803), .Z(n27798) );
  XNOR U28087 ( .A(n27804), .B(n24391), .Z(n27803) );
  XOR U28088 ( .A(n27805), .B(n27787), .Z(n24391) );
  ANDN U28089 ( .B(n27806), .A(n27634), .Z(n27805) );
  XOR U28090 ( .A(n27807), .B(n27782), .Z(n25897) );
  AND U28091 ( .A(n27617), .B(n27808), .Z(n27807) );
  XOR U28092 ( .A(n27809), .B(n27810), .Z(n25512) );
  XOR U28093 ( .A(n27811), .B(n25664), .Z(n27810) );
  XNOR U28094 ( .A(n27812), .B(n27813), .Z(n25664) );
  ANDN U28095 ( .B(n27814), .A(n27815), .Z(n27812) );
  XOR U28096 ( .A(n25139), .B(n27816), .Z(n27809) );
  XOR U28097 ( .A(n24631), .B(n24597), .Z(n27816) );
  XNOR U28098 ( .A(n27817), .B(n27818), .Z(n24597) );
  NOR U28099 ( .A(n27531), .B(n27819), .Z(n27817) );
  XNOR U28100 ( .A(n27820), .B(n27821), .Z(n24631) );
  NOR U28101 ( .A(n27822), .B(n27517), .Z(n27820) );
  XNOR U28102 ( .A(n27823), .B(n27824), .Z(n25139) );
  ANDN U28103 ( .B(n27527), .A(n27825), .Z(n27823) );
  XNOR U28104 ( .A(n27826), .B(n20626), .Z(n18041) );
  XNOR U28105 ( .A(n27827), .B(n21368), .Z(n20626) );
  XNOR U28106 ( .A(n27828), .B(n27829), .Z(n27728) );
  XNOR U28107 ( .A(n26729), .B(n24757), .Z(n27829) );
  XNOR U28108 ( .A(n27830), .B(n26742), .Z(n24757) );
  ANDN U28109 ( .B(n26743), .A(n27831), .Z(n27830) );
  XNOR U28110 ( .A(n27832), .B(n27833), .Z(n26729) );
  NOR U28111 ( .A(n27834), .B(n27835), .Z(n27832) );
  XNOR U28112 ( .A(n25670), .B(n27836), .Z(n27828) );
  XOR U28113 ( .A(n24628), .B(n24606), .Z(n27836) );
  XNOR U28114 ( .A(n27837), .B(n27838), .Z(n24606) );
  AND U28115 ( .A(n27839), .B(n27840), .Z(n27837) );
  XNOR U28116 ( .A(n27841), .B(n26737), .Z(n24628) );
  NOR U28117 ( .A(n26736), .B(n27842), .Z(n27841) );
  IV U28118 ( .A(n27843), .Z(n26736) );
  XNOR U28119 ( .A(n27844), .B(n26746), .Z(n25670) );
  ANDN U28120 ( .B(n26747), .A(n27845), .Z(n27844) );
  ANDN U28121 ( .B(n23799), .A(n24500), .Z(n27826) );
  XOR U28122 ( .A(n22213), .B(n27847), .Z(n24500) );
  XOR U28123 ( .A(n27848), .B(n27849), .Z(n22213) );
  IV U28124 ( .A(n21808), .Z(n23799) );
  XOR U28125 ( .A(n27850), .B(n25766), .Z(n21808) );
  IV U28126 ( .A(n25776), .Z(n25766) );
  XOR U28127 ( .A(n26420), .B(n27851), .Z(n25776) );
  XOR U28128 ( .A(n27852), .B(n27853), .Z(n26420) );
  XOR U28129 ( .A(n24834), .B(n25354), .Z(n27853) );
  XOR U28130 ( .A(n27854), .B(n27855), .Z(n25354) );
  ANDN U28131 ( .B(n27856), .A(n27857), .Z(n27854) );
  XOR U28132 ( .A(n27858), .B(n27859), .Z(n24834) );
  NOR U28133 ( .A(n27860), .B(n27861), .Z(n27858) );
  XOR U28134 ( .A(n27862), .B(n27863), .Z(n27852) );
  XOR U28135 ( .A(n25666), .B(n25081), .Z(n27863) );
  XNOR U28136 ( .A(n27864), .B(n27772), .Z(n25081) );
  XOR U28137 ( .A(n27867), .B(n27767), .Z(n25666) );
  ANDN U28138 ( .B(n27868), .A(n27869), .Z(n27867) );
  XOR U28139 ( .A(n27870), .B(n20617), .Z(n21183) );
  XOR U28140 ( .A(n27871), .B(n22943), .Z(n20617) );
  NOR U28141 ( .A(n21810), .B(n21811), .Z(n27870) );
  XOR U28142 ( .A(n22641), .B(n27872), .Z(n21811) );
  XOR U28143 ( .A(n27874), .B(n27875), .Z(n24379) );
  XOR U28144 ( .A(n11227), .B(n27876), .Z(n26664) );
  XOR U28145 ( .A(n11113), .B(n14181), .Z(n27876) );
  XNOR U28146 ( .A(n27877), .B(n16210), .Z(n14181) );
  XNOR U28147 ( .A(n24204), .B(n16531), .Z(n16210) );
  XOR U28148 ( .A(n20134), .B(n20077), .Z(n16531) );
  XNOR U28149 ( .A(n27878), .B(n27879), .Z(n20077) );
  XOR U28150 ( .A(n19511), .B(n16601), .Z(n27879) );
  XOR U28151 ( .A(n27880), .B(n21102), .Z(n16601) );
  ANDN U28152 ( .B(n19619), .A(n21101), .Z(n27880) );
  XOR U28153 ( .A(n25916), .B(n27881), .Z(n21101) );
  XOR U28154 ( .A(n26089), .B(n27882), .Z(n19619) );
  XOR U28155 ( .A(n27883), .B(n21106), .Z(n19511) );
  ANDN U28156 ( .B(n21472), .A(n21470), .Z(n27883) );
  XOR U28157 ( .A(n23422), .B(n25524), .Z(n21470) );
  XOR U28158 ( .A(n27884), .B(n27255), .Z(n25524) );
  ANDN U28159 ( .B(n27885), .A(n27886), .Z(n27884) );
  XOR U28160 ( .A(n26886), .B(n26579), .Z(n21472) );
  XNOR U28161 ( .A(n27889), .B(n27890), .Z(n26579) );
  XOR U28162 ( .A(n27891), .B(n27892), .Z(n26886) );
  ANDN U28163 ( .B(n27182), .A(n27893), .Z(n27891) );
  XNOR U28164 ( .A(n18446), .B(n27894), .Z(n27878) );
  XNOR U28165 ( .A(n18527), .B(n19762), .Z(n27894) );
  XNOR U28166 ( .A(n27895), .B(n21147), .Z(n19762) );
  AND U28167 ( .A(n19843), .B(n21148), .Z(n27895) );
  XOR U28168 ( .A(n27896), .B(n22536), .Z(n21148) );
  IV U28169 ( .A(n25551), .Z(n22536) );
  XOR U28170 ( .A(n27899), .B(n24150), .Z(n19843) );
  IV U28171 ( .A(n22517), .Z(n24150) );
  XOR U28172 ( .A(n27902), .B(n27903), .Z(n18527) );
  XNOR U28173 ( .A(n25362), .B(n27904), .Z(n19626) );
  XOR U28174 ( .A(n27905), .B(n21112), .Z(n18446) );
  NOR U28175 ( .A(n20022), .B(n21111), .Z(n27905) );
  XOR U28176 ( .A(n24623), .B(n27906), .Z(n21111) );
  XOR U28177 ( .A(n27907), .B(n27908), .Z(n24623) );
  XNOR U28178 ( .A(n25282), .B(n27909), .Z(n20022) );
  IV U28179 ( .A(n25986), .Z(n25282) );
  XOR U28180 ( .A(n27910), .B(n27911), .Z(n20134) );
  XNOR U28181 ( .A(n19548), .B(n18101), .Z(n27911) );
  XNOR U28182 ( .A(n27912), .B(n22765), .Z(n18101) );
  NOR U28183 ( .A(n21047), .B(n22764), .Z(n27912) );
  XOR U28184 ( .A(n27913), .B(n24193), .Z(n22764) );
  XOR U28185 ( .A(n27313), .B(n23825), .Z(n21047) );
  IV U28186 ( .A(n25974), .Z(n23825) );
  XNOR U28187 ( .A(n27914), .B(n27915), .Z(n27313) );
  NOR U28188 ( .A(n27916), .B(n27917), .Z(n27914) );
  XNOR U28189 ( .A(n27918), .B(n22772), .Z(n19548) );
  ANDN U28190 ( .B(n21056), .A(n22773), .Z(n27918) );
  XOR U28191 ( .A(n27919), .B(n24296), .Z(n22773) );
  XOR U28192 ( .A(n23489), .B(n27920), .Z(n21056) );
  XOR U28193 ( .A(n18883), .B(n27921), .Z(n27910) );
  XOR U28194 ( .A(n21096), .B(n19384), .Z(n27921) );
  XNOR U28195 ( .A(n27922), .B(n22769), .Z(n19384) );
  XOR U28196 ( .A(n27525), .B(n21725), .Z(n21051) );
  XNOR U28197 ( .A(n27924), .B(n27925), .Z(n26518) );
  XOR U28198 ( .A(n24171), .B(n24817), .Z(n27925) );
  XOR U28199 ( .A(n27926), .B(n27927), .Z(n24817) );
  XOR U28200 ( .A(n27928), .B(n27929), .Z(n27627) );
  XNOR U28201 ( .A(n27930), .B(n27931), .Z(n24171) );
  ANDN U28202 ( .B(n27630), .A(n27632), .Z(n27930) );
  XOR U28203 ( .A(n24194), .B(n27934), .Z(n27924) );
  XOR U28204 ( .A(n26670), .B(n26630), .Z(n27934) );
  XNOR U28205 ( .A(n27935), .B(n27802), .Z(n26630) );
  XOR U28206 ( .A(n27938), .B(n27939), .Z(n27623) );
  XNOR U28207 ( .A(n27940), .B(n27806), .Z(n26670) );
  AND U28208 ( .A(n27634), .B(n27636), .Z(n27940) );
  XOR U28209 ( .A(n27941), .B(n27942), .Z(n27636) );
  XNOR U28210 ( .A(n27943), .B(n27944), .Z(n27634) );
  XNOR U28211 ( .A(n27945), .B(n27808), .Z(n24194) );
  NOR U28212 ( .A(n27617), .B(n27618), .Z(n27945) );
  XOR U28213 ( .A(n27946), .B(n27947), .Z(n27618) );
  XOR U28214 ( .A(n27948), .B(n27949), .Z(n27617) );
  XOR U28215 ( .A(n27950), .B(n27814), .Z(n27525) );
  NOR U28216 ( .A(n27951), .B(n27952), .Z(n27950) );
  XOR U28217 ( .A(n22829), .B(n27953), .Z(n22770) );
  XOR U28218 ( .A(n27954), .B(n27955), .Z(n22829) );
  XNOR U28219 ( .A(n27956), .B(n22761), .Z(n21096) );
  AND U28220 ( .A(n22762), .B(n21060), .Z(n27956) );
  XOR U28221 ( .A(n24278), .B(n27957), .Z(n21060) );
  XNOR U28222 ( .A(n27958), .B(n27959), .Z(n24278) );
  XOR U28223 ( .A(n27960), .B(n23250), .Z(n22762) );
  XNOR U28224 ( .A(n27961), .B(n22777), .Z(n18883) );
  NOR U28225 ( .A(n21064), .B(n22776), .Z(n27961) );
  XOR U28226 ( .A(n27962), .B(n22776), .Z(n24204) );
  XNOR U28227 ( .A(n22944), .B(n27963), .Z(n22776) );
  XOR U28228 ( .A(n27964), .B(n26258), .Z(n22944) );
  XOR U28229 ( .A(n27965), .B(n27966), .Z(n26258) );
  XOR U28230 ( .A(n27735), .B(n27967), .Z(n27966) );
  XNOR U28231 ( .A(n27968), .B(n27969), .Z(n27735) );
  ANDN U28232 ( .B(n27970), .A(n27971), .Z(n27968) );
  XOR U28233 ( .A(n27722), .B(n27972), .Z(n27965) );
  XNOR U28234 ( .A(n25456), .B(n27973), .Z(n27972) );
  XNOR U28235 ( .A(n27974), .B(n27975), .Z(n25456) );
  NOR U28236 ( .A(n27976), .B(n27977), .Z(n27974) );
  XOR U28237 ( .A(n27978), .B(n27979), .Z(n27722) );
  NOR U28238 ( .A(n27980), .B(n27981), .Z(n27978) );
  ANDN U28239 ( .B(n21064), .A(n27982), .Z(n27962) );
  XNOR U28240 ( .A(n27983), .B(n24857), .Z(n21064) );
  XNOR U28241 ( .A(n27984), .B(n26866), .Z(n24857) );
  XNOR U28242 ( .A(n27985), .B(n27986), .Z(n26866) );
  XNOR U28243 ( .A(n27987), .B(n27988), .Z(n27986) );
  XNOR U28244 ( .A(n25378), .B(n27989), .Z(n27985) );
  XNOR U28245 ( .A(n26284), .B(n23067), .Z(n27989) );
  XNOR U28246 ( .A(n27990), .B(n27991), .Z(n23067) );
  ANDN U28247 ( .B(n27992), .A(n27993), .Z(n27990) );
  ANDN U28248 ( .B(n27996), .A(n27997), .Z(n27994) );
  XOR U28249 ( .A(n27998), .B(n27999), .Z(n25378) );
  XOR U28250 ( .A(n18530), .B(n22456), .Z(n13502) );
  XNOR U28251 ( .A(n28002), .B(n25639), .Z(n22456) );
  IV U28252 ( .A(n28003), .Z(n25639) );
  NOR U28253 ( .A(n23208), .B(n23206), .Z(n28002) );
  IV U28254 ( .A(n16753), .Z(n18530) );
  XOR U28255 ( .A(n22911), .B(n21253), .Z(n16753) );
  XOR U28256 ( .A(n28004), .B(n28005), .Z(n21253) );
  XOR U28257 ( .A(n18038), .B(n22208), .Z(n28005) );
  XOR U28258 ( .A(n28006), .B(n26033), .Z(n22208) );
  XOR U28259 ( .A(n24778), .B(n28007), .Z(n26033) );
  IV U28260 ( .A(n23905), .Z(n24778) );
  XOR U28261 ( .A(n28008), .B(n28009), .Z(n23905) );
  ANDN U28262 ( .B(n22478), .A(n22476), .Z(n28006) );
  IV U28263 ( .A(n26047), .Z(n22476) );
  XOR U28264 ( .A(n25016), .B(n28010), .Z(n26047) );
  XNOR U28265 ( .A(n25476), .B(n28011), .Z(n22478) );
  XOR U28266 ( .A(n28012), .B(n26373), .Z(n25476) );
  XNOR U28267 ( .A(n28013), .B(n28014), .Z(n26373) );
  XOR U28268 ( .A(n21583), .B(n28015), .Z(n28014) );
  XNOR U28269 ( .A(n28016), .B(n28017), .Z(n21583) );
  ANDN U28270 ( .B(n28018), .A(n28019), .Z(n28016) );
  XOR U28271 ( .A(n23069), .B(n28020), .Z(n28013) );
  XOR U28272 ( .A(n25510), .B(n26193), .Z(n28020) );
  XNOR U28273 ( .A(n28021), .B(n28022), .Z(n26193) );
  NOR U28274 ( .A(n28023), .B(n28024), .Z(n28021) );
  XNOR U28275 ( .A(n28025), .B(n28026), .Z(n25510) );
  NOR U28276 ( .A(n28027), .B(n28028), .Z(n28025) );
  XNOR U28277 ( .A(n28029), .B(n28030), .Z(n23069) );
  ANDN U28278 ( .B(n28031), .A(n28032), .Z(n28029) );
  XOR U28279 ( .A(n28033), .B(n22250), .Z(n18038) );
  XNOR U28280 ( .A(n26568), .B(n27569), .Z(n22250) );
  XNOR U28281 ( .A(n28034), .B(n28035), .Z(n27569) );
  NOR U28282 ( .A(n28036), .B(n28037), .Z(n28034) );
  ANDN U28283 ( .B(n22251), .A(n22484), .Z(n28033) );
  XOR U28284 ( .A(n28038), .B(n24525), .Z(n22484) );
  IV U28285 ( .A(n24846), .Z(n24525) );
  XOR U28286 ( .A(n28039), .B(n26153), .Z(n24846) );
  XNOR U28287 ( .A(n28040), .B(n28041), .Z(n26153) );
  XNOR U28288 ( .A(n24026), .B(n25256), .Z(n28041) );
  XOR U28289 ( .A(n28042), .B(n27368), .Z(n25256) );
  ANDN U28290 ( .B(n28043), .A(n27367), .Z(n28042) );
  XNOR U28291 ( .A(n28044), .B(n28045), .Z(n24026) );
  XOR U28292 ( .A(n26415), .B(n28047), .Z(n28040) );
  XNOR U28293 ( .A(n24245), .B(n27361), .Z(n28047) );
  XNOR U28294 ( .A(n28048), .B(n27377), .Z(n27361) );
  ANDN U28295 ( .B(n28049), .A(n28050), .Z(n28048) );
  XNOR U28296 ( .A(n28051), .B(n28052), .Z(n24245) );
  ANDN U28297 ( .B(n28053), .A(n27611), .Z(n28051) );
  XNOR U28298 ( .A(n28054), .B(n27381), .Z(n26415) );
  XOR U28299 ( .A(n28056), .B(n24366), .Z(n22251) );
  XOR U28300 ( .A(n19520), .B(n28057), .Z(n28004) );
  XOR U28301 ( .A(n17748), .B(n17600), .Z(n28057) );
  XOR U28302 ( .A(n28058), .B(n22246), .Z(n17600) );
  XOR U28303 ( .A(n28059), .B(n23855), .Z(n22246) );
  IV U28304 ( .A(n27678), .Z(n23855) );
  XOR U28305 ( .A(n28060), .B(n28061), .Z(n27678) );
  ANDN U28306 ( .B(n22247), .A(n22472), .Z(n28058) );
  XOR U28307 ( .A(n26656), .B(n25942), .Z(n22472) );
  XNOR U28308 ( .A(n28062), .B(n28063), .Z(n26656) );
  ANDN U28309 ( .B(n28064), .A(n28065), .Z(n28062) );
  XOR U28310 ( .A(n22409), .B(n28066), .Z(n22247) );
  IV U28311 ( .A(n25916), .Z(n22409) );
  XOR U28312 ( .A(n27959), .B(n26541), .Z(n25916) );
  XNOR U28313 ( .A(n28067), .B(n28068), .Z(n26541) );
  XOR U28314 ( .A(n26392), .B(n24378), .Z(n28068) );
  XNOR U28315 ( .A(n28069), .B(n28070), .Z(n24378) );
  ANDN U28316 ( .B(n28071), .A(n28072), .Z(n28069) );
  XNOR U28317 ( .A(n28073), .B(n28074), .Z(n26392) );
  ANDN U28318 ( .B(n28075), .A(n28076), .Z(n28073) );
  XOR U28319 ( .A(n26339), .B(n28077), .Z(n28067) );
  XNOR U28320 ( .A(n27873), .B(n24956), .Z(n28077) );
  XNOR U28321 ( .A(n28078), .B(n28079), .Z(n24956) );
  ANDN U28322 ( .B(n28080), .A(n28081), .Z(n28078) );
  XNOR U28323 ( .A(n28082), .B(n28083), .Z(n27873) );
  NOR U28324 ( .A(n28084), .B(n28085), .Z(n28082) );
  XOR U28325 ( .A(n28086), .B(n28087), .Z(n26339) );
  ANDN U28326 ( .B(n28088), .A(n28089), .Z(n28086) );
  XNOR U28327 ( .A(n28090), .B(n28091), .Z(n27959) );
  XOR U28328 ( .A(n28056), .B(n28092), .Z(n28091) );
  XNOR U28329 ( .A(n28093), .B(n28094), .Z(n28056) );
  ANDN U28330 ( .B(n28095), .A(n28096), .Z(n28093) );
  XNOR U28331 ( .A(n24365), .B(n28097), .Z(n28090) );
  XNOR U28332 ( .A(n28098), .B(n26906), .Z(n28097) );
  XOR U28333 ( .A(n28099), .B(n28100), .Z(n26906) );
  ANDN U28334 ( .B(n28101), .A(n28102), .Z(n28099) );
  XNOR U28335 ( .A(n28103), .B(n28104), .Z(n24365) );
  ANDN U28336 ( .B(n28105), .A(n28106), .Z(n28103) );
  XNOR U28337 ( .A(n28107), .B(n22240), .Z(n17748) );
  XOR U28338 ( .A(n28108), .B(n25996), .Z(n22240) );
  IV U28339 ( .A(n23250), .Z(n25996) );
  AND U28340 ( .A(n22481), .B(n22241), .Z(n28107) );
  XOR U28341 ( .A(n27691), .B(n25032), .Z(n22241) );
  XNOR U28342 ( .A(n28110), .B(n28111), .Z(n26863) );
  XOR U28343 ( .A(n28112), .B(n24230), .Z(n28111) );
  XOR U28344 ( .A(n28113), .B(n28114), .Z(n24230) );
  ANDN U28345 ( .B(n27685), .A(n27683), .Z(n28113) );
  IV U28346 ( .A(n28115), .Z(n27683) );
  XOR U28347 ( .A(n26923), .B(n28116), .Z(n28110) );
  XOR U28348 ( .A(n27001), .B(n26223), .Z(n28116) );
  XNOR U28349 ( .A(n28117), .B(n28118), .Z(n26223) );
  XNOR U28350 ( .A(n28121), .B(n28122), .Z(n27001) );
  NOR U28351 ( .A(n28123), .B(n27694), .Z(n28121) );
  XOR U28352 ( .A(n28124), .B(n28125), .Z(n26923) );
  NOR U28353 ( .A(n27697), .B(n27698), .Z(n28124) );
  XNOR U28354 ( .A(n28126), .B(n28120), .Z(n27691) );
  ANDN U28355 ( .B(n28119), .A(n28127), .Z(n28126) );
  XOR U28356 ( .A(n27116), .B(n25182), .Z(n22481) );
  XNOR U28357 ( .A(n28128), .B(n28129), .Z(n27116) );
  ANDN U28358 ( .B(n28130), .A(n28131), .Z(n28128) );
  XNOR U28359 ( .A(n28132), .B(n26040), .Z(n19520) );
  IV U28360 ( .A(n22236), .Z(n26040) );
  XOR U28361 ( .A(n26924), .B(n28133), .Z(n22236) );
  XNOR U28362 ( .A(n23725), .B(n28134), .Z(n22470) );
  XOR U28363 ( .A(n28135), .B(n26812), .Z(n23725) );
  XNOR U28364 ( .A(n28136), .B(n28137), .Z(n26812) );
  XNOR U28365 ( .A(n26920), .B(n27485), .Z(n28137) );
  XOR U28366 ( .A(n28138), .B(n28139), .Z(n27485) );
  NOR U28367 ( .A(n28140), .B(n28141), .Z(n28138) );
  XOR U28368 ( .A(n28142), .B(n28143), .Z(n26920) );
  ANDN U28369 ( .B(n26800), .A(n28144), .Z(n28142) );
  XNOR U28370 ( .A(n24721), .B(n28145), .Z(n28136) );
  XOR U28371 ( .A(n26077), .B(n24181), .Z(n28145) );
  XNOR U28372 ( .A(n28146), .B(n28147), .Z(n24181) );
  ANDN U28373 ( .B(n28148), .A(n28149), .Z(n28146) );
  XNOR U28374 ( .A(n28150), .B(n28151), .Z(n26077) );
  NOR U28375 ( .A(n26807), .B(n28152), .Z(n28150) );
  XNOR U28376 ( .A(n28153), .B(n28154), .Z(n24721) );
  NOR U28377 ( .A(n28155), .B(n28156), .Z(n28153) );
  XNOR U28378 ( .A(n28157), .B(n24946), .Z(n22237) );
  IV U28379 ( .A(n25805), .Z(n24946) );
  XOR U28380 ( .A(n28158), .B(n28159), .Z(n25805) );
  XOR U28381 ( .A(n28160), .B(n28161), .Z(n22911) );
  XOR U28382 ( .A(n17130), .B(n20067), .Z(n28161) );
  XOR U28383 ( .A(n28162), .B(n25633), .Z(n20067) );
  NOR U28384 ( .A(n22454), .B(n22453), .Z(n28162) );
  XOR U28385 ( .A(n26831), .B(n28163), .Z(n22453) );
  XNOR U28386 ( .A(n28164), .B(n28165), .Z(n26831) );
  ANDN U28387 ( .B(n28166), .A(n28167), .Z(n28164) );
  XOR U28388 ( .A(n28098), .B(n24366), .Z(n22454) );
  XNOR U28389 ( .A(n28168), .B(n28169), .Z(n28098) );
  NOR U28390 ( .A(n28170), .B(n28171), .Z(n28168) );
  XNOR U28391 ( .A(n28172), .B(n25635), .Z(n17130) );
  ANDN U28392 ( .B(n22463), .A(n22464), .Z(n28172) );
  XNOR U28393 ( .A(n26533), .B(n26620), .Z(n22464) );
  XOR U28394 ( .A(n28173), .B(n27558), .Z(n26533) );
  NOR U28395 ( .A(n28174), .B(n28175), .Z(n28173) );
  XOR U28396 ( .A(n25577), .B(n28176), .Z(n22463) );
  XNOR U28397 ( .A(n28039), .B(n26264), .Z(n25577) );
  XNOR U28398 ( .A(n28177), .B(n28178), .Z(n26264) );
  XNOR U28399 ( .A(n26509), .B(n25806), .Z(n28178) );
  XNOR U28400 ( .A(n28179), .B(n28180), .Z(n25806) );
  ANDN U28401 ( .B(n26303), .A(n28181), .Z(n28179) );
  XNOR U28402 ( .A(n28182), .B(n28183), .Z(n26509) );
  ANDN U28403 ( .B(n28184), .A(n26309), .Z(n28182) );
  IV U28404 ( .A(n28185), .Z(n26309) );
  XOR U28405 ( .A(n25279), .B(n28186), .Z(n28177) );
  XNOR U28406 ( .A(n24771), .B(n25052), .Z(n28186) );
  XNOR U28407 ( .A(n28187), .B(n28188), .Z(n25052) );
  XNOR U28408 ( .A(n28190), .B(n28191), .Z(n24771) );
  ANDN U28409 ( .B(n28192), .A(n28193), .Z(n28190) );
  XNOR U28410 ( .A(n28194), .B(n28195), .Z(n25279) );
  ANDN U28411 ( .B(n26299), .A(n28196), .Z(n28194) );
  XOR U28412 ( .A(n28197), .B(n28198), .Z(n28039) );
  XOR U28413 ( .A(n28199), .B(n26068), .Z(n28198) );
  XNOR U28414 ( .A(n28200), .B(n28201), .Z(n26068) );
  XOR U28415 ( .A(n23046), .B(n28204), .Z(n28197) );
  XNOR U28416 ( .A(n27871), .B(n22942), .Z(n28204) );
  XOR U28417 ( .A(n28205), .B(n27604), .Z(n22942) );
  ANDN U28418 ( .B(n28206), .A(n28207), .Z(n28205) );
  XNOR U28419 ( .A(n28208), .B(n27599), .Z(n27871) );
  NOR U28420 ( .A(n28209), .B(n28210), .Z(n28208) );
  XNOR U28421 ( .A(n28211), .B(n27591), .Z(n23046) );
  NOR U28422 ( .A(n28212), .B(n28213), .Z(n28211) );
  XOR U28423 ( .A(n17307), .B(n28214), .Z(n28160) );
  XNOR U28424 ( .A(n21502), .B(n17551), .Z(n28214) );
  XOR U28425 ( .A(n28215), .B(n25644), .Z(n17551) );
  NOR U28426 ( .A(n25645), .B(n22460), .Z(n28215) );
  XNOR U28427 ( .A(n24930), .B(n28216), .Z(n22460) );
  XOR U28428 ( .A(n28217), .B(n24397), .Z(n25645) );
  IV U28429 ( .A(n24281), .Z(n24397) );
  XNOR U28430 ( .A(n27486), .B(n27052), .Z(n24281) );
  XNOR U28431 ( .A(n28218), .B(n28219), .Z(n27052) );
  XNOR U28432 ( .A(n25283), .B(n27909), .Z(n28219) );
  XNOR U28433 ( .A(n28220), .B(n28221), .Z(n27909) );
  ANDN U28434 ( .B(n28222), .A(n28223), .Z(n28220) );
  XNOR U28435 ( .A(n28224), .B(n28225), .Z(n25283) );
  ANDN U28436 ( .B(n28226), .A(n28227), .Z(n28224) );
  XOR U28437 ( .A(n28228), .B(n28229), .Z(n28218) );
  XNOR U28438 ( .A(n25987), .B(n28230), .Z(n28229) );
  XOR U28439 ( .A(n28231), .B(n28232), .Z(n25987) );
  XOR U28440 ( .A(n28235), .B(n28236), .Z(n27486) );
  XOR U28441 ( .A(n26554), .B(n28237), .Z(n28236) );
  XNOR U28442 ( .A(n28238), .B(n28239), .Z(n26554) );
  AND U28443 ( .A(n28139), .B(n28141), .Z(n28238) );
  XNOR U28444 ( .A(n26002), .B(n28240), .Z(n28235) );
  XOR U28445 ( .A(n22819), .B(n28241), .Z(n28240) );
  XOR U28446 ( .A(n28242), .B(n26809), .Z(n22819) );
  AND U28447 ( .A(n28152), .B(n28151), .Z(n28242) );
  XOR U28448 ( .A(n28243), .B(n28244), .Z(n26002) );
  AND U28449 ( .A(n28154), .B(n28156), .Z(n28243) );
  XNOR U28450 ( .A(n28245), .B(n25638), .Z(n21502) );
  ANDN U28451 ( .B(n23206), .A(n28003), .Z(n28245) );
  XOR U28452 ( .A(n28246), .B(n22506), .Z(n28003) );
  IV U28453 ( .A(n25865), .Z(n22506) );
  XNOR U28454 ( .A(n28247), .B(n28248), .Z(n25968) );
  XOR U28455 ( .A(n24667), .B(n23722), .Z(n28248) );
  XOR U28456 ( .A(n28249), .B(n28250), .Z(n23722) );
  ANDN U28457 ( .B(n28251), .A(n28252), .Z(n28249) );
  XNOR U28458 ( .A(n28253), .B(n28254), .Z(n24667) );
  NOR U28459 ( .A(n28255), .B(n28256), .Z(n28253) );
  XOR U28460 ( .A(n26690), .B(n28257), .Z(n28247) );
  XNOR U28461 ( .A(n26767), .B(n23709), .Z(n28257) );
  XNOR U28462 ( .A(n28258), .B(n28259), .Z(n23709) );
  ANDN U28463 ( .B(n28260), .A(n28261), .Z(n28258) );
  XNOR U28464 ( .A(n28262), .B(n28263), .Z(n26767) );
  ANDN U28465 ( .B(n28264), .A(n28265), .Z(n28262) );
  XNOR U28466 ( .A(n28266), .B(n28267), .Z(n26690) );
  ANDN U28467 ( .B(n28268), .A(n28269), .Z(n28266) );
  XNOR U28468 ( .A(n27118), .B(n23029), .Z(n23206) );
  IV U28469 ( .A(n25182), .Z(n23029) );
  XOR U28470 ( .A(n28272), .B(n28273), .Z(n26350) );
  XNOR U28471 ( .A(n26635), .B(n28274), .Z(n28273) );
  XOR U28472 ( .A(n28275), .B(n28276), .Z(n26635) );
  ANDN U28473 ( .B(n27122), .A(n27120), .Z(n28275) );
  XOR U28474 ( .A(n24723), .B(n28277), .Z(n28272) );
  XNOR U28475 ( .A(n23999), .B(n26142), .Z(n28277) );
  XNOR U28476 ( .A(n28278), .B(n28279), .Z(n26142) );
  AND U28477 ( .A(n27109), .B(n27111), .Z(n28278) );
  XNOR U28478 ( .A(n28280), .B(n28281), .Z(n23999) );
  ANDN U28479 ( .B(n27113), .A(n27114), .Z(n28280) );
  XNOR U28480 ( .A(n28282), .B(n28283), .Z(n24723) );
  ANDN U28481 ( .B(n28129), .A(n28130), .Z(n28282) );
  XOR U28482 ( .A(n28284), .B(n28285), .Z(n27118) );
  NOR U28483 ( .A(n28286), .B(n28287), .Z(n28284) );
  XNOR U28484 ( .A(n28288), .B(n25641), .Z(n17307) );
  NOR U28485 ( .A(n22449), .B(n22450), .Z(n28288) );
  IV U28486 ( .A(n25642), .Z(n22449) );
  XOR U28487 ( .A(n26658), .B(n25942), .Z(n25642) );
  IV U28488 ( .A(n23019), .Z(n25942) );
  XNOR U28489 ( .A(n28292), .B(n28293), .Z(n26658) );
  ANDN U28490 ( .B(n28294), .A(n28295), .Z(n28292) );
  XOR U28491 ( .A(n17659), .B(n22750), .Z(n13501) );
  XNOR U28492 ( .A(n28296), .B(n21075), .Z(n22750) );
  ANDN U28493 ( .B(n22780), .A(n22779), .Z(n28296) );
  XNOR U28494 ( .A(n28297), .B(n23584), .Z(n22780) );
  XOR U28495 ( .A(n25875), .B(n21894), .Z(n17659) );
  XOR U28496 ( .A(n28298), .B(n28299), .Z(n21894) );
  XNOR U28497 ( .A(n18588), .B(n19029), .Z(n28299) );
  XNOR U28498 ( .A(n28300), .B(n21057), .Z(n19029) );
  XOR U28499 ( .A(n28301), .B(n23566), .Z(n21057) );
  XNOR U28500 ( .A(n28302), .B(n28012), .Z(n23566) );
  XOR U28501 ( .A(n28303), .B(n28304), .Z(n28012) );
  XNOR U28502 ( .A(n25492), .B(n25870), .Z(n28304) );
  XOR U28503 ( .A(n28305), .B(n28306), .Z(n25870) );
  ANDN U28504 ( .B(n28307), .A(n28308), .Z(n28305) );
  XNOR U28505 ( .A(n28309), .B(n28310), .Z(n25492) );
  ANDN U28506 ( .B(n28311), .A(n28312), .Z(n28309) );
  XOR U28507 ( .A(n28313), .B(n28314), .Z(n28303) );
  XNOR U28508 ( .A(n24394), .B(n25800), .Z(n28314) );
  XOR U28509 ( .A(n28315), .B(n28316), .Z(n25800) );
  NOR U28510 ( .A(n28317), .B(n28318), .Z(n28315) );
  XOR U28511 ( .A(n28319), .B(n28320), .Z(n24394) );
  ANDN U28512 ( .B(n28321), .A(n28322), .Z(n28319) );
  AND U28513 ( .A(n22772), .B(n21058), .Z(n28300) );
  XNOR U28514 ( .A(n28323), .B(n27796), .Z(n21058) );
  XOR U28515 ( .A(n28324), .B(n24408), .Z(n22772) );
  IV U28516 ( .A(n25170), .Z(n24408) );
  XNOR U28517 ( .A(n28325), .B(n28326), .Z(n27778) );
  XNOR U28518 ( .A(n28327), .B(n25541), .Z(n28326) );
  XNOR U28519 ( .A(n28328), .B(n27713), .Z(n25541) );
  ANDN U28520 ( .B(n28329), .A(n26686), .Z(n28328) );
  XNOR U28521 ( .A(n24210), .B(n28330), .Z(n28325) );
  XOR U28522 ( .A(n26134), .B(n28331), .Z(n28330) );
  ANDN U28523 ( .B(n26676), .A(n28333), .Z(n28332) );
  XOR U28524 ( .A(n28334), .B(n27710), .Z(n24210) );
  XOR U28525 ( .A(n28336), .B(n28337), .Z(n27202) );
  XNOR U28526 ( .A(n27872), .B(n28338), .Z(n28337) );
  XOR U28527 ( .A(n28339), .B(n28340), .Z(n27872) );
  ANDN U28528 ( .B(n28341), .A(n28342), .Z(n28339) );
  XOR U28529 ( .A(n25121), .B(n28343), .Z(n28336) );
  XOR U28530 ( .A(n22640), .B(n24820), .Z(n28343) );
  XNOR U28531 ( .A(n28344), .B(n28345), .Z(n24820) );
  AND U28532 ( .A(n28346), .B(n28347), .Z(n28344) );
  XNOR U28533 ( .A(n28348), .B(n28349), .Z(n22640) );
  XNOR U28534 ( .A(n28352), .B(n28353), .Z(n25121) );
  ANDN U28535 ( .B(n28354), .A(n28355), .Z(n28352) );
  XNOR U28536 ( .A(n28356), .B(n21049), .Z(n18588) );
  XOR U28537 ( .A(n24250), .B(n28357), .Z(n21049) );
  IV U28538 ( .A(n25490), .Z(n24250) );
  ANDN U28539 ( .B(n22765), .A(n21048), .Z(n28356) );
  XNOR U28540 ( .A(n25986), .B(n28228), .Z(n22765) );
  XNOR U28541 ( .A(n28359), .B(n28360), .Z(n28228) );
  NOR U28542 ( .A(n28361), .B(n28362), .Z(n28359) );
  XOR U28543 ( .A(n18922), .B(n28363), .Z(n28298) );
  XOR U28544 ( .A(n19613), .B(n15890), .Z(n28363) );
  XNOR U28545 ( .A(n28364), .B(n21061), .Z(n15890) );
  IV U28546 ( .A(n24207), .Z(n21061) );
  XOR U28547 ( .A(n28365), .B(n22960), .Z(n24207) );
  ANDN U28548 ( .B(n21062), .A(n22761), .Z(n28364) );
  XNOR U28549 ( .A(n28366), .B(n26280), .Z(n22761) );
  XNOR U28550 ( .A(n28367), .B(n28368), .Z(n27060) );
  XNOR U28551 ( .A(n23142), .B(n24184), .Z(n28368) );
  XNOR U28552 ( .A(n28369), .B(n28370), .Z(n24184) );
  XNOR U28553 ( .A(n28371), .B(n28372), .Z(n23142) );
  ANDN U28554 ( .B(n26598), .A(n26596), .Z(n28371) );
  XOR U28555 ( .A(n26095), .B(n28373), .Z(n28367) );
  XOR U28556 ( .A(n25955), .B(n28374), .Z(n28373) );
  XOR U28557 ( .A(n28375), .B(n28376), .Z(n25955) );
  ANDN U28558 ( .B(n26606), .A(n26607), .Z(n28375) );
  XNOR U28559 ( .A(n28377), .B(n28378), .Z(n26095) );
  ANDN U28560 ( .B(n27062), .A(n28379), .Z(n28377) );
  XOR U28561 ( .A(n28380), .B(n28381), .Z(n26119) );
  XOR U28562 ( .A(n26505), .B(n25723), .Z(n28381) );
  XOR U28563 ( .A(n28382), .B(n28383), .Z(n25723) );
  NOR U28564 ( .A(n27494), .B(n28384), .Z(n28382) );
  XOR U28565 ( .A(n28385), .B(n28386), .Z(n26505) );
  ANDN U28566 ( .B(n27490), .A(n28387), .Z(n28385) );
  XOR U28567 ( .A(n25406), .B(n28388), .Z(n28380) );
  XOR U28568 ( .A(n21220), .B(n25096), .Z(n28388) );
  XNOR U28569 ( .A(n28389), .B(n28390), .Z(n25096) );
  XNOR U28570 ( .A(n28392), .B(n28393), .Z(n21220) );
  ANDN U28571 ( .B(n28394), .A(n27499), .Z(n28392) );
  XOR U28572 ( .A(n28395), .B(n28396), .Z(n25406) );
  ANDN U28573 ( .B(n27507), .A(n28397), .Z(n28395) );
  XOR U28574 ( .A(n28015), .B(n21584), .Z(n21062) );
  XOR U28575 ( .A(n28398), .B(n26879), .Z(n21584) );
  XNOR U28576 ( .A(n28399), .B(n28400), .Z(n26879) );
  XNOR U28577 ( .A(n21386), .B(n28401), .Z(n28400) );
  XNOR U28578 ( .A(n28402), .B(n28403), .Z(n21386) );
  ANDN U28579 ( .B(n28404), .A(n28405), .Z(n28402) );
  XNOR U28580 ( .A(n26480), .B(n28406), .Z(n28399) );
  XOR U28581 ( .A(n28407), .B(n23516), .Z(n28406) );
  XNOR U28582 ( .A(n28408), .B(n28409), .Z(n23516) );
  ANDN U28583 ( .B(n28024), .A(n28022), .Z(n28408) );
  XOR U28584 ( .A(n28410), .B(n28411), .Z(n26480) );
  XNOR U28585 ( .A(n28412), .B(n28404), .Z(n28015) );
  ANDN U28586 ( .B(n28405), .A(n28413), .Z(n28412) );
  XOR U28587 ( .A(n28414), .B(n21052), .Z(n19613) );
  XNOR U28588 ( .A(n22495), .B(n28415), .Z(n21052) );
  ANDN U28589 ( .B(n22769), .A(n22768), .Z(n28414) );
  XOR U28590 ( .A(n26824), .B(n28163), .Z(n22768) );
  IV U28591 ( .A(n23869), .Z(n28163) );
  XNOR U28592 ( .A(n28418), .B(n28419), .Z(n26257) );
  XNOR U28593 ( .A(n26229), .B(n23857), .Z(n28419) );
  XOR U28594 ( .A(n28420), .B(n27893), .Z(n23857) );
  ANDN U28595 ( .B(n27184), .A(n27182), .Z(n28420) );
  XOR U28596 ( .A(n28421), .B(n28422), .Z(n27182) );
  XNOR U28597 ( .A(n28423), .B(n26903), .Z(n26229) );
  ANDN U28598 ( .B(n27180), .A(n26902), .Z(n28423) );
  XOR U28599 ( .A(n28424), .B(n28425), .Z(n26902) );
  XOR U28600 ( .A(n23874), .B(n28426), .Z(n28418) );
  XNOR U28601 ( .A(n24787), .B(n24252), .Z(n28426) );
  XOR U28602 ( .A(n28427), .B(n26898), .Z(n24252) );
  AND U28603 ( .A(n27188), .B(n26899), .Z(n28427) );
  XOR U28604 ( .A(n28428), .B(n28429), .Z(n26899) );
  XNOR U28605 ( .A(n28430), .B(n26889), .Z(n24787) );
  NOR U28606 ( .A(n26890), .B(n27193), .Z(n28430) );
  XOR U28607 ( .A(n28431), .B(n28432), .Z(n26890) );
  XNOR U28608 ( .A(n28433), .B(n28434), .Z(n23874) );
  ANDN U28609 ( .B(n27191), .A(n26894), .Z(n28433) );
  XOR U28610 ( .A(n28435), .B(n28436), .Z(n26894) );
  XNOR U28611 ( .A(n28437), .B(n28438), .Z(n27101) );
  XNOR U28612 ( .A(n25212), .B(n23716), .Z(n28438) );
  XNOR U28613 ( .A(n28439), .B(n28440), .Z(n23716) );
  NOR U28614 ( .A(n26834), .B(n26833), .Z(n28439) );
  XNOR U28615 ( .A(n28441), .B(n28442), .Z(n25212) );
  ANDN U28616 ( .B(n28443), .A(n28444), .Z(n28441) );
  XNOR U28617 ( .A(n26882), .B(n28445), .Z(n28437) );
  XOR U28618 ( .A(n25585), .B(n22226), .Z(n28445) );
  XOR U28619 ( .A(n28446), .B(n28447), .Z(n22226) );
  ANDN U28620 ( .B(n26828), .A(n26826), .Z(n28446) );
  XOR U28621 ( .A(n28448), .B(n28449), .Z(n25585) );
  XNOR U28622 ( .A(n28450), .B(n28451), .Z(n26882) );
  ANDN U28623 ( .B(n27332), .A(n28452), .Z(n28450) );
  XNOR U28624 ( .A(n28453), .B(n28443), .Z(n26824) );
  XNOR U28625 ( .A(n28374), .B(n24185), .Z(n22769) );
  XOR U28626 ( .A(n28455), .B(n26507), .Z(n24185) );
  XNOR U28627 ( .A(n28456), .B(n28457), .Z(n26507) );
  XNOR U28628 ( .A(n28458), .B(n27701), .Z(n28457) );
  XNOR U28629 ( .A(n28459), .B(n28460), .Z(n27701) );
  NOR U28630 ( .A(n28378), .B(n27062), .Z(n28459) );
  XNOR U28631 ( .A(n28461), .B(n28462), .Z(n27062) );
  IV U28632 ( .A(n28463), .Z(n28378) );
  XNOR U28633 ( .A(n26905), .B(n28464), .Z(n28456) );
  XOR U28634 ( .A(n28465), .B(n25290), .Z(n28464) );
  XOR U28635 ( .A(n28466), .B(n28467), .Z(n25290) );
  NOR U28636 ( .A(n26592), .B(n28370), .Z(n28466) );
  XOR U28637 ( .A(n28468), .B(n28469), .Z(n26592) );
  XNOR U28638 ( .A(n28470), .B(n28471), .Z(n26905) );
  ANDN U28639 ( .B(n26596), .A(n28372), .Z(n28470) );
  XOR U28640 ( .A(n28472), .B(n28473), .Z(n26596) );
  XOR U28641 ( .A(n28474), .B(n28475), .Z(n28374) );
  NOR U28642 ( .A(n26602), .B(n26603), .Z(n28474) );
  XNOR U28643 ( .A(n28476), .B(n21066), .Z(n18922) );
  IV U28644 ( .A(n27982), .Z(n21066) );
  XNOR U28645 ( .A(n28477), .B(n25424), .Z(n27982) );
  ANDN U28646 ( .B(n22777), .A(n21065), .Z(n28476) );
  IV U28647 ( .A(n22775), .Z(n21065) );
  XNOR U28648 ( .A(n28478), .B(n23708), .Z(n22775) );
  XOR U28649 ( .A(n28135), .B(n28479), .Z(n23708) );
  XOR U28650 ( .A(n28480), .B(n28481), .Z(n28135) );
  XNOR U28651 ( .A(n24396), .B(n25156), .Z(n28481) );
  XNOR U28652 ( .A(n28482), .B(n28483), .Z(n25156) );
  NOR U28653 ( .A(n28484), .B(n28485), .Z(n28482) );
  XNOR U28654 ( .A(n28486), .B(n28361), .Z(n24396) );
  ANDN U28655 ( .B(n28362), .A(n28487), .Z(n28486) );
  XOR U28656 ( .A(n25518), .B(n28488), .Z(n28480) );
  XNOR U28657 ( .A(n28217), .B(n24280), .Z(n28488) );
  XNOR U28658 ( .A(n28489), .B(n28234), .Z(n24280) );
  ANDN U28659 ( .B(n28490), .A(n28233), .Z(n28489) );
  XOR U28660 ( .A(n28491), .B(n28227), .Z(n28217) );
  NOR U28661 ( .A(n28492), .B(n28226), .Z(n28491) );
  XNOR U28662 ( .A(n28493), .B(n28222), .Z(n25518) );
  ANDN U28663 ( .B(n28223), .A(n28494), .Z(n28493) );
  XOR U28664 ( .A(n28495), .B(n24146), .Z(n22777) );
  XOR U28665 ( .A(n28496), .B(n28497), .Z(n25875) );
  XOR U28666 ( .A(n16619), .B(n17482), .Z(n28497) );
  XNOR U28667 ( .A(n28498), .B(n21072), .Z(n17482) );
  XNOR U28668 ( .A(n28499), .B(n24515), .Z(n21072) );
  IV U28669 ( .A(n23941), .Z(n24515) );
  XOR U28670 ( .A(n25967), .B(n25198), .Z(n23941) );
  XNOR U28671 ( .A(n28500), .B(n28501), .Z(n25198) );
  XOR U28672 ( .A(n26761), .B(n22957), .Z(n28501) );
  XOR U28673 ( .A(n28502), .B(n28503), .Z(n22957) );
  NOR U28674 ( .A(n28504), .B(n28505), .Z(n28502) );
  XOR U28675 ( .A(n28506), .B(n27480), .Z(n26761) );
  ANDN U28676 ( .B(n28507), .A(n28508), .Z(n28506) );
  XNOR U28677 ( .A(n25314), .B(n28509), .Z(n28500) );
  XNOR U28678 ( .A(n22403), .B(n28510), .Z(n28509) );
  XOR U28679 ( .A(n28511), .B(n27484), .Z(n22403) );
  ANDN U28680 ( .B(n28512), .A(n28513), .Z(n28511) );
  XOR U28681 ( .A(n28514), .B(n27476), .Z(n25314) );
  ANDN U28682 ( .B(n28515), .A(n28516), .Z(n28514) );
  XOR U28683 ( .A(n28517), .B(n28518), .Z(n25967) );
  XNOR U28684 ( .A(n25288), .B(n27734), .Z(n28518) );
  XNOR U28685 ( .A(n28519), .B(n28520), .Z(n27734) );
  ANDN U28686 ( .B(n28521), .A(n28522), .Z(n28519) );
  XNOR U28687 ( .A(n28523), .B(n28524), .Z(n25288) );
  XOR U28688 ( .A(n28216), .B(n28527), .Z(n28517) );
  XNOR U28689 ( .A(n28528), .B(n24931), .Z(n28527) );
  XOR U28690 ( .A(n28529), .B(n28530), .Z(n24931) );
  ANDN U28691 ( .B(n28531), .A(n28532), .Z(n28529) );
  XNOR U28692 ( .A(n28533), .B(n28534), .Z(n28216) );
  ANDN U28693 ( .B(n28535), .A(n28536), .Z(n28533) );
  NOR U28694 ( .A(n21122), .B(n21071), .Z(n28498) );
  XOR U28695 ( .A(n28537), .B(n28538), .Z(n21071) );
  XOR U28696 ( .A(n28539), .B(n21372), .Z(n21122) );
  XNOR U28697 ( .A(n28540), .B(n24190), .Z(n16619) );
  XOR U28698 ( .A(n24755), .B(n28541), .Z(n24190) );
  IV U28699 ( .A(n23737), .Z(n24755) );
  XOR U28700 ( .A(n28542), .B(n28543), .Z(n23737) );
  ANDN U28701 ( .B(n22779), .A(n21075), .Z(n28540) );
  XOR U28702 ( .A(n27295), .B(n25043), .Z(n21075) );
  IV U28703 ( .A(n25079), .Z(n25043) );
  XNOR U28704 ( .A(n28544), .B(n28545), .Z(n26378) );
  XNOR U28705 ( .A(n27260), .B(n23947), .Z(n28545) );
  XOR U28706 ( .A(n28546), .B(n28547), .Z(n23947) );
  XNOR U28707 ( .A(n28548), .B(n28549), .Z(n27260) );
  ANDN U28708 ( .B(n27291), .A(n27293), .Z(n28548) );
  XNOR U28709 ( .A(n26626), .B(n28550), .Z(n28544) );
  XNOR U28710 ( .A(n24789), .B(n27512), .Z(n28550) );
  XNOR U28711 ( .A(n28551), .B(n28552), .Z(n27512) );
  NOR U28712 ( .A(n28553), .B(n28554), .Z(n28551) );
  XOR U28713 ( .A(n28555), .B(n28556), .Z(n24789) );
  ANDN U28714 ( .B(n27289), .A(n28557), .Z(n28555) );
  IV U28715 ( .A(n28558), .Z(n27289) );
  XNOR U28716 ( .A(n28559), .B(n28560), .Z(n26626) );
  ANDN U28717 ( .B(n27301), .A(n27302), .Z(n28559) );
  XOR U28718 ( .A(n28561), .B(n28562), .Z(n26342) );
  XOR U28719 ( .A(n25482), .B(n24810), .Z(n28562) );
  XOR U28720 ( .A(n28563), .B(n27952), .Z(n24810) );
  XNOR U28721 ( .A(n28564), .B(n28565), .Z(n25482) );
  NOR U28722 ( .A(n27818), .B(n27532), .Z(n28564) );
  IV U28723 ( .A(n28566), .Z(n27818) );
  XOR U28724 ( .A(n25899), .B(n28567), .Z(n28561) );
  XOR U28725 ( .A(n26762), .B(n23863), .Z(n28567) );
  XNOR U28726 ( .A(n28568), .B(n27519), .Z(n23863) );
  NOR U28727 ( .A(n27821), .B(n27518), .Z(n28568) );
  XNOR U28728 ( .A(n28569), .B(n27522), .Z(n26762) );
  ANDN U28729 ( .B(n28570), .A(n27523), .Z(n28569) );
  XOR U28730 ( .A(n28571), .B(n27529), .Z(n25899) );
  ANDN U28731 ( .B(n27528), .A(n27824), .Z(n28571) );
  XNOR U28732 ( .A(n28572), .B(n28553), .Z(n27295) );
  AND U28733 ( .A(n28573), .B(n28554), .Z(n28572) );
  XOR U28734 ( .A(n28574), .B(n21606), .Z(n22779) );
  XOR U28735 ( .A(n28575), .B(n28576), .Z(n27240) );
  XOR U28736 ( .A(n23726), .B(n24746), .Z(n28576) );
  XOR U28737 ( .A(n28577), .B(n28578), .Z(n24746) );
  ANDN U28738 ( .B(n28579), .A(n27275), .Z(n28577) );
  XNOR U28739 ( .A(n28580), .B(n28581), .Z(n23726) );
  AND U28740 ( .A(n27269), .B(n28582), .Z(n28580) );
  XOR U28741 ( .A(n28583), .B(n28584), .Z(n28575) );
  XOR U28742 ( .A(n25483), .B(n26131), .Z(n28584) );
  XNOR U28743 ( .A(n28585), .B(n28586), .Z(n26131) );
  ANDN U28744 ( .B(n27279), .A(n28587), .Z(n28585) );
  XNOR U28745 ( .A(n28588), .B(n28589), .Z(n25483) );
  ANDN U28746 ( .B(n28590), .A(n27671), .Z(n28588) );
  IV U28747 ( .A(n28591), .Z(n27671) );
  XOR U28748 ( .A(n28592), .B(n28593), .Z(n27955) );
  XNOR U28749 ( .A(n21832), .B(n22310), .Z(n28593) );
  XNOR U28750 ( .A(n28594), .B(n27093), .Z(n22310) );
  AND U28751 ( .A(n27094), .B(n28595), .Z(n28594) );
  XNOR U28752 ( .A(n28596), .B(n27081), .Z(n21832) );
  AND U28753 ( .A(n28597), .B(n27080), .Z(n28596) );
  XOR U28754 ( .A(n26003), .B(n28598), .Z(n28592) );
  XNOR U28755 ( .A(n23331), .B(n25665), .Z(n28598) );
  XOR U28756 ( .A(n28599), .B(n27090), .Z(n25665) );
  ANDN U28757 ( .B(n28600), .A(n27089), .Z(n28599) );
  XNOR U28758 ( .A(n28601), .B(n28602), .Z(n23331) );
  ANDN U28759 ( .B(n28603), .A(n28604), .Z(n28601) );
  XOR U28760 ( .A(n28605), .B(n27085), .Z(n26003) );
  XNOR U28761 ( .A(n16514), .B(n28607), .Z(n28496) );
  XNOR U28762 ( .A(n16109), .B(n21043), .Z(n28607) );
  XNOR U28763 ( .A(n28608), .B(n21082), .Z(n21043) );
  XNOR U28764 ( .A(n28092), .B(n24366), .Z(n21082) );
  IV U28765 ( .A(n26907), .Z(n24366) );
  XNOR U28766 ( .A(n26290), .B(n27875), .Z(n26907) );
  XNOR U28767 ( .A(n28609), .B(n28610), .Z(n27875) );
  XOR U28768 ( .A(n26023), .B(n25162), .Z(n28610) );
  XNOR U28769 ( .A(n28611), .B(n28612), .Z(n25162) );
  AND U28770 ( .A(n28613), .B(n28614), .Z(n28611) );
  XNOR U28771 ( .A(n28615), .B(n28616), .Z(n26023) );
  ANDN U28772 ( .B(n28094), .A(n28095), .Z(n28615) );
  XNOR U28773 ( .A(n26266), .B(n28617), .Z(n28609) );
  XOR U28774 ( .A(n23828), .B(n28618), .Z(n28617) );
  XOR U28775 ( .A(n28619), .B(n28620), .Z(n23828) );
  ANDN U28776 ( .B(n28171), .A(n28621), .Z(n28619) );
  XNOR U28777 ( .A(n28622), .B(n28623), .Z(n26266) );
  ANDN U28778 ( .B(n28104), .A(n28105), .Z(n28622) );
  XOR U28779 ( .A(n28624), .B(n28625), .Z(n26290) );
  XNOR U28780 ( .A(n28626), .B(n24038), .Z(n28625) );
  XOR U28781 ( .A(n28627), .B(n28628), .Z(n24038) );
  XOR U28782 ( .A(n22353), .B(n28631), .Z(n28624) );
  XOR U28783 ( .A(n26148), .B(n27383), .Z(n28631) );
  XNOR U28784 ( .A(n28632), .B(n28633), .Z(n27383) );
  ANDN U28785 ( .B(n28634), .A(n28635), .Z(n28632) );
  XNOR U28786 ( .A(n28636), .B(n28637), .Z(n26148) );
  AND U28787 ( .A(n28638), .B(n28639), .Z(n28636) );
  XNOR U28788 ( .A(n28640), .B(n28641), .Z(n22353) );
  ANDN U28789 ( .B(n28642), .A(n28643), .Z(n28640) );
  XNOR U28790 ( .A(n28644), .B(n28614), .Z(n28092) );
  NOR U28791 ( .A(n28645), .B(n28613), .Z(n28644) );
  ANDN U28792 ( .B(n21081), .A(n21127), .Z(n28608) );
  XOR U28793 ( .A(n27967), .B(n27723), .Z(n21127) );
  XNOR U28794 ( .A(n28646), .B(n28647), .Z(n27967) );
  NOR U28795 ( .A(n28648), .B(n28649), .Z(n28646) );
  XOR U28796 ( .A(n25414), .B(n28650), .Z(n21081) );
  XOR U28797 ( .A(n28651), .B(n28652), .Z(n25414) );
  XNOR U28798 ( .A(n28653), .B(n21086), .Z(n16109) );
  XNOR U28799 ( .A(n27144), .B(n23050), .Z(n21086) );
  XOR U28800 ( .A(n28008), .B(n28654), .Z(n23050) );
  XOR U28801 ( .A(n28655), .B(n28656), .Z(n28008) );
  XOR U28802 ( .A(n26973), .B(n27197), .Z(n28656) );
  XOR U28803 ( .A(n28657), .B(n28658), .Z(n27197) );
  NOR U28804 ( .A(n27161), .B(n27159), .Z(n28657) );
  XNOR U28805 ( .A(n28659), .B(n28660), .Z(n26973) );
  ANDN U28806 ( .B(n27156), .A(n28661), .Z(n28659) );
  XNOR U28807 ( .A(n24961), .B(n28662), .Z(n28655) );
  XOR U28808 ( .A(n26058), .B(n24760), .Z(n28662) );
  XNOR U28809 ( .A(n28663), .B(n28664), .Z(n24760) );
  NOR U28810 ( .A(n28665), .B(n27152), .Z(n28663) );
  XNOR U28811 ( .A(n28666), .B(n28667), .Z(n26058) );
  ANDN U28812 ( .B(n27147), .A(n27146), .Z(n28666) );
  XNOR U28813 ( .A(n28668), .B(n28669), .Z(n24961) );
  ANDN U28814 ( .B(n28670), .A(n28671), .Z(n28668) );
  XNOR U28815 ( .A(n28672), .B(n28673), .Z(n27144) );
  NOR U28816 ( .A(n28670), .B(n28674), .Z(n28672) );
  ANDN U28817 ( .B(n21119), .A(n21085), .Z(n28653) );
  XOR U28818 ( .A(n28675), .B(n24798), .Z(n21085) );
  XOR U28819 ( .A(n28416), .B(n27408), .Z(n24798) );
  XNOR U28820 ( .A(n28676), .B(n28677), .Z(n27408) );
  XNOR U28821 ( .A(n28678), .B(n25838), .Z(n28677) );
  XNOR U28822 ( .A(n28679), .B(n28680), .Z(n25838) );
  ANDN U28823 ( .B(n28681), .A(n28682), .Z(n28679) );
  XOR U28824 ( .A(n25221), .B(n28683), .Z(n28676) );
  XOR U28825 ( .A(n27009), .B(n26696), .Z(n28683) );
  XNOR U28826 ( .A(n28684), .B(n28685), .Z(n26696) );
  NOR U28827 ( .A(n28686), .B(n28687), .Z(n28684) );
  XNOR U28828 ( .A(n28688), .B(n28689), .Z(n27009) );
  ANDN U28829 ( .B(n28690), .A(n28691), .Z(n28688) );
  XNOR U28830 ( .A(n28692), .B(n28693), .Z(n25221) );
  ANDN U28831 ( .B(n28694), .A(n28695), .Z(n28692) );
  XOR U28832 ( .A(n28696), .B(n28697), .Z(n28416) );
  XOR U28833 ( .A(n23481), .B(n24276), .Z(n28697) );
  XNOR U28834 ( .A(n28698), .B(n25534), .Z(n24276) );
  AND U28835 ( .A(n27257), .B(n25535), .Z(n28698) );
  XOR U28836 ( .A(n28699), .B(n28700), .Z(n23481) );
  NOR U28837 ( .A(n27330), .B(n27249), .Z(n28699) );
  XOR U28838 ( .A(n25520), .B(n28701), .Z(n28696) );
  XOR U28839 ( .A(n23706), .B(n25058), .Z(n28701) );
  XNOR U28840 ( .A(n28702), .B(n27885), .Z(n25058) );
  ANDN U28841 ( .B(n27886), .A(n27253), .Z(n28702) );
  IV U28842 ( .A(n28703), .Z(n27253) );
  XNOR U28843 ( .A(n28704), .B(n26990), .Z(n23706) );
  ANDN U28844 ( .B(n26991), .A(n27245), .Z(n28704) );
  XNOR U28845 ( .A(n28705), .B(n25531), .Z(n25520) );
  NOR U28846 ( .A(n28706), .B(n25530), .Z(n28705) );
  XOR U28847 ( .A(n28707), .B(n23333), .Z(n21119) );
  IV U28848 ( .A(n23839), .Z(n23333) );
  XNOR U28849 ( .A(n28708), .B(n24198), .Z(n16514) );
  XNOR U28850 ( .A(n28709), .B(n28710), .Z(n24198) );
  NOR U28851 ( .A(n21130), .B(n22757), .Z(n28708) );
  XOR U28852 ( .A(n28711), .B(n23810), .Z(n22757) );
  XOR U28853 ( .A(n28712), .B(n23250), .Z(n21130) );
  XNOR U28854 ( .A(n28715), .B(n14724), .Z(n11113) );
  XOR U28855 ( .A(n20363), .B(n18326), .Z(n14724) );
  XOR U28856 ( .A(n22258), .B(n20481), .Z(n18326) );
  XOR U28857 ( .A(n28716), .B(n28717), .Z(n20481) );
  XNOR U28858 ( .A(n14171), .B(n18304), .Z(n28717) );
  XNOR U28859 ( .A(n28718), .B(n22933), .Z(n18304) );
  XOR U28860 ( .A(n28719), .B(n27228), .Z(n22933) );
  NOR U28861 ( .A(n18849), .B(n20753), .Z(n28718) );
  XOR U28862 ( .A(n24288), .B(n27648), .Z(n20753) );
  XNOR U28863 ( .A(n28720), .B(n28721), .Z(n27648) );
  AND U28864 ( .A(n27137), .B(n27665), .Z(n28720) );
  XOR U28865 ( .A(n28722), .B(n28723), .Z(n27137) );
  IV U28866 ( .A(n25488), .Z(n24288) );
  XNOR U28867 ( .A(n28724), .B(n24374), .Z(n18849) );
  IV U28868 ( .A(n28725), .Z(n24374) );
  XNOR U28869 ( .A(n28726), .B(n20188), .Z(n14171) );
  XOR U28870 ( .A(n26803), .B(n24998), .Z(n20188) );
  XNOR U28871 ( .A(n28727), .B(n28728), .Z(n26803) );
  ANDN U28872 ( .B(n28729), .A(n28244), .Z(n28727) );
  AND U28873 ( .A(n20187), .B(n20748), .Z(n28726) );
  XOR U28874 ( .A(n24836), .B(n28730), .Z(n20748) );
  XNOR U28875 ( .A(n28731), .B(n26543), .Z(n24836) );
  XNOR U28876 ( .A(n28732), .B(n28733), .Z(n26543) );
  XNOR U28877 ( .A(n26250), .B(n25729), .Z(n28733) );
  XNOR U28878 ( .A(n28734), .B(n26603), .Z(n25729) );
  XOR U28879 ( .A(n28735), .B(n28736), .Z(n26603) );
  XOR U28880 ( .A(n28738), .B(n26598), .Z(n26250) );
  XOR U28881 ( .A(n28739), .B(n28740), .Z(n26598) );
  ANDN U28882 ( .B(n26597), .A(n28471), .Z(n28738) );
  XOR U28883 ( .A(n24612), .B(n28741), .Z(n28732) );
  XOR U28884 ( .A(n25576), .B(n24073), .Z(n28741) );
  XOR U28885 ( .A(n28742), .B(n26593), .Z(n24073) );
  XNOR U28886 ( .A(n28743), .B(n28744), .Z(n26593) );
  XNOR U28887 ( .A(n28745), .B(n28379), .Z(n25576) );
  IV U28888 ( .A(n27064), .Z(n28379) );
  XOR U28889 ( .A(n28746), .B(n28747), .Z(n27064) );
  NOR U28890 ( .A(n27063), .B(n28460), .Z(n28745) );
  XNOR U28891 ( .A(n28748), .B(n26607), .Z(n24612) );
  XOR U28892 ( .A(n28749), .B(n28750), .Z(n26607) );
  ANDN U28893 ( .B(n26608), .A(n28751), .Z(n28748) );
  XOR U28894 ( .A(n28752), .B(n24709), .Z(n20187) );
  IV U28895 ( .A(n23983), .Z(n24709) );
  XOR U28896 ( .A(n28753), .B(n27890), .Z(n23983) );
  XNOR U28897 ( .A(n28754), .B(n28755), .Z(n27890) );
  XNOR U28898 ( .A(n22007), .B(n28756), .Z(n28755) );
  XOR U28899 ( .A(n28757), .B(n27183), .Z(n22007) );
  AND U28900 ( .A(n27893), .B(n27892), .Z(n28757) );
  XOR U28901 ( .A(n28758), .B(n28759), .Z(n27893) );
  XNOR U28902 ( .A(n28709), .B(n28760), .Z(n28754) );
  XNOR U28903 ( .A(n26750), .B(n25417), .Z(n28760) );
  XOR U28904 ( .A(n28761), .B(n27194), .Z(n25417) );
  NOR U28905 ( .A(n26888), .B(n26889), .Z(n28761) );
  XOR U28906 ( .A(n28762), .B(n28763), .Z(n26889) );
  XNOR U28907 ( .A(n28764), .B(n27187), .Z(n26750) );
  ANDN U28908 ( .B(n26897), .A(n26898), .Z(n28764) );
  XOR U28909 ( .A(n28765), .B(n28766), .Z(n26898) );
  XNOR U28910 ( .A(n28767), .B(n27179), .Z(n28709) );
  ANDN U28911 ( .B(n26901), .A(n26903), .Z(n28767) );
  XOR U28912 ( .A(n28768), .B(n28769), .Z(n26903) );
  XOR U28913 ( .A(n17435), .B(n28770), .Z(n28716) );
  XOR U28914 ( .A(n17949), .B(n18341), .Z(n28770) );
  XNOR U28915 ( .A(n28771), .B(n20178), .Z(n18341) );
  XOR U28916 ( .A(n24484), .B(n28772), .Z(n20178) );
  ANDN U28917 ( .B(n20177), .A(n18910), .Z(n28771) );
  XNOR U28918 ( .A(n21385), .B(n28401), .Z(n18910) );
  XOR U28919 ( .A(n28773), .B(n28774), .Z(n28401) );
  AND U28920 ( .A(n28026), .B(n28028), .Z(n28773) );
  XOR U28921 ( .A(n26733), .B(n22988), .Z(n20177) );
  XNOR U28922 ( .A(n28775), .B(n28776), .Z(n26733) );
  ANDN U28923 ( .B(n27835), .A(n27833), .Z(n28775) );
  XNOR U28924 ( .A(n28777), .B(n20184), .Z(n17949) );
  XNOR U28925 ( .A(n28778), .B(n26749), .Z(n20184) );
  IV U28926 ( .A(n24411), .Z(n26749) );
  XOR U28927 ( .A(n28779), .B(n28780), .Z(n24411) );
  NOR U28928 ( .A(n18845), .B(n20183), .Z(n28777) );
  XNOR U28929 ( .A(n26089), .B(n28781), .Z(n20183) );
  XOR U28930 ( .A(n22636), .B(n27273), .Z(n18845) );
  XNOR U28931 ( .A(n28782), .B(n28783), .Z(n27273) );
  ANDN U28932 ( .B(n28784), .A(n28785), .Z(n28782) );
  IV U28933 ( .A(n26454), .Z(n22636) );
  XOR U28934 ( .A(n28786), .B(n27888), .Z(n26454) );
  XOR U28935 ( .A(n28787), .B(n28788), .Z(n27888) );
  XNOR U28936 ( .A(n23851), .B(n24419), .Z(n28788) );
  XNOR U28937 ( .A(n28789), .B(n27254), .Z(n24419) );
  ANDN U28938 ( .B(n27255), .A(n27885), .Z(n28789) );
  XOR U28939 ( .A(n28790), .B(n28791), .Z(n27885) );
  XOR U28940 ( .A(n28792), .B(n28793), .Z(n27255) );
  XNOR U28941 ( .A(n28794), .B(n27246), .Z(n23851) );
  ANDN U28942 ( .B(n26989), .A(n26990), .Z(n28794) );
  XOR U28943 ( .A(n28795), .B(n28796), .Z(n26990) );
  XOR U28944 ( .A(n28797), .B(n28798), .Z(n26989) );
  XNOR U28945 ( .A(n24591), .B(n28799), .Z(n28787) );
  XNOR U28946 ( .A(n25313), .B(n26615), .Z(n28799) );
  XOR U28947 ( .A(n28800), .B(n27258), .Z(n26615) );
  NOR U28948 ( .A(n25534), .B(n25533), .Z(n28800) );
  XOR U28949 ( .A(n28801), .B(n28802), .Z(n25533) );
  XOR U28950 ( .A(n28803), .B(n28804), .Z(n25534) );
  XNOR U28951 ( .A(n28805), .B(n28806), .Z(n25313) );
  XOR U28952 ( .A(n28807), .B(n28808), .Z(n25531) );
  XOR U28953 ( .A(n28809), .B(n27251), .Z(n24591) );
  IV U28954 ( .A(n28810), .Z(n27251) );
  NOR U28955 ( .A(n27329), .B(n27250), .Z(n28809) );
  XNOR U28956 ( .A(n28811), .B(n28812), .Z(n27250) );
  IV U28957 ( .A(n28700), .Z(n27329) );
  XOR U28958 ( .A(n28813), .B(n28814), .Z(n28700) );
  XNOR U28959 ( .A(n28815), .B(n20175), .Z(n17435) );
  XOR U28960 ( .A(n28816), .B(n24228), .Z(n20175) );
  XOR U28961 ( .A(n25812), .B(n26693), .Z(n24228) );
  XNOR U28962 ( .A(n28817), .B(n28818), .Z(n26693) );
  XNOR U28963 ( .A(n26759), .B(n25475), .Z(n28818) );
  XNOR U28964 ( .A(n28819), .B(n28405), .Z(n25475) );
  XOR U28965 ( .A(n28820), .B(n28821), .Z(n28405) );
  XOR U28966 ( .A(n28823), .B(n28024), .Z(n26759) );
  XNOR U28967 ( .A(n28824), .B(n28825), .Z(n28024) );
  AND U28968 ( .A(n28023), .B(n28826), .Z(n28823) );
  XOR U28969 ( .A(n25818), .B(n28827), .Z(n28817) );
  XNOR U28970 ( .A(n25717), .B(n28011), .Z(n28827) );
  XOR U28971 ( .A(n28828), .B(n28032), .Z(n28011) );
  ANDN U28972 ( .B(n28829), .A(n28031), .Z(n28828) );
  XOR U28973 ( .A(n28830), .B(n28028), .Z(n25717) );
  XNOR U28974 ( .A(n28831), .B(n28832), .Z(n28028) );
  AND U28975 ( .A(n28027), .B(n28833), .Z(n28830) );
  XNOR U28976 ( .A(n28834), .B(n28019), .Z(n25818) );
  XOR U28977 ( .A(n28835), .B(n28836), .Z(n28019) );
  NOR U28978 ( .A(n28018), .B(n28837), .Z(n28834) );
  XOR U28979 ( .A(n28838), .B(n28839), .Z(n25812) );
  XOR U28980 ( .A(n26070), .B(n21226), .Z(n28839) );
  XNOR U28981 ( .A(n28840), .B(n28841), .Z(n21226) );
  ANDN U28982 ( .B(n28842), .A(n28843), .Z(n28840) );
  XNOR U28983 ( .A(n28844), .B(n28845), .Z(n26070) );
  NOR U28984 ( .A(n28846), .B(n28847), .Z(n28844) );
  XNOR U28985 ( .A(n26371), .B(n28848), .Z(n28838) );
  XOR U28986 ( .A(n24413), .B(n25772), .Z(n28848) );
  XNOR U28987 ( .A(n28849), .B(n28850), .Z(n25772) );
  NOR U28988 ( .A(n28851), .B(n28852), .Z(n28849) );
  XNOR U28989 ( .A(n28853), .B(n28854), .Z(n24413) );
  ANDN U28990 ( .B(n28855), .A(n28856), .Z(n28853) );
  XNOR U28991 ( .A(n28857), .B(n28858), .Z(n26371) );
  ANDN U28992 ( .B(n28859), .A(n28860), .Z(n28857) );
  ANDN U28993 ( .B(n19729), .A(n20174), .Z(n28815) );
  XOR U28994 ( .A(n26568), .B(n27567), .Z(n20174) );
  XNOR U28995 ( .A(n28861), .B(n28862), .Z(n27567) );
  ANDN U28996 ( .B(n28863), .A(n28864), .Z(n28861) );
  XOR U28997 ( .A(n28865), .B(n24506), .Z(n19729) );
  XOR U28998 ( .A(n28866), .B(n28867), .Z(n22258) );
  XNOR U28999 ( .A(n18891), .B(n18259), .Z(n28867) );
  XNOR U29000 ( .A(n28868), .B(n21233), .Z(n18259) );
  XOR U29001 ( .A(n23695), .B(n26844), .Z(n21233) );
  XOR U29002 ( .A(n28869), .B(n26106), .Z(n26844) );
  XNOR U29003 ( .A(n28870), .B(n26719), .Z(n23695) );
  XNOR U29004 ( .A(n28871), .B(n28872), .Z(n26719) );
  XNOR U29005 ( .A(n24818), .B(n24559), .Z(n28872) );
  XOR U29006 ( .A(n28873), .B(n25862), .Z(n24559) );
  NOR U29007 ( .A(n27457), .B(n25861), .Z(n28873) );
  XNOR U29008 ( .A(n28874), .B(n28875), .Z(n25861) );
  XOR U29009 ( .A(n28876), .B(n28759), .Z(n27457) );
  XNOR U29010 ( .A(n28877), .B(n26105), .Z(n24818) );
  ANDN U29011 ( .B(n26106), .A(n27461), .Z(n28877) );
  XOR U29012 ( .A(n28878), .B(n28879), .Z(n27461) );
  XNOR U29013 ( .A(n28880), .B(n28881), .Z(n26106) );
  XOR U29014 ( .A(n22222), .B(n28882), .Z(n28871) );
  XOR U29015 ( .A(n24781), .B(n25197), .Z(n28882) );
  XNOR U29016 ( .A(n28883), .B(n25857), .Z(n25197) );
  NOR U29017 ( .A(n26850), .B(n26852), .Z(n28883) );
  XNOR U29018 ( .A(n28884), .B(n28885), .Z(n26852) );
  XNOR U29019 ( .A(n28886), .B(n28887), .Z(n26850) );
  XNOR U29020 ( .A(n28888), .B(n25847), .Z(n24781) );
  ANDN U29021 ( .B(n26859), .A(n26857), .Z(n28888) );
  IV U29022 ( .A(n25848), .Z(n26857) );
  XNOR U29023 ( .A(n28889), .B(n28890), .Z(n25848) );
  XNOR U29024 ( .A(n28891), .B(n28892), .Z(n26859) );
  XNOR U29025 ( .A(n28893), .B(n25852), .Z(n22222) );
  NOR U29026 ( .A(n26847), .B(n25851), .Z(n28893) );
  XOR U29027 ( .A(n28894), .B(n28895), .Z(n25851) );
  XOR U29028 ( .A(n28896), .B(n28897), .Z(n26847) );
  ANDN U29029 ( .B(n19885), .A(n21237), .Z(n28868) );
  XNOR U29030 ( .A(n28898), .B(n20169), .Z(n18891) );
  XOR U29031 ( .A(n28899), .B(n28900), .Z(n20169) );
  ANDN U29032 ( .B(n19898), .A(n20365), .Z(n28898) );
  IV U29033 ( .A(n20170), .Z(n20365) );
  XOR U29034 ( .A(n25001), .B(n28901), .Z(n20170) );
  XNOR U29035 ( .A(n27035), .B(n28902), .Z(n25001) );
  XOR U29036 ( .A(n28903), .B(n28904), .Z(n27035) );
  XOR U29037 ( .A(n25284), .B(n23693), .Z(n28904) );
  XNOR U29038 ( .A(n28905), .B(n28906), .Z(n23693) );
  NOR U29039 ( .A(n28907), .B(n28908), .Z(n28905) );
  XOR U29040 ( .A(n28909), .B(n28910), .Z(n25284) );
  NOR U29041 ( .A(n28911), .B(n28912), .Z(n28909) );
  XOR U29042 ( .A(n23621), .B(n28913), .Z(n28903) );
  XNOR U29043 ( .A(n23012), .B(n28914), .Z(n28913) );
  XOR U29044 ( .A(n28915), .B(n28916), .Z(n23012) );
  ANDN U29045 ( .B(n28917), .A(n28918), .Z(n28915) );
  XOR U29046 ( .A(n28919), .B(n28920), .Z(n23621) );
  ANDN U29047 ( .B(n28921), .A(n28922), .Z(n28919) );
  XOR U29048 ( .A(n28923), .B(n22825), .Z(n19898) );
  XOR U29049 ( .A(n27198), .B(n27580), .Z(n22825) );
  XNOR U29050 ( .A(n28924), .B(n28925), .Z(n27580) );
  XNOR U29051 ( .A(n23058), .B(n28926), .Z(n28925) );
  XNOR U29052 ( .A(n28927), .B(n28928), .Z(n23058) );
  NOR U29053 ( .A(n28929), .B(n28930), .Z(n28927) );
  XOR U29054 ( .A(n24866), .B(n28931), .Z(n28924) );
  XOR U29055 ( .A(n26087), .B(n26234), .Z(n28931) );
  XNOR U29056 ( .A(n28932), .B(n28933), .Z(n26234) );
  NOR U29057 ( .A(n28934), .B(n28935), .Z(n28932) );
  XNOR U29058 ( .A(n28936), .B(n28937), .Z(n26087) );
  NOR U29059 ( .A(n28938), .B(n28939), .Z(n28936) );
  XNOR U29060 ( .A(n28940), .B(n28941), .Z(n24866) );
  XOR U29061 ( .A(n28944), .B(n28945), .Z(n27198) );
  XNOR U29062 ( .A(n28946), .B(n27919), .Z(n28945) );
  XOR U29063 ( .A(n28947), .B(n27839), .Z(n27919) );
  ANDN U29064 ( .B(n28948), .A(n28949), .Z(n28947) );
  XOR U29065 ( .A(n24401), .B(n28950), .Z(n28944) );
  XNOR U29066 ( .A(n24295), .B(n27033), .Z(n28950) );
  XOR U29067 ( .A(n28951), .B(n28952), .Z(n27033) );
  NOR U29068 ( .A(n28953), .B(n26745), .Z(n28951) );
  XNOR U29069 ( .A(n28954), .B(n27842), .Z(n24295) );
  AND U29070 ( .A(n28955), .B(n26735), .Z(n28954) );
  XNOR U29071 ( .A(n28956), .B(n27834), .Z(n24401) );
  ANDN U29072 ( .B(n28957), .A(n28776), .Z(n28956) );
  XOR U29073 ( .A(n17794), .B(n28958), .Z(n28866) );
  XOR U29074 ( .A(n20156), .B(n19067), .Z(n28958) );
  XNOR U29075 ( .A(n28959), .B(n21141), .Z(n19067) );
  XOR U29076 ( .A(n26955), .B(n22951), .Z(n21141) );
  IV U29077 ( .A(n25305), .Z(n22951) );
  XOR U29078 ( .A(n28960), .B(n26408), .Z(n25305) );
  XNOR U29079 ( .A(n28961), .B(n28962), .Z(n26408) );
  XNOR U29080 ( .A(n24920), .B(n25894), .Z(n28962) );
  XNOR U29081 ( .A(n28963), .B(n28175), .Z(n25894) );
  ANDN U29082 ( .B(n27559), .A(n27557), .Z(n28963) );
  XOR U29083 ( .A(n28964), .B(n28965), .Z(n24920) );
  XOR U29084 ( .A(n26814), .B(n28966), .Z(n28961) );
  XOR U29085 ( .A(n24460), .B(n24627), .Z(n28966) );
  XNOR U29086 ( .A(n28967), .B(n26624), .Z(n24627) );
  IV U29087 ( .A(n28968), .Z(n26624) );
  XOR U29088 ( .A(n28969), .B(n28970), .Z(n24460) );
  ANDN U29089 ( .B(n27550), .A(n27552), .Z(n28969) );
  XNOR U29090 ( .A(n28971), .B(n26995), .Z(n26814) );
  AND U29091 ( .A(n27543), .B(n27542), .Z(n28971) );
  XOR U29092 ( .A(n28972), .B(n28973), .Z(n26955) );
  ANDN U29093 ( .B(n28974), .A(n28975), .Z(n28972) );
  ANDN U29094 ( .B(n20369), .A(n19894), .Z(n28959) );
  XOR U29095 ( .A(n23712), .B(n28976), .Z(n19894) );
  XNOR U29096 ( .A(n27907), .B(n27585), .Z(n23712) );
  XNOR U29097 ( .A(n28977), .B(n28978), .Z(n27585) );
  XNOR U29098 ( .A(n23789), .B(n28979), .Z(n28978) );
  XNOR U29099 ( .A(n28980), .B(n28981), .Z(n23789) );
  AND U29100 ( .A(n27368), .B(n27366), .Z(n28980) );
  XOR U29101 ( .A(n28982), .B(n28983), .Z(n27368) );
  XNOR U29102 ( .A(n26071), .B(n28984), .Z(n28977) );
  XNOR U29103 ( .A(n24770), .B(n24376), .Z(n28984) );
  XOR U29104 ( .A(n28985), .B(n28986), .Z(n24376) );
  ANDN U29105 ( .B(n27376), .A(n27377), .Z(n28985) );
  XOR U29106 ( .A(n28987), .B(n28988), .Z(n27377) );
  XNOR U29107 ( .A(n28989), .B(n28990), .Z(n24770) );
  ANDN U29108 ( .B(n27610), .A(n28052), .Z(n28989) );
  IV U29109 ( .A(n27612), .Z(n28052) );
  XOR U29110 ( .A(n28991), .B(n28992), .Z(n27612) );
  XOR U29111 ( .A(n28993), .B(n28994), .Z(n26071) );
  ANDN U29112 ( .B(n27370), .A(n28045), .Z(n28993) );
  IV U29113 ( .A(n27372), .Z(n28045) );
  XOR U29114 ( .A(n28995), .B(n28996), .Z(n27372) );
  XOR U29115 ( .A(n28997), .B(n28998), .Z(n27907) );
  XOR U29116 ( .A(n25257), .B(n26479), .Z(n28998) );
  XNOR U29117 ( .A(n28999), .B(n29000), .Z(n26479) );
  NOR U29118 ( .A(n26170), .B(n29001), .Z(n28999) );
  XOR U29119 ( .A(n29002), .B(n29003), .Z(n25257) );
  ANDN U29120 ( .B(n29004), .A(n26161), .Z(n29002) );
  XOR U29121 ( .A(n29005), .B(n29006), .Z(n28997) );
  XOR U29122 ( .A(n25044), .B(n25782), .Z(n29006) );
  XNOR U29123 ( .A(n29007), .B(n29008), .Z(n25782) );
  NOR U29124 ( .A(n26166), .B(n29009), .Z(n29007) );
  XNOR U29125 ( .A(n29010), .B(n29011), .Z(n25044) );
  ANDN U29126 ( .B(n26157), .A(n29012), .Z(n29010) );
  XNOR U29127 ( .A(n28510), .B(n22958), .Z(n20369) );
  IV U29128 ( .A(n22404), .Z(n22958) );
  XOR U29129 ( .A(n26108), .B(n29013), .Z(n22404) );
  XOR U29130 ( .A(n29014), .B(n29015), .Z(n26108) );
  XNOR U29131 ( .A(n25421), .B(n24568), .Z(n29015) );
  XOR U29132 ( .A(n29016), .B(n29017), .Z(n24568) );
  AND U29133 ( .A(n28503), .B(n28504), .Z(n29016) );
  XNOR U29134 ( .A(n29018), .B(n27479), .Z(n25421) );
  XOR U29135 ( .A(n29019), .B(n29020), .Z(n27480) );
  XOR U29136 ( .A(n24459), .B(n29021), .Z(n29014) );
  XOR U29137 ( .A(n25588), .B(n24793), .Z(n29021) );
  XOR U29138 ( .A(n29022), .B(n27483), .Z(n24793) );
  ANDN U29139 ( .B(n27484), .A(n28512), .Z(n29022) );
  XOR U29140 ( .A(n29023), .B(n29024), .Z(n27484) );
  XNOR U29141 ( .A(n29025), .B(n27475), .Z(n25588) );
  XOR U29142 ( .A(n29026), .B(n29027), .Z(n27476) );
  XNOR U29143 ( .A(n29028), .B(n27470), .Z(n24459) );
  ANDN U29144 ( .B(n27471), .A(n29029), .Z(n29028) );
  XOR U29145 ( .A(n29030), .B(n27471), .Z(n28510) );
  XOR U29146 ( .A(n29031), .B(n29032), .Z(n27471) );
  XNOR U29147 ( .A(n29034), .B(n20160), .Z(n20156) );
  XOR U29148 ( .A(n29035), .B(n25958), .Z(n20160) );
  IV U29149 ( .A(n27228), .Z(n25958) );
  NOR U29150 ( .A(n23556), .B(n19881), .Z(n29034) );
  XNOR U29151 ( .A(n22641), .B(n28338), .Z(n19881) );
  XNOR U29152 ( .A(n29036), .B(n29037), .Z(n28338) );
  ANDN U29153 ( .B(n29038), .A(n29039), .Z(n29036) );
  XOR U29154 ( .A(n29040), .B(n29041), .Z(n22641) );
  IV U29155 ( .A(n20161), .Z(n23556) );
  XOR U29156 ( .A(n28756), .B(n22008), .Z(n20161) );
  IV U29157 ( .A(n28710), .Z(n22008) );
  XNOR U29158 ( .A(n26584), .B(n26711), .Z(n28710) );
  XNOR U29159 ( .A(n29042), .B(n29043), .Z(n26711) );
  XOR U29160 ( .A(n23802), .B(n23075), .Z(n29043) );
  XNOR U29161 ( .A(n29044), .B(n27193), .Z(n23075) );
  XNOR U29162 ( .A(n29045), .B(n29046), .Z(n27193) );
  XNOR U29163 ( .A(n29047), .B(n29048), .Z(n27194) );
  XOR U29164 ( .A(n29049), .B(n29050), .Z(n26888) );
  XOR U29165 ( .A(n29051), .B(n27180), .Z(n23802) );
  XOR U29166 ( .A(n29052), .B(n29053), .Z(n27180) );
  NOR U29167 ( .A(n27179), .B(n26901), .Z(n29051) );
  XOR U29168 ( .A(n29054), .B(n29055), .Z(n26901) );
  XNOR U29169 ( .A(n29056), .B(n29057), .Z(n27179) );
  XOR U29170 ( .A(n27174), .B(n29058), .Z(n29042) );
  XOR U29171 ( .A(n26874), .B(n23702), .Z(n29058) );
  XOR U29172 ( .A(n29059), .B(n27191), .Z(n23702) );
  XOR U29173 ( .A(n29060), .B(n29061), .Z(n27191) );
  NOR U29174 ( .A(n29062), .B(n26893), .Z(n29059) );
  XOR U29175 ( .A(n29063), .B(n27188), .Z(n26874) );
  XNOR U29176 ( .A(n29064), .B(n29065), .Z(n27188) );
  NOR U29177 ( .A(n26897), .B(n27187), .Z(n29063) );
  XOR U29178 ( .A(n29066), .B(n29067), .Z(n27187) );
  XOR U29179 ( .A(n29068), .B(n27933), .Z(n26897) );
  XOR U29180 ( .A(n29069), .B(n27184), .Z(n27174) );
  XOR U29181 ( .A(n29070), .B(n29071), .Z(n27184) );
  XOR U29182 ( .A(n29072), .B(n29073), .Z(n27892) );
  XOR U29183 ( .A(n29074), .B(n29075), .Z(n27183) );
  XOR U29184 ( .A(n29076), .B(n29077), .Z(n26584) );
  XOR U29185 ( .A(n25948), .B(n25306), .Z(n29077) );
  XOR U29186 ( .A(n29078), .B(n27981), .Z(n25306) );
  AND U29187 ( .A(n29079), .B(n29080), .Z(n29078) );
  XNOR U29188 ( .A(n29081), .B(n29082), .Z(n25948) );
  ANDN U29189 ( .B(n29083), .A(n29084), .Z(n29081) );
  XNOR U29190 ( .A(n23836), .B(n29085), .Z(n29076) );
  XNOR U29191 ( .A(n29086), .B(n25431), .Z(n29085) );
  XNOR U29192 ( .A(n29087), .B(n28649), .Z(n25431) );
  NOR U29193 ( .A(n29088), .B(n29089), .Z(n29087) );
  XOR U29194 ( .A(n29090), .B(n27976), .Z(n23836) );
  ANDN U29195 ( .B(n29091), .A(n29092), .Z(n29090) );
  XNOR U29196 ( .A(n29093), .B(n29062), .Z(n28756) );
  IV U29197 ( .A(n27190), .Z(n29062) );
  XOR U29198 ( .A(n29094), .B(n29095), .Z(n27190) );
  ANDN U29199 ( .B(n26893), .A(n28434), .Z(n29093) );
  IV U29200 ( .A(n26895), .Z(n28434) );
  XNOR U29201 ( .A(n29096), .B(n28887), .Z(n26895) );
  XOR U29202 ( .A(n29097), .B(n29098), .Z(n26893) );
  XNOR U29203 ( .A(n29099), .B(n20164), .Z(n17794) );
  XOR U29204 ( .A(n24528), .B(n29100), .Z(n20164) );
  XNOR U29205 ( .A(n26616), .B(n25872), .Z(n24528) );
  XNOR U29206 ( .A(n29101), .B(n29102), .Z(n25872) );
  XOR U29207 ( .A(n29103), .B(n24064), .Z(n29102) );
  XNOR U29208 ( .A(n29104), .B(n27418), .Z(n24064) );
  ANDN U29209 ( .B(n29105), .A(n29106), .Z(n29104) );
  XNOR U29210 ( .A(n25320), .B(n29107), .Z(n29101) );
  XOR U29211 ( .A(n22642), .B(n24886), .Z(n29107) );
  XNOR U29212 ( .A(n29108), .B(n27422), .Z(n24886) );
  IV U29213 ( .A(n29109), .Z(n27422) );
  ANDN U29214 ( .B(n29110), .A(n29111), .Z(n29108) );
  XNOR U29215 ( .A(n29112), .B(n27413), .Z(n22642) );
  IV U29216 ( .A(n29113), .Z(n27413) );
  AND U29217 ( .A(n29114), .B(n29115), .Z(n29112) );
  XOR U29218 ( .A(n29116), .B(n27431), .Z(n25320) );
  ANDN U29219 ( .B(n29117), .A(n29118), .Z(n29116) );
  XOR U29220 ( .A(n29119), .B(n29120), .Z(n26616) );
  XOR U29221 ( .A(n25464), .B(n24033), .Z(n29120) );
  XNOR U29222 ( .A(n29121), .B(n29122), .Z(n24033) );
  AND U29223 ( .A(n29123), .B(n29124), .Z(n29121) );
  XNOR U29224 ( .A(n29125), .B(n28681), .Z(n25464) );
  ANDN U29225 ( .B(n29126), .A(n29127), .Z(n29125) );
  XNOR U29226 ( .A(n23984), .B(n29128), .Z(n29119) );
  XNOR U29227 ( .A(n29129), .B(n29130), .Z(n29128) );
  XOR U29228 ( .A(n29131), .B(n28695), .Z(n23984) );
  AND U29229 ( .A(n29132), .B(n29133), .Z(n29131) );
  ANDN U29230 ( .B(n19890), .A(n20163), .Z(n29099) );
  XNOR U29231 ( .A(n28914), .B(n23013), .Z(n20163) );
  XOR U29232 ( .A(n28060), .B(n29134), .Z(n23013) );
  XOR U29233 ( .A(n29135), .B(n29136), .Z(n28060) );
  XOR U29234 ( .A(n22940), .B(n26072), .Z(n29136) );
  XNOR U29235 ( .A(n29137), .B(n29138), .Z(n26072) );
  ANDN U29236 ( .B(n28920), .A(n28921), .Z(n29137) );
  XNOR U29237 ( .A(n29139), .B(n29140), .Z(n22940) );
  AND U29238 ( .A(n29141), .B(n29142), .Z(n29139) );
  XOR U29239 ( .A(n24933), .B(n29143), .Z(n29135) );
  XOR U29240 ( .A(n23986), .B(n26219), .Z(n29143) );
  XOR U29241 ( .A(n29144), .B(n29145), .Z(n26219) );
  ANDN U29242 ( .B(n28908), .A(n29146), .Z(n29144) );
  XOR U29243 ( .A(n29147), .B(n29148), .Z(n23986) );
  ANDN U29244 ( .B(n28912), .A(n28910), .Z(n29147) );
  XNOR U29245 ( .A(n29149), .B(n29150), .Z(n24933) );
  NOR U29246 ( .A(n28916), .B(n28917), .Z(n29149) );
  IV U29247 ( .A(n29151), .Z(n28916) );
  XNOR U29248 ( .A(n29152), .B(n29141), .Z(n28914) );
  NOR U29249 ( .A(n29153), .B(n29142), .Z(n29152) );
  XNOR U29250 ( .A(n25986), .B(n28230), .Z(n19890) );
  XOR U29251 ( .A(n29154), .B(n29155), .Z(n28230) );
  XNOR U29252 ( .A(n26781), .B(n29156), .Z(n25986) );
  XOR U29253 ( .A(n29157), .B(n29158), .Z(n26781) );
  XOR U29254 ( .A(n24422), .B(n25470), .Z(n29158) );
  XNOR U29255 ( .A(n29159), .B(n29160), .Z(n25470) );
  NOR U29256 ( .A(n28221), .B(n28222), .Z(n29159) );
  XOR U29257 ( .A(n29161), .B(n29162), .Z(n28222) );
  XNOR U29258 ( .A(n29163), .B(n29164), .Z(n24422) );
  ANDN U29259 ( .B(n28232), .A(n28234), .Z(n29163) );
  XOR U29260 ( .A(n29165), .B(n29166), .Z(n28234) );
  XNOR U29261 ( .A(n26794), .B(n29167), .Z(n29157) );
  XOR U29262 ( .A(n26639), .B(n23841), .Z(n29167) );
  XNOR U29263 ( .A(n29168), .B(n29169), .Z(n23841) );
  ANDN U29264 ( .B(n28227), .A(n28225), .Z(n29168) );
  XOR U29265 ( .A(n29170), .B(n29171), .Z(n28227) );
  XNOR U29266 ( .A(n29172), .B(n29173), .Z(n26639) );
  ANDN U29267 ( .B(n29155), .A(n28483), .Z(n29172) );
  XOR U29268 ( .A(n29174), .B(n29175), .Z(n28483) );
  XNOR U29269 ( .A(n29176), .B(n29177), .Z(n26794) );
  ANDN U29270 ( .B(n28361), .A(n28360), .Z(n29176) );
  XOR U29271 ( .A(n29178), .B(n29179), .Z(n28361) );
  XNOR U29272 ( .A(n29180), .B(n21237), .Z(n20363) );
  XOR U29273 ( .A(n27973), .B(n27723), .Z(n21237) );
  XOR U29274 ( .A(n26231), .B(n26645), .Z(n27723) );
  XNOR U29275 ( .A(n29181), .B(n29182), .Z(n26645) );
  XOR U29276 ( .A(n22510), .B(n25148), .Z(n29182) );
  XNOR U29277 ( .A(n29183), .B(n29184), .Z(n25148) );
  ANDN U29278 ( .B(n29185), .A(n29186), .Z(n29183) );
  XNOR U29279 ( .A(n29187), .B(n29188), .Z(n22510) );
  ANDN U29280 ( .B(n29189), .A(n29190), .Z(n29187) );
  XNOR U29281 ( .A(n29191), .B(n29192), .Z(n29181) );
  XOR U29282 ( .A(n25826), .B(n21828), .Z(n29192) );
  XNOR U29283 ( .A(n29193), .B(n29194), .Z(n21828) );
  ANDN U29284 ( .B(n29195), .A(n29196), .Z(n29193) );
  XNOR U29285 ( .A(n29197), .B(n29198), .Z(n25826) );
  ANDN U29286 ( .B(n29199), .A(n29200), .Z(n29197) );
  XOR U29287 ( .A(n29201), .B(n29202), .Z(n26231) );
  XOR U29288 ( .A(n26370), .B(n25799), .Z(n29202) );
  XOR U29289 ( .A(n29203), .B(n29080), .Z(n25799) );
  ANDN U29290 ( .B(n27980), .A(n27979), .Z(n29203) );
  XNOR U29291 ( .A(n29204), .B(n29083), .Z(n26370) );
  ANDN U29292 ( .B(n29205), .A(n29206), .Z(n29204) );
  XOR U29293 ( .A(n25246), .B(n29207), .Z(n29201) );
  XNOR U29294 ( .A(n29208), .B(n29209), .Z(n29207) );
  XNOR U29295 ( .A(n29210), .B(n29088), .Z(n25246) );
  ANDN U29296 ( .B(n28648), .A(n28647), .Z(n29210) );
  XOR U29297 ( .A(n29211), .B(n29206), .Z(n27973) );
  NOR U29298 ( .A(n29205), .B(n29082), .Z(n29211) );
  NOR U29299 ( .A(n21232), .B(n19885), .Z(n29180) );
  XNOR U29300 ( .A(n29212), .B(n24262), .Z(n19885) );
  XNOR U29301 ( .A(n29213), .B(n29214), .Z(n26727) );
  XOR U29302 ( .A(n24900), .B(n29215), .Z(n29214) );
  XNOR U29303 ( .A(n29216), .B(n29217), .Z(n24900) );
  AND U29304 ( .A(n29218), .B(n29219), .Z(n29216) );
  XOR U29305 ( .A(n25615), .B(n29220), .Z(n29213) );
  XNOR U29306 ( .A(n29221), .B(n27055), .Z(n29220) );
  XOR U29307 ( .A(n29222), .B(n28847), .Z(n27055) );
  XNOR U29308 ( .A(n29225), .B(n28855), .Z(n25615) );
  NOR U29309 ( .A(n29226), .B(n29227), .Z(n29225) );
  XNOR U29310 ( .A(n29228), .B(n29229), .Z(n25873) );
  XNOR U29311 ( .A(n24823), .B(n22816), .Z(n29229) );
  XNOR U29312 ( .A(n29230), .B(n29231), .Z(n22816) );
  AND U29313 ( .A(n29232), .B(n29233), .Z(n29230) );
  XNOR U29314 ( .A(n29234), .B(n29235), .Z(n24823) );
  ANDN U29315 ( .B(n29236), .A(n29237), .Z(n29234) );
  XOR U29316 ( .A(n25767), .B(n29238), .Z(n29228) );
  XOR U29317 ( .A(n25934), .B(n26054), .Z(n29238) );
  XOR U29318 ( .A(n29239), .B(n26206), .Z(n26054) );
  NOR U29319 ( .A(n29240), .B(n29241), .Z(n29239) );
  XOR U29320 ( .A(n29242), .B(n26211), .Z(n25934) );
  ANDN U29321 ( .B(n29243), .A(n29244), .Z(n29242) );
  XNOR U29322 ( .A(n29245), .B(n26216), .Z(n25767) );
  AND U29323 ( .A(n29246), .B(n29247), .Z(n29245) );
  IV U29324 ( .A(n19887), .Z(n21232) );
  XNOR U29325 ( .A(n26537), .B(n26620), .Z(n19887) );
  XNOR U29326 ( .A(n29248), .B(n27547), .Z(n26537) );
  NOR U29327 ( .A(n29249), .B(n28965), .Z(n29248) );
  ANDN U29328 ( .B(n13505), .A(n16724), .Z(n28715) );
  IV U29329 ( .A(n13507), .Z(n16724) );
  XNOR U29330 ( .A(n22107), .B(n17630), .Z(n13507) );
  XNOR U29331 ( .A(n23424), .B(n23519), .Z(n17630) );
  XOR U29332 ( .A(n29250), .B(n29251), .Z(n23519) );
  XOR U29333 ( .A(n17957), .B(n18592), .Z(n29251) );
  XOR U29334 ( .A(n29252), .B(n23102), .Z(n18592) );
  XNOR U29335 ( .A(n25362), .B(n29253), .Z(n23102) );
  XOR U29336 ( .A(n29254), .B(n29255), .Z(n26768) );
  XNOR U29337 ( .A(n25685), .B(n25467), .Z(n29255) );
  XNOR U29338 ( .A(n29256), .B(n28908), .Z(n25467) );
  XOR U29339 ( .A(n29257), .B(n29258), .Z(n28908) );
  XNOR U29340 ( .A(n29260), .B(n28912), .Z(n25685) );
  XOR U29341 ( .A(n29261), .B(n29262), .Z(n28912) );
  ANDN U29342 ( .B(n28911), .A(n29263), .Z(n29260) );
  XOR U29343 ( .A(n21589), .B(n29264), .Z(n29254) );
  XNOR U29344 ( .A(n26046), .B(n27034), .Z(n29264) );
  XNOR U29345 ( .A(n29265), .B(n29142), .Z(n27034) );
  XOR U29346 ( .A(n29266), .B(n29267), .Z(n29142) );
  ANDN U29347 ( .B(n29153), .A(n29268), .Z(n29265) );
  IV U29348 ( .A(n29269), .Z(n29153) );
  XOR U29349 ( .A(n29270), .B(n28917), .Z(n26046) );
  XOR U29350 ( .A(n29271), .B(n29272), .Z(n28917) );
  ANDN U29351 ( .B(n28918), .A(n29273), .Z(n29270) );
  XNOR U29352 ( .A(n29274), .B(n28921), .Z(n21589) );
  XNOR U29353 ( .A(n29275), .B(n29071), .Z(n28921) );
  XOR U29354 ( .A(n29278), .B(n26030), .Z(n21923) );
  XOR U29355 ( .A(n28946), .B(n24296), .Z(n21924) );
  IV U29356 ( .A(n24402), .Z(n24296) );
  XOR U29357 ( .A(n29280), .B(n29281), .Z(n26015) );
  XOR U29358 ( .A(n25028), .B(n27827), .Z(n29281) );
  XNOR U29359 ( .A(n29282), .B(n26747), .Z(n27827) );
  XOR U29360 ( .A(n29283), .B(n29284), .Z(n26747) );
  ANDN U29361 ( .B(n28953), .A(n28952), .Z(n29282) );
  IV U29362 ( .A(n27845), .Z(n28952) );
  XOR U29363 ( .A(n29285), .B(n29286), .Z(n27845) );
  XOR U29364 ( .A(n29287), .B(n27835), .Z(n25028) );
  XOR U29365 ( .A(n29288), .B(n29289), .Z(n27835) );
  ANDN U29366 ( .B(n27834), .A(n28957), .Z(n29287) );
  XOR U29367 ( .A(n29290), .B(n29291), .Z(n27834) );
  XNOR U29368 ( .A(n23325), .B(n29292), .Z(n29280) );
  XNOR U29369 ( .A(n21367), .B(n23491), .Z(n29292) );
  XOR U29370 ( .A(n29293), .B(n26743), .Z(n23491) );
  XOR U29371 ( .A(n29294), .B(n29295), .Z(n26743) );
  ANDN U29372 ( .B(n27831), .A(n29296), .Z(n29293) );
  XOR U29373 ( .A(n29297), .B(n27843), .Z(n21367) );
  XOR U29374 ( .A(n29298), .B(n29299), .Z(n27843) );
  ANDN U29375 ( .B(n27842), .A(n28955), .Z(n29297) );
  XNOR U29376 ( .A(n29300), .B(n29301), .Z(n27842) );
  XOR U29377 ( .A(n29302), .B(n27840), .Z(n23325) );
  NOR U29378 ( .A(n27839), .B(n28948), .Z(n29302) );
  XNOR U29379 ( .A(n29303), .B(n29304), .Z(n27839) );
  XNOR U29380 ( .A(n29305), .B(n27831), .Z(n28946) );
  XOR U29381 ( .A(n29306), .B(n29307), .Z(n27831) );
  ANDN U29382 ( .B(n26741), .A(n29308), .Z(n29305) );
  XNOR U29383 ( .A(n29309), .B(n23093), .Z(n17957) );
  IV U29384 ( .A(n25740), .Z(n23093) );
  XOR U29385 ( .A(n29310), .B(n23577), .Z(n25740) );
  NOR U29386 ( .A(n26137), .B(n21913), .Z(n29309) );
  XOR U29387 ( .A(n27467), .B(n24842), .Z(n21913) );
  IV U29388 ( .A(n23996), .Z(n24842) );
  XNOR U29389 ( .A(n26841), .B(n29311), .Z(n23996) );
  XOR U29390 ( .A(n29312), .B(n29313), .Z(n26841) );
  XNOR U29391 ( .A(n27195), .B(n23441), .Z(n29313) );
  XNOR U29392 ( .A(n29314), .B(n28516), .Z(n23441) );
  XOR U29393 ( .A(n29315), .B(n29316), .Z(n27475) );
  XNOR U29394 ( .A(n29317), .B(n29033), .Z(n27195) );
  NOR U29395 ( .A(n27470), .B(n27469), .Z(n29317) );
  XOR U29396 ( .A(n29318), .B(n28892), .Z(n27470) );
  XOR U29397 ( .A(n25658), .B(n29319), .Z(n29312) );
  XNOR U29398 ( .A(n23754), .B(n29320), .Z(n29319) );
  XNOR U29399 ( .A(n29321), .B(n28513), .Z(n23754) );
  XOR U29400 ( .A(n29322), .B(n27949), .Z(n27483) );
  XNOR U29401 ( .A(n29323), .B(n28508), .Z(n25658) );
  ANDN U29402 ( .B(n27478), .A(n27479), .Z(n29323) );
  XOR U29403 ( .A(n29324), .B(n29325), .Z(n27479) );
  XNOR U29404 ( .A(n29326), .B(n29327), .Z(n27467) );
  NOR U29405 ( .A(n29017), .B(n28503), .Z(n29326) );
  XOR U29406 ( .A(n29328), .B(n29329), .Z(n28503) );
  IV U29407 ( .A(n21915), .Z(n26137) );
  XOR U29408 ( .A(n24484), .B(n29330), .Z(n21915) );
  IV U29409 ( .A(n21235), .Z(n24484) );
  XOR U29410 ( .A(n27310), .B(n27846), .Z(n21235) );
  XOR U29411 ( .A(n29331), .B(n29332), .Z(n27846) );
  XNOR U29412 ( .A(n25707), .B(n29333), .Z(n29332) );
  XOR U29413 ( .A(n29334), .B(n29335), .Z(n25707) );
  NOR U29414 ( .A(n28933), .B(n29336), .Z(n29334) );
  XNOR U29415 ( .A(n23255), .B(n29337), .Z(n29331) );
  XOR U29416 ( .A(n26582), .B(n22789), .Z(n29337) );
  XNOR U29417 ( .A(n29338), .B(n29339), .Z(n22789) );
  ANDN U29418 ( .B(n29340), .A(n28937), .Z(n29338) );
  XNOR U29419 ( .A(n29341), .B(n29342), .Z(n26582) );
  ANDN U29420 ( .B(n29343), .A(n29344), .Z(n29341) );
  XOR U29421 ( .A(n29345), .B(n29346), .Z(n23255) );
  ANDN U29422 ( .B(n29347), .A(n28928), .Z(n29345) );
  XNOR U29423 ( .A(n29348), .B(n29349), .Z(n27310) );
  XOR U29424 ( .A(n25460), .B(n28289), .Z(n29349) );
  XNOR U29425 ( .A(n29350), .B(n29351), .Z(n28289) );
  ANDN U29426 ( .B(n29352), .A(n29353), .Z(n29350) );
  XNOR U29427 ( .A(n29354), .B(n29355), .Z(n25460) );
  ANDN U29428 ( .B(n29356), .A(n29357), .Z(n29354) );
  XOR U29429 ( .A(n29358), .B(n29359), .Z(n29348) );
  XOR U29430 ( .A(n26275), .B(n25360), .Z(n29359) );
  XNOR U29431 ( .A(n29360), .B(n29361), .Z(n25360) );
  ANDN U29432 ( .B(n29362), .A(n29363), .Z(n29360) );
  XNOR U29433 ( .A(n29364), .B(n29365), .Z(n26275) );
  ANDN U29434 ( .B(n29366), .A(n29367), .Z(n29364) );
  XOR U29435 ( .A(n20014), .B(n29368), .Z(n29250) );
  XOR U29436 ( .A(n23084), .B(n20080), .Z(n29368) );
  XNOR U29437 ( .A(n29369), .B(n23089), .Z(n20080) );
  XNOR U29438 ( .A(n27054), .B(n29221), .Z(n23089) );
  XNOR U29439 ( .A(n29370), .B(n28843), .Z(n29221) );
  ANDN U29440 ( .B(n29371), .A(n29372), .Z(n29370) );
  ANDN U29441 ( .B(n21921), .A(n23090), .Z(n29369) );
  XOR U29442 ( .A(n29373), .B(n24506), .Z(n23090) );
  XNOR U29443 ( .A(n29374), .B(n26771), .Z(n24506) );
  XOR U29444 ( .A(n29375), .B(n29376), .Z(n26771) );
  XNOR U29445 ( .A(n26925), .B(n28133), .Z(n29376) );
  XNOR U29446 ( .A(n29377), .B(n29378), .Z(n28133) );
  NOR U29447 ( .A(n29379), .B(n27321), .Z(n29377) );
  XNOR U29448 ( .A(n29380), .B(n29381), .Z(n26925) );
  ANDN U29449 ( .B(n29382), .A(n27915), .Z(n29380) );
  XNOR U29450 ( .A(n29383), .B(n29384), .Z(n29375) );
  XNOR U29451 ( .A(n29385), .B(n25069), .Z(n29384) );
  XNOR U29452 ( .A(n29386), .B(n29387), .Z(n25069) );
  NOR U29453 ( .A(n29388), .B(n27325), .Z(n29386) );
  XOR U29454 ( .A(n29389), .B(n23139), .Z(n21921) );
  XNOR U29455 ( .A(n29391), .B(n29392), .Z(n27199) );
  XOR U29456 ( .A(n25584), .B(n25168), .Z(n29392) );
  XOR U29457 ( .A(n29393), .B(n29394), .Z(n25168) );
  ANDN U29458 ( .B(n29395), .A(n27151), .Z(n29393) );
  IV U29459 ( .A(n28665), .Z(n27151) );
  XNOR U29460 ( .A(n29396), .B(n29397), .Z(n28665) );
  XNOR U29461 ( .A(n29398), .B(n29399), .Z(n25584) );
  NOR U29462 ( .A(n27155), .B(n28660), .Z(n29398) );
  IV U29463 ( .A(n28661), .Z(n27155) );
  XOR U29464 ( .A(n29400), .B(n29401), .Z(n28661) );
  XNOR U29465 ( .A(n25416), .B(n29402), .Z(n29391) );
  XNOR U29466 ( .A(n23601), .B(n26013), .Z(n29402) );
  XNOR U29467 ( .A(n29403), .B(n29404), .Z(n26013) );
  ANDN U29468 ( .B(n27146), .A(n28667), .Z(n29403) );
  XNOR U29469 ( .A(n29405), .B(n29032), .Z(n27146) );
  XOR U29470 ( .A(n29406), .B(n29407), .Z(n23601) );
  ANDN U29471 ( .B(n27159), .A(n28658), .Z(n29406) );
  XNOR U29472 ( .A(n29408), .B(n29409), .Z(n27159) );
  XOR U29473 ( .A(n29410), .B(n29411), .Z(n25416) );
  NOR U29474 ( .A(n28673), .B(n28669), .Z(n29410) );
  IV U29475 ( .A(n28671), .Z(n28673) );
  XOR U29476 ( .A(n29412), .B(n29413), .Z(n28671) );
  XNOR U29477 ( .A(n29414), .B(n25701), .Z(n23084) );
  XOR U29478 ( .A(n23742), .B(n29415), .Z(n25701) );
  IV U29479 ( .A(n24446), .Z(n23742) );
  XNOR U29480 ( .A(n26510), .B(n25842), .Z(n24446) );
  XNOR U29481 ( .A(n29416), .B(n29417), .Z(n25842) );
  XOR U29482 ( .A(n24491), .B(n25143), .Z(n29417) );
  XOR U29483 ( .A(n29418), .B(n27345), .Z(n25143) );
  XNOR U29484 ( .A(n29420), .B(n27353), .Z(n24491) );
  ANDN U29485 ( .B(n29421), .A(n29422), .Z(n29420) );
  XOR U29486 ( .A(n26817), .B(n29423), .Z(n29416) );
  XOR U29487 ( .A(n29424), .B(n25473), .Z(n29423) );
  XOR U29488 ( .A(n29425), .B(n27351), .Z(n25473) );
  ANDN U29489 ( .B(n26499), .A(n29426), .Z(n29425) );
  XNOR U29490 ( .A(n29427), .B(n27343), .Z(n26817) );
  ANDN U29491 ( .B(n26488), .A(n29428), .Z(n29427) );
  XOR U29492 ( .A(n29429), .B(n29430), .Z(n26510) );
  XNOR U29493 ( .A(n26476), .B(n25151), .Z(n29430) );
  XOR U29494 ( .A(n29431), .B(n26337), .Z(n25151) );
  AND U29495 ( .A(n29432), .B(n29433), .Z(n29431) );
  XNOR U29496 ( .A(n29434), .B(n26333), .Z(n26476) );
  AND U29497 ( .A(n29435), .B(n29436), .Z(n29434) );
  XOR U29498 ( .A(n29437), .B(n29438), .Z(n29429) );
  XNOR U29499 ( .A(n26519), .B(n25536), .Z(n29438) );
  XNOR U29500 ( .A(n29439), .B(n26321), .Z(n25536) );
  ANDN U29501 ( .B(n29440), .A(n29441), .Z(n29439) );
  XNOR U29502 ( .A(n29442), .B(n26330), .Z(n26519) );
  ANDN U29503 ( .B(n21909), .A(n21910), .Z(n29414) );
  XNOR U29504 ( .A(n28237), .B(n22820), .Z(n21910) );
  XNOR U29505 ( .A(n29445), .B(n29446), .Z(n28237) );
  XNOR U29506 ( .A(n29447), .B(n24146), .Z(n21909) );
  XNOR U29507 ( .A(n29448), .B(n29449), .Z(n25262) );
  XNOR U29508 ( .A(n26526), .B(n29450), .Z(n29449) );
  XOR U29509 ( .A(n29451), .B(n28355), .Z(n26526) );
  ANDN U29510 ( .B(n29452), .A(n29453), .Z(n29451) );
  XOR U29511 ( .A(n26380), .B(n29454), .Z(n29448) );
  XNOR U29512 ( .A(n29455), .B(n25832), .Z(n29454) );
  XOR U29513 ( .A(n29456), .B(n28347), .Z(n25832) );
  AND U29514 ( .A(n29457), .B(n29458), .Z(n29456) );
  XNOR U29515 ( .A(n29459), .B(n29039), .Z(n26380) );
  ANDN U29516 ( .B(n29460), .A(n29461), .Z(n29459) );
  XNOR U29517 ( .A(n29462), .B(n29463), .Z(n28780) );
  XOR U29518 ( .A(n26460), .B(n24978), .Z(n29463) );
  XNOR U29519 ( .A(n29464), .B(n29465), .Z(n24978) );
  AND U29520 ( .A(n29466), .B(n29467), .Z(n29464) );
  XNOR U29521 ( .A(n29468), .B(n29469), .Z(n26460) );
  XNOR U29522 ( .A(n24791), .B(n29472), .Z(n29462) );
  XNOR U29523 ( .A(n23992), .B(n25669), .Z(n29472) );
  XOR U29524 ( .A(n29473), .B(n29474), .Z(n25669) );
  XNOR U29525 ( .A(n29477), .B(n29478), .Z(n23992) );
  ANDN U29526 ( .B(n29479), .A(n29480), .Z(n29477) );
  XOR U29527 ( .A(n29481), .B(n29482), .Z(n24791) );
  ANDN U29528 ( .B(n29483), .A(n29484), .Z(n29481) );
  XNOR U29529 ( .A(n29485), .B(n23099), .Z(n20014) );
  XNOR U29530 ( .A(n25659), .B(n29486), .Z(n23099) );
  IV U29531 ( .A(n23335), .Z(n25659) );
  XNOR U29532 ( .A(n29487), .B(n28753), .Z(n23335) );
  XNOR U29533 ( .A(n29488), .B(n29489), .Z(n28753) );
  XOR U29534 ( .A(n25943), .B(n26710), .Z(n29489) );
  XNOR U29535 ( .A(n29490), .B(n27333), .Z(n26710) );
  ANDN U29536 ( .B(n28451), .A(n29491), .Z(n29490) );
  XOR U29537 ( .A(n29492), .B(n26835), .Z(n25943) );
  ANDN U29538 ( .B(n28440), .A(n29493), .Z(n29492) );
  XNOR U29539 ( .A(n22808), .B(n29494), .Z(n29488) );
  XNOR U29540 ( .A(n26066), .B(n26406), .Z(n29494) );
  XNOR U29541 ( .A(n29495), .B(n28166), .Z(n26406) );
  ANDN U29542 ( .B(n29496), .A(n28449), .Z(n29495) );
  XOR U29543 ( .A(n29497), .B(n28454), .Z(n26066) );
  ANDN U29544 ( .B(n28442), .A(n29498), .Z(n29497) );
  XNOR U29545 ( .A(n29499), .B(n26827), .Z(n22808) );
  ANDN U29546 ( .B(n29500), .A(n28447), .Z(n29499) );
  ANDN U29547 ( .B(n23098), .A(n23522), .Z(n29485) );
  XOR U29548 ( .A(n29501), .B(n22394), .Z(n23522) );
  XNOR U29549 ( .A(n29502), .B(n26813), .Z(n22394) );
  XNOR U29550 ( .A(n29503), .B(n29504), .Z(n26813) );
  XNOR U29551 ( .A(n26094), .B(n26414), .Z(n29504) );
  XNOR U29552 ( .A(n29505), .B(n27492), .Z(n26414) );
  NOR U29553 ( .A(n28386), .B(n27491), .Z(n29505) );
  XNOR U29554 ( .A(n29506), .B(n27505), .Z(n26094) );
  ANDN U29555 ( .B(n28390), .A(n27504), .Z(n29506) );
  XNOR U29556 ( .A(n23052), .B(n29507), .Z(n29503) );
  XNOR U29557 ( .A(n26542), .B(n26447), .Z(n29507) );
  XOR U29558 ( .A(n29508), .B(n29509), .Z(n26447) );
  ANDN U29559 ( .B(n28383), .A(n27495), .Z(n29508) );
  XNOR U29560 ( .A(n29510), .B(n27500), .Z(n26542) );
  ANDN U29561 ( .B(n27501), .A(n28393), .Z(n29510) );
  XNOR U29562 ( .A(n29511), .B(n27509), .Z(n23052) );
  AND U29563 ( .A(n27508), .B(n28396), .Z(n29511) );
  XOR U29564 ( .A(n23998), .B(n28274), .Z(n23098) );
  XOR U29565 ( .A(n29512), .B(n29513), .Z(n28274) );
  ANDN U29566 ( .B(n28287), .A(n28285), .Z(n29512) );
  XOR U29567 ( .A(n27141), .B(n27663), .Z(n23998) );
  XOR U29568 ( .A(n29514), .B(n29515), .Z(n27663) );
  XNOR U29569 ( .A(n26274), .B(n25359), .Z(n29515) );
  XOR U29570 ( .A(n29516), .B(n29517), .Z(n25359) );
  XOR U29571 ( .A(n29518), .B(n29519), .Z(n27109) );
  XOR U29572 ( .A(n29520), .B(n29521), .Z(n26274) );
  NOR U29573 ( .A(n28281), .B(n27113), .Z(n29520) );
  XNOR U29574 ( .A(n28831), .B(n29522), .Z(n27113) );
  IV U29575 ( .A(n29523), .Z(n28281) );
  XOR U29576 ( .A(n24428), .B(n29524), .Z(n29514) );
  XOR U29577 ( .A(n24441), .B(n29525), .Z(n29524) );
  XNOR U29578 ( .A(n29526), .B(n29527), .Z(n24441) );
  ANDN U29579 ( .B(n28283), .A(n28129), .Z(n29526) );
  XOR U29580 ( .A(n29528), .B(n29529), .Z(n28129) );
  XOR U29581 ( .A(n29530), .B(n29531), .Z(n24428) );
  ANDN U29582 ( .B(n27120), .A(n28276), .Z(n29530) );
  XOR U29583 ( .A(n29532), .B(n29533), .Z(n27120) );
  XOR U29584 ( .A(n29534), .B(n29535), .Z(n27141) );
  XOR U29585 ( .A(n26009), .B(n23906), .Z(n29535) );
  XNOR U29586 ( .A(n29536), .B(n29537), .Z(n23906) );
  NOR U29587 ( .A(n29538), .B(n29539), .Z(n29536) );
  XOR U29588 ( .A(n29540), .B(n29541), .Z(n26009) );
  ANDN U29589 ( .B(n29542), .A(n29543), .Z(n29540) );
  XOR U29590 ( .A(n28007), .B(n29544), .Z(n29534) );
  XOR U29591 ( .A(n24777), .B(n25867), .Z(n29544) );
  XNOR U29592 ( .A(n29545), .B(n29546), .Z(n25867) );
  ANDN U29593 ( .B(n29547), .A(n29548), .Z(n29545) );
  XNOR U29594 ( .A(n29549), .B(n29550), .Z(n24777) );
  ANDN U29595 ( .B(n29551), .A(n29552), .Z(n29549) );
  XNOR U29596 ( .A(n29553), .B(n29554), .Z(n28007) );
  NOR U29597 ( .A(n29555), .B(n29556), .Z(n29553) );
  XOR U29598 ( .A(n29557), .B(n29558), .Z(n23424) );
  XOR U29599 ( .A(n17041), .B(n16997), .Z(n29558) );
  XNOR U29600 ( .A(n29559), .B(n20882), .Z(n16997) );
  XNOR U29601 ( .A(n28528), .B(n24930), .Z(n20882) );
  XNOR U29602 ( .A(n29560), .B(n29561), .Z(n29013) );
  XOR U29603 ( .A(n29562), .B(n27259), .Z(n29561) );
  XNOR U29604 ( .A(n29563), .B(n29564), .Z(n27259) );
  ANDN U29605 ( .B(n28520), .A(n28521), .Z(n29563) );
  XOR U29606 ( .A(n24192), .B(n29565), .Z(n29560) );
  XNOR U29607 ( .A(n24372), .B(n27913), .Z(n29565) );
  XOR U29608 ( .A(n29566), .B(n29567), .Z(n27913) );
  NOR U29609 ( .A(n29568), .B(n29569), .Z(n29566) );
  XOR U29610 ( .A(n29570), .B(n29571), .Z(n24372) );
  XNOR U29611 ( .A(n29572), .B(n29573), .Z(n24192) );
  NOR U29612 ( .A(n28534), .B(n28535), .Z(n29572) );
  IV U29613 ( .A(n29574), .Z(n28534) );
  XOR U29614 ( .A(n29575), .B(n29576), .Z(n26769) );
  XNOR U29615 ( .A(n28901), .B(n25000), .Z(n29576) );
  XNOR U29616 ( .A(n29577), .B(n29578), .Z(n25000) );
  ANDN U29617 ( .B(n28267), .A(n29579), .Z(n29577) );
  ANDN U29618 ( .B(n28259), .A(n29582), .Z(n29580) );
  XNOR U29619 ( .A(n25661), .B(n29583), .Z(n29575) );
  XNOR U29620 ( .A(n23502), .B(n24235), .Z(n29583) );
  XNOR U29621 ( .A(n29584), .B(n29585), .Z(n24235) );
  ANDN U29622 ( .B(n28250), .A(n28251), .Z(n29584) );
  XNOR U29623 ( .A(n29586), .B(n29587), .Z(n23502) );
  ANDN U29624 ( .B(n28254), .A(n29588), .Z(n29586) );
  XNOR U29625 ( .A(n29589), .B(n29590), .Z(n25661) );
  ANDN U29626 ( .B(n28263), .A(n28264), .Z(n29589) );
  XNOR U29627 ( .A(n29591), .B(n29592), .Z(n28528) );
  ANDN U29628 ( .B(n29569), .A(n29593), .Z(n29591) );
  ANDN U29629 ( .B(n21670), .A(n26115), .Z(n29559) );
  XOR U29630 ( .A(n29594), .B(n25810), .Z(n26115) );
  IV U29631 ( .A(n24949), .Z(n25810) );
  XOR U29632 ( .A(n27100), .B(n27901), .Z(n24949) );
  XNOR U29633 ( .A(n29595), .B(n29596), .Z(n27901) );
  XOR U29634 ( .A(n25835), .B(n25886), .Z(n29596) );
  XOR U29635 ( .A(n29597), .B(n29598), .Z(n25886) );
  NOR U29636 ( .A(n29599), .B(n29600), .Z(n29597) );
  XNOR U29637 ( .A(n29601), .B(n29602), .Z(n25835) );
  ANDN U29638 ( .B(n29603), .A(n29604), .Z(n29601) );
  XOR U29639 ( .A(n25420), .B(n29605), .Z(n29595) );
  XOR U29640 ( .A(n22390), .B(n23339), .Z(n29605) );
  XNOR U29641 ( .A(n29606), .B(n29607), .Z(n23339) );
  ANDN U29642 ( .B(n29608), .A(n29609), .Z(n29606) );
  XNOR U29643 ( .A(n29610), .B(n29611), .Z(n22390) );
  AND U29644 ( .A(n29612), .B(n29613), .Z(n29610) );
  XNOR U29645 ( .A(n29614), .B(n29615), .Z(n25420) );
  ANDN U29646 ( .B(n29616), .A(n29617), .Z(n29614) );
  XOR U29647 ( .A(n29618), .B(n29619), .Z(n27100) );
  XOR U29648 ( .A(n26571), .B(n22620), .Z(n29619) );
  XOR U29649 ( .A(n29620), .B(n29621), .Z(n22620) );
  ANDN U29650 ( .B(n29622), .A(n29623), .Z(n29620) );
  XNOR U29651 ( .A(n29624), .B(n29625), .Z(n26571) );
  ANDN U29652 ( .B(n29626), .A(n29627), .Z(n29624) );
  XOR U29653 ( .A(n24240), .B(n29628), .Z(n29618) );
  XNOR U29654 ( .A(n25956), .B(n29629), .Z(n29628) );
  XOR U29655 ( .A(n29630), .B(n29631), .Z(n25956) );
  ANDN U29656 ( .B(n29632), .A(n29633), .Z(n29630) );
  XNOR U29657 ( .A(n29634), .B(n29635), .Z(n24240) );
  ANDN U29658 ( .B(n29636), .A(n29637), .Z(n29634) );
  XOR U29659 ( .A(n29638), .B(n22982), .Z(n21670) );
  XNOR U29660 ( .A(n29639), .B(n29640), .Z(n27579) );
  XNOR U29661 ( .A(n28538), .B(n29641), .Z(n29640) );
  XOR U29662 ( .A(n29642), .B(n29357), .Z(n28538) );
  NOR U29663 ( .A(n29643), .B(n29644), .Z(n29642) );
  XOR U29664 ( .A(n25604), .B(n29645), .Z(n29639) );
  XOR U29665 ( .A(n25914), .B(n26643), .Z(n29645) );
  XOR U29666 ( .A(n29646), .B(n29363), .Z(n26643) );
  NOR U29667 ( .A(n29647), .B(n29648), .Z(n29646) );
  XNOR U29668 ( .A(n29649), .B(n29353), .Z(n25914) );
  XOR U29669 ( .A(n29652), .B(n29653), .Z(n25604) );
  NOR U29670 ( .A(n29654), .B(n29655), .Z(n29652) );
  XNOR U29671 ( .A(n29657), .B(n20878), .Z(n17041) );
  XNOR U29672 ( .A(n28313), .B(n25801), .Z(n20878) );
  IV U29673 ( .A(n24395), .Z(n25801) );
  XOR U29674 ( .A(n28398), .B(n26987), .Z(n24395) );
  XNOR U29675 ( .A(n29658), .B(n29659), .Z(n26987) );
  XOR U29676 ( .A(n24258), .B(n23958), .Z(n29659) );
  XNOR U29677 ( .A(n29660), .B(n29608), .Z(n23958) );
  ANDN U29678 ( .B(n29661), .A(n29662), .Z(n29660) );
  XOR U29679 ( .A(n29663), .B(n29604), .Z(n24258) );
  ANDN U29680 ( .B(n29664), .A(n29665), .Z(n29663) );
  XNOR U29681 ( .A(n29666), .B(n29667), .Z(n29658) );
  XOR U29682 ( .A(n25583), .B(n26611), .Z(n29667) );
  XNOR U29683 ( .A(n29668), .B(n29669), .Z(n26611) );
  ANDN U29684 ( .B(n29670), .A(n29671), .Z(n29668) );
  XNOR U29685 ( .A(n29672), .B(n29616), .Z(n25583) );
  AND U29686 ( .A(n29673), .B(n29674), .Z(n29672) );
  XOR U29687 ( .A(n29675), .B(n29676), .Z(n28398) );
  XNOR U29688 ( .A(n23014), .B(n26790), .Z(n29676) );
  XNOR U29689 ( .A(n29677), .B(n29678), .Z(n26790) );
  ANDN U29690 ( .B(n28308), .A(n28306), .Z(n29677) );
  XOR U29691 ( .A(n29679), .B(n29680), .Z(n23014) );
  ANDN U29692 ( .B(n28310), .A(n28311), .Z(n29679) );
  XNOR U29693 ( .A(n26018), .B(n29681), .Z(n29675) );
  XNOR U29694 ( .A(n24229), .B(n24953), .Z(n29681) );
  XNOR U29695 ( .A(n29682), .B(n29683), .Z(n24953) );
  ANDN U29696 ( .B(n28317), .A(n28316), .Z(n29682) );
  XNOR U29697 ( .A(n29684), .B(n29685), .Z(n24229) );
  ANDN U29698 ( .B(n28322), .A(n28320), .Z(n29684) );
  XOR U29699 ( .A(n29686), .B(n29687), .Z(n26018) );
  XNOR U29700 ( .A(n29690), .B(n29688), .Z(n28313) );
  NOR U29701 ( .A(n29689), .B(n29691), .Z(n29690) );
  XOR U29702 ( .A(n29692), .B(n27796), .Z(n22109) );
  XNOR U29703 ( .A(n29693), .B(n23839), .Z(n21677) );
  XNOR U29704 ( .A(n29694), .B(n29695), .Z(n27900) );
  XOR U29705 ( .A(n29696), .B(n23060), .Z(n29695) );
  XOR U29706 ( .A(n29697), .B(n28321), .Z(n23060) );
  ANDN U29707 ( .B(n29685), .A(n29698), .Z(n29697) );
  XOR U29708 ( .A(n21604), .B(n29699), .Z(n29694) );
  XNOR U29709 ( .A(n24002), .B(n29700), .Z(n29699) );
  XNOR U29710 ( .A(n29701), .B(n28312), .Z(n24002) );
  NOR U29711 ( .A(n29680), .B(n29702), .Z(n29701) );
  XOR U29712 ( .A(n29703), .B(n28318), .Z(n21604) );
  XOR U29713 ( .A(n21665), .B(n29706), .Z(n29557) );
  XOR U29714 ( .A(n18547), .B(n17521), .Z(n29706) );
  XNOR U29715 ( .A(n29707), .B(n21674), .Z(n17521) );
  XOR U29716 ( .A(n25149), .B(n29708), .Z(n21674) );
  IV U29717 ( .A(n21713), .Z(n25149) );
  XNOR U29718 ( .A(n28786), .B(n28158), .Z(n21713) );
  XOR U29719 ( .A(n29709), .B(n29710), .Z(n28158) );
  XOR U29720 ( .A(n25419), .B(n22938), .Z(n29710) );
  XOR U29721 ( .A(n29711), .B(n27089), .Z(n22938) );
  XOR U29722 ( .A(n29712), .B(n29713), .Z(n27089) );
  NOR U29723 ( .A(n29714), .B(n28600), .Z(n29711) );
  XNOR U29724 ( .A(n29715), .B(n27086), .Z(n25419) );
  XNOR U29725 ( .A(n29716), .B(n29717), .Z(n27086) );
  ANDN U29726 ( .B(n29718), .A(n28606), .Z(n29715) );
  XOR U29727 ( .A(n21605), .B(n29719), .Z(n29709) );
  XOR U29728 ( .A(n28574), .B(n25357), .Z(n29719) );
  XNOR U29729 ( .A(n29720), .B(n27080), .Z(n25357) );
  XNOR U29730 ( .A(n29721), .B(n29722), .Z(n27080) );
  NOR U29731 ( .A(n29723), .B(n28597), .Z(n29720) );
  XNOR U29732 ( .A(n29724), .B(n27094), .Z(n28574) );
  XNOR U29733 ( .A(n29725), .B(n29413), .Z(n27094) );
  ANDN U29734 ( .B(n29726), .A(n28595), .Z(n29724) );
  XNOR U29735 ( .A(n29727), .B(n28603), .Z(n21605) );
  ANDN U29736 ( .B(n29728), .A(n29729), .Z(n29727) );
  XOR U29737 ( .A(n29730), .B(n29731), .Z(n28786) );
  XNOR U29738 ( .A(n26877), .B(n25506), .Z(n29731) );
  XOR U29739 ( .A(n29732), .B(n28582), .Z(n25506) );
  NOR U29740 ( .A(n27270), .B(n27269), .Z(n29732) );
  XOR U29741 ( .A(n29733), .B(n29734), .Z(n27269) );
  XNOR U29742 ( .A(n29735), .B(n28590), .Z(n26877) );
  ANDN U29743 ( .B(n27673), .A(n28591), .Z(n29735) );
  XOR U29744 ( .A(n29736), .B(n29737), .Z(n28591) );
  XOR U29745 ( .A(n23791), .B(n29738), .Z(n29730) );
  XOR U29746 ( .A(n27239), .B(n25203), .Z(n29738) );
  XNOR U29747 ( .A(n29739), .B(n28579), .Z(n25203) );
  XOR U29748 ( .A(n29740), .B(n29741), .Z(n27275) );
  XOR U29749 ( .A(n29742), .B(n29743), .Z(n27239) );
  ANDN U29750 ( .B(n28785), .A(n29744), .Z(n29742) );
  XNOR U29751 ( .A(n29745), .B(n28587), .Z(n23791) );
  ANDN U29752 ( .B(n27281), .A(n27279), .Z(n29745) );
  XNOR U29753 ( .A(n29746), .B(n29747), .Z(n27279) );
  ANDN U29754 ( .B(n26112), .A(n21673), .Z(n29707) );
  XOR U29755 ( .A(n29748), .B(n21680), .Z(n18547) );
  XOR U29756 ( .A(n27804), .B(n24390), .Z(n21680) );
  XNOR U29757 ( .A(n29749), .B(n27789), .Z(n27804) );
  NOR U29758 ( .A(n27931), .B(n27630), .Z(n29749) );
  XOR U29759 ( .A(n29750), .B(n29519), .Z(n27630) );
  IV U29760 ( .A(n29751), .Z(n27931) );
  AND U29761 ( .A(n22103), .B(n21681), .Z(n29748) );
  XNOR U29762 ( .A(n29130), .B(n25465), .Z(n21681) );
  IV U29763 ( .A(n23985), .Z(n25465) );
  XNOR U29764 ( .A(n29752), .B(n29753), .Z(n29130) );
  ANDN U29765 ( .B(n29754), .A(n29755), .Z(n29752) );
  XOR U29766 ( .A(n29756), .B(n23079), .Z(n22103) );
  XOR U29767 ( .A(n26564), .B(n26880), .Z(n23079) );
  XNOR U29768 ( .A(n29757), .B(n29758), .Z(n26880) );
  XOR U29769 ( .A(n26405), .B(n26725), .Z(n29758) );
  XOR U29770 ( .A(n29759), .B(n29223), .Z(n26725) );
  ANDN U29771 ( .B(n28845), .A(n29224), .Z(n29759) );
  XOR U29772 ( .A(n29760), .B(n29227), .Z(n26405) );
  XOR U29773 ( .A(n25074), .B(n29761), .Z(n29757) );
  XOR U29774 ( .A(n25049), .B(n26713), .Z(n29761) );
  XNOR U29775 ( .A(n29762), .B(n29218), .Z(n26713) );
  XOR U29776 ( .A(n29763), .B(n29372), .Z(n25049) );
  ANDN U29777 ( .B(n28841), .A(n29371), .Z(n29763) );
  XNOR U29778 ( .A(n29764), .B(n29765), .Z(n25074) );
  ANDN U29779 ( .B(n28858), .A(n29766), .Z(n29764) );
  XOR U29780 ( .A(n29767), .B(n29768), .Z(n26564) );
  XNOR U29781 ( .A(n25879), .B(n25779), .Z(n29768) );
  XNOR U29782 ( .A(n29769), .B(n29246), .Z(n25779) );
  ANDN U29783 ( .B(n26214), .A(n29247), .Z(n29769) );
  XNOR U29784 ( .A(n29770), .B(n29244), .Z(n25879) );
  ANDN U29785 ( .B(n26210), .A(n29243), .Z(n29770) );
  XNOR U29786 ( .A(n29212), .B(n29771), .Z(n29767) );
  XOR U29787 ( .A(n21729), .B(n24261), .Z(n29771) );
  XNOR U29788 ( .A(n29772), .B(n29773), .Z(n24261) );
  ANDN U29789 ( .B(n29774), .A(n29236), .Z(n29772) );
  XNOR U29790 ( .A(n29775), .B(n29233), .Z(n21729) );
  ANDN U29791 ( .B(n29776), .A(n29232), .Z(n29775) );
  XOR U29792 ( .A(n29777), .B(n29241), .Z(n29212) );
  XNOR U29793 ( .A(n29778), .B(n20872), .Z(n21665) );
  IV U29794 ( .A(n21683), .Z(n20872) );
  XOR U29795 ( .A(n26010), .B(n29779), .Z(n21683) );
  IV U29796 ( .A(n24633), .Z(n26010) );
  XNOR U29797 ( .A(n27874), .B(n29780), .Z(n24633) );
  XOR U29798 ( .A(n29781), .B(n29782), .Z(n27874) );
  XNOR U29799 ( .A(n21598), .B(n26467), .Z(n29782) );
  XNOR U29800 ( .A(n29783), .B(n29784), .Z(n26467) );
  ANDN U29801 ( .B(n28084), .A(n28083), .Z(n29783) );
  XNOR U29802 ( .A(n29785), .B(n29786), .Z(n21598) );
  ANDN U29803 ( .B(n28089), .A(n28087), .Z(n29785) );
  XOR U29804 ( .A(n23860), .B(n29787), .Z(n29781) );
  XOR U29805 ( .A(n25796), .B(n24975), .Z(n29787) );
  XNOR U29806 ( .A(n29788), .B(n29789), .Z(n24975) );
  NOR U29807 ( .A(n29790), .B(n28071), .Z(n29788) );
  XNOR U29808 ( .A(n29791), .B(n29792), .Z(n25796) );
  NOR U29809 ( .A(n29793), .B(n28079), .Z(n29791) );
  XOR U29810 ( .A(n29794), .B(n29795), .Z(n23860) );
  ANDN U29811 ( .B(n28076), .A(n28074), .Z(n29794) );
  AND U29812 ( .A(n21684), .B(n22105), .Z(n29778) );
  XOR U29813 ( .A(n21718), .B(n29796), .Z(n22105) );
  IV U29814 ( .A(n23322), .Z(n21718) );
  XNOR U29815 ( .A(n29797), .B(n22401), .Z(n21684) );
  IV U29816 ( .A(n25227), .Z(n22401) );
  XNOR U29817 ( .A(n29798), .B(n29799), .Z(n26782) );
  XOR U29818 ( .A(n23963), .B(n24392), .Z(n29799) );
  XOR U29819 ( .A(n29800), .B(n29801), .Z(n24392) );
  ANDN U29820 ( .B(n29802), .A(n29803), .Z(n29800) );
  XNOR U29821 ( .A(n29804), .B(n29805), .Z(n23963) );
  ANDN U29822 ( .B(n29806), .A(n29807), .Z(n29804) );
  XOR U29823 ( .A(n29808), .B(n29809), .Z(n29798) );
  XNOR U29824 ( .A(n24021), .B(n26374), .Z(n29809) );
  XOR U29825 ( .A(n29810), .B(n29811), .Z(n26374) );
  NOR U29826 ( .A(n29812), .B(n29813), .Z(n29810) );
  XNOR U29827 ( .A(n29814), .B(n29815), .Z(n24021) );
  ANDN U29828 ( .B(n29816), .A(n29817), .Z(n29814) );
  XOR U29829 ( .A(n29818), .B(n29819), .Z(n26530) );
  XNOR U29830 ( .A(n23844), .B(n24197), .Z(n29819) );
  XNOR U29831 ( .A(n29820), .B(n28037), .Z(n24197) );
  ANDN U29832 ( .B(n29821), .A(n29822), .Z(n29820) );
  XNOR U29833 ( .A(n29823), .B(n28864), .Z(n23844) );
  NOR U29834 ( .A(n29824), .B(n29825), .Z(n29823) );
  XOR U29835 ( .A(n25883), .B(n29826), .Z(n29818) );
  XOR U29836 ( .A(n24003), .B(n27581), .Z(n29826) );
  XNOR U29837 ( .A(n29827), .B(n27573), .Z(n27581) );
  XNOR U29838 ( .A(n29830), .B(n29831), .Z(n24003) );
  AND U29839 ( .A(n29832), .B(n29833), .Z(n29830) );
  XNOR U29840 ( .A(n29834), .B(n29835), .Z(n25883) );
  ANDN U29841 ( .B(n29836), .A(n29837), .Z(n29834) );
  XOR U29842 ( .A(n29838), .B(n21673), .Z(n22107) );
  XOR U29843 ( .A(n29839), .B(n25424), .Z(n21673) );
  ANDN U29844 ( .B(n24466), .A(n26112), .Z(n29838) );
  XOR U29845 ( .A(n24571), .B(n26306), .Z(n26112) );
  XNOR U29846 ( .A(n29840), .B(n28192), .Z(n26306) );
  NOR U29847 ( .A(n29841), .B(n29842), .Z(n29840) );
  IV U29848 ( .A(n24432), .Z(n24571) );
  XOR U29849 ( .A(n25709), .B(n29843), .Z(n24432) );
  XOR U29850 ( .A(n29844), .B(n29845), .Z(n25709) );
  XOR U29851 ( .A(n27162), .B(n29846), .Z(n29845) );
  XOR U29852 ( .A(n29847), .B(n29848), .Z(n27162) );
  AND U29853 ( .A(n26325), .B(n26323), .Z(n29847) );
  XNOR U29854 ( .A(n26974), .B(n29849), .Z(n29844) );
  XOR U29855 ( .A(n24873), .B(n27010), .Z(n29849) );
  XOR U29856 ( .A(n29850), .B(n29443), .Z(n27010) );
  ANDN U29857 ( .B(n26329), .A(n26328), .Z(n29850) );
  IV U29858 ( .A(n29851), .Z(n26328) );
  XNOR U29859 ( .A(n29852), .B(n29440), .Z(n24873) );
  ANDN U29860 ( .B(n26319), .A(n26320), .Z(n29852) );
  XNOR U29861 ( .A(n29853), .B(n29432), .Z(n26974) );
  AND U29862 ( .A(n26336), .B(n26338), .Z(n29853) );
  XOR U29863 ( .A(n26135), .B(n28331), .Z(n24466) );
  XOR U29864 ( .A(n29854), .B(n27716), .Z(n28331) );
  ANDN U29865 ( .B(n29855), .A(n29856), .Z(n29854) );
  XNOR U29866 ( .A(n23168), .B(n17699), .Z(n13505) );
  XOR U29867 ( .A(n26144), .B(n22856), .Z(n17699) );
  XNOR U29868 ( .A(n29857), .B(n29858), .Z(n22856) );
  XNOR U29869 ( .A(n19400), .B(n22033), .Z(n29858) );
  XNOR U29870 ( .A(n29859), .B(n23274), .Z(n22033) );
  XOR U29871 ( .A(n28678), .B(n25839), .Z(n23274) );
  XNOR U29872 ( .A(n29860), .B(n29861), .Z(n25521) );
  XOR U29873 ( .A(n27920), .B(n24750), .Z(n29861) );
  XNOR U29874 ( .A(n29862), .B(n29126), .Z(n24750) );
  ANDN U29875 ( .B(n28682), .A(n28680), .Z(n29862) );
  XNOR U29876 ( .A(n29863), .B(n29755), .Z(n27920) );
  ANDN U29877 ( .B(n29864), .A(n29865), .Z(n29863) );
  XNOR U29878 ( .A(n29866), .B(n29867), .Z(n29860) );
  XNOR U29879 ( .A(n23488), .B(n26186), .Z(n29867) );
  XOR U29880 ( .A(n29868), .B(n29869), .Z(n26186) );
  XNOR U29881 ( .A(n29870), .B(n29123), .Z(n23488) );
  AND U29882 ( .A(n28687), .B(n28685), .Z(n29870) );
  XNOR U29883 ( .A(n29871), .B(n29872), .Z(n26779) );
  XNOR U29884 ( .A(n24984), .B(n26563), .Z(n29872) );
  XNOR U29885 ( .A(n29873), .B(n29105), .Z(n26563) );
  ANDN U29886 ( .B(n29874), .A(n27417), .Z(n29873) );
  XNOR U29887 ( .A(n29875), .B(n29117), .Z(n24984) );
  NOR U29888 ( .A(n27429), .B(n27430), .Z(n29875) );
  XOR U29889 ( .A(n24041), .B(n29876), .Z(n29871) );
  XOR U29890 ( .A(n23732), .B(n24813), .Z(n29876) );
  XNOR U29891 ( .A(n29877), .B(n29878), .Z(n24813) );
  ANDN U29892 ( .B(n27425), .A(n27426), .Z(n29877) );
  XNOR U29893 ( .A(n29879), .B(n29111), .Z(n23732) );
  AND U29894 ( .A(n27421), .B(n27423), .Z(n29879) );
  XOR U29895 ( .A(n29880), .B(n29115), .Z(n24041) );
  ANDN U29896 ( .B(n27414), .A(n27412), .Z(n29880) );
  XNOR U29897 ( .A(n29881), .B(n29864), .Z(n28678) );
  ANDN U29898 ( .B(n29865), .A(n29882), .Z(n29881) );
  ANDN U29899 ( .B(n24084), .A(n25318), .Z(n29859) );
  XNOR U29900 ( .A(n27216), .B(n23878), .Z(n25318) );
  XNOR U29901 ( .A(n27908), .B(n29883), .Z(n23878) );
  XOR U29902 ( .A(n29884), .B(n29885), .Z(n27908) );
  XNOR U29903 ( .A(n22214), .B(n27358), .Z(n29885) );
  XNOR U29904 ( .A(n29886), .B(n29887), .Z(n27358) );
  ANDN U29905 ( .B(n29888), .A(n29889), .Z(n29886) );
  XOR U29906 ( .A(n29890), .B(n29891), .Z(n22214) );
  NOR U29907 ( .A(n29892), .B(n29893), .Z(n29890) );
  XOR U29908 ( .A(n25240), .B(n29894), .Z(n29884) );
  XOR U29909 ( .A(n25594), .B(n27847), .Z(n29894) );
  XNOR U29910 ( .A(n29895), .B(n29896), .Z(n27847) );
  ANDN U29911 ( .B(n29897), .A(n29898), .Z(n29895) );
  XOR U29912 ( .A(n29899), .B(n29900), .Z(n25594) );
  XNOR U29913 ( .A(n29903), .B(n29904), .Z(n25240) );
  ANDN U29914 ( .B(n29905), .A(n29906), .Z(n29903) );
  XOR U29915 ( .A(n29907), .B(n29908), .Z(n27216) );
  ANDN U29916 ( .B(n29909), .A(n29910), .Z(n29907) );
  XOR U29917 ( .A(n29424), .B(n24492), .Z(n24084) );
  IV U29918 ( .A(n25144), .Z(n24492) );
  XOR U29919 ( .A(n26107), .B(n29911), .Z(n25144) );
  XOR U29920 ( .A(n29912), .B(n29913), .Z(n26107) );
  XOR U29921 ( .A(n24694), .B(n25084), .Z(n29913) );
  XOR U29922 ( .A(n29914), .B(n26858), .Z(n25084) );
  XOR U29923 ( .A(n29915), .B(n29916), .Z(n26858) );
  XNOR U29924 ( .A(n28739), .B(n29917), .Z(n25847) );
  XOR U29925 ( .A(n29918), .B(n29919), .Z(n25846) );
  XNOR U29926 ( .A(n29921), .B(n29922), .Z(n26854) );
  NOR U29927 ( .A(n29923), .B(n25860), .Z(n29920) );
  XOR U29928 ( .A(n29924), .B(n29925), .Z(n25860) );
  IV U29929 ( .A(n25862), .Z(n29923) );
  XOR U29930 ( .A(n25680), .B(n29928), .Z(n29912) );
  XNOR U29931 ( .A(n27453), .B(n26227), .Z(n29928) );
  XOR U29932 ( .A(n29929), .B(n27462), .Z(n26227) );
  XOR U29933 ( .A(n29930), .B(n29931), .Z(n27462) );
  ANDN U29934 ( .B(n26104), .A(n26105), .Z(n29929) );
  XNOR U29935 ( .A(n29932), .B(n28432), .Z(n26105) );
  XNOR U29936 ( .A(n29933), .B(n29934), .Z(n26104) );
  XOR U29937 ( .A(n29935), .B(n26851), .Z(n27453) );
  XOR U29938 ( .A(n29936), .B(n29937), .Z(n26851) );
  NOR U29939 ( .A(n25857), .B(n25856), .Z(n29935) );
  XOR U29940 ( .A(n29938), .B(n29939), .Z(n25856) );
  XOR U29941 ( .A(n29940), .B(n29941), .Z(n25857) );
  XNOR U29942 ( .A(n29942), .B(n26846), .Z(n25680) );
  XNOR U29943 ( .A(n29943), .B(n29944), .Z(n26846) );
  XOR U29944 ( .A(n29945), .B(n29946), .Z(n25852) );
  XNOR U29945 ( .A(n29947), .B(n29948), .Z(n25850) );
  XNOR U29946 ( .A(n29949), .B(n27348), .Z(n29424) );
  ANDN U29947 ( .B(n26722), .A(n29950), .Z(n29949) );
  XNOR U29948 ( .A(n29951), .B(n23286), .Z(n19400) );
  XOR U29949 ( .A(n29952), .B(n27796), .Z(n23286) );
  ANDN U29950 ( .B(n24093), .A(n24865), .Z(n29951) );
  XOR U29951 ( .A(n29953), .B(n25177), .Z(n24865) );
  IV U29952 ( .A(n21819), .Z(n25177) );
  XOR U29953 ( .A(n29955), .B(n29956), .Z(n29843) );
  XOR U29954 ( .A(n25785), .B(n24165), .Z(n29956) );
  XOR U29955 ( .A(n29957), .B(n28181), .Z(n24165) );
  ANDN U29956 ( .B(n26305), .A(n26303), .Z(n29957) );
  XOR U29957 ( .A(n29924), .B(n29958), .Z(n26303) );
  IV U29958 ( .A(n29959), .Z(n29924) );
  XNOR U29959 ( .A(n29960), .B(n28184), .Z(n25785) );
  ANDN U29960 ( .B(n26311), .A(n28185), .Z(n29960) );
  XOR U29961 ( .A(n29961), .B(n29962), .Z(n28185) );
  XOR U29962 ( .A(n26262), .B(n29963), .Z(n29955) );
  XNOR U29963 ( .A(n25758), .B(n25251), .Z(n29963) );
  XOR U29964 ( .A(n29964), .B(n28193), .Z(n25251) );
  ANDN U29965 ( .B(n29842), .A(n28192), .Z(n29964) );
  XOR U29966 ( .A(n29965), .B(n29966), .Z(n28192) );
  XNOR U29967 ( .A(n29967), .B(n28189), .Z(n25758) );
  ANDN U29968 ( .B(n26314), .A(n26313), .Z(n29967) );
  XOR U29969 ( .A(n29968), .B(n29969), .Z(n26313) );
  XOR U29970 ( .A(n29970), .B(n28196), .Z(n26262) );
  ANDN U29971 ( .B(n26301), .A(n26299), .Z(n29970) );
  XOR U29972 ( .A(n29971), .B(n29067), .Z(n26299) );
  XOR U29973 ( .A(n27314), .B(n25974), .Z(n24093) );
  XNOR U29974 ( .A(n29972), .B(n29973), .Z(n25974) );
  XOR U29975 ( .A(n29974), .B(n29975), .Z(n27314) );
  NOR U29976 ( .A(n29976), .B(n29977), .Z(n29974) );
  XNOR U29977 ( .A(n22361), .B(n29978), .Z(n29857) );
  XOR U29978 ( .A(n19280), .B(n21622), .Z(n29978) );
  XNOR U29979 ( .A(n29979), .B(n23267), .Z(n21622) );
  XOR U29980 ( .A(n29980), .B(n28725), .Z(n23267) );
  XNOR U29981 ( .A(n29981), .B(n29982), .Z(n28271) );
  XOR U29982 ( .A(n25449), .B(n27140), .Z(n29982) );
  XNOR U29983 ( .A(n29983), .B(n29548), .Z(n27140) );
  NOR U29984 ( .A(n29984), .B(n29547), .Z(n29983) );
  XOR U29985 ( .A(n29985), .B(n29551), .Z(n25449) );
  NOR U29986 ( .A(n29986), .B(n29987), .Z(n29985) );
  XNOR U29987 ( .A(n25165), .B(n29988), .Z(n29981) );
  XNOR U29988 ( .A(n25795), .B(n25947), .Z(n29988) );
  XNOR U29989 ( .A(n29989), .B(n29555), .Z(n25947) );
  ANDN U29990 ( .B(n29556), .A(n29990), .Z(n29989) );
  XOR U29991 ( .A(n29991), .B(n29542), .Z(n25795) );
  NOR U29992 ( .A(n29992), .B(n29993), .Z(n29991) );
  XNOR U29993 ( .A(n29994), .B(n29539), .Z(n25165) );
  ANDN U29994 ( .B(n29995), .A(n29996), .Z(n29994) );
  XNOR U29995 ( .A(n29997), .B(n29998), .Z(n27729) );
  XNOR U29996 ( .A(n24382), .B(n23691), .Z(n29998) );
  XNOR U29997 ( .A(n29999), .B(n28670), .Z(n23691) );
  XOR U29998 ( .A(n30000), .B(n30001), .Z(n28670) );
  XOR U29999 ( .A(n30002), .B(n27152), .Z(n24382) );
  XNOR U30000 ( .A(n30003), .B(n30004), .Z(n27152) );
  ANDN U30001 ( .B(n27153), .A(n29394), .Z(n30002) );
  XOR U30002 ( .A(n25115), .B(n30005), .Z(n29997) );
  XNOR U30003 ( .A(n23744), .B(n25076), .Z(n30005) );
  XNOR U30004 ( .A(n30006), .B(n27147), .Z(n25076) );
  XOR U30005 ( .A(n30007), .B(n28473), .Z(n27147) );
  ANDN U30006 ( .B(n27148), .A(n29404), .Z(n30006) );
  XOR U30007 ( .A(n30008), .B(n27161), .Z(n23744) );
  XNOR U30008 ( .A(n30009), .B(n30010), .Z(n27161) );
  NOR U30009 ( .A(n30011), .B(n27160), .Z(n30008) );
  XNOR U30010 ( .A(n30012), .B(n27156), .Z(n25115) );
  XOR U30011 ( .A(n30013), .B(n30014), .Z(n27156) );
  ANDN U30012 ( .B(n27157), .A(n29399), .Z(n30012) );
  ANDN U30013 ( .B(n24859), .A(n24082), .Z(n29979) );
  XNOR U30014 ( .A(n22635), .B(n26208), .Z(n24082) );
  XNOR U30015 ( .A(n30015), .B(n29776), .Z(n26208) );
  ANDN U30016 ( .B(n30016), .A(n29231), .Z(n30015) );
  XNOR U30017 ( .A(n29455), .B(n26381), .Z(n24859) );
  XNOR U30018 ( .A(n30017), .B(n28350), .Z(n29455) );
  AND U30019 ( .A(n30018), .B(n30019), .Z(n30017) );
  XNOR U30020 ( .A(n30020), .B(n23278), .Z(n19280) );
  XOR U30021 ( .A(n30021), .B(n23346), .Z(n23278) );
  ANDN U30022 ( .B(n24855), .A(n25324), .Z(n30020) );
  XOR U30023 ( .A(n30022), .B(n25757), .Z(n25324) );
  XNOR U30024 ( .A(n30023), .B(n30024), .Z(n25937) );
  XOR U30025 ( .A(n28976), .B(n26379), .Z(n30024) );
  XNOR U30026 ( .A(n30025), .B(n29004), .Z(n26379) );
  ANDN U30027 ( .B(n26161), .A(n26162), .Z(n30025) );
  XOR U30028 ( .A(n30026), .B(n30027), .Z(n26161) );
  XOR U30029 ( .A(n30028), .B(n30029), .Z(n28976) );
  XOR U30030 ( .A(n23713), .B(n30030), .Z(n30023) );
  XOR U30031 ( .A(n26609), .B(n27095), .Z(n30030) );
  XNOR U30032 ( .A(n30031), .B(n30032), .Z(n27095) );
  NOR U30033 ( .A(n26157), .B(n26158), .Z(n30031) );
  XNOR U30034 ( .A(n28987), .B(n30033), .Z(n26157) );
  XOR U30035 ( .A(n30034), .B(n29009), .Z(n26609) );
  ANDN U30036 ( .B(n26166), .A(n30035), .Z(n30034) );
  XOR U30037 ( .A(n30036), .B(n28897), .Z(n26166) );
  XNOR U30038 ( .A(n30037), .B(n29001), .Z(n23713) );
  ANDN U30039 ( .B(n26170), .A(n26172), .Z(n30037) );
  XOR U30040 ( .A(n30038), .B(n30039), .Z(n26170) );
  XNOR U30041 ( .A(n30040), .B(n30041), .Z(n27204) );
  XNOR U30042 ( .A(n27906), .B(n26458), .Z(n30041) );
  XOR U30043 ( .A(n30042), .B(n29902), .Z(n26458) );
  ANDN U30044 ( .B(n29901), .A(n30043), .Z(n30042) );
  XOR U30045 ( .A(n30044), .B(n29905), .Z(n27906) );
  NOR U30046 ( .A(n30045), .B(n30046), .Z(n30044) );
  XNOR U30047 ( .A(n26130), .B(n30047), .Z(n30040) );
  XNOR U30048 ( .A(n24624), .B(n27305), .Z(n30047) );
  XNOR U30049 ( .A(n30048), .B(n29888), .Z(n27305) );
  ANDN U30050 ( .B(n30049), .A(n30050), .Z(n30048) );
  XOR U30051 ( .A(n30051), .B(n29897), .Z(n24624) );
  XNOR U30052 ( .A(n30053), .B(n29892), .Z(n26130) );
  IV U30053 ( .A(n30054), .Z(n29892) );
  ANDN U30054 ( .B(n29893), .A(n30055), .Z(n30053) );
  XOR U30055 ( .A(n26932), .B(n27002), .Z(n24855) );
  IV U30056 ( .A(n25356), .Z(n27002) );
  XNOR U30057 ( .A(n30056), .B(n27449), .Z(n26932) );
  IV U30058 ( .A(n30057), .Z(n27449) );
  ANDN U30059 ( .B(n27024), .A(n30058), .Z(n30056) );
  XNOR U30060 ( .A(n30059), .B(n23283), .Z(n22361) );
  XOR U30061 ( .A(n30060), .B(n26017), .Z(n23283) );
  IV U30062 ( .A(n28900), .Z(n26017) );
  XNOR U30063 ( .A(n30061), .B(n30062), .Z(n27264) );
  XNOR U30064 ( .A(n21714), .B(n25150), .Z(n30062) );
  XOR U30065 ( .A(n30063), .B(n28606), .Z(n25150) );
  XOR U30066 ( .A(n29943), .B(n30064), .Z(n28606) );
  ANDN U30067 ( .B(n27084), .A(n29718), .Z(n30063) );
  XOR U30068 ( .A(n30065), .B(n28597), .Z(n21714) );
  XOR U30069 ( .A(n30066), .B(n30067), .Z(n28597) );
  XOR U30070 ( .A(n24881), .B(n30068), .Z(n30061) );
  XNOR U30071 ( .A(n24457), .B(n29708), .Z(n30068) );
  XNOR U30072 ( .A(n30069), .B(n29729), .Z(n29708) );
  IV U30073 ( .A(n28604), .Z(n29729) );
  XOR U30074 ( .A(n30070), .B(n30071), .Z(n28604) );
  NOR U30075 ( .A(n30072), .B(n29728), .Z(n30069) );
  XOR U30076 ( .A(n30073), .B(n28600), .Z(n24457) );
  XOR U30077 ( .A(n30074), .B(n30075), .Z(n28600) );
  ANDN U30078 ( .B(n29714), .A(n27088), .Z(n30073) );
  XOR U30079 ( .A(n30076), .B(n28595), .Z(n24881) );
  XOR U30080 ( .A(n30077), .B(n30078), .Z(n28595) );
  ANDN U30081 ( .B(n27092), .A(n29726), .Z(n30076) );
  XNOR U30082 ( .A(n30079), .B(n30080), .Z(n28543) );
  XOR U30083 ( .A(n25804), .B(n26553), .Z(n30080) );
  XOR U30084 ( .A(n30081), .B(n30082), .Z(n26553) );
  ANDN U30085 ( .B(n30083), .A(n30084), .Z(n30081) );
  XNOR U30086 ( .A(n30085), .B(n30086), .Z(n25804) );
  XNOR U30087 ( .A(n28157), .B(n30089), .Z(n30079) );
  XNOR U30088 ( .A(n24945), .B(n27452), .Z(n30089) );
  XNOR U30089 ( .A(n30090), .B(n30091), .Z(n27452) );
  NOR U30090 ( .A(n30092), .B(n30093), .Z(n30090) );
  XNOR U30091 ( .A(n30094), .B(n30095), .Z(n24945) );
  ANDN U30092 ( .B(n30096), .A(n30097), .Z(n30094) );
  XNOR U30093 ( .A(n30098), .B(n30099), .Z(n28157) );
  ANDN U30094 ( .B(n30100), .A(n30101), .Z(n30098) );
  ANDN U30095 ( .B(n24090), .A(n24868), .Z(n30059) );
  XOR U30096 ( .A(n24442), .B(n29525), .Z(n24868) );
  XOR U30097 ( .A(n30102), .B(n30103), .Z(n29525) );
  XOR U30098 ( .A(n30104), .B(n30105), .Z(n28285) );
  XOR U30099 ( .A(n30107), .B(n30108), .Z(n28009) );
  XNOR U30100 ( .A(n23138), .B(n25728), .Z(n30108) );
  XNOR U30101 ( .A(n30109), .B(n30110), .Z(n25728) );
  ANDN U30102 ( .B(n29555), .A(n29554), .Z(n30109) );
  XNOR U30103 ( .A(n30111), .B(n30112), .Z(n29555) );
  XNOR U30104 ( .A(n30113), .B(n30114), .Z(n23138) );
  NOR U30105 ( .A(n29551), .B(n29550), .Z(n30113) );
  XNOR U30106 ( .A(n30115), .B(n30116), .Z(n29551) );
  XOR U30107 ( .A(n23800), .B(n30117), .Z(n30107) );
  XNOR U30108 ( .A(n26561), .B(n29389), .Z(n30117) );
  XNOR U30109 ( .A(n30118), .B(n30119), .Z(n29389) );
  ANDN U30110 ( .B(n29539), .A(n29537), .Z(n30118) );
  XOR U30111 ( .A(n30120), .B(n30121), .Z(n29539) );
  XNOR U30112 ( .A(n30122), .B(n30123), .Z(n26561) );
  ANDN U30113 ( .B(n29548), .A(n29546), .Z(n30122) );
  XNOR U30114 ( .A(n30124), .B(n30125), .Z(n29548) );
  XNOR U30115 ( .A(n30126), .B(n30127), .Z(n23800) );
  ANDN U30116 ( .B(n29541), .A(n29542), .Z(n30126) );
  XOR U30117 ( .A(n30128), .B(n30129), .Z(n29542) );
  XOR U30118 ( .A(n28583), .B(n23727), .Z(n24090) );
  IV U30119 ( .A(n24747), .Z(n23727) );
  XNOR U30120 ( .A(n26004), .B(n30130), .Z(n24747) );
  XOR U30121 ( .A(n30131), .B(n30132), .Z(n26004) );
  XOR U30122 ( .A(n24578), .B(n22496), .Z(n30132) );
  XNOR U30123 ( .A(n30133), .B(n27271), .Z(n22496) );
  XNOR U30124 ( .A(n30134), .B(n29413), .Z(n28582) );
  XOR U30125 ( .A(n30135), .B(n27280), .Z(n24578) );
  XNOR U30126 ( .A(n30136), .B(n28881), .Z(n28587) );
  XNOR U30127 ( .A(n24368), .B(n30137), .Z(n30131) );
  XNOR U30128 ( .A(n24600), .B(n28415), .Z(n30137) );
  XOR U30129 ( .A(n30138), .B(n28784), .Z(n28415) );
  ANDN U30130 ( .B(n29743), .A(n30139), .Z(n30138) );
  XNOR U30131 ( .A(n30140), .B(n27277), .Z(n24600) );
  ANDN U30132 ( .B(n28578), .A(n28579), .Z(n30140) );
  XOR U30133 ( .A(n30141), .B(n30142), .Z(n28579) );
  XOR U30134 ( .A(n30143), .B(n27672), .Z(n24368) );
  ANDN U30135 ( .B(n28589), .A(n28590), .Z(n30143) );
  XOR U30136 ( .A(n30144), .B(n30145), .Z(n28590) );
  XOR U30137 ( .A(n30146), .B(n30139), .Z(n28583) );
  ANDN U30138 ( .B(n29744), .A(n29743), .Z(n30146) );
  XOR U30139 ( .A(n30147), .B(n30148), .Z(n29743) );
  IV U30140 ( .A(n28783), .Z(n29744) );
  XNOR U30141 ( .A(n30149), .B(n30150), .Z(n28783) );
  XNOR U30142 ( .A(n30151), .B(n30152), .Z(n26144) );
  XOR U30143 ( .A(n18617), .B(n16044), .Z(n30152) );
  XOR U30144 ( .A(n30153), .B(n23302), .Z(n16044) );
  XNOR U30145 ( .A(n27038), .B(n25706), .Z(n23302) );
  NOR U30146 ( .A(n30155), .B(n30156), .Z(n30154) );
  XOR U30147 ( .A(n30157), .B(n26030), .Z(n23161) );
  IV U30148 ( .A(n26718), .Z(n26030) );
  XNOR U30149 ( .A(n30158), .B(n21216), .Z(n23163) );
  XOR U30150 ( .A(n29390), .B(n30159), .Z(n21216) );
  XNOR U30151 ( .A(n30160), .B(n30161), .Z(n29390) );
  XNOR U30152 ( .A(n30162), .B(n25067), .Z(n30161) );
  XNOR U30153 ( .A(n30163), .B(n29995), .Z(n25067) );
  AND U30154 ( .A(n30119), .B(n29537), .Z(n30163) );
  XNOR U30155 ( .A(n30164), .B(n30165), .Z(n29537) );
  XOR U30156 ( .A(n23970), .B(n30166), .Z(n30160) );
  XNOR U30157 ( .A(n23997), .B(n25056), .Z(n30166) );
  XNOR U30158 ( .A(n30167), .B(n29990), .Z(n25056) );
  ANDN U30159 ( .B(n29554), .A(n30168), .Z(n30167) );
  XOR U30160 ( .A(n30169), .B(n30170), .Z(n29554) );
  XNOR U30161 ( .A(n30171), .B(n29993), .Z(n23997) );
  ANDN U30162 ( .B(n30127), .A(n29541), .Z(n30171) );
  XOR U30163 ( .A(n30172), .B(n30004), .Z(n29541) );
  XNOR U30164 ( .A(n30173), .B(n29984), .Z(n23970) );
  AND U30165 ( .A(n29546), .B(n30123), .Z(n30173) );
  XOR U30166 ( .A(n30174), .B(n30175), .Z(n29546) );
  XNOR U30167 ( .A(n30176), .B(n23296), .Z(n18617) );
  XOR U30168 ( .A(n27759), .B(n23974), .Z(n23296) );
  XOR U30169 ( .A(n30177), .B(n25102), .Z(n23974) );
  XNOR U30170 ( .A(n30178), .B(n30179), .Z(n25102) );
  XNOR U30171 ( .A(n21595), .B(n30180), .Z(n30179) );
  XNOR U30172 ( .A(n30181), .B(n26426), .Z(n21595) );
  NOR U30173 ( .A(n27755), .B(n27756), .Z(n30181) );
  XOR U30174 ( .A(n22895), .B(n30182), .Z(n30178) );
  XNOR U30175 ( .A(n26184), .B(n22324), .Z(n30182) );
  XNOR U30176 ( .A(n30183), .B(n26434), .Z(n22324) );
  IV U30177 ( .A(n30184), .Z(n26434) );
  ANDN U30178 ( .B(n27750), .A(n27749), .Z(n30183) );
  XOR U30179 ( .A(n30185), .B(n30186), .Z(n26184) );
  NOR U30180 ( .A(n30187), .B(n27752), .Z(n30185) );
  XNOR U30181 ( .A(n30188), .B(n26430), .Z(n22895) );
  ANDN U30182 ( .B(n27746), .A(n27745), .Z(n30188) );
  IV U30183 ( .A(n30189), .Z(n27746) );
  XNOR U30184 ( .A(n30190), .B(n30191), .Z(n27759) );
  ANDN U30185 ( .B(n23165), .A(n23166), .Z(n30176) );
  XNOR U30186 ( .A(n27243), .B(n23065), .Z(n23166) );
  XNOR U30187 ( .A(n30193), .B(n30194), .Z(n30130) );
  XNOR U30188 ( .A(n28675), .B(n25154), .Z(n30194) );
  XOR U30189 ( .A(n30195), .B(n26991), .Z(n25154) );
  XOR U30190 ( .A(n30196), .B(n29304), .Z(n26991) );
  IV U30191 ( .A(n30197), .Z(n29304) );
  XNOR U30192 ( .A(n30198), .B(n30199), .Z(n27246) );
  XOR U30193 ( .A(n30200), .B(n30201), .Z(n27245) );
  XOR U30194 ( .A(n30202), .B(n25530), .Z(n28675) );
  XOR U30195 ( .A(n30203), .B(n30204), .Z(n25530) );
  XOR U30196 ( .A(n27669), .B(n30205), .Z(n30193) );
  XNOR U30197 ( .A(n27794), .B(n24797), .Z(n30205) );
  XNOR U30198 ( .A(n30206), .B(n27330), .Z(n24797) );
  ANDN U30199 ( .B(n27249), .A(n28810), .Z(n30206) );
  XOR U30200 ( .A(n30209), .B(n30210), .Z(n28810) );
  XOR U30201 ( .A(n30211), .B(n30212), .Z(n27249) );
  XNOR U30202 ( .A(n30213), .B(n27886), .Z(n27794) );
  XNOR U30203 ( .A(n30214), .B(n30215), .Z(n27886) );
  ANDN U30204 ( .B(n27254), .A(n28703), .Z(n30213) );
  XOR U30205 ( .A(n30216), .B(n30217), .Z(n28703) );
  XOR U30206 ( .A(n30218), .B(n30219), .Z(n27254) );
  XOR U30207 ( .A(n30220), .B(n25535), .Z(n27669) );
  XOR U30208 ( .A(n30221), .B(n29329), .Z(n25535) );
  ANDN U30209 ( .B(n27258), .A(n27257), .Z(n30220) );
  XOR U30210 ( .A(n30222), .B(n30223), .Z(n27257) );
  XNOR U30211 ( .A(n30224), .B(n29948), .Z(n27258) );
  XOR U30212 ( .A(n30226), .B(n28706), .Z(n27243) );
  XOR U30213 ( .A(n30227), .B(n30228), .Z(n28706) );
  ANDN U30214 ( .B(n28806), .A(n25529), .Z(n30226) );
  XNOR U30215 ( .A(n30229), .B(n30230), .Z(n25529) );
  XNOR U30216 ( .A(n30231), .B(n30232), .Z(n28806) );
  XNOR U30217 ( .A(n24749), .B(n29866), .Z(n23165) );
  XNOR U30218 ( .A(n30233), .B(n29133), .Z(n29866) );
  ANDN U30219 ( .B(n28693), .A(n28694), .Z(n30233) );
  IV U30220 ( .A(n23489), .Z(n24749) );
  XOR U30221 ( .A(n27887), .B(n26565), .Z(n23489) );
  XNOR U30222 ( .A(n30234), .B(n30235), .Z(n26565) );
  XOR U30223 ( .A(n25344), .B(n25794), .Z(n30235) );
  XOR U30224 ( .A(n30236), .B(n29106), .Z(n25794) );
  NOR U30225 ( .A(n29874), .B(n29105), .Z(n30236) );
  XOR U30226 ( .A(n30237), .B(n30116), .Z(n29105) );
  IV U30227 ( .A(n27416), .Z(n29874) );
  XOR U30228 ( .A(n30238), .B(n30239), .Z(n27416) );
  XNOR U30229 ( .A(n30240), .B(n30241), .Z(n25344) );
  ANDN U30230 ( .B(n29878), .A(n27425), .Z(n30240) );
  XOR U30231 ( .A(n30242), .B(n30243), .Z(n27425) );
  XNOR U30232 ( .A(n25499), .B(n30244), .Z(n30234) );
  XNOR U30233 ( .A(n23039), .B(n25871), .Z(n30244) );
  XNOR U30234 ( .A(n30245), .B(n29114), .Z(n25871) );
  ANDN U30235 ( .B(n27412), .A(n29115), .Z(n30245) );
  XNOR U30236 ( .A(n30246), .B(n30247), .Z(n29115) );
  XNOR U30237 ( .A(n30248), .B(n30249), .Z(n27412) );
  XNOR U30238 ( .A(n30250), .B(n29110), .Z(n23039) );
  ANDN U30239 ( .B(n29111), .A(n27421), .Z(n30250) );
  XOR U30240 ( .A(n30251), .B(n30252), .Z(n27421) );
  XNOR U30241 ( .A(n30253), .B(n30254), .Z(n29111) );
  XOR U30242 ( .A(n30255), .B(n29118), .Z(n25499) );
  IV U30243 ( .A(n30256), .Z(n29118) );
  ANDN U30244 ( .B(n27429), .A(n29117), .Z(n30255) );
  XNOR U30245 ( .A(n30257), .B(n30258), .Z(n29117) );
  XNOR U30246 ( .A(n30259), .B(n30260), .Z(n27429) );
  XOR U30247 ( .A(n30261), .B(n30262), .Z(n27887) );
  XNOR U30248 ( .A(n24638), .B(n22347), .Z(n30262) );
  XNOR U30249 ( .A(n30263), .B(n29132), .Z(n22347) );
  NOR U30250 ( .A(n28693), .B(n29133), .Z(n30263) );
  XOR U30251 ( .A(n30264), .B(n30265), .Z(n29133) );
  XOR U30252 ( .A(n30266), .B(n30267), .Z(n28693) );
  XNOR U30253 ( .A(n30268), .B(n29754), .Z(n24638) );
  ANDN U30254 ( .B(n29755), .A(n29864), .Z(n30268) );
  XOR U30255 ( .A(n30269), .B(n30071), .Z(n29864) );
  XOR U30256 ( .A(n30270), .B(n28750), .Z(n29755) );
  XNOR U30257 ( .A(n24527), .B(n30271), .Z(n30261) );
  XOR U30258 ( .A(n22632), .B(n29100), .Z(n30271) );
  XOR U30259 ( .A(n30272), .B(n29127), .Z(n29100) );
  XNOR U30260 ( .A(n30273), .B(n28793), .Z(n29126) );
  XNOR U30261 ( .A(n30274), .B(n30275), .Z(n28680) );
  XNOR U30262 ( .A(n30276), .B(n29124), .Z(n22632) );
  NOR U30263 ( .A(n29123), .B(n28685), .Z(n30276) );
  XOR U30264 ( .A(n30277), .B(n30278), .Z(n28685) );
  XOR U30265 ( .A(n30279), .B(n29948), .Z(n29123) );
  XOR U30266 ( .A(n30280), .B(n30281), .Z(n24527) );
  AND U30267 ( .A(n28689), .B(n29869), .Z(n30280) );
  XNOR U30268 ( .A(n30282), .B(n29050), .Z(n28689) );
  XOR U30269 ( .A(n24077), .B(n30283), .Z(n30151) );
  XOR U30270 ( .A(n17938), .B(n15544), .Z(n30283) );
  XOR U30271 ( .A(n30284), .B(n23293), .Z(n15544) );
  XOR U30272 ( .A(n30285), .B(n24272), .Z(n23293) );
  IV U30273 ( .A(n26619), .Z(n24272) );
  XOR U30274 ( .A(n28960), .B(n28270), .Z(n26619) );
  XOR U30275 ( .A(n30286), .B(n30287), .Z(n28270) );
  XNOR U30276 ( .A(n25363), .B(n27645), .Z(n30287) );
  XOR U30277 ( .A(n30288), .B(n29269), .Z(n27645) );
  XOR U30278 ( .A(n30289), .B(n30290), .Z(n29269) );
  ANDN U30279 ( .B(n29140), .A(n30291), .Z(n30288) );
  XNOR U30280 ( .A(n30292), .B(n28911), .Z(n25363) );
  XOR U30281 ( .A(n30293), .B(n30294), .Z(n28911) );
  ANDN U30282 ( .B(n30295), .A(n30296), .Z(n30292) );
  XOR U30283 ( .A(n27904), .B(n30297), .Z(n30286) );
  XOR U30284 ( .A(n29253), .B(n26449), .Z(n30297) );
  XNOR U30285 ( .A(n30298), .B(n28922), .Z(n26449) );
  XOR U30286 ( .A(n30299), .B(n30300), .Z(n28922) );
  ANDN U30287 ( .B(n29138), .A(n29276), .Z(n30298) );
  XNOR U30288 ( .A(n30301), .B(n28918), .Z(n29253) );
  XNOR U30289 ( .A(n30302), .B(n30303), .Z(n28918) );
  NOR U30290 ( .A(n30304), .B(n29150), .Z(n30301) );
  XNOR U30291 ( .A(n30305), .B(n28907), .Z(n27904) );
  XNOR U30292 ( .A(n30306), .B(n30307), .Z(n28907) );
  NOR U30293 ( .A(n29259), .B(n29145), .Z(n30305) );
  XOR U30294 ( .A(n30308), .B(n30309), .Z(n28960) );
  XNOR U30295 ( .A(n22493), .B(n26368), .Z(n30309) );
  XNOR U30296 ( .A(n30310), .B(n27045), .Z(n26368) );
  IV U30297 ( .A(n30311), .Z(n27045) );
  ANDN U30298 ( .B(n26964), .A(n26962), .Z(n30310) );
  XNOR U30299 ( .A(n30312), .B(n30155), .Z(n22493) );
  ANDN U30300 ( .B(n26972), .A(n30313), .Z(n30312) );
  XOR U30301 ( .A(n23135), .B(n30314), .Z(n30308) );
  XNOR U30302 ( .A(n30315), .B(n23858), .Z(n30314) );
  XNOR U30303 ( .A(n30316), .B(n27048), .Z(n23858) );
  AND U30304 ( .A(n26968), .B(n26966), .Z(n30316) );
  XNOR U30305 ( .A(n30317), .B(n27040), .Z(n23135) );
  ANDN U30306 ( .B(n26959), .A(n26957), .Z(n30317) );
  XOR U30307 ( .A(n30318), .B(n23810), .Z(n23171) );
  XOR U30308 ( .A(n30320), .B(n30321), .Z(n26252) );
  XNOR U30309 ( .A(n24562), .B(n26217), .Z(n30321) );
  XNOR U30310 ( .A(n30322), .B(n27402), .Z(n26217) );
  ANDN U30311 ( .B(n30323), .A(n27400), .Z(n30322) );
  XOR U30312 ( .A(n30324), .B(n27406), .Z(n24562) );
  NOR U30313 ( .A(n27405), .B(n30325), .Z(n30324) );
  XOR U30314 ( .A(n24488), .B(n30326), .Z(n30320) );
  XNOR U30315 ( .A(n23076), .B(n27387), .Z(n30326) );
  XOR U30316 ( .A(n30327), .B(n30328), .Z(n27387) );
  ANDN U30317 ( .B(n27395), .A(n30329), .Z(n30327) );
  XNOR U30318 ( .A(n30330), .B(n27536), .Z(n23076) );
  NOR U30319 ( .A(n27537), .B(n30331), .Z(n30330) );
  XOR U30320 ( .A(n30332), .B(n30333), .Z(n24488) );
  NOR U30321 ( .A(n30334), .B(n30335), .Z(n30332) );
  XOR U30322 ( .A(n28112), .B(n26224), .Z(n23173) );
  IV U30323 ( .A(n24231), .Z(n26224) );
  XNOR U30324 ( .A(n29973), .B(n26540), .Z(n24231) );
  XNOR U30325 ( .A(n30336), .B(n30337), .Z(n26540) );
  XNOR U30326 ( .A(n27167), .B(n26873), .Z(n30337) );
  XNOR U30327 ( .A(n30338), .B(n30339), .Z(n26873) );
  ANDN U30328 ( .B(n30340), .A(n30341), .Z(n30338) );
  XNOR U30329 ( .A(n30342), .B(n30343), .Z(n27167) );
  NOR U30330 ( .A(n30344), .B(n30345), .Z(n30342) );
  XNOR U30331 ( .A(n26011), .B(n30346), .Z(n30336) );
  XOR U30332 ( .A(n24634), .B(n29779), .Z(n30346) );
  XNOR U30333 ( .A(n30347), .B(n30348), .Z(n29779) );
  NOR U30334 ( .A(n30349), .B(n30350), .Z(n30347) );
  XNOR U30335 ( .A(n30351), .B(n30352), .Z(n24634) );
  ANDN U30336 ( .B(n30353), .A(n30354), .Z(n30351) );
  XNOR U30337 ( .A(n30355), .B(n30356), .Z(n26011) );
  NOR U30338 ( .A(n30357), .B(n30358), .Z(n30355) );
  XNOR U30339 ( .A(n30359), .B(n30360), .Z(n29973) );
  XNOR U30340 ( .A(n30361), .B(n25228), .Z(n30360) );
  XNOR U30341 ( .A(n30362), .B(n30363), .Z(n25228) );
  AND U30342 ( .A(n28125), .B(n27697), .Z(n30362) );
  XNOR U30343 ( .A(n30364), .B(n30365), .Z(n27697) );
  XOR U30344 ( .A(n24269), .B(n30366), .Z(n30359) );
  XOR U30345 ( .A(n21371), .B(n28539), .Z(n30366) );
  XNOR U30346 ( .A(n30367), .B(n30368), .Z(n28539) );
  ANDN U30347 ( .B(n28123), .A(n30369), .Z(n30367) );
  IV U30348 ( .A(n27693), .Z(n28123) );
  XNOR U30349 ( .A(n30370), .B(n30371), .Z(n27693) );
  XOR U30350 ( .A(n30372), .B(n30373), .Z(n21371) );
  NOR U30351 ( .A(n28115), .B(n28114), .Z(n30372) );
  XOR U30352 ( .A(n30374), .B(n30375), .Z(n28115) );
  XOR U30353 ( .A(n30376), .B(n30377), .Z(n24269) );
  AND U30354 ( .A(n30378), .B(n27687), .Z(n30376) );
  XNOR U30355 ( .A(n30379), .B(n30378), .Z(n28112) );
  NOR U30356 ( .A(n27688), .B(n27687), .Z(n30379) );
  XOR U30357 ( .A(n30380), .B(n30381), .Z(n27687) );
  XOR U30358 ( .A(n30382), .B(n23300), .Z(n17938) );
  IV U30359 ( .A(n25560), .Z(n23300) );
  XOR U30360 ( .A(n26381), .B(n29450), .Z(n25560) );
  AND U30361 ( .A(n30384), .B(n30385), .Z(n30383) );
  XNOR U30362 ( .A(n30386), .B(n26461), .Z(n26381) );
  XNOR U30363 ( .A(n30387), .B(n30388), .Z(n26461) );
  XNOR U30364 ( .A(n21727), .B(n25188), .Z(n30388) );
  XOR U30365 ( .A(n30389), .B(n30390), .Z(n25188) );
  NOR U30366 ( .A(n29465), .B(n29467), .Z(n30389) );
  XOR U30367 ( .A(n30391), .B(n30392), .Z(n21727) );
  XOR U30368 ( .A(n22350), .B(n30393), .Z(n30387) );
  XOR U30369 ( .A(n30394), .B(n25722), .Z(n30393) );
  XNOR U30370 ( .A(n30395), .B(n30396), .Z(n25722) );
  ANDN U30371 ( .B(n29474), .A(n29476), .Z(n30395) );
  XNOR U30372 ( .A(n30397), .B(n30398), .Z(n22350) );
  NOR U30373 ( .A(n30399), .B(n29483), .Z(n30397) );
  ANDN U30374 ( .B(n23177), .A(n23175), .Z(n30382) );
  XNOR U30375 ( .A(n30400), .B(n22960), .Z(n23175) );
  XNOR U30376 ( .A(n27438), .B(n26585), .Z(n22960) );
  XNOR U30377 ( .A(n30401), .B(n30402), .Z(n26585) );
  XNOR U30378 ( .A(n26043), .B(n30403), .Z(n30402) );
  XNOR U30379 ( .A(n30404), .B(n30405), .Z(n26043) );
  AND U30380 ( .A(n29194), .B(n30406), .Z(n30404) );
  XOR U30381 ( .A(n24964), .B(n30407), .Z(n30401) );
  XNOR U30382 ( .A(n25927), .B(n25517), .Z(n30407) );
  XNOR U30383 ( .A(n30408), .B(n30409), .Z(n25517) );
  XOR U30384 ( .A(n30411), .B(n30412), .Z(n25927) );
  ANDN U30385 ( .B(n30413), .A(n29184), .Z(n30411) );
  IV U30386 ( .A(n30414), .Z(n29184) );
  XNOR U30387 ( .A(n30415), .B(n30416), .Z(n24964) );
  XOR U30388 ( .A(n30419), .B(n30420), .Z(n27438) );
  XNOR U30389 ( .A(n26445), .B(n25692), .Z(n30420) );
  XNOR U30390 ( .A(n30421), .B(n30422), .Z(n25692) );
  ANDN U30391 ( .B(n28293), .A(n30423), .Z(n30421) );
  XNOR U30392 ( .A(n30424), .B(n30425), .Z(n26445) );
  ANDN U30393 ( .B(n28063), .A(n30426), .Z(n30424) );
  XNOR U30394 ( .A(n27011), .B(n30427), .Z(n30419) );
  XOR U30395 ( .A(n25270), .B(n24744), .Z(n30427) );
  XNOR U30396 ( .A(n30428), .B(n30429), .Z(n24744) );
  ANDN U30397 ( .B(n26649), .A(n30430), .Z(n30428) );
  XNOR U30398 ( .A(n30431), .B(n30432), .Z(n25270) );
  ANDN U30399 ( .B(n26653), .A(n30433), .Z(n30431) );
  XNOR U30400 ( .A(n30434), .B(n30435), .Z(n27011) );
  ANDN U30401 ( .B(n26660), .A(n30436), .Z(n30434) );
  XNOR U30402 ( .A(n25016), .B(n30437), .Z(n23177) );
  IV U30403 ( .A(n23686), .Z(n25016) );
  XOR U30404 ( .A(n27074), .B(n26867), .Z(n23686) );
  XNOR U30405 ( .A(n30438), .B(n30439), .Z(n26867) );
  XNOR U30406 ( .A(n25830), .B(n25744), .Z(n30439) );
  XNOR U30407 ( .A(n30440), .B(n30441), .Z(n25744) );
  ANDN U30408 ( .B(n30442), .A(n30443), .Z(n30440) );
  XNOR U30409 ( .A(n30444), .B(n30445), .Z(n25830) );
  ANDN U30410 ( .B(n30446), .A(n30447), .Z(n30444) );
  XOR U30411 ( .A(n30448), .B(n30449), .Z(n30438) );
  XNOR U30412 ( .A(n25814), .B(n25427), .Z(n30449) );
  XNOR U30413 ( .A(n30450), .B(n30451), .Z(n25427) );
  ANDN U30414 ( .B(n30452), .A(n30453), .Z(n30450) );
  XOR U30415 ( .A(n30454), .B(n30455), .Z(n25814) );
  NOR U30416 ( .A(n30456), .B(n30457), .Z(n30454) );
  XNOR U30417 ( .A(n30458), .B(n30459), .Z(n27074) );
  XNOR U30418 ( .A(n23909), .B(n23428), .Z(n30459) );
  XNOR U30419 ( .A(n30460), .B(n30461), .Z(n23428) );
  NOR U30420 ( .A(n30462), .B(n30463), .Z(n30460) );
  XOR U30421 ( .A(n30464), .B(n30100), .Z(n23909) );
  ANDN U30422 ( .B(n30465), .A(n30466), .Z(n30464) );
  XOR U30423 ( .A(n26411), .B(n30467), .Z(n30458) );
  XOR U30424 ( .A(n24556), .B(n26183), .Z(n30467) );
  XOR U30425 ( .A(n30468), .B(n30083), .Z(n26183) );
  ANDN U30426 ( .B(n30469), .A(n30470), .Z(n30468) );
  XNOR U30427 ( .A(n30471), .B(n30087), .Z(n24556) );
  NOR U30428 ( .A(n30472), .B(n30473), .Z(n30471) );
  XNOR U30429 ( .A(n30474), .B(n30475), .Z(n26411) );
  NOR U30430 ( .A(n30476), .B(n30477), .Z(n30474) );
  XNOR U30431 ( .A(n30478), .B(n24889), .Z(n24077) );
  XNOR U30432 ( .A(n30180), .B(n22325), .Z(n24889) );
  XOR U30433 ( .A(n30480), .B(n30481), .Z(n26082) );
  XOR U30434 ( .A(n25330), .B(n22525), .Z(n30481) );
  XNOR U30435 ( .A(n30482), .B(n26425), .Z(n22525) );
  AND U30436 ( .A(n27755), .B(n26426), .Z(n30482) );
  XNOR U30437 ( .A(n30483), .B(n30484), .Z(n26426) );
  XNOR U30438 ( .A(n30306), .B(n30485), .Z(n27755) );
  XOR U30439 ( .A(n26438), .B(n30486), .Z(n25330) );
  XOR U30440 ( .A(n30487), .B(n21688), .Z(n30486) );
  ANDN U30441 ( .B(n27742), .A(n30488), .Z(n30487) );
  XNOR U30442 ( .A(n24509), .B(n30489), .Z(n30480) );
  XNOR U30443 ( .A(n25823), .B(n23720), .Z(n30489) );
  XNOR U30444 ( .A(n30490), .B(n26435), .Z(n23720) );
  ANDN U30445 ( .B(n27749), .A(n30184), .Z(n30490) );
  XOR U30446 ( .A(n30491), .B(n30492), .Z(n30184) );
  XOR U30447 ( .A(n30493), .B(n30494), .Z(n27749) );
  XOR U30448 ( .A(n30495), .B(n26442), .Z(n25823) );
  ANDN U30449 ( .B(n27752), .A(n30186), .Z(n30495) );
  IV U30450 ( .A(n26443), .Z(n30186) );
  XOR U30451 ( .A(n30496), .B(n28736), .Z(n26443) );
  XNOR U30452 ( .A(n30497), .B(n29166), .Z(n27752) );
  XOR U30453 ( .A(n30498), .B(n26429), .Z(n24509) );
  XOR U30454 ( .A(n30499), .B(n30500), .Z(n26430) );
  XOR U30455 ( .A(n30501), .B(n30502), .Z(n27745) );
  XNOR U30456 ( .A(n30503), .B(n26439), .Z(n30180) );
  IV U30457 ( .A(n30488), .Z(n26439) );
  XOR U30458 ( .A(n30504), .B(n30505), .Z(n30488) );
  NOR U30459 ( .A(n27743), .B(n27742), .Z(n30503) );
  XNOR U30460 ( .A(n30506), .B(n30507), .Z(n27742) );
  ANDN U30461 ( .B(n25557), .A(n24876), .Z(n30478) );
  XNOR U30462 ( .A(n30508), .B(n25557), .Z(n23168) );
  XNOR U30463 ( .A(n26738), .B(n26238), .Z(n25557) );
  IV U30464 ( .A(n22988), .Z(n26238) );
  XNOR U30465 ( .A(n30509), .B(n28654), .Z(n22988) );
  XNOR U30466 ( .A(n30510), .B(n30511), .Z(n28654) );
  XNOR U30467 ( .A(n26102), .B(n28923), .Z(n30511) );
  XOR U30468 ( .A(n30512), .B(n28948), .Z(n28923) );
  XNOR U30469 ( .A(n30513), .B(n30514), .Z(n28948) );
  AND U30470 ( .A(n28949), .B(n27838), .Z(n30512) );
  XNOR U30471 ( .A(n30515), .B(n29308), .Z(n26102) );
  IV U30472 ( .A(n29296), .Z(n29308) );
  XOR U30473 ( .A(n30516), .B(n30517), .Z(n29296) );
  NOR U30474 ( .A(n26742), .B(n26741), .Z(n30515) );
  XOR U30475 ( .A(n30518), .B(n30204), .Z(n26741) );
  XOR U30476 ( .A(n30519), .B(n30520), .Z(n26742) );
  XNOR U30477 ( .A(n27168), .B(n30521), .Z(n30510) );
  XNOR U30478 ( .A(n24386), .B(n22824), .Z(n30521) );
  XNOR U30479 ( .A(n30522), .B(n28953), .Z(n22824) );
  XNOR U30480 ( .A(n30523), .B(n30524), .Z(n28953) );
  XOR U30481 ( .A(n30525), .B(n29934), .Z(n26746) );
  XOR U30482 ( .A(n28747), .B(n30526), .Z(n26745) );
  XOR U30483 ( .A(n30527), .B(n28955), .Z(n24386) );
  XOR U30484 ( .A(n30528), .B(n30529), .Z(n28955) );
  NOR U30485 ( .A(n26737), .B(n26735), .Z(n30527) );
  XOR U30486 ( .A(n30530), .B(n30531), .Z(n26735) );
  XOR U30487 ( .A(n30532), .B(n30267), .Z(n26737) );
  XOR U30488 ( .A(n30533), .B(n28957), .Z(n27168) );
  XOR U30489 ( .A(n30534), .B(n30535), .Z(n28957) );
  XOR U30490 ( .A(n30536), .B(n30537), .Z(n27833) );
  XNOR U30491 ( .A(n30538), .B(n30539), .Z(n28776) );
  XNOR U30492 ( .A(n30540), .B(n28949), .Z(n26738) );
  XNOR U30493 ( .A(n30541), .B(n30542), .Z(n28949) );
  NOR U30494 ( .A(n27840), .B(n27838), .Z(n30540) );
  XOR U30495 ( .A(n30543), .B(n30544), .Z(n27838) );
  XOR U30496 ( .A(n30545), .B(n29032), .Z(n27840) );
  XNOR U30497 ( .A(n29562), .B(n24193), .Z(n24876) );
  XNOR U30498 ( .A(n25590), .B(n28902), .Z(n24193) );
  XNOR U30499 ( .A(n30546), .B(n30547), .Z(n28902) );
  XOR U30500 ( .A(n25747), .B(n27677), .Z(n30547) );
  XOR U30501 ( .A(n30548), .B(n30549), .Z(n27677) );
  ANDN U30502 ( .B(n29581), .A(n28259), .Z(n30548) );
  XOR U30503 ( .A(n30550), .B(n30112), .Z(n28259) );
  XNOR U30504 ( .A(n30551), .B(n30552), .Z(n25747) );
  NOR U30505 ( .A(n29590), .B(n28263), .Z(n30551) );
  XNOR U30506 ( .A(n30553), .B(n30554), .Z(n28263) );
  XOR U30507 ( .A(n28059), .B(n30555), .Z(n30546) );
  XOR U30508 ( .A(n23854), .B(n26124), .Z(n30555) );
  XOR U30509 ( .A(n30556), .B(n30557), .Z(n26124) );
  NOR U30510 ( .A(n29578), .B(n28267), .Z(n30556) );
  XNOR U30511 ( .A(n30558), .B(n30559), .Z(n28267) );
  XNOR U30512 ( .A(n30560), .B(n30561), .Z(n23854) );
  NOR U30513 ( .A(n28254), .B(n29587), .Z(n30560) );
  XNOR U30514 ( .A(n30562), .B(n30563), .Z(n28254) );
  XNOR U30515 ( .A(n30564), .B(n30565), .Z(n28059) );
  NOR U30516 ( .A(n29585), .B(n28250), .Z(n30564) );
  XOR U30517 ( .A(n30566), .B(n30567), .Z(n28250) );
  XNOR U30518 ( .A(n30568), .B(n30569), .Z(n25590) );
  XNOR U30519 ( .A(n23030), .B(n22533), .Z(n30569) );
  XNOR U30520 ( .A(n30570), .B(n30571), .Z(n22533) );
  ANDN U30521 ( .B(n30572), .A(n29574), .Z(n30570) );
  XNOR U30522 ( .A(n30573), .B(n30574), .Z(n29574) );
  XNOR U30523 ( .A(n30575), .B(n30576), .Z(n23030) );
  NOR U30524 ( .A(n28530), .B(n30577), .Z(n30575) );
  XOR U30525 ( .A(n25786), .B(n30578), .Z(n30568) );
  XNOR U30526 ( .A(n30579), .B(n22955), .Z(n30578) );
  XOR U30527 ( .A(n30580), .B(n30581), .Z(n22955) );
  NOR U30528 ( .A(n29564), .B(n28520), .Z(n30580) );
  XOR U30529 ( .A(n30582), .B(n30583), .Z(n28520) );
  XNOR U30530 ( .A(n30584), .B(n30585), .Z(n25786) );
  ANDN U30531 ( .B(n29567), .A(n29592), .Z(n30584) );
  IV U30532 ( .A(n29568), .Z(n29592) );
  XOR U30533 ( .A(n30586), .B(n30587), .Z(n29568) );
  IV U30534 ( .A(n30588), .Z(n29567) );
  XNOR U30535 ( .A(n30589), .B(n30577), .Z(n29562) );
  ANDN U30536 ( .B(n28530), .A(n28531), .Z(n30589) );
  XNOR U30537 ( .A(n30590), .B(n28814), .Z(n28530) );
  IV U30538 ( .A(n24888), .Z(n24878) );
  XOR U30539 ( .A(n25603), .B(n29641), .Z(n24888) );
  XOR U30540 ( .A(n30591), .B(n29367), .Z(n29641) );
  ANDN U30541 ( .B(n30592), .A(n30593), .Z(n30591) );
  IV U30542 ( .A(n28537), .Z(n25603) );
  XOR U30543 ( .A(n30594), .B(n27700), .Z(n28537) );
  XOR U30544 ( .A(n30595), .B(n30596), .Z(n27700) );
  XNOR U30545 ( .A(n26228), .B(n24345), .Z(n30596) );
  XNOR U30546 ( .A(n30597), .B(n27326), .Z(n24345) );
  AND U30547 ( .A(n29387), .B(n27327), .Z(n30597) );
  XNOR U30548 ( .A(n30598), .B(n27319), .Z(n26228) );
  ANDN U30549 ( .B(n30599), .A(n27318), .Z(n30598) );
  XOR U30550 ( .A(n26861), .B(n30600), .Z(n30595) );
  XNOR U30551 ( .A(n26123), .B(n26062), .Z(n30600) );
  XNOR U30552 ( .A(n30601), .B(n27323), .Z(n26062) );
  ANDN U30553 ( .B(n29378), .A(n27322), .Z(n30601) );
  XNOR U30554 ( .A(n30602), .B(n27916), .Z(n26123) );
  XNOR U30555 ( .A(n30603), .B(n29976), .Z(n26861) );
  AND U30556 ( .A(n30604), .B(n29977), .Z(n30603) );
  XNOR U30557 ( .A(n30605), .B(n16219), .Z(n11227) );
  IV U30558 ( .A(n14720), .Z(n16219) );
  XNOR U30559 ( .A(n16770), .B(n25626), .Z(n14720) );
  XNOR U30560 ( .A(n30606), .B(n23202), .Z(n25626) );
  NOR U30561 ( .A(n25647), .B(n25648), .Z(n30606) );
  XNOR U30562 ( .A(n30607), .B(n22892), .Z(n25648) );
  XOR U30563 ( .A(n26815), .B(n27051), .Z(n22892) );
  XNOR U30564 ( .A(n30608), .B(n30609), .Z(n27051) );
  XNOR U30565 ( .A(n26780), .B(n25118), .Z(n30609) );
  XNOR U30566 ( .A(n30610), .B(n30611), .Z(n25118) );
  ANDN U30567 ( .B(n30612), .A(n30613), .Z(n30610) );
  XOR U30568 ( .A(n30614), .B(n30615), .Z(n26780) );
  ANDN U30569 ( .B(n30616), .A(n29802), .Z(n30614) );
  XNOR U30570 ( .A(n23071), .B(n30617), .Z(n30608) );
  XOR U30571 ( .A(n25994), .B(n25939), .Z(n30617) );
  XOR U30572 ( .A(n30618), .B(n29806), .Z(n25939) );
  ANDN U30573 ( .B(n29807), .A(n30619), .Z(n30618) );
  XNOR U30574 ( .A(n30620), .B(n29817), .Z(n25994) );
  ANDN U30575 ( .B(n30621), .A(n29816), .Z(n30620) );
  ANDN U30576 ( .B(n29813), .A(n30623), .Z(n30622) );
  XOR U30577 ( .A(n30624), .B(n30625), .Z(n26815) );
  XOR U30578 ( .A(n29797), .B(n25338), .Z(n30625) );
  XOR U30579 ( .A(n30626), .B(n29837), .Z(n25338) );
  XOR U30580 ( .A(n30627), .B(n29825), .Z(n29797) );
  AND U30581 ( .A(n29824), .B(n28862), .Z(n30627) );
  XOR U30582 ( .A(n25226), .B(n30628), .Z(n30624) );
  XOR U30583 ( .A(n22400), .B(n25495), .Z(n30628) );
  XOR U30584 ( .A(n30629), .B(n29832), .Z(n25495) );
  ANDN U30585 ( .B(n30630), .A(n29833), .Z(n30629) );
  XNOR U30586 ( .A(n30631), .B(n29829), .Z(n22400) );
  AND U30587 ( .A(n29828), .B(n27571), .Z(n30631) );
  XNOR U30588 ( .A(n30632), .B(n29821), .Z(n25226) );
  AND U30589 ( .A(n28035), .B(n29822), .Z(n30632) );
  XOR U30590 ( .A(n22384), .B(n22998), .Z(n16770) );
  XNOR U30591 ( .A(n30633), .B(n30634), .Z(n22998) );
  XOR U30592 ( .A(n20371), .B(n16584), .Z(n30634) );
  XOR U30593 ( .A(n30635), .B(n22451), .Z(n16584) );
  XOR U30594 ( .A(n25745), .B(n30448), .Z(n22451) );
  XNOR U30595 ( .A(n30636), .B(n30637), .Z(n30448) );
  NOR U30596 ( .A(n30638), .B(n30639), .Z(n30636) );
  XOR U30597 ( .A(n30640), .B(n26413), .Z(n25745) );
  XNOR U30598 ( .A(n30641), .B(n30642), .Z(n26413) );
  XNOR U30599 ( .A(n28899), .B(n26016), .Z(n30642) );
  XNOR U30600 ( .A(n30643), .B(n30101), .Z(n26016) );
  ANDN U30601 ( .B(n30466), .A(n30100), .Z(n30643) );
  XOR U30602 ( .A(n30644), .B(n30645), .Z(n30100) );
  XOR U30603 ( .A(n30646), .B(n30088), .Z(n28899) );
  AND U30604 ( .A(n30087), .B(n30472), .Z(n30646) );
  XOR U30605 ( .A(n30647), .B(n28885), .Z(n30087) );
  XNOR U30606 ( .A(n26481), .B(n30648), .Z(n30641) );
  XOR U30607 ( .A(n26869), .B(n30060), .Z(n30648) );
  XNOR U30608 ( .A(n30649), .B(n30093), .Z(n30060) );
  ANDN U30609 ( .B(n30476), .A(n30475), .Z(n30649) );
  IV U30610 ( .A(n30092), .Z(n30475) );
  XOR U30611 ( .A(n30650), .B(n30651), .Z(n30092) );
  XNOR U30612 ( .A(n30652), .B(n30084), .Z(n26869) );
  ANDN U30613 ( .B(n30470), .A(n30083), .Z(n30652) );
  XOR U30614 ( .A(n30653), .B(n30654), .Z(n30083) );
  XOR U30615 ( .A(n30655), .B(n30096), .Z(n26481) );
  ANDN U30616 ( .B(n30462), .A(n30461), .Z(n30655) );
  IV U30617 ( .A(n30097), .Z(n30461) );
  XOR U30618 ( .A(n30227), .B(n30656), .Z(n30097) );
  IV U30619 ( .A(n30657), .Z(n30227) );
  NOR U30620 ( .A(n25641), .B(n23213), .Z(n30635) );
  XNOR U30621 ( .A(n30658), .B(n30659), .Z(n26795) );
  XOR U30622 ( .A(n25880), .B(n27164), .Z(n30659) );
  XOR U30623 ( .A(n30660), .B(n28485), .Z(n27164) );
  NOR U30624 ( .A(n29155), .B(n29173), .Z(n30660) );
  XOR U30625 ( .A(n30661), .B(n30662), .Z(n29155) );
  XNOR U30626 ( .A(n30663), .B(n28487), .Z(n25880) );
  ANDN U30627 ( .B(n28360), .A(n29177), .Z(n30663) );
  XOR U30628 ( .A(n30664), .B(n30014), .Z(n28360) );
  XOR U30629 ( .A(n25454), .B(n30665), .Z(n30658) );
  XOR U30630 ( .A(n24617), .B(n24970), .Z(n30665) );
  XNOR U30631 ( .A(n30666), .B(n28492), .Z(n24970) );
  ANDN U30632 ( .B(n28225), .A(n30667), .Z(n30666) );
  XOR U30633 ( .A(n30066), .B(n30668), .Z(n28225) );
  XNOR U30634 ( .A(n30669), .B(n28494), .Z(n24617) );
  XOR U30635 ( .A(n30670), .B(n30671), .Z(n28221) );
  XNOR U30636 ( .A(n30672), .B(n30673), .Z(n25454) );
  NOR U30637 ( .A(n28232), .B(n29164), .Z(n30672) );
  XNOR U30638 ( .A(n30674), .B(n30675), .Z(n28232) );
  XOR U30639 ( .A(n30676), .B(n30677), .Z(n27583) );
  XOR U30640 ( .A(n22020), .B(n30678), .Z(n30677) );
  XNOR U30641 ( .A(n30679), .B(n30680), .Z(n22020) );
  ANDN U30642 ( .B(n29817), .A(n29815), .Z(n30679) );
  XOR U30643 ( .A(n30681), .B(n30682), .Z(n29817) );
  XOR U30644 ( .A(n24159), .B(n30683), .Z(n30676) );
  XOR U30645 ( .A(n25082), .B(n26139), .Z(n30683) );
  XOR U30646 ( .A(n30684), .B(n30685), .Z(n26139) );
  ANDN U30647 ( .B(n29812), .A(n29811), .Z(n30684) );
  XNOR U30648 ( .A(n30686), .B(n30687), .Z(n29812) );
  XNOR U30649 ( .A(n30688), .B(n30689), .Z(n25082) );
  NOR U30650 ( .A(n30615), .B(n29801), .Z(n30688) );
  IV U30651 ( .A(n29803), .Z(n30615) );
  XOR U30652 ( .A(n30690), .B(n30691), .Z(n29803) );
  XOR U30653 ( .A(n30692), .B(n30693), .Z(n24159) );
  XNOR U30654 ( .A(n30695), .B(n30694), .Z(n29808) );
  NOR U30655 ( .A(n30611), .B(n30612), .Z(n30695) );
  XOR U30656 ( .A(n30696), .B(n30697), .Z(n30611) );
  XOR U30657 ( .A(n24702), .B(n30698), .Z(n25641) );
  XOR U30658 ( .A(n26628), .B(n30699), .Z(n24702) );
  XOR U30659 ( .A(n30700), .B(n30701), .Z(n26628) );
  XOR U30660 ( .A(n25562), .B(n25496), .Z(n30701) );
  XOR U30661 ( .A(n30702), .B(n30703), .Z(n25496) );
  NOR U30662 ( .A(n30704), .B(n30705), .Z(n30702) );
  XOR U30663 ( .A(n30706), .B(n28629), .Z(n25562) );
  ANDN U30664 ( .B(n30707), .A(n30708), .Z(n30706) );
  XOR U30665 ( .A(n23576), .B(n30709), .Z(n30700) );
  XOR U30666 ( .A(n30710), .B(n29310), .Z(n30709) );
  XOR U30667 ( .A(n30711), .B(n28638), .Z(n29310) );
  ANDN U30668 ( .B(n30712), .A(n30713), .Z(n30711) );
  XOR U30669 ( .A(n30714), .B(n28635), .Z(n23576) );
  ANDN U30670 ( .B(n30715), .A(n30716), .Z(n30714) );
  XNOR U30671 ( .A(n30717), .B(n22461), .Z(n20371) );
  XNOR U30672 ( .A(n25490), .B(n30718), .Z(n22461) );
  ANDN U30673 ( .B(n25644), .A(n23218), .Z(n30717) );
  XOR U30674 ( .A(n30719), .B(n25952), .Z(n23218) );
  XOR U30675 ( .A(n29208), .B(n25247), .Z(n25644) );
  AND U30676 ( .A(n27975), .B(n27977), .Z(n30720) );
  XOR U30677 ( .A(n22577), .B(n30721), .Z(n30633) );
  XOR U30678 ( .A(n19561), .B(n15687), .Z(n30721) );
  XNOR U30679 ( .A(n30722), .B(n23208), .Z(n15687) );
  XOR U30680 ( .A(n30723), .B(n23731), .Z(n23208) );
  IV U30681 ( .A(n22793), .Z(n23731) );
  NOR U30682 ( .A(n23207), .B(n25638), .Z(n30722) );
  XOR U30683 ( .A(n29437), .B(n25152), .Z(n25638) );
  XOR U30684 ( .A(n30727), .B(n30728), .Z(n29911) );
  XNOR U30685 ( .A(n27339), .B(n23700), .Z(n30728) );
  XNOR U30686 ( .A(n30729), .B(n26501), .Z(n23700) );
  XNOR U30687 ( .A(n29045), .B(n30730), .Z(n26501) );
  ANDN U30688 ( .B(n27351), .A(n30731), .Z(n30729) );
  XOR U30689 ( .A(n30732), .B(n30243), .Z(n27351) );
  IV U30690 ( .A(n30733), .Z(n30243) );
  XNOR U30691 ( .A(n30734), .B(n26489), .Z(n27339) );
  XNOR U30692 ( .A(n28765), .B(n30735), .Z(n26489) );
  ANDN U30693 ( .B(n27343), .A(n30736), .Z(n30734) );
  XOR U30694 ( .A(n30737), .B(n29927), .Z(n27343) );
  XOR U30695 ( .A(n23989), .B(n30738), .Z(n30727) );
  XOR U30696 ( .A(n24782), .B(n25721), .Z(n30738) );
  XNOR U30697 ( .A(n30739), .B(n26724), .Z(n25721) );
  XNOR U30698 ( .A(n30740), .B(n30687), .Z(n26724) );
  ANDN U30699 ( .B(n27348), .A(n30741), .Z(n30739) );
  XOR U30700 ( .A(n30742), .B(n30743), .Z(n27348) );
  XNOR U30701 ( .A(n30744), .B(n26549), .Z(n24782) );
  XNOR U30702 ( .A(n30745), .B(n30746), .Z(n26549) );
  NOR U30703 ( .A(n27353), .B(n29421), .Z(n30744) );
  XOR U30704 ( .A(n30747), .B(n30748), .Z(n27353) );
  XOR U30705 ( .A(n30749), .B(n26493), .Z(n23989) );
  XOR U30706 ( .A(n30750), .B(n30129), .Z(n26493) );
  NOR U30707 ( .A(n29419), .B(n27345), .Z(n30749) );
  XOR U30708 ( .A(n30751), .B(n30752), .Z(n27345) );
  XOR U30709 ( .A(n30753), .B(n26324), .Z(n29437) );
  ANDN U30710 ( .B(n30754), .A(n29848), .Z(n30753) );
  XOR U30711 ( .A(n27054), .B(n29215), .Z(n23207) );
  XNOR U30712 ( .A(n30755), .B(n28860), .Z(n29215) );
  ANDN U30713 ( .B(n29765), .A(n30756), .Z(n30755) );
  IV U30714 ( .A(n24899), .Z(n27054) );
  XOR U30715 ( .A(n30757), .B(n30758), .Z(n29705) );
  XNOR U30716 ( .A(n24318), .B(n26692), .Z(n30758) );
  XOR U30717 ( .A(n30759), .B(n28413), .Z(n26692) );
  XOR U30718 ( .A(n30760), .B(n30761), .Z(n28413) );
  ANDN U30719 ( .B(n28403), .A(n28822), .Z(n30759) );
  XNOR U30720 ( .A(n30762), .B(n28023), .Z(n24318) );
  XOR U30721 ( .A(n30763), .B(n30764), .Z(n28023) );
  NOR U30722 ( .A(n28409), .B(n28826), .Z(n30762) );
  XOR U30723 ( .A(n23435), .B(n30765), .Z(n30757) );
  XNOR U30724 ( .A(n24521), .B(n24902), .Z(n30765) );
  XOR U30725 ( .A(n30766), .B(n28018), .Z(n24902) );
  XOR U30726 ( .A(n30767), .B(n30768), .Z(n28018) );
  ANDN U30727 ( .B(n28837), .A(n28411), .Z(n30766) );
  XNOR U30728 ( .A(n30769), .B(n28027), .Z(n24521) );
  XOR U30729 ( .A(n30198), .B(n30770), .Z(n28027) );
  XOR U30730 ( .A(n30771), .B(n28031), .Z(n23435) );
  XOR U30731 ( .A(n30772), .B(n30078), .Z(n28031) );
  ANDN U30732 ( .B(n30773), .A(n28829), .Z(n30771) );
  XNOR U30733 ( .A(n30774), .B(n30775), .Z(n26056) );
  XNOR U30734 ( .A(n24179), .B(n26472), .Z(n30775) );
  XOR U30735 ( .A(n30776), .B(n28852), .Z(n26472) );
  NOR U30736 ( .A(n29217), .B(n29218), .Z(n30776) );
  XNOR U30737 ( .A(n30573), .B(n30777), .Z(n29218) );
  IV U30738 ( .A(n28851), .Z(n29217) );
  XOR U30739 ( .A(n30778), .B(n30267), .Z(n28851) );
  XNOR U30740 ( .A(n30779), .B(n30780), .Z(n24179) );
  ANDN U30741 ( .B(n28847), .A(n29223), .Z(n30779) );
  XOR U30742 ( .A(n30781), .B(n30782), .Z(n29223) );
  XOR U30743 ( .A(n30783), .B(n30784), .Z(n28847) );
  XOR U30744 ( .A(n28816), .B(n30785), .Z(n30774) );
  XOR U30745 ( .A(n25242), .B(n24227), .Z(n30785) );
  XNOR U30746 ( .A(n30786), .B(n30787), .Z(n24227) );
  ANDN U30747 ( .B(n29227), .A(n28855), .Z(n30786) );
  XOR U30748 ( .A(n29528), .B(n30788), .Z(n28855) );
  XNOR U30749 ( .A(n30789), .B(n30790), .Z(n29227) );
  XNOR U30750 ( .A(n30791), .B(n28842), .Z(n25242) );
  XOR U30751 ( .A(n30792), .B(n28469), .Z(n28843) );
  XOR U30752 ( .A(n30793), .B(n30794), .Z(n29372) );
  XNOR U30753 ( .A(n30795), .B(n28859), .Z(n28816) );
  ANDN U30754 ( .B(n28860), .A(n29765), .Z(n30795) );
  XOR U30755 ( .A(n30796), .B(n29095), .Z(n29765) );
  XOR U30756 ( .A(n30797), .B(n30798), .Z(n28860) );
  XNOR U30757 ( .A(n30799), .B(n23216), .Z(n19561) );
  XOR U30758 ( .A(n26924), .B(n29383), .Z(n23216) );
  XNOR U30759 ( .A(n30800), .B(n30599), .Z(n29383) );
  NOR U30760 ( .A(n30801), .B(n27317), .Z(n30800) );
  ANDN U30761 ( .B(n25633), .A(n23215), .Z(n30799) );
  XOR U30762 ( .A(n30802), .B(n25206), .Z(n23215) );
  XOR U30763 ( .A(n24455), .B(n30803), .Z(n25633) );
  XOR U30764 ( .A(n30804), .B(n22465), .Z(n22577) );
  XOR U30765 ( .A(n30805), .B(n25026), .Z(n22465) );
  IV U30766 ( .A(n25352), .Z(n25026) );
  NOR U30767 ( .A(n25635), .B(n23210), .Z(n30804) );
  XNOR U30768 ( .A(n29005), .B(n25045), .Z(n23210) );
  XOR U30769 ( .A(n30807), .B(n30808), .Z(n27849) );
  XOR U30770 ( .A(n27337), .B(n24341), .Z(n30808) );
  XOR U30771 ( .A(n30809), .B(n26176), .Z(n24341) );
  ANDN U30772 ( .B(n30810), .A(n30029), .Z(n30809) );
  XNOR U30773 ( .A(n30811), .B(n26167), .Z(n27337) );
  AND U30774 ( .A(n29008), .B(n29009), .Z(n30811) );
  XNOR U30775 ( .A(n30812), .B(n30781), .Z(n29009) );
  XNOR U30776 ( .A(n30813), .B(n30814), .Z(n30807) );
  XOR U30777 ( .A(n24274), .B(n27436), .Z(n30814) );
  XNOR U30778 ( .A(n30815), .B(n26171), .Z(n27436) );
  XOR U30779 ( .A(n30816), .B(n30817), .Z(n29001) );
  XOR U30780 ( .A(n30818), .B(n26163), .Z(n24274) );
  NOR U30781 ( .A(n29003), .B(n29004), .Z(n30818) );
  XOR U30782 ( .A(n30000), .B(n30819), .Z(n29004) );
  IV U30783 ( .A(n30820), .Z(n29003) );
  XNOR U30784 ( .A(n30821), .B(n30810), .Z(n29005) );
  ANDN U30785 ( .B(n30029), .A(n26174), .Z(n30821) );
  XNOR U30786 ( .A(n30822), .B(n30823), .Z(n26174) );
  XNOR U30787 ( .A(n28995), .B(n30824), .Z(n30029) );
  XOR U30788 ( .A(n22645), .B(n27391), .Z(n25635) );
  XNOR U30789 ( .A(n30825), .B(n30826), .Z(n27391) );
  ANDN U30790 ( .B(n30334), .A(n30333), .Z(n30825) );
  IV U30791 ( .A(n22608), .Z(n22645) );
  XOR U30792 ( .A(n28455), .B(n27984), .Z(n22608) );
  XOR U30793 ( .A(n30827), .B(n30828), .Z(n27984) );
  XNOR U30794 ( .A(n24437), .B(n30829), .Z(n30828) );
  XOR U30795 ( .A(n30830), .B(n30831), .Z(n24437) );
  XOR U30796 ( .A(n25275), .B(n30834), .Z(n30827) );
  XOR U30797 ( .A(n26997), .B(n24503), .Z(n30834) );
  XOR U30798 ( .A(n30835), .B(n30836), .Z(n24503) );
  ANDN U30799 ( .B(n30837), .A(n30838), .Z(n30835) );
  XNOR U30800 ( .A(n30839), .B(n30840), .Z(n26997) );
  XNOR U30801 ( .A(n30843), .B(n30844), .Z(n25275) );
  XOR U30802 ( .A(n30847), .B(n30848), .Z(n28455) );
  XOR U30803 ( .A(n24831), .B(n22024), .Z(n30848) );
  XOR U30804 ( .A(n30849), .B(n30850), .Z(n22024) );
  AND U30805 ( .A(n27404), .B(n27406), .Z(n30849) );
  XOR U30806 ( .A(n30851), .B(n30852), .Z(n27406) );
  XNOR U30807 ( .A(n30853), .B(n30854), .Z(n24831) );
  ANDN U30808 ( .B(n27535), .A(n27536), .Z(n30853) );
  XNOR U30809 ( .A(n30855), .B(n30856), .Z(n27536) );
  XOR U30810 ( .A(n25216), .B(n30857), .Z(n30847) );
  XOR U30811 ( .A(n26978), .B(n26286), .Z(n30857) );
  XNOR U30812 ( .A(n30858), .B(n30859), .Z(n26286) );
  AND U30813 ( .A(n30333), .B(n30826), .Z(n30858) );
  XOR U30814 ( .A(n30860), .B(n30861), .Z(n30333) );
  XOR U30815 ( .A(n30862), .B(n30863), .Z(n26978) );
  ANDN U30816 ( .B(n27393), .A(n27394), .Z(n30862) );
  IV U30817 ( .A(n30328), .Z(n27394) );
  XNOR U30818 ( .A(n30866), .B(n30867), .Z(n25216) );
  ANDN U30819 ( .B(n27399), .A(n27402), .Z(n30866) );
  XOR U30820 ( .A(n30868), .B(n30869), .Z(n27402) );
  XOR U30821 ( .A(n30870), .B(n30871), .Z(n22384) );
  XOR U30822 ( .A(n20223), .B(n20128), .Z(n30871) );
  XOR U30823 ( .A(n30872), .B(n23201), .Z(n20128) );
  XOR U30824 ( .A(n30873), .B(n25952), .Z(n23201) );
  IV U30825 ( .A(n26570), .Z(n25952) );
  XOR U30826 ( .A(n27964), .B(n27898), .Z(n26570) );
  XOR U30827 ( .A(n30874), .B(n30875), .Z(n27898) );
  XNOR U30828 ( .A(n24139), .B(n22218), .Z(n30875) );
  XNOR U30829 ( .A(n30876), .B(n26654), .Z(n22218) );
  ANDN U30830 ( .B(n26655), .A(n30432), .Z(n30876) );
  XNOR U30831 ( .A(n30877), .B(n28294), .Z(n24139) );
  ANDN U30832 ( .B(n28295), .A(n30422), .Z(n30877) );
  XOR U30833 ( .A(n23816), .B(n30878), .Z(n30874) );
  XOR U30834 ( .A(n25130), .B(n23337), .Z(n30878) );
  XNOR U30835 ( .A(n30879), .B(n28064), .Z(n23337) );
  NOR U30836 ( .A(n30880), .B(n30425), .Z(n30879) );
  XNOR U30837 ( .A(n30881), .B(n26661), .Z(n25130) );
  ANDN U30838 ( .B(n26662), .A(n30435), .Z(n30881) );
  XOR U30839 ( .A(n30882), .B(n26651), .Z(n23816) );
  ANDN U30840 ( .B(n26650), .A(n30429), .Z(n30882) );
  IV U30841 ( .A(n30883), .Z(n30429) );
  XOR U30842 ( .A(n30884), .B(n30885), .Z(n27964) );
  XNOR U30843 ( .A(n26093), .B(n25780), .Z(n30885) );
  XOR U30844 ( .A(n30886), .B(n30887), .Z(n25780) );
  ANDN U30845 ( .B(n30888), .A(n30416), .Z(n30886) );
  XNOR U30846 ( .A(n30889), .B(n30890), .Z(n26093) );
  ANDN U30847 ( .B(n30891), .A(n29189), .Z(n30889) );
  XOR U30848 ( .A(n26644), .B(n30892), .Z(n30884) );
  XOR U30849 ( .A(n24622), .B(n26397), .Z(n30892) );
  XOR U30850 ( .A(n30893), .B(n29186), .Z(n26397) );
  NOR U30851 ( .A(n30894), .B(n29185), .Z(n30893) );
  XOR U30852 ( .A(n30895), .B(n29200), .Z(n24622) );
  NOR U30853 ( .A(n30409), .B(n29199), .Z(n30895) );
  XNOR U30854 ( .A(n30896), .B(n30897), .Z(n26644) );
  NOR U30855 ( .A(n30405), .B(n29195), .Z(n30896) );
  XOR U30856 ( .A(n28926), .B(n23059), .Z(n23202) );
  XNOR U30857 ( .A(n30594), .B(n29279), .Z(n23059) );
  XNOR U30858 ( .A(n30898), .B(n30899), .Z(n29279) );
  XNOR U30859 ( .A(n24485), .B(n29330), .Z(n30899) );
  XNOR U30860 ( .A(n30900), .B(n29336), .Z(n29330) );
  XNOR U30861 ( .A(n30901), .B(n28750), .Z(n28933) );
  IV U30862 ( .A(n29057), .Z(n28750) );
  XNOR U30863 ( .A(n30902), .B(n29347), .Z(n24485) );
  AND U30864 ( .A(n28928), .B(n28929), .Z(n30902) );
  XOR U30865 ( .A(n30903), .B(n30904), .Z(n28928) );
  XOR U30866 ( .A(n21236), .B(n30905), .Z(n30898) );
  XNOR U30867 ( .A(n26141), .B(n28772), .Z(n30905) );
  XOR U30868 ( .A(n30906), .B(n30907), .Z(n28772) );
  ANDN U30869 ( .B(n28941), .A(n28943), .Z(n30906) );
  XNOR U30870 ( .A(n30908), .B(n29343), .Z(n26141) );
  AND U30871 ( .A(n29344), .B(n30909), .Z(n30908) );
  XNOR U30872 ( .A(n30910), .B(n29340), .Z(n21236) );
  AND U30873 ( .A(n28937), .B(n28939), .Z(n30910) );
  XNOR U30874 ( .A(n30911), .B(n30912), .Z(n28937) );
  XOR U30875 ( .A(n30913), .B(n30914), .Z(n30594) );
  XNOR U30876 ( .A(n25267), .B(n25822), .Z(n30914) );
  XNOR U30877 ( .A(n30915), .B(n29356), .Z(n25822) );
  XNOR U30878 ( .A(n30916), .B(n28890), .Z(n29357) );
  XNOR U30879 ( .A(n30917), .B(n29362), .Z(n25267) );
  AND U30880 ( .A(n29648), .B(n29363), .Z(n30917) );
  XOR U30881 ( .A(n30918), .B(n30919), .Z(n29363) );
  XOR U30882 ( .A(n27309), .B(n30920), .Z(n30913) );
  XOR U30883 ( .A(n22653), .B(n23846), .Z(n30920) );
  XNOR U30884 ( .A(n30921), .B(n29366), .Z(n23846) );
  ANDN U30885 ( .B(n29367), .A(n30592), .Z(n30921) );
  XNOR U30886 ( .A(n30922), .B(n30923), .Z(n29367) );
  XNOR U30887 ( .A(n30924), .B(n30925), .Z(n22653) );
  AND U30888 ( .A(n29655), .B(n29653), .Z(n30924) );
  XNOR U30889 ( .A(n30926), .B(n29352), .Z(n27309) );
  ANDN U30890 ( .B(n29353), .A(n29651), .Z(n30926) );
  XOR U30891 ( .A(n30927), .B(n30928), .Z(n29353) );
  XOR U30892 ( .A(n30929), .B(n29344), .Z(n28926) );
  XNOR U30893 ( .A(n30930), .B(n30559), .Z(n29344) );
  NOR U30894 ( .A(n30931), .B(n30909), .Z(n30929) );
  XNOR U30895 ( .A(n30932), .B(n22231), .Z(n25647) );
  XOR U30896 ( .A(n30933), .B(n30934), .Z(n22231) );
  XNOR U30897 ( .A(n30935), .B(n23187), .Z(n20223) );
  XNOR U30898 ( .A(n30936), .B(n23584), .Z(n23187) );
  XNOR U30899 ( .A(n26986), .B(n26712), .Z(n23584) );
  XOR U30900 ( .A(n30937), .B(n30938), .Z(n26712) );
  XOR U30901 ( .A(n25194), .B(n24932), .Z(n30938) );
  XNOR U30902 ( .A(n30939), .B(n28444), .Z(n24932) );
  XOR U30903 ( .A(n30940), .B(n30941), .Z(n28444) );
  ANDN U30904 ( .B(n29498), .A(n28454), .Z(n30939) );
  XOR U30905 ( .A(n30942), .B(n30943), .Z(n28454) );
  XOR U30906 ( .A(n30944), .B(n26828), .Z(n25194) );
  XOR U30907 ( .A(n30945), .B(n30219), .Z(n26828) );
  NOR U30908 ( .A(n29500), .B(n26827), .Z(n30944) );
  XNOR U30909 ( .A(n30946), .B(n30947), .Z(n26827) );
  XOR U30910 ( .A(n22341), .B(n30948), .Z(n30937) );
  XOR U30911 ( .A(n23570), .B(n25725), .Z(n30948) );
  XNOR U30912 ( .A(n30949), .B(n28167), .Z(n25725) );
  XOR U30913 ( .A(n30950), .B(n29289), .Z(n28167) );
  NOR U30914 ( .A(n28166), .B(n29496), .Z(n30949) );
  XOR U30915 ( .A(n28995), .B(n30951), .Z(n28166) );
  XNOR U30916 ( .A(n30952), .B(n26834), .Z(n23570) );
  XNOR U30917 ( .A(n30953), .B(n30687), .Z(n26834) );
  ANDN U30918 ( .B(n26835), .A(n30954), .Z(n30952) );
  XNOR U30919 ( .A(n30955), .B(n30956), .Z(n26835) );
  XNOR U30920 ( .A(n30957), .B(n27334), .Z(n22341) );
  IV U30921 ( .A(n28452), .Z(n27334) );
  XOR U30922 ( .A(n30958), .B(n30959), .Z(n28452) );
  NOR U30923 ( .A(n30960), .B(n27333), .Z(n30957) );
  XOR U30924 ( .A(n30961), .B(n30962), .Z(n27333) );
  XOR U30925 ( .A(n30963), .B(n30964), .Z(n26986) );
  XNOR U30926 ( .A(n26402), .B(n24006), .Z(n30964) );
  ANDN U30927 ( .B(n30966), .A(n30967), .Z(n30965) );
  IV U30928 ( .A(n30968), .Z(n30967) );
  XNOR U30929 ( .A(n30969), .B(n29633), .Z(n26402) );
  XOR U30930 ( .A(n26820), .B(n30972), .Z(n30963) );
  XNOR U30931 ( .A(n24775), .B(n26036), .Z(n30972) );
  XNOR U30932 ( .A(n30973), .B(n30974), .Z(n26036) );
  ANDN U30933 ( .B(n30975), .A(n30976), .Z(n30973) );
  XNOR U30934 ( .A(n30977), .B(n30978), .Z(n24775) );
  ANDN U30935 ( .B(n30979), .A(n30980), .Z(n30977) );
  XNOR U30936 ( .A(n30981), .B(n29622), .Z(n26820) );
  AND U30937 ( .A(n30982), .B(n30983), .Z(n30981) );
  NOR U30938 ( .A(n22925), .B(n23186), .Z(n30935) );
  XNOR U30939 ( .A(n30984), .B(n25352), .Z(n23186) );
  XOR U30940 ( .A(n26629), .B(n30985), .Z(n25352) );
  XNOR U30941 ( .A(n30986), .B(n30987), .Z(n26629) );
  XOR U30942 ( .A(n27957), .B(n27386), .Z(n30987) );
  XNOR U30943 ( .A(n30988), .B(n28171), .Z(n27386) );
  XNOR U30944 ( .A(n30989), .B(n30990), .Z(n28171) );
  ANDN U30945 ( .B(n28170), .A(n30991), .Z(n30988) );
  XOR U30946 ( .A(n30992), .B(n28105), .Z(n27957) );
  XOR U30947 ( .A(n30781), .B(n30993), .Z(n28105) );
  XNOR U30948 ( .A(n24279), .B(n30995), .Z(n30986) );
  XNOR U30949 ( .A(n24604), .B(n27733), .Z(n30995) );
  XNOR U30950 ( .A(n30996), .B(n30997), .Z(n27733) );
  ANDN U30951 ( .B(n28102), .A(n30998), .Z(n30996) );
  XOR U30952 ( .A(n30999), .B(n28095), .Z(n24604) );
  XOR U30953 ( .A(n31000), .B(n31001), .Z(n28095) );
  ANDN U30954 ( .B(n28096), .A(n31002), .Z(n30999) );
  IV U30955 ( .A(n31003), .Z(n28096) );
  XNOR U30956 ( .A(n31004), .B(n28613), .Z(n24279) );
  XNOR U30957 ( .A(n31005), .B(n31006), .Z(n28613) );
  XNOR U30958 ( .A(n29358), .B(n25361), .Z(n22925) );
  XOR U30959 ( .A(n29972), .B(n31008), .Z(n25361) );
  XOR U30960 ( .A(n31009), .B(n31010), .Z(n29972) );
  XNOR U30961 ( .A(n25693), .B(n26770), .Z(n31010) );
  XNOR U30962 ( .A(n31011), .B(n30801), .Z(n26770) );
  AND U30963 ( .A(n27317), .B(n27319), .Z(n31011) );
  XOR U30964 ( .A(n30541), .B(n31012), .Z(n27319) );
  XNOR U30965 ( .A(n31013), .B(n27937), .Z(n27317) );
  XNOR U30966 ( .A(n31014), .B(n29382), .Z(n25693) );
  XNOR U30967 ( .A(n31015), .B(n29027), .Z(n27915) );
  XOR U30968 ( .A(n31016), .B(n30928), .Z(n27916) );
  XOR U30969 ( .A(n25310), .B(n31017), .Z(n31009) );
  XNOR U30970 ( .A(n26640), .B(n24034), .Z(n31017) );
  XOR U30971 ( .A(n31018), .B(n29379), .Z(n24034) );
  AND U30972 ( .A(n27323), .B(n27321), .Z(n31018) );
  XOR U30973 ( .A(n31019), .B(n31020), .Z(n27321) );
  XNOR U30974 ( .A(n31021), .B(n31022), .Z(n27323) );
  ANDN U30975 ( .B(n29975), .A(n31025), .Z(n31023) );
  IV U30976 ( .A(n29976), .Z(n31025) );
  XNOR U30977 ( .A(n31026), .B(n31027), .Z(n29976) );
  XNOR U30978 ( .A(n31028), .B(n29388), .Z(n25310) );
  AND U30979 ( .A(n27325), .B(n27326), .Z(n31028) );
  XNOR U30980 ( .A(n31029), .B(n31030), .Z(n27326) );
  XNOR U30981 ( .A(n29266), .B(n31031), .Z(n27325) );
  XNOR U30982 ( .A(n31032), .B(n31033), .Z(n29358) );
  NOR U30983 ( .A(n30925), .B(n29653), .Z(n31032) );
  XOR U30984 ( .A(n31034), .B(n31035), .Z(n29653) );
  XOR U30985 ( .A(n23182), .B(n31036), .Z(n30870) );
  XOR U30986 ( .A(n18747), .B(n16515), .Z(n31036) );
  XNOR U30987 ( .A(n31037), .B(n26261), .Z(n16515) );
  XOR U30988 ( .A(n30579), .B(n23031), .Z(n26261) );
  IV U30989 ( .A(n22534), .Z(n23031) );
  XNOR U30990 ( .A(n31038), .B(n31039), .Z(n29311) );
  XOR U30991 ( .A(n24001), .B(n22625), .Z(n31039) );
  XNOR U30992 ( .A(n31040), .B(n29593), .Z(n22625) );
  XOR U30993 ( .A(n31041), .B(n29401), .Z(n30588) );
  XNOR U30994 ( .A(n31042), .B(n28522), .Z(n24001) );
  IV U30995 ( .A(n31043), .Z(n28522) );
  ANDN U30996 ( .B(n29564), .A(n31044), .Z(n31042) );
  XOR U30997 ( .A(n31045), .B(n31046), .Z(n29564) );
  XOR U30998 ( .A(n25617), .B(n31047), .Z(n31038) );
  XOR U30999 ( .A(n24445), .B(n27575), .Z(n31047) );
  XNOR U31000 ( .A(n31048), .B(n28532), .Z(n27575) );
  ANDN U31001 ( .B(n30577), .A(n30576), .Z(n31048) );
  XOR U31002 ( .A(n31049), .B(n31050), .Z(n30577) );
  XNOR U31003 ( .A(n31051), .B(n28536), .Z(n24445) );
  IV U31004 ( .A(n31052), .Z(n28536) );
  ANDN U31005 ( .B(n29573), .A(n31053), .Z(n31051) );
  IV U31006 ( .A(n30572), .Z(n29573) );
  XNOR U31007 ( .A(n31054), .B(n31055), .Z(n30572) );
  XNOR U31008 ( .A(n31056), .B(n28526), .Z(n25617) );
  NOR U31009 ( .A(n29571), .B(n31057), .Z(n31056) );
  XOR U31010 ( .A(n31058), .B(n31059), .Z(n28061) );
  XOR U31011 ( .A(n29952), .B(n27795), .Z(n31059) );
  XOR U31012 ( .A(n31060), .B(n28260), .Z(n27795) );
  ANDN U31013 ( .B(n30549), .A(n29581), .Z(n31060) );
  XNOR U31014 ( .A(n31061), .B(n28890), .Z(n29581) );
  XOR U31015 ( .A(n31062), .B(n28256), .Z(n29952) );
  AND U31016 ( .A(n30561), .B(n29587), .Z(n31062) );
  XNOR U31017 ( .A(n30573), .B(n31063), .Z(n29587) );
  XNOR U31018 ( .A(n28323), .B(n31064), .Z(n31058) );
  XOR U31019 ( .A(n29692), .B(n31065), .Z(n31064) );
  XOR U31020 ( .A(n31066), .B(n28265), .Z(n29692) );
  AND U31021 ( .A(n29590), .B(n30552), .Z(n31066) );
  XNOR U31022 ( .A(n31067), .B(n31068), .Z(n29590) );
  XOR U31023 ( .A(n31069), .B(n28252), .Z(n28323) );
  AND U31024 ( .A(n29585), .B(n30565), .Z(n31069) );
  XOR U31025 ( .A(n31070), .B(n28992), .Z(n29585) );
  IV U31026 ( .A(n31071), .Z(n28992) );
  XOR U31027 ( .A(n31072), .B(n31057), .Z(n30579) );
  ANDN U31028 ( .B(n29571), .A(n28524), .Z(n31072) );
  XOR U31029 ( .A(n31073), .B(n30567), .Z(n28524) );
  XOR U31030 ( .A(n31074), .B(n28802), .Z(n29571) );
  ANDN U31031 ( .B(n23198), .A(n22921), .Z(n31037) );
  XOR U31032 ( .A(n30829), .B(n25276), .Z(n22921) );
  IV U31033 ( .A(n24438), .Z(n25276) );
  XNOR U31034 ( .A(n31075), .B(n26979), .Z(n24438) );
  XNOR U31035 ( .A(n31076), .B(n31077), .Z(n26979) );
  XNOR U31036 ( .A(n26754), .B(n23750), .Z(n31077) );
  XOR U31037 ( .A(n31078), .B(n31079), .Z(n23750) );
  NOR U31038 ( .A(n30842), .B(n30840), .Z(n31078) );
  XNOR U31039 ( .A(n31080), .B(n31081), .Z(n26754) );
  ANDN U31040 ( .B(n30831), .A(n30832), .Z(n31080) );
  XNOR U31041 ( .A(n26695), .B(n31082), .Z(n31076) );
  XNOR U31042 ( .A(n26027), .B(n26240), .Z(n31082) );
  XNOR U31043 ( .A(n31083), .B(n31084), .Z(n26240) );
  ANDN U31044 ( .B(n31085), .A(n31086), .Z(n31083) );
  XNOR U31045 ( .A(n31087), .B(n31088), .Z(n26027) );
  AND U31046 ( .A(n30836), .B(n30838), .Z(n31087) );
  XNOR U31047 ( .A(n31089), .B(n31090), .Z(n26695) );
  NOR U31048 ( .A(n30844), .B(n30845), .Z(n31089) );
  XOR U31049 ( .A(n31091), .B(n31085), .Z(n30829) );
  ANDN U31050 ( .B(n31086), .A(n31092), .Z(n31091) );
  IV U31051 ( .A(n25622), .Z(n23198) );
  XOR U31052 ( .A(n31093), .B(n25206), .Z(n25622) );
  XNOR U31053 ( .A(n30159), .B(n30479), .Z(n25206) );
  XNOR U31054 ( .A(n31094), .B(n31095), .Z(n30479) );
  XNOR U31055 ( .A(n23850), .B(n23506), .Z(n31095) );
  XNOR U31056 ( .A(n31096), .B(n27139), .Z(n23506) );
  XOR U31057 ( .A(n31097), .B(n30520), .Z(n27139) );
  ANDN U31058 ( .B(n28721), .A(n27138), .Z(n31096) );
  XOR U31059 ( .A(n31098), .B(n26363), .Z(n23850) );
  XOR U31060 ( .A(n31099), .B(n31100), .Z(n26363) );
  ANDN U31061 ( .B(n27132), .A(n31101), .Z(n31098) );
  XNOR U31062 ( .A(n24387), .B(n31102), .Z(n31094) );
  XOR U31063 ( .A(n26116), .B(n27105), .Z(n31102) );
  XNOR U31064 ( .A(n31103), .B(n26948), .Z(n27105) );
  XNOR U31065 ( .A(n29396), .B(n31104), .Z(n26948) );
  ANDN U31066 ( .B(n27129), .A(n27650), .Z(n31103) );
  XNOR U31067 ( .A(n31105), .B(n26366), .Z(n26116) );
  XNOR U31068 ( .A(n31106), .B(n31107), .Z(n26366) );
  ANDN U31069 ( .B(n27656), .A(n31108), .Z(n31105) );
  XNOR U31070 ( .A(n31110), .B(n30784), .Z(n26357) );
  ANDN U31071 ( .B(n27660), .A(n31111), .Z(n31109) );
  XNOR U31072 ( .A(n31112), .B(n31113), .Z(n30159) );
  XNOR U31073 ( .A(n23048), .B(n23827), .Z(n31113) );
  XOR U31074 ( .A(n31114), .B(n27122), .Z(n23827) );
  XOR U31075 ( .A(n31115), .B(n30697), .Z(n27122) );
  IV U31076 ( .A(n31116), .Z(n30697) );
  ANDN U31077 ( .B(n29531), .A(n27121), .Z(n31114) );
  XOR U31078 ( .A(n31117), .B(n27114), .Z(n23048) );
  XOR U31079 ( .A(n31118), .B(n31119), .Z(n27114) );
  AND U31080 ( .A(n29521), .B(n27115), .Z(n31117) );
  XOR U31081 ( .A(n23920), .B(n31120), .Z(n31112) );
  XOR U31082 ( .A(n26575), .B(n23627), .Z(n31120) );
  XOR U31083 ( .A(n31121), .B(n28130), .Z(n23627) );
  XOR U31084 ( .A(n31122), .B(n31123), .Z(n28130) );
  ANDN U31085 ( .B(n28131), .A(n29527), .Z(n31121) );
  IV U31086 ( .A(n31124), .Z(n29527) );
  XOR U31087 ( .A(n31125), .B(n28287), .Z(n26575) );
  XOR U31088 ( .A(n31126), .B(n31127), .Z(n28287) );
  XOR U31089 ( .A(n31128), .B(n27111), .Z(n23920) );
  XOR U31090 ( .A(n31129), .B(n29734), .Z(n27111) );
  ANDN U31091 ( .B(n29517), .A(n31130), .Z(n31128) );
  XNOR U31092 ( .A(n31131), .B(n23194), .Z(n18747) );
  XOR U31093 ( .A(n30678), .B(n25083), .Z(n23194) );
  XNOR U31094 ( .A(n27165), .B(n27057), .Z(n25083) );
  XNOR U31095 ( .A(n31132), .B(n31133), .Z(n27057) );
  XNOR U31096 ( .A(n26641), .B(n28478), .Z(n31133) );
  XOR U31097 ( .A(n31134), .B(n30621), .Z(n28478) );
  XNOR U31098 ( .A(n31135), .B(n28887), .Z(n29815) );
  XNOR U31099 ( .A(n31136), .B(n30623), .Z(n26641) );
  ANDN U31100 ( .B(n29811), .A(n30685), .Z(n31136) );
  XOR U31101 ( .A(n31137), .B(n31138), .Z(n29811) );
  XNOR U31102 ( .A(n23707), .B(n31139), .Z(n31132) );
  XNOR U31103 ( .A(n23761), .B(n24186), .Z(n31139) );
  XOR U31104 ( .A(n31140), .B(n30616), .Z(n24186) );
  XOR U31105 ( .A(n31141), .B(n31142), .Z(n29801) );
  XOR U31106 ( .A(n31143), .B(n30619), .Z(n23761) );
  AND U31107 ( .A(n29805), .B(n31144), .Z(n31143) );
  XOR U31108 ( .A(n31145), .B(n30613), .Z(n23707) );
  IV U31109 ( .A(n31146), .Z(n30613) );
  ANDN U31110 ( .B(n30694), .A(n30693), .Z(n31145) );
  XOR U31111 ( .A(n31147), .B(n31148), .Z(n30694) );
  XOR U31112 ( .A(n31149), .B(n31150), .Z(n27165) );
  XOR U31113 ( .A(n25788), .B(n26113), .Z(n31150) );
  XNOR U31114 ( .A(n31151), .B(n28362), .Z(n26113) );
  XNOR U31115 ( .A(n31152), .B(n30559), .Z(n28362) );
  XOR U31116 ( .A(n31153), .B(n31154), .Z(n29177) );
  XOR U31117 ( .A(n31155), .B(n27939), .Z(n28487) );
  XOR U31118 ( .A(n31156), .B(n28223), .Z(n25788) );
  XNOR U31119 ( .A(n31157), .B(n29053), .Z(n28223) );
  AND U31120 ( .A(n28494), .B(n29160), .Z(n31156) );
  XOR U31121 ( .A(n31158), .B(n31159), .Z(n29160) );
  XOR U31122 ( .A(n29324), .B(n31160), .Z(n28494) );
  XNOR U31123 ( .A(n28134), .B(n31161), .Z(n31149) );
  XNOR U31124 ( .A(n23724), .B(n26278), .Z(n31161) );
  XNOR U31125 ( .A(n31162), .B(n28233), .Z(n26278) );
  XOR U31126 ( .A(n31163), .B(n31164), .Z(n28233) );
  ANDN U31127 ( .B(n29164), .A(n28490), .Z(n31162) );
  IV U31128 ( .A(n30673), .Z(n28490) );
  XOR U31129 ( .A(n31165), .B(n28887), .Z(n30673) );
  XOR U31130 ( .A(n31166), .B(n28885), .Z(n29164) );
  XOR U31131 ( .A(n31167), .B(n28226), .Z(n23724) );
  XOR U31132 ( .A(n31168), .B(n31169), .Z(n28226) );
  XOR U31133 ( .A(n30248), .B(n31170), .Z(n28492) );
  IV U31134 ( .A(n29169), .Z(n30667) );
  XNOR U31135 ( .A(n30306), .B(n31171), .Z(n29169) );
  XOR U31136 ( .A(n31172), .B(n28484), .Z(n28134) );
  XNOR U31137 ( .A(n31173), .B(n30682), .Z(n28484) );
  IV U31138 ( .A(n29946), .Z(n30682) );
  AND U31139 ( .A(n28485), .B(n29173), .Z(n31172) );
  XOR U31140 ( .A(n31174), .B(n30990), .Z(n29173) );
  XOR U31141 ( .A(n31175), .B(n30125), .Z(n28485) );
  XOR U31142 ( .A(n31176), .B(n31144), .Z(n30678) );
  NOR U31143 ( .A(n29805), .B(n29806), .Z(n31176) );
  XOR U31144 ( .A(n31179), .B(n31159), .Z(n29805) );
  ANDN U31145 ( .B(n23195), .A(n22916), .Z(n31131) );
  XOR U31146 ( .A(n30361), .B(n21372), .Z(n22916) );
  XOR U31147 ( .A(n29780), .B(n26772), .Z(n21372) );
  XNOR U31148 ( .A(n31180), .B(n31181), .Z(n26772) );
  XNOR U31149 ( .A(n31182), .B(n25054), .Z(n31181) );
  XNOR U31150 ( .A(n31183), .B(n27695), .Z(n25054) );
  ANDN U31151 ( .B(n30368), .A(n28122), .Z(n31183) );
  IV U31152 ( .A(n30369), .Z(n28122) );
  XOR U31153 ( .A(n31184), .B(n31185), .Z(n30369) );
  XOR U31154 ( .A(n25004), .B(n31186), .Z(n31180) );
  XOR U31155 ( .A(n24699), .B(n24907), .Z(n31186) );
  XNOR U31156 ( .A(n31187), .B(n28127), .Z(n24907) );
  ANDN U31157 ( .B(n28118), .A(n31188), .Z(n31187) );
  XNOR U31158 ( .A(n31189), .B(n27684), .Z(n24699) );
  ANDN U31159 ( .B(n28114), .A(n30373), .Z(n31189) );
  XOR U31160 ( .A(n31190), .B(n31191), .Z(n28114) );
  XNOR U31161 ( .A(n31192), .B(n27699), .Z(n25004) );
  ANDN U31162 ( .B(n30363), .A(n28125), .Z(n31192) );
  XOR U31163 ( .A(n31193), .B(n30748), .Z(n28125) );
  XOR U31164 ( .A(n31194), .B(n31195), .Z(n29780) );
  XOR U31165 ( .A(n30021), .B(n26233), .Z(n31195) );
  XNOR U31166 ( .A(n31196), .B(n31197), .Z(n26233) );
  ANDN U31167 ( .B(n30352), .A(n30353), .Z(n31196) );
  ANDN U31168 ( .B(n30339), .A(n30340), .Z(n31198) );
  XNOR U31169 ( .A(n26783), .B(n31200), .Z(n31194) );
  XOR U31170 ( .A(n23345), .B(n31201), .Z(n31200) );
  XNOR U31171 ( .A(n31202), .B(n31203), .Z(n23345) );
  AND U31172 ( .A(n30343), .B(n30344), .Z(n31202) );
  XOR U31173 ( .A(n31204), .B(n31205), .Z(n26783) );
  AND U31174 ( .A(n30349), .B(n30348), .Z(n31204) );
  XOR U31175 ( .A(n31206), .B(n31188), .Z(n30361) );
  NOR U31176 ( .A(n28120), .B(n28118), .Z(n31206) );
  XNOR U31177 ( .A(n31207), .B(n29050), .Z(n28118) );
  XOR U31178 ( .A(n31208), .B(n30790), .Z(n28120) );
  XOR U31179 ( .A(n29320), .B(n23442), .Z(n23195) );
  XOR U31180 ( .A(n31209), .B(n31210), .Z(n28870) );
  XOR U31181 ( .A(n27726), .B(n23940), .Z(n31210) );
  XNOR U31182 ( .A(n31211), .B(n29029), .Z(n23940) );
  AND U31183 ( .A(n27469), .B(n29033), .Z(n31211) );
  XNOR U31184 ( .A(n28982), .B(n31213), .Z(n29033) );
  XOR U31185 ( .A(n31214), .B(n29289), .Z(n27469) );
  XNOR U31186 ( .A(n31215), .B(n28507), .Z(n27726) );
  XNOR U31187 ( .A(n31216), .B(n29409), .Z(n28507) );
  ANDN U31188 ( .B(n28508), .A(n27478), .Z(n31215) );
  XOR U31189 ( .A(n29930), .B(n31217), .Z(n27478) );
  XOR U31190 ( .A(n31218), .B(n31219), .Z(n28508) );
  XNOR U31191 ( .A(n28499), .B(n31220), .Z(n31209) );
  XOR U31192 ( .A(n24514), .B(n25891), .Z(n31220) );
  XOR U31193 ( .A(n31221), .B(n28504), .Z(n25891) );
  XOR U31194 ( .A(n31222), .B(n31223), .Z(n28504) );
  ANDN U31195 ( .B(n28505), .A(n29327), .Z(n31221) );
  XNOR U31196 ( .A(n31224), .B(n28512), .Z(n24514) );
  XNOR U31197 ( .A(n31225), .B(n31226), .Z(n28512) );
  ANDN U31198 ( .B(n28513), .A(n27482), .Z(n31224) );
  XNOR U31199 ( .A(n30231), .B(n31227), .Z(n27482) );
  XOR U31200 ( .A(n31228), .B(n31229), .Z(n28513) );
  XOR U31201 ( .A(n31230), .B(n28515), .Z(n28499) );
  XOR U31202 ( .A(n31231), .B(n31127), .Z(n28515) );
  ANDN U31203 ( .B(n28516), .A(n27474), .Z(n31230) );
  XOR U31204 ( .A(n31232), .B(n31233), .Z(n27474) );
  XOR U31205 ( .A(n31234), .B(n29741), .Z(n28516) );
  XOR U31206 ( .A(n31235), .B(n31236), .Z(n27577) );
  XNOR U31207 ( .A(n23688), .B(n25966), .Z(n31236) );
  XOR U31208 ( .A(n31237), .B(n29569), .Z(n25966) );
  XOR U31209 ( .A(n31238), .B(n31239), .Z(n29569) );
  ANDN U31210 ( .B(n29593), .A(n30585), .Z(n31237) );
  XOR U31211 ( .A(n31240), .B(n31241), .Z(n30585) );
  XOR U31212 ( .A(n31242), .B(n31142), .Z(n29593) );
  XNOR U31213 ( .A(n31243), .B(n28521), .Z(n23688) );
  XOR U31214 ( .A(n28765), .B(n31244), .Z(n28521) );
  ANDN U31215 ( .B(n31044), .A(n31043), .Z(n31243) );
  XNOR U31216 ( .A(n31245), .B(n31127), .Z(n31043) );
  IV U31217 ( .A(n30581), .Z(n31044) );
  XOR U31218 ( .A(n29064), .B(n31246), .Z(n30581) );
  XNOR U31219 ( .A(n24426), .B(n31247), .Z(n31235) );
  XNOR U31220 ( .A(n25714), .B(n23596), .Z(n31247) );
  XNOR U31221 ( .A(n31248), .B(n28525), .Z(n23596) );
  XOR U31222 ( .A(n31249), .B(n31250), .Z(n28525) );
  ANDN U31223 ( .B(n31057), .A(n28526), .Z(n31248) );
  XNOR U31224 ( .A(n31251), .B(n30230), .Z(n28526) );
  XOR U31225 ( .A(n31252), .B(n31253), .Z(n31057) );
  XNOR U31226 ( .A(n31254), .B(n28535), .Z(n25714) );
  XNOR U31227 ( .A(n31255), .B(n31256), .Z(n28535) );
  ANDN U31228 ( .B(n31053), .A(n31052), .Z(n31254) );
  XOR U31229 ( .A(n31257), .B(n31258), .Z(n31052) );
  IV U31230 ( .A(n30571), .Z(n31053) );
  XOR U31231 ( .A(n30264), .B(n31259), .Z(n30571) );
  XNOR U31232 ( .A(n31260), .B(n28531), .Z(n24426) );
  XOR U31233 ( .A(n31262), .B(n30956), .Z(n28532) );
  XOR U31234 ( .A(n31263), .B(n31264), .Z(n30576) );
  XNOR U31235 ( .A(n31265), .B(n28505), .Z(n29320) );
  XOR U31236 ( .A(n31266), .B(n30258), .Z(n28505) );
  XOR U31237 ( .A(n31267), .B(n31268), .Z(n29017) );
  XNOR U31238 ( .A(n30211), .B(n31269), .Z(n29327) );
  XNOR U31239 ( .A(n31270), .B(n23191), .Z(n23182) );
  XOR U31240 ( .A(n23788), .B(n28979), .Z(n23191) );
  XNOR U31241 ( .A(n31271), .B(n31272), .Z(n28979) );
  NOR U31242 ( .A(n27380), .B(n27381), .Z(n31271) );
  XNOR U31243 ( .A(n30860), .B(n31273), .Z(n27381) );
  IV U31244 ( .A(n31274), .Z(n27380) );
  IV U31245 ( .A(n24375), .Z(n23788) );
  XNOR U31246 ( .A(n30806), .B(n25751), .Z(n24375) );
  XOR U31247 ( .A(n31275), .B(n31276), .Z(n25751) );
  XOR U31248 ( .A(n26555), .B(n24909), .Z(n31276) );
  XNOR U31249 ( .A(n31277), .B(n28213), .Z(n24909) );
  ANDN U31250 ( .B(n27589), .A(n27590), .Z(n31277) );
  XOR U31251 ( .A(n31278), .B(n28202), .Z(n26555) );
  ANDN U31252 ( .B(n27595), .A(n31279), .Z(n31278) );
  XNOR U31253 ( .A(n21818), .B(n31280), .Z(n31275) );
  XOR U31254 ( .A(n29953), .B(n25176), .Z(n31280) );
  XNOR U31255 ( .A(n31281), .B(n28210), .Z(n25176) );
  ANDN U31256 ( .B(n27598), .A(n27600), .Z(n31281) );
  NOR U31257 ( .A(n27602), .B(n27603), .Z(n31282) );
  XNOR U31258 ( .A(n31283), .B(n31284), .Z(n21818) );
  ANDN U31259 ( .B(n27606), .A(n27607), .Z(n31283) );
  XNOR U31260 ( .A(n31285), .B(n31286), .Z(n30806) );
  XOR U31261 ( .A(n27227), .B(n25957), .Z(n31286) );
  XNOR U31262 ( .A(n31287), .B(n28046), .Z(n25957) );
  ANDN U31263 ( .B(n28994), .A(n27370), .Z(n31287) );
  XNOR U31264 ( .A(n31288), .B(n31289), .Z(n27370) );
  XNOR U31265 ( .A(n31290), .B(n28055), .Z(n27227) );
  ANDN U31266 ( .B(n31272), .A(n31274), .Z(n31290) );
  XOR U31267 ( .A(n31291), .B(n31142), .Z(n31274) );
  IV U31268 ( .A(n30531), .Z(n31142) );
  XNOR U31269 ( .A(n29035), .B(n31292), .Z(n31285) );
  XNOR U31270 ( .A(n28719), .B(n31293), .Z(n31292) );
  XNOR U31271 ( .A(n31294), .B(n28043), .Z(n28719) );
  ANDN U31272 ( .B(n28981), .A(n27366), .Z(n31294) );
  XOR U31273 ( .A(n31295), .B(n31296), .Z(n27366) );
  XNOR U31274 ( .A(n31297), .B(n28049), .Z(n29035) );
  ANDN U31275 ( .B(n28986), .A(n27376), .Z(n31297) );
  XOR U31276 ( .A(n31298), .B(n31299), .Z(n27376) );
  NOR U31277 ( .A(n23190), .B(n22929), .Z(n31270) );
  XNOR U31278 ( .A(n31201), .B(n23346), .Z(n22929) );
  IV U31279 ( .A(n26784), .Z(n23346) );
  XNOR U31280 ( .A(n26468), .B(n31300), .Z(n26784) );
  XOR U31281 ( .A(n31301), .B(n31302), .Z(n26468) );
  XNOR U31282 ( .A(n27173), .B(n28650), .Z(n31302) );
  XNOR U31283 ( .A(n31303), .B(n31304), .Z(n28650) );
  AND U31284 ( .A(n29795), .B(n28074), .Z(n31303) );
  XOR U31285 ( .A(n31305), .B(n29071), .Z(n28074) );
  XOR U31286 ( .A(n31306), .B(n31307), .Z(n27173) );
  ANDN U31287 ( .B(n29789), .A(n28070), .Z(n31306) );
  IV U31288 ( .A(n29790), .Z(n28070) );
  XOR U31289 ( .A(n30657), .B(n31308), .Z(n29790) );
  XOR U31290 ( .A(n27638), .B(n31309), .Z(n31301) );
  XNOR U31291 ( .A(n25415), .B(n26138), .Z(n31309) );
  XOR U31292 ( .A(n31310), .B(n31311), .Z(n26138) );
  ANDN U31293 ( .B(n28087), .A(n31312), .Z(n31310) );
  XOR U31294 ( .A(n31313), .B(n31314), .Z(n28087) );
  XNOR U31295 ( .A(n31315), .B(n31316), .Z(n25415) );
  AND U31296 ( .A(n28079), .B(n29792), .Z(n31315) );
  XNOR U31297 ( .A(n31317), .B(n30514), .Z(n28079) );
  XNOR U31298 ( .A(n31318), .B(n31319), .Z(n27638) );
  ANDN U31299 ( .B(n28083), .A(n31320), .Z(n31318) );
  XNOR U31300 ( .A(n31321), .B(n31322), .Z(n28083) );
  XOR U31301 ( .A(n31323), .B(n31324), .Z(n31201) );
  AND U31302 ( .A(n30356), .B(n30357), .Z(n31323) );
  XOR U31303 ( .A(n30315), .B(n23136), .Z(n23190) );
  XOR U31304 ( .A(n26816), .B(n29277), .Z(n23136) );
  XNOR U31305 ( .A(n31325), .B(n31326), .Z(n29277) );
  XOR U31306 ( .A(n22314), .B(n25325), .Z(n31326) );
  XNOR U31307 ( .A(n31327), .B(n30156), .Z(n25325) );
  ANDN U31308 ( .B(n30155), .A(n26970), .Z(n31327) );
  IV U31309 ( .A(n30313), .Z(n26970) );
  XOR U31310 ( .A(n31328), .B(n29299), .Z(n30313) );
  XNOR U31311 ( .A(n31330), .B(n27049), .Z(n22314) );
  IV U31312 ( .A(n31331), .Z(n27049) );
  NOR U31313 ( .A(n27048), .B(n26966), .Z(n31330) );
  XNOR U31314 ( .A(n31332), .B(n31333), .Z(n26966) );
  XOR U31315 ( .A(n31334), .B(n29717), .Z(n27048) );
  XOR U31316 ( .A(n22338), .B(n31335), .Z(n31325) );
  XOR U31317 ( .A(n24614), .B(n25979), .Z(n31335) );
  XNOR U31318 ( .A(n31336), .B(n27041), .Z(n25979) );
  XOR U31319 ( .A(n31337), .B(n31338), .Z(n26957) );
  XOR U31320 ( .A(n31339), .B(n31340), .Z(n27040) );
  XNOR U31321 ( .A(n31341), .B(n31342), .Z(n24614) );
  NOR U31322 ( .A(n31343), .B(n28973), .Z(n31341) );
  XNOR U31323 ( .A(n31344), .B(n27046), .Z(n22338) );
  ANDN U31324 ( .B(n26962), .A(n30311), .Z(n31344) );
  XOR U31325 ( .A(n31345), .B(n31346), .Z(n30311) );
  XOR U31326 ( .A(n31347), .B(n31348), .Z(n26962) );
  XNOR U31327 ( .A(n31349), .B(n31350), .Z(n26816) );
  XNOR U31328 ( .A(n26529), .B(n22953), .Z(n31350) );
  XNOR U31329 ( .A(n31351), .B(n28174), .Z(n22953) );
  IV U31330 ( .A(n31352), .Z(n28174) );
  AND U31331 ( .A(n27557), .B(n28175), .Z(n31351) );
  XNOR U31332 ( .A(n31353), .B(n30078), .Z(n28175) );
  XOR U31333 ( .A(n31354), .B(n29307), .Z(n27557) );
  IV U31334 ( .A(n31355), .Z(n29307) );
  XNOR U31335 ( .A(n31356), .B(n31357), .Z(n26529) );
  ANDN U31336 ( .B(n28965), .A(n27545), .Z(n31356) );
  XNOR U31337 ( .A(n31358), .B(n29922), .Z(n27545) );
  XOR U31338 ( .A(n31359), .B(n31360), .Z(n28965) );
  XNOR U31339 ( .A(n24954), .B(n31361), .Z(n31349) );
  XOR U31340 ( .A(n22499), .B(n23608), .Z(n31361) );
  XNOR U31341 ( .A(n31362), .B(n26623), .Z(n23608) );
  NOR U31342 ( .A(n28968), .B(n27554), .Z(n31362) );
  XOR U31343 ( .A(n31363), .B(n30507), .Z(n27554) );
  XOR U31344 ( .A(n31364), .B(n31365), .Z(n28968) );
  XNOR U31345 ( .A(n31366), .B(n26994), .Z(n22499) );
  ANDN U31346 ( .B(n26995), .A(n27542), .Z(n31366) );
  XNOR U31347 ( .A(n31367), .B(n31264), .Z(n27542) );
  XOR U31348 ( .A(n31368), .B(n31369), .Z(n26995) );
  XOR U31349 ( .A(n31370), .B(n31371), .Z(n24954) );
  ANDN U31350 ( .B(n28970), .A(n27550), .Z(n31370) );
  XNOR U31351 ( .A(n31372), .B(n30928), .Z(n27550) );
  XOR U31352 ( .A(n31373), .B(n31374), .Z(n30315) );
  ANDN U31353 ( .B(n28973), .A(n28974), .Z(n31373) );
  XNOR U31354 ( .A(n31375), .B(n31376), .Z(n28973) );
  ANDN U31355 ( .B(n13492), .A(n16741), .Z(n30605) );
  XOR U31356 ( .A(n16957), .B(n21109), .Z(n16741) );
  XNOR U31357 ( .A(n31377), .B(n19627), .Z(n21109) );
  NOR U31358 ( .A(n21465), .B(n27903), .Z(n31377) );
  XOR U31359 ( .A(n23957), .B(n29666), .Z(n21465) );
  XNOR U31360 ( .A(n31378), .B(n29612), .Z(n29666) );
  NOR U31361 ( .A(n31379), .B(n31380), .Z(n31378) );
  IV U31362 ( .A(n24257), .Z(n23957) );
  XOR U31363 ( .A(n26821), .B(n26792), .Z(n24257) );
  XNOR U31364 ( .A(n31381), .B(n31382), .Z(n26792) );
  XNOR U31365 ( .A(n25809), .B(n24948), .Z(n31382) );
  XNOR U31366 ( .A(n31383), .B(n29609), .Z(n24948) );
  NOR U31367 ( .A(n29661), .B(n29608), .Z(n31383) );
  XNOR U31368 ( .A(n31384), .B(n29946), .Z(n29608) );
  XNOR U31369 ( .A(n31385), .B(n29600), .Z(n25809) );
  ANDN U31370 ( .B(n29599), .A(n31386), .Z(n31385) );
  IV U31371 ( .A(n29669), .Z(n29599) );
  XNOR U31372 ( .A(n30000), .B(n31387), .Z(n29669) );
  XOR U31373 ( .A(n29594), .B(n31388), .Z(n31381) );
  XOR U31374 ( .A(n25516), .B(n26126), .Z(n31388) );
  XNOR U31375 ( .A(n31389), .B(n29617), .Z(n26126) );
  NOR U31376 ( .A(n29616), .B(n29673), .Z(n31389) );
  XOR U31377 ( .A(n29097), .B(n31390), .Z(n29616) );
  XNOR U31378 ( .A(n31391), .B(n29603), .Z(n25516) );
  ANDN U31379 ( .B(n29604), .A(n29664), .Z(n31391) );
  XOR U31380 ( .A(n31392), .B(n30798), .Z(n29604) );
  XOR U31381 ( .A(n31393), .B(n29613), .Z(n29594) );
  ANDN U31382 ( .B(n31380), .A(n29612), .Z(n31393) );
  XOR U31383 ( .A(n31394), .B(n31395), .Z(n29612) );
  XOR U31384 ( .A(n31396), .B(n31397), .Z(n26821) );
  XOR U31385 ( .A(n23820), .B(n22796), .Z(n31397) );
  XOR U31386 ( .A(n31398), .B(n31399), .Z(n22796) );
  ANDN U31387 ( .B(n30978), .A(n31400), .Z(n31398) );
  XNOR U31388 ( .A(n31401), .B(n29632), .Z(n23820) );
  ANDN U31389 ( .B(n29633), .A(n30971), .Z(n31401) );
  XOR U31390 ( .A(n31402), .B(n30217), .Z(n29633) );
  XOR U31391 ( .A(n27099), .B(n31403), .Z(n31396) );
  XOR U31392 ( .A(n21218), .B(n24435), .Z(n31403) );
  XNOR U31393 ( .A(n31404), .B(n29626), .Z(n24435) );
  ANDN U31394 ( .B(n29627), .A(n30968), .Z(n31404) );
  XNOR U31395 ( .A(n31405), .B(n31406), .Z(n29627) );
  XNOR U31396 ( .A(n31407), .B(n29636), .Z(n21218) );
  NOR U31397 ( .A(n30974), .B(n30975), .Z(n31407) );
  IV U31398 ( .A(n29637), .Z(n30974) );
  XNOR U31399 ( .A(n31408), .B(n29396), .Z(n29637) );
  XNOR U31400 ( .A(n31409), .B(n31410), .Z(n27099) );
  NOR U31401 ( .A(n29622), .B(n30983), .Z(n31409) );
  XOR U31402 ( .A(n31411), .B(n31412), .Z(n29622) );
  XNOR U31403 ( .A(n19828), .B(n21895), .Z(n16957) );
  XNOR U31404 ( .A(n31413), .B(n31414), .Z(n21895) );
  XNOR U31405 ( .A(n18382), .B(n18636), .Z(n31414) );
  XOR U31406 ( .A(n31415), .B(n20023), .Z(n18636) );
  XOR U31407 ( .A(n30394), .B(n25189), .Z(n20023) );
  IV U31408 ( .A(n21728), .Z(n25189) );
  XNOR U31409 ( .A(n27201), .B(n30177), .Z(n21728) );
  XOR U31410 ( .A(n31416), .B(n31417), .Z(n30177) );
  XNOR U31411 ( .A(n25369), .B(n26080), .Z(n31417) );
  XNOR U31412 ( .A(n31418), .B(n27869), .Z(n26080) );
  ANDN U31413 ( .B(n27766), .A(n31419), .Z(n31418) );
  XNOR U31414 ( .A(n31420), .B(n27856), .Z(n25369) );
  ANDN U31415 ( .B(n30191), .A(n30192), .Z(n31420) );
  XNOR U31416 ( .A(n24922), .B(n31421), .Z(n31416) );
  XNOR U31417 ( .A(n25599), .B(n23146), .Z(n31421) );
  XNOR U31418 ( .A(n31422), .B(n27861), .Z(n23146) );
  ANDN U31419 ( .B(n27774), .A(n27775), .Z(n31422) );
  XOR U31420 ( .A(n31423), .B(n31424), .Z(n25599) );
  ANDN U31421 ( .B(n27762), .A(n27761), .Z(n31423) );
  XNOR U31422 ( .A(n31425), .B(n27866), .Z(n24922) );
  ANDN U31423 ( .B(n27770), .A(n27771), .Z(n31425) );
  XOR U31424 ( .A(n31426), .B(n31427), .Z(n27201) );
  XOR U31425 ( .A(n24805), .B(n25332), .Z(n31427) );
  XNOR U31426 ( .A(n31428), .B(n31429), .Z(n25332) );
  ANDN U31427 ( .B(n29469), .A(n31430), .Z(n31428) );
  XOR U31428 ( .A(n31431), .B(n31432), .Z(n24805) );
  XNOR U31429 ( .A(n31433), .B(n31434), .Z(n29478) );
  XOR U31430 ( .A(n25048), .B(n31435), .Z(n31426) );
  XOR U31431 ( .A(n31436), .B(n23593), .Z(n31435) );
  XNOR U31432 ( .A(n31437), .B(n31438), .Z(n23593) );
  ANDN U31433 ( .B(n29465), .A(n30390), .Z(n31437) );
  XOR U31434 ( .A(n31439), .B(n31440), .Z(n29465) );
  XNOR U31435 ( .A(n31441), .B(n31442), .Z(n25048) );
  ANDN U31436 ( .B(n30396), .A(n29474), .Z(n31441) );
  XOR U31437 ( .A(n31443), .B(n31444), .Z(n29474) );
  XNOR U31438 ( .A(n31445), .B(n31446), .Z(n30394) );
  NOR U31439 ( .A(n29471), .B(n29469), .Z(n31445) );
  XNOR U31440 ( .A(n31447), .B(n31448), .Z(n29469) );
  ANDN U31441 ( .B(n21112), .A(n20024), .Z(n31415) );
  XOR U31442 ( .A(n29191), .B(n21829), .Z(n20024) );
  XNOR U31443 ( .A(n31449), .B(n28290), .Z(n21829) );
  XNOR U31444 ( .A(n31450), .B(n31451), .Z(n28290) );
  XNOR U31445 ( .A(n26471), .B(n26344), .Z(n31451) );
  XNOR U31446 ( .A(n31452), .B(n30436), .Z(n26344) );
  NOR U31447 ( .A(n26661), .B(n26660), .Z(n31452) );
  XNOR U31448 ( .A(n31453), .B(n31454), .Z(n26660) );
  XOR U31449 ( .A(n31455), .B(n31456), .Z(n26661) );
  XNOR U31450 ( .A(n31457), .B(n31458), .Z(n26471) );
  NOR U31451 ( .A(n28064), .B(n28063), .Z(n31457) );
  XOR U31452 ( .A(n31459), .B(n31460), .Z(n28063) );
  XOR U31453 ( .A(n31461), .B(n29941), .Z(n28064) );
  XOR U31454 ( .A(n25220), .B(n31462), .Z(n31450) );
  XOR U31455 ( .A(n25975), .B(n27437), .Z(n31462) );
  XNOR U31456 ( .A(n31463), .B(n31464), .Z(n27437) );
  NOR U31457 ( .A(n28294), .B(n28293), .Z(n31463) );
  XNOR U31458 ( .A(n31240), .B(n31465), .Z(n28293) );
  XNOR U31459 ( .A(n31466), .B(n31467), .Z(n28294) );
  XNOR U31460 ( .A(n31468), .B(n31469), .Z(n25975) );
  NOR U31461 ( .A(n26654), .B(n26653), .Z(n31468) );
  XNOR U31462 ( .A(n31470), .B(n31471), .Z(n26653) );
  XNOR U31463 ( .A(n31472), .B(n29055), .Z(n26654) );
  XNOR U31464 ( .A(n31473), .B(n30430), .Z(n25220) );
  ANDN U31465 ( .B(n26651), .A(n26649), .Z(n31473) );
  XOR U31466 ( .A(n31474), .B(n30746), .Z(n26649) );
  XOR U31467 ( .A(n31475), .B(n28897), .Z(n26651) );
  XNOR U31468 ( .A(n31476), .B(n30418), .Z(n29191) );
  NOR U31469 ( .A(n31477), .B(n30888), .Z(n31476) );
  XOR U31470 ( .A(n31478), .B(n25255), .Z(n21112) );
  IV U31471 ( .A(n25350), .Z(n25255) );
  XNOR U31472 ( .A(n28542), .B(n26755), .Z(n25350) );
  XOR U31473 ( .A(n31479), .B(n31480), .Z(n26755) );
  XNOR U31474 ( .A(n23730), .B(n30723), .Z(n31480) );
  XNOR U31475 ( .A(n31481), .B(n31482), .Z(n30723) );
  XOR U31476 ( .A(n31484), .B(n31485), .Z(n23730) );
  NOR U31477 ( .A(n31486), .B(n31487), .Z(n31484) );
  XOR U31478 ( .A(n25297), .B(n31488), .Z(n31479) );
  XNOR U31479 ( .A(n22792), .B(n27721), .Z(n31488) );
  XNOR U31480 ( .A(n31489), .B(n31490), .Z(n27721) );
  XNOR U31481 ( .A(n31492), .B(n31493), .Z(n22792) );
  ANDN U31482 ( .B(n27995), .A(n31494), .Z(n31492) );
  XNOR U31483 ( .A(n31495), .B(n31496), .Z(n25297) );
  ANDN U31484 ( .B(n31497), .A(n31498), .Z(n31495) );
  XOR U31485 ( .A(n31499), .B(n31500), .Z(n28542) );
  XNOR U31486 ( .A(n25451), .B(n26393), .Z(n31500) );
  XOR U31487 ( .A(n31501), .B(n31502), .Z(n26393) );
  NOR U31488 ( .A(n31503), .B(n30445), .Z(n31501) );
  XNOR U31489 ( .A(n31504), .B(n31505), .Z(n25451) );
  ANDN U31490 ( .B(n31506), .A(n30451), .Z(n31504) );
  XOR U31491 ( .A(n25223), .B(n31507), .Z(n31499) );
  XOR U31492 ( .A(n25108), .B(n31508), .Z(n31507) );
  XNOR U31493 ( .A(n31509), .B(n31510), .Z(n25108) );
  NOR U31494 ( .A(n30455), .B(n31511), .Z(n31509) );
  IV U31495 ( .A(n31512), .Z(n30455) );
  XNOR U31496 ( .A(n31513), .B(n31514), .Z(n25223) );
  ANDN U31497 ( .B(n30637), .A(n31515), .Z(n31513) );
  XNOR U31498 ( .A(n31516), .B(n19621), .Z(n18382) );
  XOR U31499 ( .A(n26805), .B(n24998), .Z(n19621) );
  XOR U31500 ( .A(n31517), .B(n31518), .Z(n26805) );
  ANDN U31501 ( .B(n31519), .A(n31520), .Z(n31517) );
  XOR U31502 ( .A(n31182), .B(n24908), .Z(n21102) );
  XOR U31503 ( .A(n31521), .B(n31300), .Z(n24908) );
  XNOR U31504 ( .A(n31522), .B(n31523), .Z(n31300) );
  XNOR U31505 ( .A(n30718), .B(n25491), .Z(n31523) );
  XOR U31506 ( .A(n31524), .B(n31525), .Z(n25491) );
  XOR U31507 ( .A(n30148), .B(n31526), .Z(n30348) );
  XNOR U31508 ( .A(n31527), .B(n31528), .Z(n30718) );
  ANDN U31509 ( .B(n31324), .A(n30356), .Z(n31527) );
  XOR U31510 ( .A(n31529), .B(n30764), .Z(n30356) );
  XOR U31511 ( .A(n28357), .B(n31530), .Z(n31522) );
  XOR U31512 ( .A(n24251), .B(n31531), .Z(n31530) );
  XNOR U31513 ( .A(n31532), .B(n31533), .Z(n24251) );
  ANDN U31514 ( .B(n31199), .A(n30339), .Z(n31532) );
  XOR U31515 ( .A(n31534), .B(n31535), .Z(n30339) );
  XNOR U31516 ( .A(n31536), .B(n31537), .Z(n28357) );
  NOR U31517 ( .A(n30343), .B(n31203), .Z(n31536) );
  XOR U31518 ( .A(n31538), .B(n31539), .Z(n30343) );
  ANDN U31519 ( .B(n30377), .A(n30378), .Z(n31540) );
  XNOR U31520 ( .A(n31541), .B(n31542), .Z(n30378) );
  XOR U31521 ( .A(n31065), .B(n27796), .Z(n19620) );
  XNOR U31522 ( .A(n27576), .B(n26220), .Z(n27796) );
  XOR U31523 ( .A(n31543), .B(n31544), .Z(n26220) );
  XNOR U31524 ( .A(n26523), .B(n30285), .Z(n31544) );
  XNOR U31525 ( .A(n31545), .B(n30291), .Z(n30285) );
  IV U31526 ( .A(n29268), .Z(n30291) );
  XOR U31527 ( .A(n31546), .B(n31107), .Z(n29268) );
  IV U31528 ( .A(n31547), .Z(n31107) );
  XOR U31529 ( .A(n31548), .B(n31549), .Z(n29141) );
  XNOR U31530 ( .A(n31550), .B(n29027), .Z(n29140) );
  XNOR U31531 ( .A(n31551), .B(n30304), .Z(n26523) );
  IV U31532 ( .A(n29273), .Z(n30304) );
  XOR U31533 ( .A(n31552), .B(n31376), .Z(n29273) );
  ANDN U31534 ( .B(n29150), .A(n29151), .Z(n31551) );
  XOR U31535 ( .A(n31553), .B(n30733), .Z(n29151) );
  XOR U31536 ( .A(n31554), .B(n31555), .Z(n29150) );
  XOR U31537 ( .A(n24271), .B(n31556), .Z(n31543) );
  XOR U31538 ( .A(n26020), .B(n26618), .Z(n31556) );
  XNOR U31539 ( .A(n31557), .B(n30296), .Z(n26618) );
  IV U31540 ( .A(n29263), .Z(n30296) );
  XOR U31541 ( .A(n31558), .B(n29747), .Z(n29263) );
  ANDN U31542 ( .B(n28910), .A(n30295), .Z(n31557) );
  IV U31543 ( .A(n29148), .Z(n30295) );
  XOR U31544 ( .A(n31559), .B(n31560), .Z(n29148) );
  XOR U31545 ( .A(n30865), .B(n31561), .Z(n28910) );
  XNOR U31546 ( .A(n31562), .B(n29259), .Z(n26020) );
  XOR U31547 ( .A(n31563), .B(n31340), .Z(n29259) );
  ANDN U31548 ( .B(n29145), .A(n28906), .Z(n31562) );
  IV U31549 ( .A(n29146), .Z(n28906) );
  XOR U31550 ( .A(n31564), .B(n31565), .Z(n29146) );
  XOR U31551 ( .A(n31566), .B(n31567), .Z(n29145) );
  XNOR U31552 ( .A(n31568), .B(n29276), .Z(n24271) );
  XOR U31553 ( .A(n31569), .B(n31071), .Z(n29276) );
  NOR U31554 ( .A(n29138), .B(n28920), .Z(n31568) );
  XOR U31555 ( .A(n31570), .B(n31571), .Z(n28920) );
  XOR U31556 ( .A(n31572), .B(n31440), .Z(n29138) );
  XOR U31557 ( .A(n31573), .B(n31574), .Z(n27576) );
  XNOR U31558 ( .A(n25864), .B(n27007), .Z(n31574) );
  XOR U31559 ( .A(n31575), .B(n28251), .Z(n27007) );
  XNOR U31560 ( .A(n31405), .B(n31576), .Z(n28251) );
  XOR U31561 ( .A(n31577), .B(n30768), .Z(n30565) );
  XOR U31562 ( .A(n31578), .B(n31579), .Z(n28252) );
  XOR U31563 ( .A(n31580), .B(n28255), .Z(n25864) );
  IV U31564 ( .A(n29588), .Z(n28255) );
  XOR U31565 ( .A(n31581), .B(n27942), .Z(n29588) );
  ANDN U31566 ( .B(n28256), .A(n30561), .Z(n31580) );
  XNOR U31567 ( .A(n31582), .B(n30105), .Z(n30561) );
  XOR U31568 ( .A(n31583), .B(n31584), .Z(n28256) );
  XOR U31569 ( .A(n26475), .B(n31585), .Z(n31573) );
  XOR U31570 ( .A(n28246), .B(n22505), .Z(n31585) );
  XOR U31571 ( .A(n31586), .B(n28261), .Z(n22505) );
  IV U31572 ( .A(n29582), .Z(n28261) );
  XOR U31573 ( .A(n30918), .B(n31587), .Z(n29582) );
  IV U31574 ( .A(n31588), .Z(n30918) );
  NOR U31575 ( .A(n28260), .B(n30549), .Z(n31586) );
  XOR U31576 ( .A(n31589), .B(n29166), .Z(n30549) );
  XNOR U31577 ( .A(n31590), .B(n30746), .Z(n28260) );
  XNOR U31578 ( .A(n31591), .B(n28264), .Z(n28246) );
  XOR U31579 ( .A(n31592), .B(n31454), .Z(n28264) );
  ANDN U31580 ( .B(n28265), .A(n30552), .Z(n31591) );
  XNOR U31581 ( .A(n31593), .B(n31565), .Z(n30552) );
  XNOR U31582 ( .A(n31594), .B(n31595), .Z(n28265) );
  XNOR U31583 ( .A(n31596), .B(n29579), .Z(n26475) );
  IV U31584 ( .A(n28269), .Z(n29579) );
  XNOR U31585 ( .A(n31597), .B(n31598), .Z(n28269) );
  NOR U31586 ( .A(n30557), .B(n28268), .Z(n31596) );
  IV U31587 ( .A(n31599), .Z(n30557) );
  XOR U31588 ( .A(n31600), .B(n28268), .Z(n31065) );
  XOR U31589 ( .A(n31601), .B(n31549), .Z(n28268) );
  ANDN U31590 ( .B(n29578), .A(n31599), .Z(n31600) );
  XOR U31591 ( .A(n30277), .B(n31602), .Z(n31599) );
  XNOR U31592 ( .A(n31359), .B(n31603), .Z(n29578) );
  XNOR U31593 ( .A(n16400), .B(n31604), .Z(n31413) );
  XOR U31594 ( .A(n15952), .B(n17125), .Z(n31604) );
  XNOR U31595 ( .A(n31605), .B(n21471), .Z(n17125) );
  XOR U31596 ( .A(n31606), .B(n23558), .Z(n21471) );
  XOR U31597 ( .A(n28731), .B(n26756), .Z(n23558) );
  XNOR U31598 ( .A(n31607), .B(n31608), .Z(n26756) );
  XOR U31599 ( .A(n31609), .B(n25537), .Z(n31608) );
  XOR U31600 ( .A(n31610), .B(n31611), .Z(n25537) );
  ANDN U31601 ( .B(n31081), .A(n30831), .Z(n31610) );
  XOR U31602 ( .A(n31612), .B(n31613), .Z(n30831) );
  XOR U31603 ( .A(n25494), .B(n31614), .Z(n31607) );
  XNOR U31604 ( .A(n26793), .B(n24424), .Z(n31614) );
  XNOR U31605 ( .A(n31615), .B(n31616), .Z(n24424) );
  ANDN U31606 ( .B(n30840), .A(n31079), .Z(n31615) );
  XOR U31607 ( .A(n31617), .B(n31618), .Z(n30840) );
  XNOR U31608 ( .A(n31619), .B(n31620), .Z(n26793) );
  XOR U31609 ( .A(n31621), .B(n31622), .Z(n30844) );
  XNOR U31610 ( .A(n31623), .B(n31624), .Z(n25494) );
  ANDN U31611 ( .B(n31084), .A(n31085), .Z(n31623) );
  XNOR U31612 ( .A(n31625), .B(n30231), .Z(n31085) );
  XOR U31613 ( .A(n31626), .B(n31627), .Z(n28731) );
  XOR U31614 ( .A(n26457), .B(n30318), .Z(n31627) );
  XOR U31615 ( .A(n31628), .B(n27395), .Z(n30318) );
  XOR U31616 ( .A(n31629), .B(n30210), .Z(n27395) );
  AND U31617 ( .A(n30863), .B(n30329), .Z(n31628) );
  XNOR U31618 ( .A(n31630), .B(n27400), .Z(n26457) );
  XNOR U31619 ( .A(n31631), .B(n31632), .Z(n27400) );
  NOR U31620 ( .A(n30323), .B(n30867), .Z(n31630) );
  XOR U31621 ( .A(n28711), .B(n31633), .Z(n31626) );
  XOR U31622 ( .A(n25748), .B(n23809), .Z(n31633) );
  XNOR U31623 ( .A(n31634), .B(n27537), .Z(n23809) );
  XOR U31624 ( .A(n31635), .B(n31636), .Z(n27537) );
  AND U31625 ( .A(n30331), .B(n30854), .Z(n31634) );
  XNOR U31626 ( .A(n31637), .B(n27405), .Z(n25748) );
  XNOR U31627 ( .A(n31622), .B(n31638), .Z(n27405) );
  AND U31628 ( .A(n30850), .B(n30325), .Z(n31637) );
  XNOR U31629 ( .A(n31639), .B(n30334), .Z(n28711) );
  XNOR U31630 ( .A(n29271), .B(n31640), .Z(n30334) );
  AND U31631 ( .A(n21104), .B(n21106), .Z(n31605) );
  XOR U31632 ( .A(n25896), .B(n27800), .Z(n21106) );
  XOR U31633 ( .A(n31641), .B(n27784), .Z(n27800) );
  ANDN U31634 ( .B(n27927), .A(n27626), .Z(n31641) );
  XOR U31635 ( .A(n31642), .B(n31643), .Z(n27626) );
  IV U31636 ( .A(n24390), .Z(n25896) );
  XOR U31637 ( .A(n31644), .B(n31645), .Z(n24390) );
  XNOR U31638 ( .A(n23484), .B(n27077), .Z(n21104) );
  XNOR U31639 ( .A(n31646), .B(n31647), .Z(n27077) );
  ANDN U31640 ( .B(n28602), .A(n28603), .Z(n31646) );
  XOR U31641 ( .A(n31648), .B(n31649), .Z(n28603) );
  IV U31642 ( .A(n21229), .Z(n23484) );
  XOR U31643 ( .A(n26412), .B(n28417), .Z(n21229) );
  XNOR U31644 ( .A(n31650), .B(n31651), .Z(n28417) );
  XOR U31645 ( .A(n24928), .B(n24838), .Z(n31651) );
  XOR U31646 ( .A(n31652), .B(n28785), .Z(n24838) );
  XOR U31647 ( .A(n31653), .B(n31654), .Z(n28785) );
  ANDN U31648 ( .B(n30139), .A(n28784), .Z(n31652) );
  XOR U31649 ( .A(n31655), .B(n30197), .Z(n28784) );
  XNOR U31650 ( .A(n31656), .B(n31657), .Z(n30139) );
  XOR U31651 ( .A(n31658), .B(n27270), .Z(n24928) );
  XOR U31652 ( .A(n31659), .B(n31660), .Z(n27270) );
  NOR U31653 ( .A(n28581), .B(n27271), .Z(n31658) );
  XNOR U31654 ( .A(n28807), .B(n31661), .Z(n27271) );
  XOR U31655 ( .A(n31662), .B(n31663), .Z(n28581) );
  XOR U31656 ( .A(n23567), .B(n31664), .Z(n31650) );
  XOR U31657 ( .A(n25287), .B(n25401), .Z(n31664) );
  XNOR U31658 ( .A(n31666), .B(n31667), .Z(n27276) );
  ANDN U31659 ( .B(n27277), .A(n28578), .Z(n31665) );
  XNOR U31660 ( .A(n31668), .B(n30524), .Z(n28578) );
  XNOR U31661 ( .A(n31669), .B(n31670), .Z(n27277) );
  XOR U31662 ( .A(n31671), .B(n27673), .Z(n25287) );
  XOR U31663 ( .A(n29938), .B(n31672), .Z(n27673) );
  ANDN U31664 ( .B(n27672), .A(n28589), .Z(n31671) );
  XOR U31665 ( .A(n31673), .B(n31674), .Z(n28589) );
  XOR U31666 ( .A(n31675), .B(n31676), .Z(n27672) );
  XNOR U31667 ( .A(n31677), .B(n27281), .Z(n23567) );
  XOR U31668 ( .A(n31678), .B(n30208), .Z(n27281) );
  ANDN U31669 ( .B(n27280), .A(n28586), .Z(n31677) );
  XOR U31670 ( .A(n31679), .B(n31680), .Z(n28586) );
  XOR U31671 ( .A(n31681), .B(n31226), .Z(n27280) );
  XOR U31672 ( .A(n31682), .B(n31683), .Z(n26412) );
  XOR U31673 ( .A(n26912), .B(n22011), .Z(n31683) );
  XOR U31674 ( .A(n31684), .B(n29714), .Z(n22011) );
  XOR U31675 ( .A(n31685), .B(n30903), .Z(n29714) );
  ANDN U31676 ( .B(n27088), .A(n27090), .Z(n31684) );
  XOR U31677 ( .A(n31686), .B(n31687), .Z(n27090) );
  XOR U31678 ( .A(n31688), .B(n27933), .Z(n27088) );
  XOR U31679 ( .A(n31689), .B(n29723), .Z(n26912) );
  XOR U31680 ( .A(n31690), .B(n29171), .Z(n29723) );
  AND U31681 ( .A(n27081), .B(n27079), .Z(n31689) );
  XOR U31682 ( .A(n30247), .B(n31691), .Z(n27079) );
  XOR U31683 ( .A(n31692), .B(n30375), .Z(n27081) );
  XOR U31684 ( .A(n24725), .B(n31693), .Z(n31682) );
  XOR U31685 ( .A(n27263), .B(n23917), .Z(n31693) );
  XOR U31686 ( .A(n31695), .B(n31539), .Z(n29718) );
  ANDN U31687 ( .B(n27085), .A(n27084), .Z(n31694) );
  XNOR U31688 ( .A(n31696), .B(n29916), .Z(n27084) );
  XOR U31689 ( .A(n31697), .B(n31698), .Z(n27085) );
  XNOR U31690 ( .A(n31699), .B(n29726), .Z(n27263) );
  XOR U31691 ( .A(n31700), .B(n31701), .Z(n29726) );
  NOR U31692 ( .A(n27092), .B(n27093), .Z(n31699) );
  XNOR U31693 ( .A(n31702), .B(n31001), .Z(n27093) );
  XOR U31694 ( .A(n31703), .B(n30544), .Z(n27092) );
  XOR U31695 ( .A(n31704), .B(n29728), .Z(n24725) );
  XOR U31696 ( .A(n31705), .B(n29045), .Z(n29728) );
  NOR U31697 ( .A(n31647), .B(n28602), .Z(n31704) );
  XOR U31698 ( .A(n31706), .B(n31707), .Z(n28602) );
  IV U31699 ( .A(n30072), .Z(n31647) );
  XOR U31700 ( .A(n31708), .B(n31709), .Z(n30072) );
  XNOR U31701 ( .A(n19845), .B(n31710), .Z(n15952) );
  XOR U31702 ( .A(n31711), .B(n31712), .Z(n31710) );
  NANDN U31703 ( .A(n19844), .B(n21147), .Z(n31712) );
  XNOR U31704 ( .A(n28626), .B(n22354), .Z(n21147) );
  XOR U31705 ( .A(n31714), .B(n31715), .Z(n29883) );
  XNOR U31706 ( .A(n24991), .B(n23832), .Z(n31715) );
  XNOR U31707 ( .A(n31716), .B(n31717), .Z(n23832) );
  ANDN U31708 ( .B(n27220), .A(n27218), .Z(n31716) );
  XNOR U31709 ( .A(n31718), .B(n31719), .Z(n24991) );
  ANDN U31710 ( .B(n27212), .A(n27213), .Z(n31718) );
  XOR U31711 ( .A(n31720), .B(n31721), .Z(n31714) );
  XOR U31712 ( .A(n24451), .B(n23990), .Z(n31721) );
  XNOR U31713 ( .A(n31722), .B(n31723), .Z(n23990) );
  XNOR U31714 ( .A(n31724), .B(n31725), .Z(n24451) );
  NOR U31715 ( .A(n31726), .B(n29909), .Z(n31724) );
  XNOR U31716 ( .A(n31727), .B(n31728), .Z(n28626) );
  AND U31717 ( .A(n30703), .B(n31729), .Z(n31727) );
  XNOR U31718 ( .A(n31730), .B(n25424), .Z(n19844) );
  XOR U31719 ( .A(n31731), .B(n24314), .Z(n25424) );
  XOR U31720 ( .A(n31732), .B(n31733), .Z(n24314) );
  XNOR U31721 ( .A(n26401), .B(n26551), .Z(n31733) );
  XNOR U31722 ( .A(n31734), .B(n29898), .Z(n26551) );
  XNOR U31723 ( .A(n31735), .B(n29717), .Z(n29898) );
  ANDN U31724 ( .B(n31736), .A(n30052), .Z(n31734) );
  XNOR U31725 ( .A(n31737), .B(n29893), .Z(n26401) );
  XOR U31726 ( .A(n31738), .B(n31739), .Z(n29893) );
  ANDN U31727 ( .B(n30055), .A(n31740), .Z(n31737) );
  XNOR U31728 ( .A(n26249), .B(n31741), .Z(n31732) );
  XNOR U31729 ( .A(n30022), .B(n25756), .Z(n31741) );
  XOR U31730 ( .A(n31742), .B(n30050), .Z(n25756) );
  IV U31731 ( .A(n29889), .Z(n30050) );
  XOR U31732 ( .A(n28762), .B(n31743), .Z(n29889) );
  NOR U31733 ( .A(n31744), .B(n30049), .Z(n31742) );
  XNOR U31734 ( .A(n31745), .B(n30045), .Z(n30022) );
  IV U31735 ( .A(n29906), .Z(n30045) );
  XOR U31736 ( .A(n31746), .B(n30258), .Z(n29906) );
  ANDN U31737 ( .B(n30046), .A(n31747), .Z(n31745) );
  XNOR U31738 ( .A(n31748), .B(n29901), .Z(n26249) );
  XNOR U31739 ( .A(n31749), .B(n31659), .Z(n29901) );
  NOR U31740 ( .A(n31750), .B(n31751), .Z(n31748) );
  XOR U31741 ( .A(n25289), .B(n28458), .Z(n19845) );
  XOR U31742 ( .A(n28737), .B(n31752), .Z(n28458) );
  XOR U31743 ( .A(n31753), .B(n4407), .Z(n31752) );
  XOR U31744 ( .A(n31754), .B(n31755), .Z(n26602) );
  XNOR U31745 ( .A(n31756), .B(n19628), .Z(n16400) );
  XNOR U31746 ( .A(n31757), .B(n23513), .Z(n19628) );
  XNOR U31747 ( .A(n31758), .B(n31759), .Z(n27704) );
  XOR U31748 ( .A(n26396), .B(n24145), .Z(n31759) );
  XOR U31749 ( .A(n31760), .B(n29458), .Z(n24145) );
  NOR U31750 ( .A(n28345), .B(n29457), .Z(n31760) );
  IV U31751 ( .A(n31761), .Z(n28345) );
  XOR U31752 ( .A(n31762), .B(n29453), .Z(n26396) );
  NOR U31753 ( .A(n29452), .B(n28353), .Z(n31762) );
  XOR U31754 ( .A(n24263), .B(n31763), .Z(n31758) );
  XNOR U31755 ( .A(n29447), .B(n28495), .Z(n31763) );
  XNOR U31756 ( .A(n31764), .B(n30384), .Z(n28495) );
  NOR U31757 ( .A(n28340), .B(n30385), .Z(n31764) );
  XNOR U31758 ( .A(n31765), .B(n30019), .Z(n29447) );
  NOR U31759 ( .A(n28349), .B(n30018), .Z(n31765) );
  XNOR U31760 ( .A(n31766), .B(n31767), .Z(n24263) );
  NOR U31761 ( .A(n29460), .B(n29037), .Z(n31766) );
  XOR U31762 ( .A(n31768), .B(n31769), .Z(n27851) );
  XOR U31763 ( .A(n27674), .B(n28778), .Z(n31769) );
  XOR U31764 ( .A(n31770), .B(n29483), .Z(n28778) );
  XOR U31765 ( .A(n31771), .B(n30520), .Z(n29483) );
  IV U31766 ( .A(n31772), .Z(n30520) );
  ANDN U31767 ( .B(n31773), .A(n31774), .Z(n31770) );
  XNOR U31768 ( .A(n29471), .B(n31775), .Z(n27674) );
  XOR U31769 ( .A(n31776), .B(n21688), .Z(n31775) );
  NANDN U31770 ( .A(rc_i[1]), .B(n4549), .Z(n21688) );
  NOR U31771 ( .A(n29470), .B(n31429), .Z(n31776) );
  XOR U31772 ( .A(n31777), .B(n30733), .Z(n29471) );
  XNOR U31773 ( .A(n27262), .B(n31778), .Z(n31768) );
  XNOR U31774 ( .A(n26748), .B(n24410), .Z(n31778) );
  XNOR U31775 ( .A(n31779), .B(n29467), .Z(n24410) );
  XOR U31776 ( .A(n31780), .B(n30514), .Z(n29467) );
  ANDN U31777 ( .B(n31438), .A(n29466), .Z(n31779) );
  XNOR U31778 ( .A(n31781), .B(n29476), .Z(n26748) );
  XOR U31779 ( .A(n31782), .B(n31783), .Z(n29476) );
  NOR U31780 ( .A(n31442), .B(n29475), .Z(n31781) );
  XOR U31781 ( .A(n31784), .B(n29480), .Z(n27262) );
  XOR U31782 ( .A(n31785), .B(n31786), .Z(n29480) );
  ANDN U31783 ( .B(n31432), .A(n29479), .Z(n31784) );
  XNOR U31784 ( .A(n29333), .B(n22790), .Z(n19627) );
  XNOR U31785 ( .A(n31787), .B(n31788), .Z(n31008) );
  XNOR U31786 ( .A(n23056), .B(n25713), .Z(n31788) );
  XNOR U31787 ( .A(n31789), .B(n29654), .Z(n25713) );
  IV U31788 ( .A(n31790), .Z(n29654) );
  XOR U31789 ( .A(n31618), .B(n31791), .Z(n30925) );
  XNOR U31790 ( .A(n31792), .B(n29647), .Z(n23056) );
  ANDN U31791 ( .B(n29361), .A(n29362), .Z(n31792) );
  XOR U31792 ( .A(n31793), .B(n31794), .Z(n29362) );
  XNOR U31793 ( .A(n24505), .B(n31795), .Z(n31787) );
  XNOR U31794 ( .A(n29373), .B(n28865), .Z(n31795) );
  XNOR U31795 ( .A(n31796), .B(n31797), .Z(n28865) );
  NOR U31796 ( .A(n29366), .B(n29365), .Z(n31796) );
  XOR U31797 ( .A(n30277), .B(n31798), .Z(n29366) );
  ANDN U31798 ( .B(n29351), .A(n29352), .Z(n31799) );
  XNOR U31799 ( .A(n31137), .B(n31800), .Z(n29352) );
  XNOR U31800 ( .A(n31801), .B(n29644), .Z(n24505) );
  NOR U31801 ( .A(n29356), .B(n29355), .Z(n31801) );
  XOR U31802 ( .A(n31802), .B(n27933), .Z(n29356) );
  XOR U31803 ( .A(n31803), .B(n31804), .Z(n26730) );
  XNOR U31804 ( .A(n26860), .B(n26151), .Z(n31804) );
  XNOR U31805 ( .A(n31805), .B(n28938), .Z(n26151) );
  NOR U31806 ( .A(n29339), .B(n29340), .Z(n31805) );
  XOR U31807 ( .A(n31806), .B(n31807), .Z(n29340) );
  IV U31808 ( .A(n31808), .Z(n29339) );
  XOR U31809 ( .A(n31809), .B(n28930), .Z(n26860) );
  ANDN U31810 ( .B(n29346), .A(n29347), .Z(n31809) );
  XOR U31811 ( .A(n31810), .B(n31811), .Z(n29347) );
  XOR U31812 ( .A(n23587), .B(n31812), .Z(n31803) );
  XOR U31813 ( .A(n22647), .B(n31813), .Z(n31812) );
  XNOR U31814 ( .A(n31814), .B(n28935), .Z(n22647) );
  XOR U31815 ( .A(n31815), .B(n30544), .Z(n29336) );
  NOR U31816 ( .A(n30907), .B(n31817), .Z(n31816) );
  XNOR U31817 ( .A(n31818), .B(n31817), .Z(n29333) );
  ANDN U31818 ( .B(n30907), .A(n28941), .Z(n31818) );
  XOR U31819 ( .A(n31819), .B(n31820), .Z(n28941) );
  XOR U31820 ( .A(n31821), .B(n31822), .Z(n30907) );
  XOR U31821 ( .A(n24063), .B(n29103), .Z(n27903) );
  XNOR U31822 ( .A(n31823), .B(n27427), .Z(n29103) );
  ANDN U31823 ( .B(n30241), .A(n29878), .Z(n31823) );
  IV U31824 ( .A(n22643), .Z(n24063) );
  XNOR U31825 ( .A(n31825), .B(n26055), .Z(n22643) );
  XOR U31826 ( .A(n31826), .B(n31827), .Z(n26055) );
  XNOR U31827 ( .A(n25019), .B(n24358), .Z(n31827) );
  XNOR U31828 ( .A(n31828), .B(n31829), .Z(n24358) );
  ANDN U31829 ( .B(n29235), .A(n29773), .Z(n31828) );
  IV U31830 ( .A(n29237), .Z(n29773) );
  XOR U31831 ( .A(n31830), .B(n31333), .Z(n29237) );
  XNOR U31832 ( .A(n31831), .B(n30016), .Z(n25019) );
  ANDN U31833 ( .B(n29231), .A(n29233), .Z(n31831) );
  XOR U31834 ( .A(n31833), .B(n31834), .Z(n29231) );
  XOR U31835 ( .A(n25811), .B(n31835), .Z(n31826) );
  XOR U31836 ( .A(n24161), .B(n25656), .Z(n31835) );
  XOR U31837 ( .A(n31836), .B(n26212), .Z(n25656) );
  ANDN U31838 ( .B(n29244), .A(n26211), .Z(n31836) );
  XNOR U31839 ( .A(n31837), .B(n29959), .Z(n26211) );
  XNOR U31840 ( .A(n31838), .B(n29528), .Z(n29244) );
  XNOR U31841 ( .A(n31839), .B(n26205), .Z(n24161) );
  AND U31842 ( .A(n26206), .B(n29241), .Z(n31839) );
  XNOR U31843 ( .A(n31840), .B(n31841), .Z(n29241) );
  XOR U31844 ( .A(n30573), .B(n31842), .Z(n26206) );
  XNOR U31845 ( .A(n31843), .B(n26215), .Z(n25811) );
  ANDN U31846 ( .B(n26216), .A(n29246), .Z(n31843) );
  XOR U31847 ( .A(n31844), .B(n31845), .Z(n29246) );
  XNOR U31848 ( .A(n29736), .B(n31846), .Z(n26216) );
  XOR U31849 ( .A(n31847), .B(n31848), .Z(n19828) );
  XOR U31850 ( .A(n18418), .B(n24799), .Z(n31848) );
  XNOR U31851 ( .A(n31849), .B(n25386), .Z(n24799) );
  XNOR U31852 ( .A(n31850), .B(n24518), .Z(n25386) );
  XNOR U31853 ( .A(n31851), .B(n31852), .Z(n28109) );
  XOR U31854 ( .A(n26539), .B(n26502), .Z(n31852) );
  XNOR U31855 ( .A(n31853), .B(n30349), .Z(n26502) );
  AND U31856 ( .A(n31525), .B(n30350), .Z(n31853) );
  XOR U31857 ( .A(n31856), .B(n30353), .Z(n26539) );
  XOR U31858 ( .A(n31857), .B(n31858), .Z(n30353) );
  ANDN U31859 ( .B(n30354), .A(n31859), .Z(n31856) );
  XOR U31860 ( .A(n24935), .B(n31860), .Z(n31851) );
  XNOR U31861 ( .A(n25946), .B(n24905), .Z(n31860) );
  XNOR U31862 ( .A(n31861), .B(n30357), .Z(n24905) );
  ANDN U31863 ( .B(n30358), .A(n31528), .Z(n31861) );
  XNOR U31864 ( .A(n31863), .B(n30344), .Z(n25946) );
  XOR U31865 ( .A(n31864), .B(n31865), .Z(n30344) );
  ANDN U31866 ( .B(n30345), .A(n31537), .Z(n31863) );
  XOR U31867 ( .A(n31866), .B(n30340), .Z(n24935) );
  XNOR U31868 ( .A(n31867), .B(n30275), .Z(n30340) );
  ANDN U31869 ( .B(n30341), .A(n31533), .Z(n31866) );
  XOR U31870 ( .A(n31868), .B(n31869), .Z(n30985) );
  XOR U31871 ( .A(n28066), .B(n24169), .Z(n31869) );
  XNOR U31872 ( .A(n31870), .B(n28089), .Z(n24169) );
  XOR U31873 ( .A(n31871), .B(n31872), .Z(n28089) );
  ANDN U31874 ( .B(n31311), .A(n28088), .Z(n31870) );
  XNOR U31875 ( .A(n31873), .B(n28081), .Z(n28066) );
  IV U31876 ( .A(n29793), .Z(n28081) );
  XNOR U31877 ( .A(n31874), .B(n28744), .Z(n29793) );
  NOR U31878 ( .A(n28080), .B(n31316), .Z(n31873) );
  XNOR U31879 ( .A(n27881), .B(n31875), .Z(n31868) );
  XOR U31880 ( .A(n25917), .B(n22410), .Z(n31875) );
  XNOR U31881 ( .A(n31876), .B(n28076), .Z(n22410) );
  XOR U31882 ( .A(n31877), .B(n29175), .Z(n28076) );
  NOR U31883 ( .A(n31304), .B(n28075), .Z(n31876) );
  XNOR U31884 ( .A(n31878), .B(n28084), .Z(n25917) );
  XOR U31885 ( .A(n31879), .B(n31880), .Z(n28084) );
  ANDN U31886 ( .B(n28085), .A(n31319), .Z(n31878) );
  XOR U31887 ( .A(n31881), .B(n28071), .Z(n27881) );
  XOR U31888 ( .A(n31882), .B(n30583), .Z(n28071) );
  ANDN U31889 ( .B(n28072), .A(n31307), .Z(n31881) );
  ANDN U31890 ( .B(n21861), .A(n24322), .Z(n31849) );
  XOR U31891 ( .A(n28618), .B(n25163), .Z(n24322) );
  XOR U31892 ( .A(n31713), .B(n26469), .Z(n25163) );
  XNOR U31893 ( .A(n31883), .B(n31884), .Z(n26469) );
  XNOR U31894 ( .A(n26181), .B(n21719), .Z(n31884) );
  XOR U31895 ( .A(n31885), .B(n30994), .Z(n21719) );
  NOR U31896 ( .A(n28623), .B(n28104), .Z(n31885) );
  XOR U31897 ( .A(n31886), .B(n31887), .Z(n28104) );
  XNOR U31898 ( .A(n31888), .B(n30991), .Z(n26181) );
  ANDN U31899 ( .B(n28620), .A(n28169), .Z(n31888) );
  IV U31900 ( .A(n28621), .Z(n28169) );
  XOR U31901 ( .A(n30657), .B(n31889), .Z(n28621) );
  XOR U31902 ( .A(n29796), .B(n31890), .Z(n31883) );
  XOR U31903 ( .A(n31891), .B(n23323), .Z(n31890) );
  XNOR U31904 ( .A(n31892), .B(n31002), .Z(n23323) );
  NOR U31905 ( .A(n28616), .B(n28094), .Z(n31892) );
  XNOR U31906 ( .A(n31893), .B(n31894), .Z(n28094) );
  XNOR U31907 ( .A(n31895), .B(n30998), .Z(n29796) );
  IV U31908 ( .A(n31896), .Z(n30998) );
  ANDN U31909 ( .B(n31897), .A(n28100), .Z(n31895) );
  IV U31910 ( .A(n31898), .Z(n28100) );
  XOR U31911 ( .A(n31899), .B(n31900), .Z(n31713) );
  XNOR U31912 ( .A(n25995), .B(n27960), .Z(n31900) );
  XNOR U31913 ( .A(n31901), .B(n31902), .Z(n27960) );
  ANDN U31914 ( .B(n28641), .A(n31903), .Z(n31901) );
  XNOR U31915 ( .A(n31904), .B(n31905), .Z(n25995) );
  NOR U31916 ( .A(n28634), .B(n28633), .Z(n31904) );
  XNOR U31917 ( .A(n23249), .B(n31906), .Z(n31899) );
  XOR U31918 ( .A(n28108), .B(n28712), .Z(n31906) );
  XNOR U31919 ( .A(n31907), .B(n31908), .Z(n28712) );
  NOR U31920 ( .A(n28639), .B(n28637), .Z(n31907) );
  XNOR U31921 ( .A(n31909), .B(n30708), .Z(n28108) );
  ANDN U31922 ( .B(n28628), .A(n28630), .Z(n31909) );
  XOR U31923 ( .A(n31910), .B(n31911), .Z(n23249) );
  NOR U31924 ( .A(n31729), .B(n31728), .Z(n31910) );
  XNOR U31925 ( .A(n31912), .B(n31897), .Z(n28618) );
  ANDN U31926 ( .B(n30997), .A(n31898), .Z(n31912) );
  IV U31927 ( .A(n28101), .Z(n30997) );
  XOR U31928 ( .A(n31914), .B(n30208), .Z(n28101) );
  XOR U31929 ( .A(n26283), .B(n27988), .Z(n21861) );
  XNOR U31930 ( .A(n31915), .B(n31487), .Z(n27988) );
  ANDN U31931 ( .B(n31916), .A(n31917), .Z(n31915) );
  XNOR U31932 ( .A(n31918), .B(n26453), .Z(n18418) );
  XOR U31933 ( .A(n26135), .B(n28327), .Z(n26453) );
  XOR U31934 ( .A(n31919), .B(n27719), .Z(n28327) );
  ANDN U31935 ( .B(n31920), .A(n31921), .Z(n31919) );
  XOR U31936 ( .A(n29040), .B(n27637), .Z(n26135) );
  XNOR U31937 ( .A(n31922), .B(n31923), .Z(n27637) );
  XOR U31938 ( .A(n25300), .B(n27703), .Z(n31923) );
  XNOR U31939 ( .A(n31924), .B(n27231), .Z(n27703) );
  XOR U31940 ( .A(n31925), .B(n31663), .Z(n27231) );
  ANDN U31941 ( .B(n27710), .A(n28335), .Z(n31924) );
  XNOR U31942 ( .A(n31926), .B(n31565), .Z(n27710) );
  XNOR U31943 ( .A(n31927), .B(n27720), .Z(n25300) );
  NOR U31944 ( .A(n27719), .B(n31920), .Z(n31927) );
  XNOR U31945 ( .A(n31928), .B(n31657), .Z(n27719) );
  XOR U31946 ( .A(n26063), .B(n31929), .Z(n31922) );
  XNOR U31947 ( .A(n23020), .B(n25553), .Z(n31929) );
  XNOR U31948 ( .A(n31930), .B(n26683), .Z(n25553) );
  XNOR U31949 ( .A(n31026), .B(n31931), .Z(n26683) );
  NOR U31950 ( .A(n29855), .B(n27716), .Z(n31930) );
  XNOR U31951 ( .A(n31932), .B(n28462), .Z(n27716) );
  XNOR U31952 ( .A(n31933), .B(n26687), .Z(n23020) );
  XOR U31953 ( .A(n31934), .B(n29291), .Z(n26687) );
  IV U31954 ( .A(n31549), .Z(n29291) );
  XNOR U31955 ( .A(n31935), .B(n30535), .Z(n27713) );
  XNOR U31956 ( .A(n31936), .B(n26678), .Z(n26063) );
  XOR U31957 ( .A(n31937), .B(n31333), .Z(n26678) );
  IV U31958 ( .A(n28879), .Z(n31333) );
  ANDN U31959 ( .B(n28333), .A(n27708), .Z(n31936) );
  XOR U31960 ( .A(n30066), .B(n31938), .Z(n27708) );
  XOR U31961 ( .A(n31939), .B(n31940), .Z(n29040) );
  XOR U31962 ( .A(n25196), .B(n25816), .Z(n31940) );
  XOR U31963 ( .A(n31941), .B(n30018), .Z(n25816) );
  XOR U31964 ( .A(n31942), .B(n31943), .Z(n30018) );
  ANDN U31965 ( .B(n28349), .A(n28351), .Z(n31941) );
  XOR U31966 ( .A(n30253), .B(n31944), .Z(n28349) );
  XNOR U31967 ( .A(n31945), .B(n29460), .Z(n25196) );
  XNOR U31968 ( .A(n28762), .B(n31946), .Z(n29460) );
  ANDN U31969 ( .B(n29037), .A(n29038), .Z(n31945) );
  XNOR U31970 ( .A(n31947), .B(n31948), .Z(n29037) );
  XOR U31971 ( .A(n25950), .B(n31949), .Z(n31939) );
  XNOR U31972 ( .A(n23512), .B(n31757), .Z(n31949) );
  XNOR U31973 ( .A(n31950), .B(n30385), .Z(n31757) );
  XOR U31974 ( .A(n31951), .B(n31952), .Z(n30385) );
  ANDN U31975 ( .B(n28340), .A(n28341), .Z(n31950) );
  XOR U31976 ( .A(n31953), .B(n30554), .Z(n28340) );
  XNOR U31977 ( .A(n31954), .B(n29452), .Z(n23512) );
  XOR U31978 ( .A(n31955), .B(n31956), .Z(n29452) );
  ANDN U31979 ( .B(n28353), .A(n28354), .Z(n31954) );
  XOR U31980 ( .A(n31957), .B(n28428), .Z(n28353) );
  XNOR U31981 ( .A(n31958), .B(n29457), .Z(n25950) );
  XOR U31982 ( .A(n31959), .B(n31960), .Z(n29457) );
  NOR U31983 ( .A(n31761), .B(n28346), .Z(n31958) );
  XNOR U31984 ( .A(n30000), .B(n31961), .Z(n31761) );
  ANDN U31985 ( .B(n24326), .A(n24324), .Z(n31918) );
  IV U31986 ( .A(n25389), .Z(n24324) );
  XOR U31987 ( .A(n29129), .B(n23985), .Z(n25389) );
  XOR U31988 ( .A(n31825), .B(n30225), .Z(n23985) );
  XNOR U31989 ( .A(n31962), .B(n31963), .Z(n30225) );
  XNOR U31990 ( .A(n24293), .B(n23977), .Z(n31963) );
  XNOR U31991 ( .A(n31964), .B(n28691), .Z(n23977) );
  XNOR U31992 ( .A(n28762), .B(n31965), .Z(n28691) );
  NOR U31993 ( .A(n28690), .B(n30281), .Z(n31964) );
  XOR U31994 ( .A(n31967), .B(n31968), .Z(n28682) );
  ANDN U31995 ( .B(n29127), .A(n28681), .Z(n31966) );
  XOR U31996 ( .A(n27661), .B(n31969), .Z(n28681) );
  XOR U31997 ( .A(n31970), .B(n30303), .Z(n29127) );
  XOR U31998 ( .A(n25977), .B(n31971), .Z(n31962) );
  XNOR U31999 ( .A(n26521), .B(n27407), .Z(n31971) );
  XOR U32000 ( .A(n31972), .B(n28687), .Z(n27407) );
  XOR U32001 ( .A(n31190), .B(n31973), .Z(n28687) );
  NOR U32002 ( .A(n29122), .B(n29124), .Z(n31972) );
  XOR U32003 ( .A(n31974), .B(n30105), .Z(n29124) );
  IV U32004 ( .A(n28686), .Z(n29122) );
  XOR U32005 ( .A(n31975), .B(n31178), .Z(n28686) );
  XNOR U32006 ( .A(n31976), .B(n29865), .Z(n26521) );
  XOR U32007 ( .A(n31977), .B(n30990), .Z(n29865) );
  NOR U32008 ( .A(n29753), .B(n29754), .Z(n31976) );
  XOR U32009 ( .A(n31978), .B(n28798), .Z(n29754) );
  IV U32010 ( .A(n29882), .Z(n29753) );
  XOR U32011 ( .A(n31979), .B(n30554), .Z(n29882) );
  XNOR U32012 ( .A(n31980), .B(n28694), .Z(n25977) );
  XOR U32013 ( .A(n29930), .B(n31981), .Z(n28694) );
  ANDN U32014 ( .B(n28695), .A(n29132), .Z(n31980) );
  XNOR U32015 ( .A(n31982), .B(n31983), .Z(n29132) );
  XNOR U32016 ( .A(n31984), .B(n31595), .Z(n28695) );
  XOR U32017 ( .A(n31985), .B(n31986), .Z(n31825) );
  XOR U32018 ( .A(n25613), .B(n26198), .Z(n31986) );
  XOR U32019 ( .A(n31987), .B(n27430), .Z(n26198) );
  XOR U32020 ( .A(n28987), .B(n31988), .Z(n27430) );
  ANDN U32021 ( .B(n27431), .A(n30256), .Z(n31987) );
  XOR U32022 ( .A(n31989), .B(n28836), .Z(n30256) );
  XNOR U32023 ( .A(n31990), .B(n31405), .Z(n27431) );
  XNOR U32024 ( .A(n31991), .B(n27414), .Z(n25613) );
  XNOR U32025 ( .A(n31992), .B(n29747), .Z(n27414) );
  NOR U32026 ( .A(n29113), .B(n29114), .Z(n31991) );
  XNOR U32027 ( .A(n31993), .B(n31071), .Z(n29114) );
  XNOR U32028 ( .A(n31994), .B(n29930), .Z(n29113) );
  XOR U32029 ( .A(n25200), .B(n31995), .Z(n31985) );
  XNOR U32030 ( .A(n22948), .B(n24385), .Z(n31995) );
  XOR U32031 ( .A(n31996), .B(n27423), .Z(n24385) );
  XOR U32032 ( .A(n31997), .B(n31998), .Z(n27423) );
  NOR U32033 ( .A(n29109), .B(n29110), .Z(n31996) );
  XOR U32034 ( .A(n31999), .B(n32000), .Z(n29110) );
  XOR U32035 ( .A(n32001), .B(n31434), .Z(n29109) );
  XOR U32036 ( .A(n32002), .B(n27417), .Z(n22948) );
  XOR U32037 ( .A(n31840), .B(n32003), .Z(n27417) );
  AND U32038 ( .A(n29106), .B(n27418), .Z(n32002) );
  XOR U32039 ( .A(n32004), .B(n31535), .Z(n27418) );
  XOR U32040 ( .A(n32005), .B(n32006), .Z(n29106) );
  XNOR U32041 ( .A(n32007), .B(n27426), .Z(n25200) );
  XOR U32042 ( .A(n32008), .B(n32009), .Z(n27426) );
  NOR U32043 ( .A(n27427), .B(n30241), .Z(n32007) );
  XNOR U32044 ( .A(n32010), .B(n32011), .Z(n30241) );
  XOR U32045 ( .A(n29072), .B(n32012), .Z(n27427) );
  XOR U32046 ( .A(n32014), .B(n32015), .Z(n28690) );
  ANDN U32047 ( .B(n30281), .A(n29869), .Z(n32013) );
  XOR U32048 ( .A(n31005), .B(n32016), .Z(n29869) );
  XOR U32049 ( .A(n32017), .B(n32018), .Z(n30281) );
  XOR U32050 ( .A(n29086), .B(n23837), .Z(n24326) );
  XOR U32051 ( .A(n32019), .B(n27175), .Z(n23837) );
  XNOR U32052 ( .A(n32020), .B(n32021), .Z(n27175) );
  XNOR U32053 ( .A(n25540), .B(n22945), .Z(n32021) );
  XOR U32054 ( .A(n32023), .B(n30078), .Z(n29205) );
  AND U32055 ( .A(n29084), .B(n29082), .Z(n32022) );
  XNOR U32056 ( .A(n30860), .B(n32024), .Z(n29082) );
  XNOR U32057 ( .A(n32025), .B(n32026), .Z(n25540) );
  ANDN U32058 ( .B(n32027), .A(n27970), .Z(n32025) );
  XNOR U32059 ( .A(n27963), .B(n32028), .Z(n32020) );
  XOR U32060 ( .A(n27435), .B(n23026), .Z(n32028) );
  XNOR U32061 ( .A(n32029), .B(n28648), .Z(n23026) );
  XOR U32062 ( .A(n31045), .B(n32030), .Z(n28648) );
  AND U32063 ( .A(n29089), .B(n28649), .Z(n32029) );
  XOR U32064 ( .A(n32031), .B(n32032), .Z(n28649) );
  XOR U32065 ( .A(n32033), .B(n27977), .Z(n27435) );
  XOR U32066 ( .A(n32034), .B(n32035), .Z(n27977) );
  XOR U32067 ( .A(n32036), .B(n32000), .Z(n27976) );
  XNOR U32068 ( .A(n32037), .B(n27980), .Z(n27963) );
  XOR U32069 ( .A(n32038), .B(n32039), .Z(n27980) );
  ANDN U32070 ( .B(n27981), .A(n29079), .Z(n32037) );
  XOR U32071 ( .A(n32040), .B(n32041), .Z(n27981) );
  XNOR U32072 ( .A(n32043), .B(n32044), .Z(n27970) );
  ANDN U32073 ( .B(n32045), .A(n32027), .Z(n32042) );
  XOR U32074 ( .A(n19357), .B(n32046), .Z(n31847) );
  XNOR U32075 ( .A(n19437), .B(n25365), .Z(n32046) );
  XOR U32076 ( .A(n32047), .B(n25393), .Z(n25365) );
  XOR U32077 ( .A(n32048), .B(n24031), .Z(n25393) );
  IV U32078 ( .A(n24884), .Z(n24031) );
  XOR U32079 ( .A(n30699), .B(n27070), .Z(n24884) );
  XNOR U32080 ( .A(n32049), .B(n32050), .Z(n27070) );
  XOR U32081 ( .A(n23823), .B(n22887), .Z(n32050) );
  XOR U32082 ( .A(n32051), .B(n30055), .Z(n22887) );
  XOR U32083 ( .A(n32052), .B(n32053), .Z(n30055) );
  XNOR U32084 ( .A(n32054), .B(n30046), .Z(n23823) );
  XNOR U32085 ( .A(n32055), .B(n30956), .Z(n30046) );
  ANDN U32086 ( .B(n31747), .A(n29904), .Z(n32054) );
  IV U32087 ( .A(n32056), .Z(n29904) );
  XNOR U32088 ( .A(n23739), .B(n32057), .Z(n32049) );
  XOR U32089 ( .A(n24313), .B(n23696), .Z(n32057) );
  XNOR U32090 ( .A(n32058), .B(n31750), .Z(n23696) );
  IV U32091 ( .A(n30043), .Z(n31750) );
  XNOR U32092 ( .A(n31642), .B(n32059), .Z(n30043) );
  AND U32093 ( .A(n31751), .B(n29900), .Z(n32058) );
  XNOR U32094 ( .A(n32060), .B(n30049), .Z(n24313) );
  XNOR U32095 ( .A(n32061), .B(n30252), .Z(n30049) );
  ANDN U32096 ( .B(n31744), .A(n29887), .Z(n32060) );
  XNOR U32097 ( .A(n32062), .B(n30052), .Z(n23739) );
  XOR U32098 ( .A(n32063), .B(n32064), .Z(n30052) );
  ANDN U32099 ( .B(n29896), .A(n31736), .Z(n32062) );
  XNOR U32100 ( .A(n32065), .B(n32066), .Z(n30699) );
  XOR U32101 ( .A(n25423), .B(n31730), .Z(n32066) );
  XOR U32102 ( .A(n32067), .B(n27223), .Z(n31730) );
  ANDN U32103 ( .B(n32068), .A(n31723), .Z(n32067) );
  XOR U32104 ( .A(n32069), .B(n27219), .Z(n25423) );
  IV U32105 ( .A(n32070), .Z(n27219) );
  ANDN U32106 ( .B(n32071), .A(n31717), .Z(n32069) );
  XNOR U32107 ( .A(n29839), .B(n32072), .Z(n32065) );
  XOR U32108 ( .A(n26008), .B(n28477), .Z(n32072) );
  XOR U32109 ( .A(n32073), .B(n27210), .Z(n28477) );
  ANDN U32110 ( .B(n32074), .A(n32075), .Z(n32073) );
  XOR U32111 ( .A(n32076), .B(n29910), .Z(n26008) );
  XOR U32112 ( .A(n32078), .B(n27214), .Z(n29839) );
  IV U32113 ( .A(n32079), .Z(n27214) );
  ANDN U32114 ( .B(n32080), .A(n31719), .Z(n32078) );
  NOR U32115 ( .A(n22874), .B(n24333), .Z(n32047) );
  XNOR U32116 ( .A(n26933), .B(n25356), .Z(n24333) );
  XNOR U32117 ( .A(n32081), .B(n32082), .Z(n28291) );
  XOR U32118 ( .A(n25411), .B(n25094), .Z(n32082) );
  XNOR U32119 ( .A(n32083), .B(n27444), .Z(n25094) );
  ANDN U32120 ( .B(n27006), .A(n27004), .Z(n32083) );
  XOR U32121 ( .A(n32084), .B(n28432), .Z(n27004) );
  XNOR U32122 ( .A(n32085), .B(n27030), .Z(n25411) );
  XOR U32123 ( .A(n32086), .B(n31565), .Z(n27030) );
  IV U32124 ( .A(n32041), .Z(n31565) );
  XNOR U32125 ( .A(n32087), .B(n32088), .Z(n32041) );
  NOR U32126 ( .A(n26937), .B(n26938), .Z(n32085) );
  XOR U32127 ( .A(n31405), .B(n32089), .Z(n26937) );
  XOR U32128 ( .A(n27282), .B(n32090), .Z(n32081) );
  XOR U32129 ( .A(n23572), .B(n25193), .Z(n32090) );
  XNOR U32130 ( .A(n32091), .B(n27022), .Z(n25193) );
  XOR U32131 ( .A(n32092), .B(n29927), .Z(n27022) );
  NOR U32132 ( .A(n32093), .B(n27447), .Z(n32091) );
  XNOR U32133 ( .A(n32094), .B(n27017), .Z(n23572) );
  XOR U32134 ( .A(n32095), .B(n31676), .Z(n27017) );
  ANDN U32135 ( .B(n26941), .A(n32096), .Z(n32094) );
  XOR U32136 ( .A(n32097), .B(n32098), .Z(n26941) );
  XNOR U32137 ( .A(n32099), .B(n27025), .Z(n27282) );
  XNOR U32138 ( .A(n32100), .B(n29409), .Z(n27025) );
  ANDN U32139 ( .B(n30058), .A(n30057), .Z(n32099) );
  XNOR U32140 ( .A(n32101), .B(n32102), .Z(n30057) );
  XOR U32141 ( .A(n32103), .B(n32104), .Z(n25513) );
  XNOR U32142 ( .A(n25233), .B(n26515), .Z(n32104) );
  XOR U32143 ( .A(n32105), .B(n28554), .Z(n26515) );
  XNOR U32144 ( .A(n32106), .B(n28744), .Z(n28554) );
  NOR U32145 ( .A(n28573), .B(n32107), .Z(n32105) );
  XNOR U32146 ( .A(n32108), .B(n27302), .Z(n25233) );
  XNOR U32147 ( .A(n32109), .B(n32110), .Z(n27302) );
  ANDN U32148 ( .B(n27303), .A(n32111), .Z(n32108) );
  XOR U32149 ( .A(n26909), .B(n32112), .Z(n32103) );
  XOR U32150 ( .A(n22630), .B(n24937), .Z(n32112) );
  XNOR U32151 ( .A(n32113), .B(n28558), .Z(n24937) );
  XNOR U32152 ( .A(n32114), .B(n31264), .Z(n28558) );
  NOR U32153 ( .A(n32115), .B(n27288), .Z(n32113) );
  XNOR U32154 ( .A(n32116), .B(n27293), .Z(n22630) );
  XOR U32155 ( .A(n32117), .B(n32118), .Z(n27293) );
  NOR U32156 ( .A(n32119), .B(n27292), .Z(n32116) );
  XOR U32157 ( .A(n32120), .B(n27298), .Z(n26909) );
  XOR U32158 ( .A(n32121), .B(n30959), .Z(n27298) );
  NOR U32159 ( .A(n32122), .B(n32123), .Z(n32120) );
  XOR U32160 ( .A(n32124), .B(n27447), .Z(n26933) );
  XOR U32161 ( .A(n32125), .B(n28723), .Z(n27447) );
  ANDN U32162 ( .B(n27020), .A(n32126), .Z(n32124) );
  XNOR U32163 ( .A(n25183), .B(n32127), .Z(n22874) );
  IV U32164 ( .A(n24455), .Z(n25183) );
  XNOR U32165 ( .A(n28302), .B(n29487), .Z(n24455) );
  XOR U32166 ( .A(n32128), .B(n32129), .Z(n29487) );
  XNOR U32167 ( .A(n25690), .B(n28297), .Z(n32129) );
  XNOR U32168 ( .A(n32130), .B(n30971), .Z(n28297) );
  XOR U32169 ( .A(n32131), .B(n32132), .Z(n30971) );
  NOR U32170 ( .A(n29631), .B(n30970), .Z(n32130) );
  XNOR U32171 ( .A(n32133), .B(n30975), .Z(n25690) );
  XNOR U32172 ( .A(n30149), .B(n32134), .Z(n30975) );
  XOR U32173 ( .A(n24602), .B(n32135), .Z(n32128) );
  XNOR U32174 ( .A(n30936), .B(n23583), .Z(n32135) );
  XNOR U32175 ( .A(n30968), .B(n32136), .Z(n23583) );
  XNOR U32176 ( .A(n11417), .B(n32137), .Z(n32136) );
  XNOR U32177 ( .A(n32138), .B(n32139), .Z(n30968) );
  XOR U32178 ( .A(n32140), .B(n30980), .Z(n30936) );
  IV U32179 ( .A(n31400), .Z(n30980) );
  XOR U32180 ( .A(n32141), .B(n32142), .Z(n31400) );
  NOR U32181 ( .A(n32143), .B(n30979), .Z(n32140) );
  XNOR U32182 ( .A(n32144), .B(n30983), .Z(n24602) );
  XNOR U32183 ( .A(n32145), .B(n29937), .Z(n30983) );
  NOR U32184 ( .A(n30982), .B(n29621), .Z(n32144) );
  XOR U32185 ( .A(n32146), .B(n32147), .Z(n28302) );
  XOR U32186 ( .A(n25924), .B(n26985), .Z(n32147) );
  XOR U32187 ( .A(n32148), .B(n31380), .Z(n26985) );
  XOR U32188 ( .A(n32149), .B(n30129), .Z(n31380) );
  NOR U32189 ( .A(n32150), .B(n29611), .Z(n32148) );
  XNOR U32190 ( .A(n32151), .B(n31386), .Z(n25924) );
  IV U32191 ( .A(n29671), .Z(n31386) );
  XNOR U32192 ( .A(n32152), .B(n29027), .Z(n29671) );
  ANDN U32193 ( .B(n29598), .A(n29670), .Z(n32151) );
  XNOR U32194 ( .A(n25095), .B(n32153), .Z(n32146) );
  XNOR U32195 ( .A(n23149), .B(n24576), .Z(n32153) );
  XNOR U32196 ( .A(n32154), .B(n29661), .Z(n24576) );
  XOR U32197 ( .A(n28803), .B(n32155), .Z(n29661) );
  ANDN U32198 ( .B(n29662), .A(n29607), .Z(n32154) );
  XOR U32199 ( .A(n32157), .B(n31178), .Z(n29664) );
  ANDN U32200 ( .B(n29602), .A(n32158), .Z(n32156) );
  IV U32201 ( .A(n29665), .Z(n32158) );
  XNOR U32202 ( .A(n32159), .B(n29673), .Z(n25095) );
  XOR U32203 ( .A(n32160), .B(n32161), .Z(n29673) );
  ANDN U32204 ( .B(n29615), .A(n29674), .Z(n32159) );
  XNOR U32205 ( .A(n32162), .B(n26388), .Z(n19437) );
  XNOR U32206 ( .A(n22635), .B(n26202), .Z(n26388) );
  XNOR U32207 ( .A(n32163), .B(n29774), .Z(n26202) );
  NOR U32208 ( .A(n32164), .B(n29235), .Z(n32163) );
  XNOR U32209 ( .A(n32165), .B(n32166), .Z(n29235) );
  XOR U32210 ( .A(n26778), .B(n26372), .Z(n22635) );
  XNOR U32211 ( .A(n32167), .B(n32168), .Z(n26372) );
  XOR U32212 ( .A(n23243), .B(n24918), .Z(n32168) );
  XNOR U32213 ( .A(n32169), .B(n29224), .Z(n24918) );
  XOR U32214 ( .A(n32170), .B(n27652), .Z(n29224) );
  NOR U32215 ( .A(n30780), .B(n28845), .Z(n32169) );
  XOR U32216 ( .A(n32171), .B(n29289), .Z(n28845) );
  IV U32217 ( .A(n32172), .Z(n29289) );
  IV U32218 ( .A(n28846), .Z(n30780) );
  XOR U32219 ( .A(n32173), .B(n30004), .Z(n28846) );
  IV U32220 ( .A(n28825), .Z(n30004) );
  XNOR U32221 ( .A(n32174), .B(n29226), .Z(n23243) );
  XOR U32222 ( .A(n32175), .B(n32176), .Z(n29226) );
  ANDN U32223 ( .B(n28856), .A(n28854), .Z(n32174) );
  XOR U32224 ( .A(n32177), .B(n29717), .Z(n28854) );
  IV U32225 ( .A(n30787), .Z(n28856) );
  XOR U32226 ( .A(n32178), .B(n31223), .Z(n30787) );
  XOR U32227 ( .A(n25207), .B(n32179), .Z(n32167) );
  XOR U32228 ( .A(n26878), .B(n24942), .Z(n32179) );
  XNOR U32229 ( .A(n32180), .B(n29219), .Z(n24942) );
  XNOR U32230 ( .A(n32181), .B(n32182), .Z(n29219) );
  ANDN U32231 ( .B(n28852), .A(n28850), .Z(n32180) );
  XOR U32232 ( .A(n30657), .B(n32183), .Z(n28850) );
  XNOR U32233 ( .A(n32184), .B(n32185), .Z(n30657) );
  XOR U32234 ( .A(n29045), .B(n32186), .Z(n28852) );
  XNOR U32235 ( .A(n32187), .B(n29371), .Z(n26878) );
  XNOR U32236 ( .A(n32188), .B(n32189), .Z(n29371) );
  NOR U32237 ( .A(n28842), .B(n28841), .Z(n32187) );
  XOR U32238 ( .A(n32190), .B(n32191), .Z(n28841) );
  XOR U32239 ( .A(n32192), .B(n32193), .Z(n28842) );
  XNOR U32240 ( .A(n32194), .B(n29766), .Z(n25207) );
  IV U32241 ( .A(n30756), .Z(n29766) );
  XOR U32242 ( .A(n32195), .B(n31164), .Z(n30756) );
  IV U32243 ( .A(n32196), .Z(n31164) );
  NOR U32244 ( .A(n28858), .B(n28859), .Z(n32194) );
  XNOR U32245 ( .A(n32197), .B(n30507), .Z(n28859) );
  XOR U32246 ( .A(n32198), .B(n30768), .Z(n28858) );
  XOR U32247 ( .A(n32199), .B(n32200), .Z(n26778) );
  XOR U32248 ( .A(n26689), .B(n26260), .Z(n32200) );
  XNOR U32249 ( .A(n32201), .B(n29240), .Z(n26260) );
  XOR U32250 ( .A(n32202), .B(n32203), .Z(n29240) );
  NOR U32251 ( .A(n26205), .B(n26204), .Z(n32201) );
  XNOR U32252 ( .A(n32204), .B(n32205), .Z(n26204) );
  XOR U32253 ( .A(n31137), .B(n32206), .Z(n26205) );
  XNOR U32254 ( .A(n32207), .B(n29247), .Z(n26689) );
  XOR U32255 ( .A(n32208), .B(n30223), .Z(n29247) );
  NOR U32256 ( .A(n26215), .B(n26214), .Z(n32207) );
  XNOR U32257 ( .A(n32209), .B(n30258), .Z(n26214) );
  XOR U32258 ( .A(n32210), .B(n32211), .Z(n30258) );
  XOR U32259 ( .A(n32212), .B(n31566), .Z(n26215) );
  XNOR U32260 ( .A(n24794), .B(n32213), .Z(n32199) );
  XNOR U32261 ( .A(n23078), .B(n29756), .Z(n32213) );
  XNOR U32262 ( .A(n32214), .B(n29232), .Z(n29756) );
  XOR U32263 ( .A(n32215), .B(n32216), .Z(n29232) );
  NOR U32264 ( .A(n30016), .B(n29776), .Z(n32214) );
  XOR U32265 ( .A(n32217), .B(n31289), .Z(n29776) );
  IV U32266 ( .A(n31687), .Z(n31289) );
  XOR U32267 ( .A(n32218), .B(n31855), .Z(n30016) );
  XOR U32268 ( .A(n32219), .B(n29243), .Z(n23078) );
  XNOR U32269 ( .A(n32220), .B(n30507), .Z(n29243) );
  ANDN U32270 ( .B(n26212), .A(n26210), .Z(n32219) );
  XOR U32271 ( .A(n32221), .B(n30252), .Z(n26210) );
  XOR U32272 ( .A(n30483), .B(n32222), .Z(n26212) );
  XNOR U32273 ( .A(n32223), .B(n29236), .Z(n24794) );
  XOR U32274 ( .A(n32224), .B(n32225), .Z(n29236) );
  NOR U32275 ( .A(n31829), .B(n29774), .Z(n32223) );
  XOR U32276 ( .A(n32226), .B(n32044), .Z(n29774) );
  IV U32277 ( .A(n32164), .Z(n31829) );
  XNOR U32278 ( .A(n28803), .B(n32227), .Z(n32164) );
  ANDN U32279 ( .B(n21867), .A(n24329), .Z(n32162) );
  XNOR U32280 ( .A(n29629), .B(n22621), .Z(n24329) );
  XNOR U32281 ( .A(n25888), .B(n26883), .Z(n22621) );
  XNOR U32282 ( .A(n32228), .B(n32229), .Z(n26883) );
  XOR U32283 ( .A(n24708), .B(n25033), .Z(n32229) );
  XOR U32284 ( .A(n32230), .B(n29496), .Z(n25033) );
  XOR U32285 ( .A(n32231), .B(n29032), .Z(n29496) );
  ANDN U32286 ( .B(n28449), .A(n28165), .Z(n32230) );
  XOR U32287 ( .A(n32232), .B(n32233), .Z(n28165) );
  XOR U32288 ( .A(n32234), .B(n28759), .Z(n28449) );
  IV U32289 ( .A(n32235), .Z(n28759) );
  XNOR U32290 ( .A(n32236), .B(n29498), .Z(n24708) );
  XOR U32291 ( .A(n32237), .B(n31598), .Z(n29498) );
  NOR U32292 ( .A(n28442), .B(n28443), .Z(n32236) );
  XOR U32293 ( .A(n32238), .B(n29057), .Z(n28443) );
  XNOR U32294 ( .A(n32239), .B(n32240), .Z(n29057) );
  XOR U32295 ( .A(n32241), .B(n29050), .Z(n28442) );
  XOR U32296 ( .A(n24716), .B(n32242), .Z(n32228) );
  XOR U32297 ( .A(n28752), .B(n23982), .Z(n32242) );
  XNOR U32298 ( .A(n32243), .B(n30954), .Z(n23982) );
  IV U32299 ( .A(n29493), .Z(n30954) );
  XOR U32300 ( .A(n28987), .B(n32244), .Z(n29493) );
  IV U32301 ( .A(n32245), .Z(n28987) );
  ANDN U32302 ( .B(n26833), .A(n28440), .Z(n32243) );
  XOR U32303 ( .A(n32246), .B(n32205), .Z(n28440) );
  XOR U32304 ( .A(n32247), .B(n32248), .Z(n26833) );
  XNOR U32305 ( .A(n32249), .B(n29500), .Z(n28752) );
  XNOR U32306 ( .A(n32250), .B(n32251), .Z(n29500) );
  AND U32307 ( .A(n28447), .B(n26826), .Z(n32249) );
  XOR U32308 ( .A(n32252), .B(n31794), .Z(n26826) );
  XOR U32309 ( .A(n32253), .B(n31355), .Z(n28447) );
  XNOR U32310 ( .A(n32254), .B(n30960), .Z(n24716) );
  IV U32311 ( .A(n29491), .Z(n30960) );
  XNOR U32312 ( .A(n32255), .B(n28887), .Z(n29491) );
  NOR U32313 ( .A(n28451), .B(n27332), .Z(n32254) );
  XOR U32314 ( .A(n32258), .B(n31229), .Z(n27332) );
  XOR U32315 ( .A(n32259), .B(n30204), .Z(n28451) );
  XNOR U32316 ( .A(n32260), .B(n32261), .Z(n25888) );
  XNOR U32317 ( .A(n23336), .B(n24645), .Z(n32261) );
  XOR U32318 ( .A(n32262), .B(n30976), .Z(n24645) );
  XNOR U32319 ( .A(n32263), .B(n31654), .Z(n30976) );
  ANDN U32320 ( .B(n29635), .A(n29636), .Z(n32262) );
  XNOR U32321 ( .A(n29968), .B(n32264), .Z(n29636) );
  XOR U32322 ( .A(n32265), .B(n32266), .Z(n29635) );
  XNOR U32323 ( .A(n32267), .B(n30966), .Z(n23336) );
  XOR U32324 ( .A(n32268), .B(n32269), .Z(n30966) );
  NOR U32325 ( .A(n29625), .B(n29626), .Z(n32267) );
  XOR U32326 ( .A(n32175), .B(n32270), .Z(n29626) );
  XNOR U32327 ( .A(n29324), .B(n32271), .Z(n29625) );
  XNOR U32328 ( .A(n24259), .B(n32272), .Z(n32260) );
  XNOR U32329 ( .A(n29486), .B(n25660), .Z(n32272) );
  XNOR U32330 ( .A(n32273), .B(n30970), .Z(n25660) );
  XOR U32331 ( .A(n32274), .B(n32275), .Z(n30970) );
  ANDN U32332 ( .B(n29631), .A(n29632), .Z(n32273) );
  XOR U32333 ( .A(n32276), .B(n31240), .Z(n29632) );
  XOR U32334 ( .A(n32277), .B(n30514), .Z(n29631) );
  XNOR U32335 ( .A(n32278), .B(n30979), .Z(n29486) );
  XNOR U32336 ( .A(n29959), .B(n32279), .Z(n30979) );
  ANDN U32337 ( .B(n32143), .A(n31399), .Z(n32278) );
  XNOR U32338 ( .A(n32280), .B(n30982), .Z(n24259) );
  XOR U32339 ( .A(n32281), .B(n32018), .Z(n30982) );
  ANDN U32340 ( .B(n29621), .A(n31410), .Z(n32280) );
  IV U32341 ( .A(n29623), .Z(n31410) );
  XOR U32342 ( .A(n32282), .B(n30687), .Z(n29623) );
  XNOR U32343 ( .A(n30860), .B(n32283), .Z(n29621) );
  XNOR U32344 ( .A(n32284), .B(n32143), .Z(n29629) );
  XNOR U32345 ( .A(n31642), .B(n32285), .Z(n32143) );
  ANDN U32346 ( .B(n31399), .A(n30978), .Z(n32284) );
  XOR U32347 ( .A(n32286), .B(n30941), .Z(n30978) );
  IV U32348 ( .A(n30752), .Z(n30941) );
  XOR U32349 ( .A(n32287), .B(n28875), .Z(n31399) );
  XNOR U32350 ( .A(n27042), .B(n25706), .Z(n21867) );
  XNOR U32351 ( .A(n32288), .B(n32289), .Z(n29134) );
  XOR U32352 ( .A(n25668), .B(n26819), .Z(n32289) );
  XOR U32353 ( .A(n32290), .B(n28974), .Z(n26819) );
  XOR U32354 ( .A(n32291), .B(n29095), .Z(n28974) );
  XOR U32355 ( .A(n32292), .B(n26959), .Z(n25668) );
  XOR U32356 ( .A(n29178), .B(n32293), .Z(n26959) );
  IV U32357 ( .A(n31238), .Z(n29178) );
  AND U32358 ( .A(n26958), .B(n27041), .Z(n32292) );
  XNOR U32359 ( .A(n32294), .B(n31185), .Z(n27041) );
  XOR U32360 ( .A(n31026), .B(n32295), .Z(n26958) );
  XNOR U32361 ( .A(n26951), .B(n32296), .Z(n32288) );
  XNOR U32362 ( .A(n25438), .B(n24557), .Z(n32296) );
  XNOR U32363 ( .A(n32297), .B(n26964), .Z(n24557) );
  XNOR U32364 ( .A(n32298), .B(n32299), .Z(n26964) );
  AND U32365 ( .A(n26963), .B(n27046), .Z(n32297) );
  XNOR U32366 ( .A(n32300), .B(n32301), .Z(n27046) );
  XOR U32367 ( .A(n32302), .B(n32303), .Z(n26963) );
  XNOR U32368 ( .A(n32304), .B(n26968), .Z(n25438) );
  XOR U32369 ( .A(n30852), .B(n32305), .Z(n26968) );
  NOR U32370 ( .A(n31331), .B(n26967), .Z(n32304) );
  XOR U32371 ( .A(n32306), .B(n32307), .Z(n26967) );
  XOR U32372 ( .A(n32308), .B(n32309), .Z(n31331) );
  XNOR U32373 ( .A(n32310), .B(n26972), .Z(n26951) );
  XNOR U32374 ( .A(n32311), .B(n31022), .Z(n26972) );
  ANDN U32375 ( .B(n30156), .A(n26971), .Z(n32310) );
  XOR U32376 ( .A(n32312), .B(n32313), .Z(n26971) );
  XOR U32377 ( .A(n32314), .B(n32315), .Z(n30156) );
  XNOR U32378 ( .A(n32317), .B(n28975), .Z(n27042) );
  XNOR U32379 ( .A(n29396), .B(n32318), .Z(n28975) );
  ANDN U32380 ( .B(n31343), .A(n31342), .Z(n32317) );
  XOR U32381 ( .A(n29965), .B(n32319), .Z(n31342) );
  IV U32382 ( .A(n31374), .Z(n31343) );
  XOR U32383 ( .A(n32320), .B(n32182), .Z(n31374) );
  XNOR U32384 ( .A(n32321), .B(n26444), .Z(n19357) );
  XOR U32385 ( .A(n32322), .B(n24825), .Z(n26444) );
  XNOR U32386 ( .A(n27954), .B(n30934), .Z(n24825) );
  XNOR U32387 ( .A(n32323), .B(n32324), .Z(n30934) );
  XNOR U32388 ( .A(n25773), .B(n25017), .Z(n32324) );
  XNOR U32389 ( .A(n32325), .B(n30442), .Z(n25017) );
  ANDN U32390 ( .B(n32326), .A(n32327), .Z(n32325) );
  XNOR U32391 ( .A(n32328), .B(n30456), .Z(n25773) );
  ANDN U32392 ( .B(n30457), .A(n31510), .Z(n32328) );
  XNOR U32393 ( .A(n30437), .B(n32329), .Z(n32323) );
  XNOR U32394 ( .A(n23687), .B(n28010), .Z(n32329) );
  XNOR U32395 ( .A(n32330), .B(n30638), .Z(n28010) );
  ANDN U32396 ( .B(n30639), .A(n31514), .Z(n32330) );
  XOR U32397 ( .A(n32331), .B(n30446), .Z(n23687) );
  ANDN U32398 ( .B(n30447), .A(n31502), .Z(n32331) );
  XOR U32399 ( .A(n32332), .B(n30452), .Z(n30437) );
  ANDN U32400 ( .B(n30453), .A(n31505), .Z(n32332) );
  XOR U32401 ( .A(n32333), .B(n32334), .Z(n27954) );
  XNOR U32402 ( .A(n26949), .B(n25214), .Z(n32334) );
  XNOR U32403 ( .A(n32335), .B(n30472), .Z(n25214) );
  XOR U32404 ( .A(n32336), .B(n30539), .Z(n30472) );
  ANDN U32405 ( .B(n30473), .A(n30086), .Z(n32335) );
  XNOR U32406 ( .A(n32337), .B(n30476), .Z(n26949) );
  XNOR U32407 ( .A(n32338), .B(n28821), .Z(n30476) );
  ANDN U32408 ( .B(n30477), .A(n30091), .Z(n32337) );
  XNOR U32409 ( .A(n27073), .B(n32339), .Z(n32333) );
  XNOR U32410 ( .A(n23814), .B(n25498), .Z(n32339) );
  XNOR U32411 ( .A(n32340), .B(n30466), .Z(n25498) );
  XNOR U32412 ( .A(n32341), .B(n30371), .Z(n30466) );
  NOR U32413 ( .A(n30099), .B(n30465), .Z(n32340) );
  XNOR U32414 ( .A(n32342), .B(n30470), .Z(n23814) );
  XOR U32415 ( .A(n32343), .B(n28744), .Z(n30470) );
  ANDN U32416 ( .B(n30082), .A(n30469), .Z(n32342) );
  XNOR U32417 ( .A(n32344), .B(n30462), .Z(n27073) );
  XOR U32418 ( .A(n31844), .B(n32345), .Z(n30462) );
  ANDN U32419 ( .B(n30463), .A(n30095), .Z(n32344) );
  ANDN U32420 ( .B(n21871), .A(n24331), .Z(n32321) );
  IV U32421 ( .A(n25396), .Z(n24331) );
  XOR U32422 ( .A(n30813), .B(n24275), .Z(n25396) );
  XOR U32423 ( .A(n32346), .B(n27071), .Z(n24275) );
  XNOR U32424 ( .A(n32347), .B(n32348), .Z(n27071) );
  XOR U32425 ( .A(n24022), .B(n22612), .Z(n32348) );
  XNOR U32426 ( .A(n32349), .B(n26175), .Z(n22612) );
  XOR U32427 ( .A(n32350), .B(n29067), .Z(n26175) );
  ANDN U32428 ( .B(n26176), .A(n30810), .Z(n32349) );
  XOR U32429 ( .A(n32351), .B(n30198), .Z(n30810) );
  XOR U32430 ( .A(n32352), .B(n29922), .Z(n26176) );
  XOR U32431 ( .A(n32353), .B(n30035), .Z(n24022) );
  IV U32432 ( .A(n26168), .Z(n30035) );
  XOR U32433 ( .A(n32354), .B(n31434), .Z(n26168) );
  NOR U32434 ( .A(n26167), .B(n29008), .Z(n32353) );
  XOR U32435 ( .A(n30253), .B(n32355), .Z(n29008) );
  XNOR U32436 ( .A(n32356), .B(n31642), .Z(n26167) );
  XOR U32437 ( .A(n25404), .B(n32357), .Z(n32347) );
  XOR U32438 ( .A(n26152), .B(n25507), .Z(n32357) );
  XOR U32439 ( .A(n32358), .B(n26158), .Z(n25507) );
  XOR U32440 ( .A(n32359), .B(n32360), .Z(n26158) );
  XNOR U32441 ( .A(n32361), .B(n26172), .Z(n26152) );
  XOR U32442 ( .A(n32362), .B(n32363), .Z(n26172) );
  NOR U32443 ( .A(n29000), .B(n26171), .Z(n32361) );
  XOR U32444 ( .A(n31982), .B(n32364), .Z(n26171) );
  IV U32445 ( .A(n32175), .Z(n31982) );
  XOR U32446 ( .A(n32365), .B(n32366), .Z(n29000) );
  XOR U32447 ( .A(n32367), .B(n26162), .Z(n25404) );
  XOR U32448 ( .A(n32368), .B(n32369), .Z(n26162) );
  ANDN U32449 ( .B(n26163), .A(n30820), .Z(n32367) );
  XNOR U32450 ( .A(n32274), .B(n32370), .Z(n30820) );
  XOR U32451 ( .A(n32371), .B(n31255), .Z(n26163) );
  IV U32452 ( .A(n30277), .Z(n31255) );
  XOR U32453 ( .A(n32372), .B(n32373), .Z(n30277) );
  XOR U32454 ( .A(n32374), .B(n26159), .Z(n30813) );
  XOR U32455 ( .A(n32375), .B(n29097), .Z(n26159) );
  IV U32456 ( .A(n32376), .Z(n29097) );
  IV U32457 ( .A(n29012), .Z(n30032) );
  XOR U32458 ( .A(n32377), .B(n28435), .Z(n29012) );
  XNOR U32459 ( .A(n32378), .B(n30573), .Z(n29011) );
  XNOR U32460 ( .A(n32379), .B(n32380), .Z(n30573) );
  XNOR U32461 ( .A(n26798), .B(n24998), .Z(n21871) );
  XNOR U32462 ( .A(n27166), .B(n26506), .Z(n24998) );
  XNOR U32463 ( .A(n32381), .B(n32382), .Z(n26506) );
  XOR U32464 ( .A(n24759), .B(n25440), .Z(n32382) );
  XNOR U32465 ( .A(n32383), .B(n27501), .Z(n25440) );
  XNOR U32466 ( .A(n32384), .B(n30204), .Z(n27501) );
  IV U32467 ( .A(n32132), .Z(n30204) );
  XOR U32468 ( .A(n32385), .B(n32386), .Z(n32132) );
  ANDN U32469 ( .B(n28393), .A(n28394), .Z(n32383) );
  XNOR U32470 ( .A(n31947), .B(n32387), .Z(n28393) );
  XOR U32471 ( .A(n32388), .B(n27491), .Z(n24759) );
  XOR U32472 ( .A(n32389), .B(n32390), .Z(n27491) );
  AND U32473 ( .A(n28387), .B(n28386), .Z(n32388) );
  XOR U32474 ( .A(n32391), .B(n31454), .Z(n28386) );
  XOR U32475 ( .A(n24768), .B(n32392), .Z(n32381) );
  XNOR U32476 ( .A(n22393), .B(n29501), .Z(n32392) );
  XNOR U32477 ( .A(n32393), .B(n27495), .Z(n29501) );
  XOR U32478 ( .A(n32394), .B(n32395), .Z(n27495) );
  ANDN U32479 ( .B(n28384), .A(n28383), .Z(n32393) );
  XOR U32480 ( .A(n32396), .B(n31348), .Z(n28383) );
  XOR U32481 ( .A(n32397), .B(n27504), .Z(n22393) );
  XOR U32482 ( .A(n32398), .B(n32315), .Z(n27504) );
  NOR U32483 ( .A(n28390), .B(n28391), .Z(n32397) );
  XOR U32484 ( .A(n32399), .B(n31858), .Z(n28390) );
  XNOR U32485 ( .A(n32400), .B(n27508), .Z(n24768) );
  XOR U32486 ( .A(n32401), .B(n32402), .Z(n27508) );
  ANDN U32487 ( .B(n28397), .A(n28396), .Z(n32400) );
  XOR U32488 ( .A(n32403), .B(n30956), .Z(n28396) );
  XOR U32489 ( .A(n32404), .B(n32405), .Z(n27166) );
  XNOR U32490 ( .A(n23509), .B(n26811), .Z(n32405) );
  XOR U32491 ( .A(n32406), .B(n28141), .Z(n26811) );
  XOR U32492 ( .A(n32407), .B(n31169), .Z(n28141) );
  XNOR U32493 ( .A(n32409), .B(n28144), .Z(n23509) );
  NOR U32494 ( .A(n26800), .B(n26801), .Z(n32409) );
  XOR U32495 ( .A(n32410), .B(n32411), .Z(n26800) );
  XNOR U32496 ( .A(n25983), .B(n32412), .Z(n32404) );
  XOR U32497 ( .A(n26663), .B(n25889), .Z(n32412) );
  XNOR U32498 ( .A(n32413), .B(n28149), .Z(n25889) );
  XOR U32499 ( .A(n32414), .B(n29175), .Z(n28149) );
  IV U32500 ( .A(n32415), .Z(n29175) );
  NOR U32501 ( .A(n28148), .B(n31519), .Z(n32413) );
  IV U32502 ( .A(n31518), .Z(n28148) );
  XNOR U32503 ( .A(n32416), .B(n30535), .Z(n31518) );
  XOR U32504 ( .A(n32417), .B(n28152), .Z(n26663) );
  XOR U32505 ( .A(n29396), .B(n32418), .Z(n28152) );
  XNOR U32506 ( .A(n32419), .B(n32184), .Z(n29396) );
  XOR U32507 ( .A(n32420), .B(n32421), .Z(n32184) );
  XOR U32508 ( .A(n32422), .B(n31928), .Z(n32421) );
  XOR U32509 ( .A(n32423), .B(n32424), .Z(n31928) );
  ANDN U32510 ( .B(n32425), .A(n32426), .Z(n32423) );
  XNOR U32511 ( .A(n32427), .B(n32428), .Z(n32420) );
  XNOR U32512 ( .A(n32429), .B(n31656), .Z(n32428) );
  XNOR U32513 ( .A(n32430), .B(n32431), .Z(n31656) );
  ANDN U32514 ( .B(n32432), .A(n32433), .Z(n32430) );
  XOR U32515 ( .A(n32434), .B(n31674), .Z(n26807) );
  XNOR U32516 ( .A(n32435), .B(n28156), .Z(n25983) );
  XOR U32517 ( .A(n32436), .B(n31068), .Z(n28156) );
  NOR U32518 ( .A(n28728), .B(n28729), .Z(n32435) );
  IV U32519 ( .A(n28155), .Z(n28728) );
  XOR U32520 ( .A(n32437), .B(n31632), .Z(n28155) );
  XNOR U32521 ( .A(n32438), .B(n28140), .Z(n26798) );
  XOR U32522 ( .A(n32439), .B(n31998), .Z(n28140) );
  IV U32523 ( .A(n30959), .Z(n31998) );
  ANDN U32524 ( .B(n32408), .A(n28239), .Z(n32438) );
  XNOR U32525 ( .A(n25905), .B(n17853), .Z(n13492) );
  XOR U32526 ( .A(n23805), .B(n21383), .Z(n17853) );
  XOR U32527 ( .A(n32440), .B(n32441), .Z(n21383) );
  XNOR U32528 ( .A(n17238), .B(n20147), .Z(n32441) );
  XNOR U32529 ( .A(n32442), .B(n23466), .Z(n20147) );
  XOR U32530 ( .A(n25490), .B(n31531), .Z(n23466) );
  XNOR U32531 ( .A(n32443), .B(n31859), .Z(n31531) );
  NOR U32532 ( .A(n31197), .B(n30352), .Z(n32443) );
  XOR U32533 ( .A(n30869), .B(n32444), .Z(n30352) );
  XNOR U32534 ( .A(n32445), .B(n32446), .Z(n26703) );
  XNOR U32535 ( .A(n31850), .B(n24517), .Z(n32446) );
  XNOR U32536 ( .A(n32447), .B(n30345), .Z(n24517) );
  XNOR U32537 ( .A(n29736), .B(n32448), .Z(n30345) );
  AND U32538 ( .A(n31203), .B(n31537), .Z(n32447) );
  XOR U32539 ( .A(n32449), .B(n32450), .Z(n31537) );
  XNOR U32540 ( .A(n32451), .B(n32452), .Z(n31203) );
  XNOR U32541 ( .A(n32453), .B(n30341), .Z(n31850) );
  XOR U32542 ( .A(n32454), .B(n31598), .Z(n30341) );
  ANDN U32543 ( .B(n31533), .A(n31199), .Z(n32453) );
  XNOR U32544 ( .A(n32455), .B(n32456), .Z(n31199) );
  XOR U32545 ( .A(n32457), .B(n31154), .Z(n31533) );
  XOR U32546 ( .A(n26067), .B(n32458), .Z(n32445) );
  XOR U32547 ( .A(n27233), .B(n25807), .Z(n32458) );
  XNOR U32548 ( .A(n32459), .B(n30358), .Z(n25807) );
  XNOR U32549 ( .A(n30000), .B(n32460), .Z(n30358) );
  XOR U32550 ( .A(n32210), .B(n32461), .Z(n30000) );
  XOR U32551 ( .A(n32462), .B(n32463), .Z(n32210) );
  XNOR U32552 ( .A(n31061), .B(n32464), .Z(n32463) );
  XNOR U32553 ( .A(n32465), .B(n32466), .Z(n31061) );
  NOR U32554 ( .A(n32467), .B(n32468), .Z(n32465) );
  XOR U32555 ( .A(n28889), .B(n32469), .Z(n32462) );
  XOR U32556 ( .A(n30916), .B(n32470), .Z(n32469) );
  XNOR U32557 ( .A(n32471), .B(n32472), .Z(n30916) );
  ANDN U32558 ( .B(n32473), .A(n32474), .Z(n32471) );
  XNOR U32559 ( .A(n32475), .B(n32476), .Z(n28889) );
  NOR U32560 ( .A(n32477), .B(n32478), .Z(n32475) );
  ANDN U32561 ( .B(n31528), .A(n31324), .Z(n32459) );
  XOR U32562 ( .A(n32479), .B(n32000), .Z(n31324) );
  XNOR U32563 ( .A(n32480), .B(n32481), .Z(n31528) );
  XOR U32564 ( .A(n32482), .B(n30354), .Z(n27233) );
  XOR U32565 ( .A(n32483), .B(n32415), .Z(n30354) );
  XOR U32566 ( .A(n30247), .B(n32484), .Z(n31197) );
  XOR U32567 ( .A(n32485), .B(n31314), .Z(n31859) );
  XNOR U32568 ( .A(n32486), .B(n30350), .Z(n26067) );
  XOR U32569 ( .A(n32487), .B(n28723), .Z(n30350) );
  IV U32570 ( .A(n31369), .Z(n28723) );
  NOR U32571 ( .A(n31205), .B(n31525), .Z(n32486) );
  XOR U32572 ( .A(n32193), .B(n32488), .Z(n31525) );
  XNOR U32573 ( .A(n32489), .B(n28897), .Z(n31205) );
  XOR U32574 ( .A(n32490), .B(n32491), .Z(n28652) );
  XOR U32575 ( .A(n25351), .B(n30984), .Z(n32491) );
  XOR U32576 ( .A(n32492), .B(n28085), .Z(n30984) );
  XNOR U32577 ( .A(n29736), .B(n32493), .Z(n28085) );
  ANDN U32578 ( .B(n31319), .A(n29784), .Z(n32492) );
  IV U32579 ( .A(n31320), .Z(n29784) );
  XOR U32580 ( .A(n32376), .B(n32494), .Z(n31320) );
  XNOR U32581 ( .A(n30231), .B(n32495), .Z(n31319) );
  XNOR U32582 ( .A(n32496), .B(n28075), .Z(n25351) );
  XNOR U32583 ( .A(n32497), .B(n32498), .Z(n28075) );
  ANDN U32584 ( .B(n31304), .A(n29795), .Z(n32496) );
  XNOR U32585 ( .A(n32499), .B(n29295), .Z(n29795) );
  IV U32586 ( .A(n32006), .Z(n29295) );
  XNOR U32587 ( .A(n32500), .B(n30252), .Z(n31304) );
  IV U32588 ( .A(n31030), .Z(n30252) );
  XOR U32589 ( .A(n26872), .B(n32503), .Z(n32490) );
  XOR U32590 ( .A(n25025), .B(n30805), .Z(n32503) );
  XOR U32591 ( .A(n32504), .B(n28080), .Z(n30805) );
  XOR U32592 ( .A(n32505), .B(n31855), .Z(n28080) );
  ANDN U32593 ( .B(n31316), .A(n29792), .Z(n32504) );
  XOR U32594 ( .A(n32506), .B(n29413), .Z(n29792) );
  XOR U32595 ( .A(n32109), .B(n32507), .Z(n31316) );
  XOR U32596 ( .A(n32509), .B(n28836), .Z(n28072) );
  ANDN U32597 ( .B(n31307), .A(n29789), .Z(n32508) );
  XNOR U32598 ( .A(n32510), .B(n32511), .Z(n29789) );
  XOR U32599 ( .A(n32512), .B(n31707), .Z(n31307) );
  XOR U32600 ( .A(n32513), .B(n28088), .Z(n26872) );
  XNOR U32601 ( .A(n32514), .B(n29409), .Z(n28088) );
  ANDN U32602 ( .B(n31312), .A(n31311), .Z(n32513) );
  XOR U32603 ( .A(n32515), .B(n30215), .Z(n31311) );
  IV U32604 ( .A(n29786), .Z(n31312) );
  XOR U32605 ( .A(n32516), .B(n32189), .Z(n29786) );
  IV U32606 ( .A(n31894), .Z(n32189) );
  XNOR U32607 ( .A(n32517), .B(n23457), .Z(n17238) );
  XOR U32608 ( .A(n24632), .B(n27811), .Z(n23457) );
  XNOR U32609 ( .A(n32518), .B(n32519), .Z(n27811) );
  NOR U32610 ( .A(n32520), .B(n27521), .Z(n32518) );
  IV U32611 ( .A(n24596), .Z(n24632) );
  XOR U32612 ( .A(n26910), .B(n31645), .Z(n24596) );
  XNOR U32613 ( .A(n32521), .B(n32522), .Z(n31645) );
  XNOR U32614 ( .A(n25264), .B(n27777), .Z(n32522) );
  XOR U32615 ( .A(n32523), .B(n27619), .Z(n27777) );
  XOR U32616 ( .A(n32524), .B(n30075), .Z(n27619) );
  ANDN U32617 ( .B(n27782), .A(n27808), .Z(n32523) );
  XOR U32618 ( .A(n32525), .B(n28469), .Z(n27808) );
  XNOR U32619 ( .A(n32526), .B(n30567), .Z(n27782) );
  IV U32620 ( .A(n29055), .Z(n30567) );
  XOR U32621 ( .A(n32527), .B(n32528), .Z(n29055) );
  XNOR U32622 ( .A(n32529), .B(n27628), .Z(n25264) );
  XOR U32623 ( .A(n32530), .B(n32531), .Z(n27628) );
  ANDN U32624 ( .B(n27784), .A(n27927), .Z(n32529) );
  XNOR U32625 ( .A(n30148), .B(n32532), .Z(n27927) );
  XNOR U32626 ( .A(n32533), .B(n30078), .Z(n27784) );
  XOR U32627 ( .A(n32534), .B(n32535), .Z(n30078) );
  XOR U32628 ( .A(n24988), .B(n32536), .Z(n32521) );
  XOR U32629 ( .A(n26757), .B(n26187), .Z(n32536) );
  XOR U32630 ( .A(n32537), .B(n27635), .Z(n26187) );
  XOR U32631 ( .A(n32538), .B(n32539), .Z(n27635) );
  ANDN U32632 ( .B(n27787), .A(n27806), .Z(n32537) );
  XNOR U32633 ( .A(n28995), .B(n32540), .Z(n27806) );
  XOR U32634 ( .A(n30491), .B(n32541), .Z(n27787) );
  XOR U32635 ( .A(n32543), .B(n29401), .Z(n27622) );
  IV U32636 ( .A(n30112), .Z(n29401) );
  XNOR U32637 ( .A(n32544), .B(n32545), .Z(n30112) );
  NOR U32638 ( .A(n27802), .B(n27791), .Z(n32542) );
  XOR U32639 ( .A(n32546), .B(n30014), .Z(n27791) );
  XNOR U32640 ( .A(n32547), .B(n29262), .Z(n27802) );
  XOR U32641 ( .A(n32548), .B(n27631), .Z(n24988) );
  XNOR U32642 ( .A(n32549), .B(n30733), .Z(n27631) );
  XOR U32643 ( .A(n32550), .B(n32551), .Z(n30733) );
  ANDN U32644 ( .B(n27789), .A(n29751), .Z(n32548) );
  XNOR U32645 ( .A(n32552), .B(n31654), .Z(n29751) );
  XOR U32646 ( .A(n32553), .B(n30651), .Z(n27789) );
  XOR U32647 ( .A(n32554), .B(n32555), .Z(n26910) );
  XNOR U32648 ( .A(n26340), .B(n25159), .Z(n32555) );
  XNOR U32649 ( .A(n32556), .B(n27523), .Z(n25159) );
  XOR U32650 ( .A(n32557), .B(n31654), .Z(n27523) );
  ANDN U32651 ( .B(n32520), .A(n28570), .Z(n32556) );
  IV U32652 ( .A(n32519), .Z(n28570) );
  XNOR U32653 ( .A(n32558), .B(n31264), .Z(n32519) );
  XNOR U32654 ( .A(n32559), .B(n27951), .Z(n26340) );
  XOR U32655 ( .A(n32117), .B(n32560), .Z(n27951) );
  AND U32656 ( .A(n27815), .B(n27813), .Z(n32559) );
  XNOR U32657 ( .A(n32561), .B(n30129), .Z(n27813) );
  XOR U32658 ( .A(n24452), .B(n32562), .Z(n32554) );
  XOR U32659 ( .A(n25755), .B(n25110), .Z(n32562) );
  XOR U32660 ( .A(n32563), .B(n27528), .Z(n25110) );
  XOR U32661 ( .A(n32564), .B(n29722), .Z(n27528) );
  XNOR U32662 ( .A(n31613), .B(n32565), .Z(n27824) );
  XNOR U32663 ( .A(n32566), .B(n27518), .Z(n25755) );
  XOR U32664 ( .A(n32567), .B(n27652), .Z(n27518) );
  IV U32665 ( .A(n31035), .Z(n27652) );
  XOR U32666 ( .A(n32568), .B(n32299), .Z(n27821) );
  XNOR U32667 ( .A(n32569), .B(n27532), .Z(n24452) );
  XNOR U32668 ( .A(n32570), .B(n31159), .Z(n27532) );
  ANDN U32669 ( .B(n27819), .A(n28566), .Z(n32569) );
  XOR U32670 ( .A(n32571), .B(n32572), .Z(n28566) );
  AND U32671 ( .A(n25910), .B(n23458), .Z(n32517) );
  XOR U32672 ( .A(n24963), .B(n30403), .Z(n23458) );
  XNOR U32673 ( .A(n32573), .B(n30891), .Z(n30403) );
  ANDN U32674 ( .B(n29188), .A(n32574), .Z(n32573) );
  IV U32675 ( .A(n25928), .Z(n24963) );
  XOR U32676 ( .A(n32019), .B(n27031), .Z(n25928) );
  XNOR U32677 ( .A(n32575), .B(n32576), .Z(n27031) );
  XOR U32678 ( .A(n25550), .B(n27896), .Z(n32576) );
  XOR U32679 ( .A(n32577), .B(n28295), .Z(n27896) );
  XNOR U32680 ( .A(n32578), .B(n30500), .Z(n28295) );
  ANDN U32681 ( .B(n30422), .A(n31464), .Z(n32577) );
  IV U32682 ( .A(n30423), .Z(n31464) );
  XNOR U32683 ( .A(n32579), .B(n30275), .Z(n30423) );
  XOR U32684 ( .A(n32580), .B(n28895), .Z(n30422) );
  XNOR U32685 ( .A(n32581), .B(n26650), .Z(n25550) );
  XNOR U32686 ( .A(n32582), .B(n32583), .Z(n26650) );
  ANDN U32687 ( .B(n30430), .A(n30883), .Z(n32581) );
  XOR U32688 ( .A(n32584), .B(n32585), .Z(n30883) );
  XNOR U32689 ( .A(n32586), .B(n32587), .Z(n30430) );
  XOR U32690 ( .A(n24869), .B(n32588), .Z(n32575) );
  XOR U32691 ( .A(n25015), .B(n22535), .Z(n32588) );
  XOR U32692 ( .A(n32589), .B(n26662), .Z(n22535) );
  XOR U32693 ( .A(n30946), .B(n32590), .Z(n26662) );
  AND U32694 ( .A(n30436), .B(n30435), .Z(n32589) );
  XOR U32695 ( .A(n28790), .B(n32591), .Z(n30435) );
  XOR U32696 ( .A(n32592), .B(n28425), .Z(n30436) );
  XOR U32697 ( .A(n32593), .B(n26655), .Z(n25015) );
  XNOR U32698 ( .A(n30264), .B(n32594), .Z(n26655) );
  IV U32699 ( .A(n32595), .Z(n30264) );
  ANDN U32700 ( .B(n30432), .A(n31469), .Z(n32593) );
  IV U32701 ( .A(n30433), .Z(n31469) );
  XOR U32702 ( .A(n32596), .B(n31894), .Z(n30433) );
  XOR U32703 ( .A(n32597), .B(n31820), .Z(n30432) );
  XNOR U32704 ( .A(n32598), .B(n30880), .Z(n24869) );
  IV U32705 ( .A(n28065), .Z(n30880) );
  XNOR U32706 ( .A(n29271), .B(n32599), .Z(n28065) );
  ANDN U32707 ( .B(n30425), .A(n31458), .Z(n32598) );
  IV U32708 ( .A(n30426), .Z(n31458) );
  XOR U32709 ( .A(n32308), .B(n32600), .Z(n30426) );
  XOR U32710 ( .A(n32601), .B(n30790), .Z(n30425) );
  IV U32711 ( .A(n32602), .Z(n30790) );
  XOR U32712 ( .A(n32603), .B(n32604), .Z(n32019) );
  XOR U32713 ( .A(n26753), .B(n26569), .Z(n32604) );
  XOR U32714 ( .A(n32605), .B(n29185), .Z(n26569) );
  XOR U32715 ( .A(n31045), .B(n32606), .Z(n29185) );
  NOR U32716 ( .A(n30412), .B(n30413), .Z(n32605) );
  IV U32717 ( .A(n30894), .Z(n30412) );
  XNOR U32718 ( .A(n32607), .B(n30748), .Z(n30894) );
  XNOR U32719 ( .A(n32608), .B(n29195), .Z(n26753) );
  XNOR U32720 ( .A(n32609), .B(n31834), .Z(n29195) );
  XOR U32721 ( .A(n32610), .B(n31229), .Z(n30405) );
  XOR U32722 ( .A(n30719), .B(n32611), .Z(n32603) );
  XNOR U32723 ( .A(n30873), .B(n25951), .Z(n32611) );
  XNOR U32724 ( .A(n32612), .B(n29189), .Z(n25951) );
  XOR U32725 ( .A(n32613), .B(n31253), .Z(n29189) );
  ANDN U32726 ( .B(n32574), .A(n30891), .Z(n32612) );
  XOR U32727 ( .A(n31337), .B(n32614), .Z(n30891) );
  XNOR U32728 ( .A(n32615), .B(n29199), .Z(n30873) );
  XOR U32729 ( .A(n32616), .B(n29027), .Z(n29199) );
  XNOR U32730 ( .A(n32617), .B(n32618), .Z(n29027) );
  XOR U32731 ( .A(n32619), .B(n32620), .Z(n30409) );
  XNOR U32732 ( .A(n32621), .B(n30888), .Z(n30719) );
  XOR U32733 ( .A(n32622), .B(n32623), .Z(n30888) );
  ANDN U32734 ( .B(n30416), .A(n30417), .Z(n32621) );
  XOR U32735 ( .A(n32624), .B(n32625), .Z(n30416) );
  XOR U32736 ( .A(n21385), .B(n28407), .Z(n25910) );
  XOR U32737 ( .A(n32626), .B(n30773), .Z(n28407) );
  ANDN U32738 ( .B(n28032), .A(n28030), .Z(n32626) );
  IV U32739 ( .A(n32627), .Z(n28030) );
  XOR U32740 ( .A(n32628), .B(n32266), .Z(n28032) );
  IV U32741 ( .A(n23515), .Z(n21385) );
  XOR U32742 ( .A(n26726), .B(n26791), .Z(n23515) );
  XNOR U32743 ( .A(n32629), .B(n32630), .Z(n26791) );
  XNOR U32744 ( .A(n22516), .B(n24149), .Z(n32630) );
  XNOR U32745 ( .A(n32631), .B(n29698), .Z(n24149) );
  ANDN U32746 ( .B(n28320), .A(n29685), .Z(n32631) );
  XOR U32747 ( .A(n31951), .B(n32632), .Z(n29685) );
  XOR U32748 ( .A(n32633), .B(n31968), .Z(n28320) );
  XNOR U32749 ( .A(n32634), .B(n32635), .Z(n22516) );
  ANDN U32750 ( .B(n29687), .A(n29688), .Z(n32634) );
  XOR U32751 ( .A(n32427), .B(n31657), .Z(n29688) );
  ANDN U32752 ( .B(n32638), .A(n32639), .Z(n32636) );
  XOR U32753 ( .A(n24552), .B(n32640), .Z(n32629) );
  XNOR U32754 ( .A(n26247), .B(n27899), .Z(n32640) );
  XNOR U32755 ( .A(n32641), .B(n32642), .Z(n27899) );
  ANDN U32756 ( .B(n28306), .A(n29678), .Z(n32641) );
  XOR U32757 ( .A(n32643), .B(n32644), .Z(n28306) );
  XNOR U32758 ( .A(n32645), .B(n29702), .Z(n26247) );
  ANDN U32759 ( .B(n29680), .A(n28310), .Z(n32645) );
  XOR U32760 ( .A(n32109), .B(n32646), .Z(n28310) );
  XOR U32761 ( .A(n32647), .B(n32648), .Z(n29680) );
  XNOR U32762 ( .A(n32649), .B(n29704), .Z(n24552) );
  ANDN U32763 ( .B(n28316), .A(n29683), .Z(n32649) );
  XNOR U32764 ( .A(n31137), .B(n32650), .Z(n29683) );
  XNOR U32765 ( .A(n32240), .B(n32651), .Z(n31137) );
  XNOR U32766 ( .A(n32652), .B(n32653), .Z(n32240) );
  XOR U32767 ( .A(n32647), .B(n30516), .Z(n32653) );
  XOR U32768 ( .A(n32654), .B(n32655), .Z(n30516) );
  ANDN U32769 ( .B(n32656), .A(n32657), .Z(n32654) );
  XNOR U32770 ( .A(n32658), .B(n32659), .Z(n32647) );
  ANDN U32771 ( .B(n32660), .A(n32661), .Z(n32658) );
  XOR U32772 ( .A(n32662), .B(n32663), .Z(n32652) );
  XOR U32773 ( .A(n32664), .B(n32665), .Z(n32663) );
  XOR U32774 ( .A(n32666), .B(n31340), .Z(n28316) );
  XOR U32775 ( .A(n32667), .B(n32668), .Z(n26726) );
  XOR U32776 ( .A(n29693), .B(n23838), .Z(n32668) );
  XNOR U32777 ( .A(n32669), .B(n28822), .Z(n23838) );
  XOR U32778 ( .A(n32670), .B(n27937), .Z(n28822) );
  NOR U32779 ( .A(n28403), .B(n28404), .Z(n32669) );
  XOR U32780 ( .A(n32664), .B(n32648), .Z(n28404) );
  IV U32781 ( .A(n30517), .Z(n32648) );
  XOR U32782 ( .A(n32671), .B(n32672), .Z(n32664) );
  NOR U32783 ( .A(n32673), .B(n32674), .Z(n32671) );
  XNOR U32784 ( .A(n28765), .B(n32675), .Z(n28403) );
  XOR U32785 ( .A(n32676), .B(n28826), .Z(n29693) );
  XNOR U32786 ( .A(n32245), .B(n32677), .Z(n28826) );
  XNOR U32787 ( .A(n32678), .B(n32679), .Z(n32245) );
  XOR U32788 ( .A(n31054), .B(n32680), .Z(n28022) );
  XOR U32789 ( .A(n32365), .B(n32681), .Z(n28409) );
  XNOR U32790 ( .A(n25180), .B(n32682), .Z(n32667) );
  XOR U32791 ( .A(n28707), .B(n23332), .Z(n32682) );
  XOR U32792 ( .A(n32683), .B(n28837), .Z(n23332) );
  XOR U32793 ( .A(n32684), .B(n32511), .Z(n28837) );
  ANDN U32794 ( .B(n28411), .A(n28017), .Z(n32683) );
  XOR U32795 ( .A(n32685), .B(n28881), .Z(n28017) );
  XOR U32796 ( .A(n32686), .B(n30071), .Z(n28411) );
  XNOR U32797 ( .A(n32687), .B(n28833), .Z(n28707) );
  XOR U32798 ( .A(n32688), .B(n32585), .Z(n28833) );
  NOR U32799 ( .A(n28774), .B(n28026), .Z(n32687) );
  XNOR U32800 ( .A(n32689), .B(n31872), .Z(n28026) );
  XOR U32801 ( .A(n32690), .B(n29962), .Z(n28774) );
  IV U32802 ( .A(n32691), .Z(n29962) );
  XNOR U32803 ( .A(n32692), .B(n28829), .Z(n25180) );
  XOR U32804 ( .A(n32693), .B(n32139), .Z(n28829) );
  NOR U32805 ( .A(n32627), .B(n30773), .Z(n32692) );
  XNOR U32806 ( .A(n32695), .B(n30784), .Z(n32627) );
  XNOR U32807 ( .A(n23219), .B(n32696), .Z(n32440) );
  XOR U32808 ( .A(n18054), .B(n19326), .Z(n32696) );
  XNOR U32809 ( .A(n32697), .B(n23462), .Z(n19326) );
  IV U32810 ( .A(n26288), .Z(n23462) );
  XOR U32811 ( .A(n23586), .B(n31813), .Z(n26288) );
  XNOR U32812 ( .A(n32698), .B(n32699), .Z(n31813) );
  NOR U32813 ( .A(n29342), .B(n29343), .Z(n32698) );
  XOR U32814 ( .A(n32700), .B(n31698), .Z(n29343) );
  XNOR U32815 ( .A(n29374), .B(n30509), .Z(n23586) );
  XNOR U32816 ( .A(n32701), .B(n32702), .Z(n30509) );
  XNOR U32817 ( .A(n23023), .B(n23493), .Z(n32702) );
  XNOR U32818 ( .A(n32703), .B(n28934), .Z(n23493) );
  XOR U32819 ( .A(n30856), .B(n32704), .Z(n28934) );
  IV U32820 ( .A(n32705), .Z(n30856) );
  ANDN U32821 ( .B(n28935), .A(n29335), .Z(n32703) );
  XNOR U32822 ( .A(n32706), .B(n29047), .Z(n29335) );
  XNOR U32823 ( .A(n30483), .B(n32707), .Z(n28935) );
  XNOR U32824 ( .A(n32708), .B(n28929), .Z(n23023) );
  XNOR U32825 ( .A(n32709), .B(n32232), .Z(n28929) );
  ANDN U32826 ( .B(n28930), .A(n29346), .Z(n32708) );
  XNOR U32827 ( .A(n32710), .B(n29299), .Z(n29346) );
  XOR U32828 ( .A(n32711), .B(n28765), .Z(n28930) );
  XOR U32829 ( .A(n32712), .B(n32713), .Z(n28765) );
  XNOR U32830 ( .A(n27384), .B(n32714), .Z(n32701) );
  XNOR U32831 ( .A(n24921), .B(n27578), .Z(n32714) );
  XNOR U32832 ( .A(n32715), .B(n30909), .Z(n27578) );
  XNOR U32833 ( .A(n32716), .B(n28836), .Z(n30909) );
  ANDN U32834 ( .B(n29342), .A(n32699), .Z(n32715) );
  IV U32835 ( .A(n30931), .Z(n32699) );
  XNOR U32836 ( .A(n32302), .B(n32717), .Z(n30931) );
  XOR U32837 ( .A(n32718), .B(n31588), .Z(n29342) );
  XNOR U32838 ( .A(n32719), .B(n28939), .Z(n24921) );
  XNOR U32839 ( .A(n30586), .B(n32720), .Z(n28939) );
  ANDN U32840 ( .B(n28938), .A(n31808), .Z(n32719) );
  XOR U32841 ( .A(n32721), .B(n31584), .Z(n31808) );
  XOR U32842 ( .A(n31666), .B(n32722), .Z(n28938) );
  XOR U32843 ( .A(n32723), .B(n28943), .Z(n27384) );
  XNOR U32844 ( .A(n30149), .B(n32724), .Z(n28943) );
  ANDN U32845 ( .B(n31817), .A(n28942), .Z(n32723) );
  XOR U32846 ( .A(n32725), .B(n29064), .Z(n28942) );
  XOR U32847 ( .A(n32726), .B(n30381), .Z(n31817) );
  XOR U32848 ( .A(n32727), .B(n32728), .Z(n29374) );
  XNOR U32849 ( .A(n26463), .B(n22981), .Z(n32728) );
  XNOR U32850 ( .A(n32729), .B(n29655), .Z(n22981) );
  XOR U32851 ( .A(n32034), .B(n32730), .Z(n29655) );
  NOR U32852 ( .A(n31790), .B(n31033), .Z(n32729) );
  XOR U32853 ( .A(n32038), .B(n32731), .Z(n31033) );
  XOR U32854 ( .A(n32732), .B(n30149), .Z(n31790) );
  XNOR U32855 ( .A(n32733), .B(n29648), .Z(n26463) );
  XOR U32856 ( .A(n32734), .B(n32015), .Z(n29648) );
  ANDN U32857 ( .B(n29647), .A(n29361), .Z(n32733) );
  XOR U32858 ( .A(n32735), .B(n32389), .Z(n29361) );
  XNOR U32859 ( .A(n28421), .B(n32736), .Z(n29647) );
  XOR U32860 ( .A(n29638), .B(n32737), .Z(n32727) );
  XOR U32861 ( .A(n25953), .B(n25029), .Z(n32737) );
  XOR U32862 ( .A(n32738), .B(n30592), .Z(n25029) );
  XOR U32863 ( .A(n32739), .B(n30293), .Z(n30592) );
  IV U32864 ( .A(n32538), .Z(n30293) );
  ANDN U32865 ( .B(n29365), .A(n31797), .Z(n32738) );
  IV U32866 ( .A(n30593), .Z(n31797) );
  XOR U32867 ( .A(n32740), .B(n31709), .Z(n30593) );
  IV U32868 ( .A(n30105), .Z(n31709) );
  XOR U32869 ( .A(n32741), .B(n32742), .Z(n30105) );
  XOR U32870 ( .A(n32743), .B(n32744), .Z(n29365) );
  XOR U32871 ( .A(n32745), .B(n29651), .Z(n25953) );
  XOR U32872 ( .A(n32746), .B(n32747), .Z(n29651) );
  NOR U32873 ( .A(n29650), .B(n29351), .Z(n32745) );
  XOR U32874 ( .A(n32748), .B(n31570), .Z(n29351) );
  XNOR U32875 ( .A(n32749), .B(n31666), .Z(n29650) );
  XNOR U32876 ( .A(n32750), .B(n29643), .Z(n29638) );
  XNOR U32877 ( .A(n32751), .B(n32302), .Z(n29643) );
  AND U32878 ( .A(n29355), .B(n29644), .Z(n32750) );
  XOR U32879 ( .A(n31754), .B(n32752), .Z(n29644) );
  XOR U32880 ( .A(n32753), .B(n29413), .Z(n29355) );
  XNOR U32881 ( .A(n32754), .B(n32755), .Z(n29413) );
  ANDN U32882 ( .B(n23463), .A(n23671), .Z(n32697) );
  XOR U32883 ( .A(n26089), .B(n32756), .Z(n23671) );
  XNOR U32884 ( .A(n30933), .B(n27388), .Z(n26089) );
  XOR U32885 ( .A(n32757), .B(n32758), .Z(n27388) );
  XNOR U32886 ( .A(n25376), .B(n24856), .Z(n32758) );
  XNOR U32887 ( .A(n32759), .B(n30845), .Z(n24856) );
  XNOR U32888 ( .A(n32760), .B(n31190), .Z(n30845) );
  NOR U32889 ( .A(n30846), .B(n31620), .Z(n32759) );
  XNOR U32890 ( .A(n32761), .B(n31086), .Z(n25376) );
  XOR U32891 ( .A(n27983), .B(n32763), .Z(n32757) );
  XOR U32892 ( .A(n26522), .B(n27102), .Z(n32763) );
  XNOR U32893 ( .A(n32764), .B(n30842), .Z(n27102) );
  XOR U32894 ( .A(n32765), .B(n32595), .Z(n30842) );
  XNOR U32895 ( .A(n32766), .B(n30832), .Z(n26522) );
  XNOR U32896 ( .A(n32767), .B(n32768), .Z(n30832) );
  ANDN U32897 ( .B(n32769), .A(n30833), .Z(n32766) );
  XOR U32898 ( .A(n32770), .B(n30838), .Z(n27983) );
  XOR U32899 ( .A(n32097), .B(n32771), .Z(n30838) );
  IV U32900 ( .A(n30852), .Z(n32097) );
  XOR U32901 ( .A(n32773), .B(n32774), .Z(n30933) );
  XNOR U32902 ( .A(n25107), .B(n25167), .Z(n32774) );
  XNOR U32903 ( .A(n32775), .B(n32776), .Z(n25167) );
  ANDN U32904 ( .B(n31485), .A(n31916), .Z(n32775) );
  XNOR U32905 ( .A(n32777), .B(n27992), .Z(n25107) );
  NOR U32906 ( .A(n32778), .B(n31490), .Z(n32777) );
  XOR U32907 ( .A(n26865), .B(n32779), .Z(n32773) );
  XNOR U32908 ( .A(n23966), .B(n23913), .Z(n32779) );
  XOR U32909 ( .A(n32780), .B(n28000), .Z(n23913) );
  ANDN U32910 ( .B(n28001), .A(n31482), .Z(n32780) );
  XNOR U32911 ( .A(n32781), .B(n27996), .Z(n23966) );
  ANDN U32912 ( .B(n27997), .A(n32782), .Z(n32781) );
  XNOR U32913 ( .A(n32783), .B(n32784), .Z(n26865) );
  ANDN U32914 ( .B(n32785), .A(n31496), .Z(n32783) );
  IV U32915 ( .A(n32786), .Z(n31496) );
  XOR U32916 ( .A(n27014), .B(n22017), .Z(n23463) );
  IV U32917 ( .A(n21586), .Z(n22017) );
  XOR U32918 ( .A(n27513), .B(n27897), .Z(n21586) );
  XNOR U32919 ( .A(n32787), .B(n32788), .Z(n27897) );
  XNOR U32920 ( .A(n24338), .B(n25311), .Z(n32788) );
  XNOR U32921 ( .A(n32789), .B(n26938), .Z(n25311) );
  XOR U32922 ( .A(n32389), .B(n32790), .Z(n26938) );
  NOR U32923 ( .A(n27028), .B(n27029), .Z(n32789) );
  XOR U32924 ( .A(n32791), .B(n32691), .Z(n27029) );
  IV U32925 ( .A(n26939), .Z(n27028) );
  XOR U32926 ( .A(n32792), .B(n32585), .Z(n26939) );
  XNOR U32927 ( .A(n32793), .B(n26943), .Z(n24338) );
  IV U32928 ( .A(n32096), .Z(n26943) );
  XOR U32929 ( .A(n32794), .B(n32587), .Z(n32096) );
  IV U32930 ( .A(n30764), .Z(n32587) );
  NOR U32931 ( .A(n26942), .B(n27016), .Z(n32793) );
  XOR U32932 ( .A(n32795), .B(n31448), .Z(n27016) );
  XOR U32933 ( .A(n32796), .B(n32531), .Z(n26942) );
  XOR U32934 ( .A(n26928), .B(n32797), .Z(n32787) );
  XOR U32935 ( .A(n24070), .B(n25674), .Z(n32797) );
  XNOR U32936 ( .A(n32798), .B(n32093), .Z(n25674) );
  IV U32937 ( .A(n32126), .Z(n32093) );
  XOR U32938 ( .A(n32799), .B(n32313), .Z(n32126) );
  NOR U32939 ( .A(n27020), .B(n27021), .Z(n32798) );
  XOR U32940 ( .A(n32800), .B(n31598), .Z(n27021) );
  XOR U32941 ( .A(n32801), .B(n32006), .Z(n27020) );
  XOR U32942 ( .A(n32802), .B(n30058), .Z(n24070) );
  XOR U32943 ( .A(n32803), .B(n32804), .Z(n30058) );
  NOR U32944 ( .A(n27024), .B(n27026), .Z(n32802) );
  XOR U32945 ( .A(n32805), .B(n30290), .Z(n27026) );
  XOR U32946 ( .A(n32806), .B(n32807), .Z(n27024) );
  XOR U32947 ( .A(n32808), .B(n27006), .Z(n26928) );
  XNOR U32948 ( .A(n32809), .B(n32018), .Z(n27006) );
  NOR U32949 ( .A(n27443), .B(n27005), .Z(n32808) );
  XOR U32950 ( .A(n32810), .B(n32811), .Z(n27513) );
  XNOR U32951 ( .A(n32812), .B(n25409), .Z(n32811) );
  XNOR U32952 ( .A(n32813), .B(n32111), .Z(n25409) );
  IV U32953 ( .A(n32814), .Z(n32111) );
  NOR U32954 ( .A(n28560), .B(n27301), .Z(n32813) );
  XOR U32955 ( .A(n31613), .B(n32815), .Z(n27301) );
  XNOR U32956 ( .A(n25688), .B(n32816), .Z(n32810) );
  XOR U32957 ( .A(n21381), .B(n25434), .Z(n32816) );
  XNOR U32958 ( .A(n32817), .B(n32115), .Z(n25434) );
  ANDN U32959 ( .B(n28556), .A(n27287), .Z(n32817) );
  IV U32960 ( .A(n28557), .Z(n27287) );
  XOR U32961 ( .A(n32818), .B(n32819), .Z(n28557) );
  XNOR U32962 ( .A(n32820), .B(n32119), .Z(n21381) );
  IV U32963 ( .A(n32821), .Z(n32119) );
  NOR U32964 ( .A(n27291), .B(n28549), .Z(n32820) );
  XNOR U32965 ( .A(n32822), .B(n30027), .Z(n27291) );
  XNOR U32966 ( .A(n32823), .B(n32107), .Z(n25688) );
  ANDN U32967 ( .B(n28553), .A(n28552), .Z(n32823) );
  IV U32968 ( .A(n32824), .Z(n28552) );
  XOR U32969 ( .A(n32825), .B(n29258), .Z(n28553) );
  IV U32970 ( .A(n32205), .Z(n29258) );
  XNOR U32971 ( .A(n32826), .B(n27005), .Z(n27014) );
  XNOR U32972 ( .A(n32827), .B(n32064), .Z(n27005) );
  ANDN U32973 ( .B(n27443), .A(n27444), .Z(n32826) );
  XOR U32974 ( .A(n32828), .B(n32829), .Z(n27444) );
  XNOR U32975 ( .A(n29271), .B(n32830), .Z(n27443) );
  XNOR U32976 ( .A(n32831), .B(n23470), .Z(n18054) );
  XNOR U32977 ( .A(n29209), .B(n25247), .Z(n23470) );
  XNOR U32978 ( .A(n27889), .B(n31449), .Z(n25247) );
  XOR U32979 ( .A(n32832), .B(n32833), .Z(n31449) );
  XOR U32980 ( .A(n26190), .B(n28365), .Z(n32833) );
  XNOR U32981 ( .A(n32834), .B(n30410), .Z(n28365) );
  XNOR U32982 ( .A(n29266), .B(n32835), .Z(n30410) );
  IV U32983 ( .A(n32747), .Z(n29266) );
  ANDN U32984 ( .B(n29200), .A(n29198), .Z(n32834) );
  XNOR U32985 ( .A(n32836), .B(n30746), .Z(n29198) );
  XNOR U32986 ( .A(n30120), .B(n32837), .Z(n29200) );
  XNOR U32987 ( .A(n32838), .B(n30413), .Z(n26190) );
  XOR U32988 ( .A(n32839), .B(n27939), .Z(n30413) );
  ANDN U32989 ( .B(n29186), .A(n30414), .Z(n32838) );
  XOR U32990 ( .A(n32840), .B(n31894), .Z(n30414) );
  XOR U32991 ( .A(n32841), .B(n32842), .Z(n31894) );
  XNOR U32992 ( .A(n32843), .B(n32602), .Z(n29186) );
  XOR U32993 ( .A(n22959), .B(n32844), .Z(n32832) );
  XNOR U32994 ( .A(n26981), .B(n30400), .Z(n32844) );
  XNOR U32995 ( .A(n32845), .B(n30417), .Z(n30400) );
  XOR U32996 ( .A(n32846), .B(n31454), .Z(n30417) );
  ANDN U32997 ( .B(n31477), .A(n30418), .Z(n32845) );
  XOR U32998 ( .A(n32847), .B(n32044), .Z(n30418) );
  IV U32999 ( .A(n30887), .Z(n31477) );
  XOR U33000 ( .A(n32848), .B(n31376), .Z(n30887) );
  XNOR U33001 ( .A(n32849), .B(n30406), .Z(n26981) );
  XOR U33002 ( .A(n32850), .B(n29329), .Z(n30406) );
  NOR U33003 ( .A(n30897), .B(n29194), .Z(n32849) );
  XOR U33004 ( .A(n30541), .B(n32851), .Z(n29194) );
  IV U33005 ( .A(n29196), .Z(n30897) );
  XOR U33006 ( .A(n32852), .B(n31855), .Z(n29196) );
  XNOR U33007 ( .A(n32853), .B(n32574), .Z(n22959) );
  XOR U33008 ( .A(n32854), .B(n32266), .Z(n32574) );
  NOR U33009 ( .A(n30890), .B(n29188), .Z(n32853) );
  XOR U33010 ( .A(n32429), .B(n31657), .Z(n29188) );
  XOR U33011 ( .A(n32855), .B(n32856), .Z(n32429) );
  AND U33012 ( .A(n32857), .B(n32858), .Z(n32855) );
  IV U33013 ( .A(n29190), .Z(n30890) );
  XOR U33014 ( .A(n30961), .B(n32859), .Z(n29190) );
  XOR U33015 ( .A(n32860), .B(n32861), .Z(n27889) );
  XOR U33016 ( .A(n25595), .B(n26557), .Z(n32861) );
  XNOR U33017 ( .A(n32862), .B(n32027), .Z(n26557) );
  XOR U33018 ( .A(n32863), .B(n29067), .Z(n32027) );
  XOR U33019 ( .A(n32864), .B(n32865), .Z(n29067) );
  NOR U33020 ( .A(n32045), .B(n27969), .Z(n32862) );
  XOR U33021 ( .A(n32866), .B(n29092), .Z(n25595) );
  XNOR U33022 ( .A(n30253), .B(n32867), .Z(n29092) );
  NOR U33023 ( .A(n29091), .B(n27975), .Z(n32866) );
  XOR U33024 ( .A(n32868), .B(n28881), .Z(n27975) );
  XOR U33025 ( .A(n32869), .B(n29937), .Z(n29091) );
  IV U33026 ( .A(n31268), .Z(n29937) );
  XOR U33027 ( .A(n26255), .B(n32870), .Z(n32860) );
  XOR U33028 ( .A(n22411), .B(n26583), .Z(n32870) );
  XOR U33029 ( .A(n32871), .B(n29084), .Z(n26583) );
  XOR U33030 ( .A(n32872), .B(n29053), .Z(n29084) );
  ANDN U33031 ( .B(n29206), .A(n29083), .Z(n32871) );
  XOR U33032 ( .A(n30865), .B(n32873), .Z(n29083) );
  XOR U33033 ( .A(n32874), .B(n32875), .Z(n29206) );
  XOR U33034 ( .A(n32876), .B(n29089), .Z(n22411) );
  XOR U33035 ( .A(n32464), .B(n28890), .Z(n29089) );
  NOR U33036 ( .A(n32879), .B(n32880), .Z(n32877) );
  XOR U33037 ( .A(n31588), .B(n32881), .Z(n28647) );
  XOR U33038 ( .A(n31943), .B(n32882), .Z(n29088) );
  XNOR U33039 ( .A(n32883), .B(n29079), .Z(n26255) );
  XOR U33040 ( .A(n32884), .B(n28469), .Z(n29079) );
  IV U33041 ( .A(n32885), .Z(n28469) );
  ANDN U33042 ( .B(n27979), .A(n29080), .Z(n32883) );
  XNOR U33043 ( .A(n32886), .B(n32887), .Z(n29080) );
  XOR U33044 ( .A(n32888), .B(n31253), .Z(n27979) );
  XOR U33045 ( .A(n32889), .B(n32045), .Z(n29209) );
  XOR U33046 ( .A(n32890), .B(n32891), .Z(n32045) );
  ANDN U33047 ( .B(n27969), .A(n32026), .Z(n32889) );
  IV U33048 ( .A(n27971), .Z(n32026) );
  XOR U33049 ( .A(n32892), .B(n31855), .Z(n27971) );
  XNOR U33050 ( .A(n32893), .B(n32894), .Z(n31855) );
  XOR U33051 ( .A(n32895), .B(n30691), .Z(n27969) );
  XOR U33052 ( .A(n23322), .B(n31891), .Z(n23668) );
  XOR U33053 ( .A(n32896), .B(n31007), .Z(n31891) );
  NOR U33054 ( .A(n28612), .B(n28614), .Z(n32896) );
  XNOR U33055 ( .A(n32897), .B(n31050), .Z(n28614) );
  XNOR U33056 ( .A(n28651), .B(n28713), .Z(n23322) );
  XNOR U33057 ( .A(n32898), .B(n32899), .Z(n28713) );
  XNOR U33058 ( .A(n30698), .B(n25192), .Z(n32899) );
  XNOR U33059 ( .A(n32900), .B(n32901), .Z(n25192) );
  NOR U33060 ( .A(n31902), .B(n28641), .Z(n32900) );
  XNOR U33061 ( .A(n32902), .B(n31434), .Z(n28641) );
  IV U33062 ( .A(n32903), .Z(n31902) );
  XNOR U33063 ( .A(n32904), .B(n30705), .Z(n30698) );
  ANDN U33064 ( .B(n31728), .A(n31911), .Z(n32904) );
  IV U33065 ( .A(n30704), .Z(n31911) );
  XOR U33066 ( .A(n32905), .B(n29916), .Z(n30704) );
  XOR U33067 ( .A(n30760), .B(n32906), .Z(n31728) );
  XOR U33068 ( .A(n26394), .B(n32907), .Z(n32898) );
  XOR U33069 ( .A(n25408), .B(n24703), .Z(n32907) );
  XOR U33070 ( .A(n32908), .B(n30707), .Z(n24703) );
  ANDN U33071 ( .B(n30708), .A(n28628), .Z(n32908) );
  XOR U33072 ( .A(n32909), .B(n31068), .Z(n28628) );
  XNOR U33073 ( .A(n32910), .B(n30071), .Z(n30708) );
  XNOR U33074 ( .A(n32911), .B(n30715), .Z(n25408) );
  ANDN U33075 ( .B(n28633), .A(n31905), .Z(n32911) );
  IV U33076 ( .A(n30716), .Z(n31905) );
  XOR U33077 ( .A(n32912), .B(n32585), .Z(n30716) );
  XOR U33078 ( .A(n32913), .B(n31654), .Z(n28633) );
  XOR U33079 ( .A(n32914), .B(n32915), .Z(n31654) );
  XOR U33080 ( .A(n32916), .B(n30712), .Z(n26394) );
  ANDN U33081 ( .B(n28637), .A(n31908), .Z(n32916) );
  IV U33082 ( .A(n30713), .Z(n31908) );
  XOR U33083 ( .A(n32917), .B(n32196), .Z(n30713) );
  XOR U33084 ( .A(n32918), .B(n29948), .Z(n28637) );
  XOR U33085 ( .A(n32919), .B(n32920), .Z(n28651) );
  XOR U33086 ( .A(n24832), .B(n24569), .Z(n32920) );
  XNOR U33087 ( .A(n32921), .B(n28645), .Z(n24569) );
  XOR U33088 ( .A(n32923), .B(n32924), .Z(n32585) );
  AND U33089 ( .A(n28612), .B(n31007), .Z(n32921) );
  XOR U33090 ( .A(n32925), .B(n31880), .Z(n31007) );
  XOR U33091 ( .A(n32926), .B(n32927), .Z(n28612) );
  XNOR U33092 ( .A(n32928), .B(n28170), .Z(n24832) );
  XNOR U33093 ( .A(n30860), .B(n32929), .Z(n28170) );
  XOR U33094 ( .A(n32930), .B(n32931), .Z(n30860) );
  ANDN U33095 ( .B(n30991), .A(n28620), .Z(n32928) );
  XNOR U33096 ( .A(n32932), .B(n30014), .Z(n28620) );
  XOR U33097 ( .A(n32933), .B(n32402), .Z(n30991) );
  XOR U33098 ( .A(n26627), .B(n32934), .Z(n32919) );
  XOR U33099 ( .A(n24959), .B(n26385), .Z(n32934) );
  XNOR U33100 ( .A(n32935), .B(n28102), .Z(n26385) );
  XNOR U33101 ( .A(n32936), .B(n31148), .Z(n28102) );
  NOR U33102 ( .A(n31896), .B(n31897), .Z(n32935) );
  XNOR U33103 ( .A(n32937), .B(n29166), .Z(n31897) );
  XOR U33104 ( .A(n32938), .B(n30071), .Z(n31896) );
  XNOR U33105 ( .A(n32939), .B(n32940), .Z(n30071) );
  XOR U33106 ( .A(n32941), .B(n31003), .Z(n24959) );
  XOR U33107 ( .A(n32942), .B(n30197), .Z(n31003) );
  AND U33108 ( .A(n31002), .B(n28616), .Z(n32941) );
  XNOR U33109 ( .A(n30364), .B(n32943), .Z(n28616) );
  XOR U33110 ( .A(n32944), .B(n31822), .Z(n31002) );
  XNOR U33111 ( .A(n32945), .B(n28106), .Z(n26627) );
  XNOR U33112 ( .A(n30483), .B(n32946), .Z(n28106) );
  ANDN U33113 ( .B(n28623), .A(n30994), .Z(n32945) );
  XOR U33114 ( .A(n32947), .B(n30691), .Z(n30994) );
  IV U33115 ( .A(n32299), .Z(n30691) );
  XOR U33116 ( .A(n32948), .B(n32949), .Z(n32299) );
  XNOR U33117 ( .A(n32950), .B(n31322), .Z(n28623) );
  XOR U33118 ( .A(n29846), .B(n26975), .Z(n23471) );
  IV U33119 ( .A(n24874), .Z(n26975) );
  XOR U33120 ( .A(n26263), .B(n26720), .Z(n24874) );
  XNOR U33121 ( .A(n32951), .B(n32952), .Z(n26720) );
  XOR U33122 ( .A(n24242), .B(n25841), .Z(n32952) );
  XNOR U33123 ( .A(n32953), .B(n29421), .Z(n25841) );
  XNOR U33124 ( .A(n30644), .B(n32954), .Z(n29421) );
  NOR U33125 ( .A(n26547), .B(n26548), .Z(n32953) );
  XOR U33126 ( .A(n32955), .B(n32956), .Z(n26548) );
  IV U33127 ( .A(n29422), .Z(n26547) );
  XOR U33128 ( .A(n32957), .B(n30208), .Z(n29422) );
  XNOR U33129 ( .A(n32958), .B(n30731), .Z(n24242) );
  IV U33130 ( .A(n29426), .Z(n30731) );
  XOR U33131 ( .A(n32959), .B(n29948), .Z(n29426) );
  XNOR U33132 ( .A(n32960), .B(n32961), .Z(n29948) );
  NOR U33133 ( .A(n27350), .B(n26499), .Z(n32958) );
  XOR U33134 ( .A(n32962), .B(n29916), .Z(n26499) );
  IV U33135 ( .A(n26500), .Z(n27350) );
  XOR U33136 ( .A(n32963), .B(n32964), .Z(n26500) );
  XNOR U33137 ( .A(n25114), .B(n32965), .Z(n32951) );
  XNOR U33138 ( .A(n24616), .B(n25339), .Z(n32965) );
  XNOR U33139 ( .A(n32966), .B(n30736), .Z(n25339) );
  IV U33140 ( .A(n29428), .Z(n30736) );
  XOR U33141 ( .A(n32967), .B(n31887), .Z(n29428) );
  ANDN U33142 ( .B(n26490), .A(n26488), .Z(n32966) );
  XOR U33143 ( .A(n32968), .B(n31264), .Z(n26488) );
  XNOR U33144 ( .A(n32969), .B(n32970), .Z(n31264) );
  XOR U33145 ( .A(n32971), .B(n32315), .Z(n26490) );
  IV U33146 ( .A(n32972), .Z(n32315) );
  XNOR U33147 ( .A(n32973), .B(n30741), .Z(n24616) );
  IV U33148 ( .A(n29950), .Z(n30741) );
  XOR U33149 ( .A(n32974), .B(n28432), .Z(n29950) );
  IV U33150 ( .A(n32975), .Z(n28432) );
  NOR U33151 ( .A(n26722), .B(n26723), .Z(n32973) );
  XNOR U33152 ( .A(n32976), .B(n30817), .Z(n26723) );
  IV U33153 ( .A(n32625), .Z(n30817) );
  XNOR U33154 ( .A(n32977), .B(n30375), .Z(n26722) );
  XNOR U33155 ( .A(n32978), .B(n29419), .Z(n25114) );
  XOR U33156 ( .A(n31026), .B(n32979), .Z(n29419) );
  ANDN U33157 ( .B(n26494), .A(n26492), .Z(n32978) );
  XNOR U33158 ( .A(n32980), .B(n30116), .Z(n26492) );
  XOR U33159 ( .A(n32981), .B(n31467), .Z(n26494) );
  XNOR U33160 ( .A(n32982), .B(n32983), .Z(n26263) );
  XOR U33161 ( .A(n25190), .B(n23743), .Z(n32983) );
  XOR U33162 ( .A(n32984), .B(n29444), .Z(n23743) );
  ANDN U33163 ( .B(n29443), .A(n29851), .Z(n32984) );
  XOR U33164 ( .A(n32985), .B(n30208), .Z(n29851) );
  XNOR U33165 ( .A(n32986), .B(n32987), .Z(n30208) );
  XOR U33166 ( .A(n32988), .B(n30554), .Z(n29443) );
  XNOR U33167 ( .A(n32989), .B(n30754), .Z(n25190) );
  ANDN U33168 ( .B(n29848), .A(n26323), .Z(n32989) );
  XNOR U33169 ( .A(n32990), .B(n32991), .Z(n26323) );
  XOR U33170 ( .A(n32992), .B(n32993), .Z(n29848) );
  XOR U33171 ( .A(n29415), .B(n32994), .Z(n32982) );
  XOR U33172 ( .A(n24447), .B(n24608), .Z(n32994) );
  XOR U33173 ( .A(n32995), .B(n29433), .Z(n24608) );
  NOR U33174 ( .A(n26336), .B(n29432), .Z(n32995) );
  XOR U33175 ( .A(n32996), .B(n31467), .Z(n29432) );
  XOR U33176 ( .A(n32997), .B(n29533), .Z(n26336) );
  IV U33177 ( .A(n32498), .Z(n29533) );
  XNOR U33178 ( .A(n32998), .B(n29435), .Z(n24447) );
  NOR U33179 ( .A(n32999), .B(n29436), .Z(n32998) );
  XNOR U33180 ( .A(n33000), .B(n29441), .Z(n29415) );
  NOR U33181 ( .A(n29440), .B(n26319), .Z(n33000) );
  XNOR U33182 ( .A(n32963), .B(n33001), .Z(n26319) );
  IV U33183 ( .A(n30946), .Z(n32963) );
  XNOR U33184 ( .A(n33002), .B(n32829), .Z(n29440) );
  XOR U33185 ( .A(n33003), .B(n29436), .Z(n29846) );
  XOR U33186 ( .A(n32274), .B(n33004), .Z(n29436) );
  ANDN U33187 ( .B(n26334), .A(n26332), .Z(n33003) );
  IV U33188 ( .A(n32999), .Z(n26332) );
  XOR U33189 ( .A(n32538), .B(n33005), .Z(n32999) );
  XNOR U33190 ( .A(n33006), .B(n23453), .Z(n23219) );
  XNOR U33191 ( .A(n21603), .B(n29696), .Z(n23453) );
  XNOR U33192 ( .A(n33007), .B(n28307), .Z(n29696) );
  ANDN U33193 ( .B(n29678), .A(n32642), .Z(n33007) );
  XOR U33194 ( .A(n33008), .B(n33009), .Z(n29678) );
  ANDN U33195 ( .B(n23676), .A(n23454), .Z(n33006) );
  XOR U33196 ( .A(n33010), .B(n26718), .Z(n23454) );
  XOR U33197 ( .A(n30726), .B(n25999), .Z(n26718) );
  XNOR U33198 ( .A(n33011), .B(n33012), .Z(n25999) );
  XNOR U33199 ( .A(n26180), .B(n26295), .Z(n33012) );
  XNOR U33200 ( .A(n33013), .B(n26311), .Z(n26295) );
  XOR U33201 ( .A(n32926), .B(n33014), .Z(n26311) );
  ANDN U33202 ( .B(n26310), .A(n28183), .Z(n33013) );
  XOR U33203 ( .A(n33015), .B(n29842), .Z(n26180) );
  XNOR U33204 ( .A(n31455), .B(n33016), .Z(n29842) );
  AND U33205 ( .A(n28191), .B(n29841), .Z(n33015) );
  XNOR U33206 ( .A(n22512), .B(n33017), .Z(n33011) );
  XOR U33207 ( .A(n25100), .B(n22529), .Z(n33017) );
  XOR U33208 ( .A(n33018), .B(n26305), .Z(n22529) );
  XOR U33209 ( .A(n33019), .B(n32620), .Z(n26305) );
  ANDN U33210 ( .B(n33020), .A(n33021), .Z(n33018) );
  XNOR U33211 ( .A(n33022), .B(n26301), .Z(n25100) );
  XOR U33212 ( .A(n28421), .B(n33023), .Z(n26301) );
  ANDN U33213 ( .B(n28195), .A(n26300), .Z(n33022) );
  XNOR U33214 ( .A(n33024), .B(n26314), .Z(n22512) );
  XNOR U33215 ( .A(n33025), .B(n30230), .Z(n26314) );
  AND U33216 ( .A(n28188), .B(n26315), .Z(n33024) );
  XOR U33217 ( .A(n33026), .B(n33027), .Z(n30726) );
  XOR U33218 ( .A(n25066), .B(n21594), .Z(n33027) );
  XNOR U33219 ( .A(n33028), .B(n26334), .Z(n21594) );
  XNOR U33220 ( .A(n33029), .B(n31119), .Z(n26334) );
  IV U33221 ( .A(n31968), .Z(n31119) );
  ANDN U33222 ( .B(n26333), .A(n29435), .Z(n33028) );
  XNOR U33223 ( .A(n33030), .B(n33031), .Z(n29435) );
  XNOR U33224 ( .A(n33032), .B(n32620), .Z(n26333) );
  IV U33225 ( .A(n31444), .Z(n32620) );
  XNOR U33226 ( .A(n33033), .B(n26329), .Z(n25066) );
  XOR U33227 ( .A(n33034), .B(n30175), .Z(n26329) );
  ANDN U33228 ( .B(n29444), .A(n26330), .Z(n33033) );
  XOR U33229 ( .A(n33035), .B(n33036), .Z(n26330) );
  XOR U33230 ( .A(n32250), .B(n33037), .Z(n29444) );
  XOR U33231 ( .A(n25579), .B(n33038), .Z(n33026) );
  XNOR U33232 ( .A(n24957), .B(n25296), .Z(n33038) );
  XNOR U33233 ( .A(n33039), .B(n26325), .Z(n25296) );
  XOR U33234 ( .A(n33040), .B(n30142), .Z(n26325) );
  IV U33235 ( .A(n31707), .Z(n30142) );
  ANDN U33236 ( .B(n26324), .A(n30754), .Z(n33039) );
  XOR U33237 ( .A(n31295), .B(n33041), .Z(n30754) );
  IV U33238 ( .A(n31045), .Z(n31295) );
  XOR U33239 ( .A(n33042), .B(n33043), .Z(n31045) );
  XOR U33240 ( .A(n33045), .B(n26338), .Z(n24957) );
  XOR U33241 ( .A(n33046), .B(n32313), .Z(n26338) );
  ANDN U33242 ( .B(n26337), .A(n29433), .Z(n33045) );
  XOR U33243 ( .A(n33047), .B(n32172), .Z(n29433) );
  XNOR U33244 ( .A(n33048), .B(n33049), .Z(n32172) );
  XOR U33245 ( .A(n33050), .B(n31547), .Z(n26337) );
  XOR U33246 ( .A(n33051), .B(n26320), .Z(n25579) );
  XOR U33247 ( .A(n33052), .B(n33053), .Z(n26320) );
  AND U33248 ( .A(n29441), .B(n26321), .Z(n33051) );
  XOR U33249 ( .A(n33054), .B(n32064), .Z(n26321) );
  XOR U33250 ( .A(n32268), .B(n33055), .Z(n29441) );
  XNOR U33251 ( .A(n26538), .B(n26620), .Z(n23676) );
  XNOR U33252 ( .A(n27582), .B(n32316), .Z(n26620) );
  XOR U33253 ( .A(n33056), .B(n33057), .Z(n32316) );
  XNOR U33254 ( .A(n24826), .B(n25348), .Z(n33057) );
  XOR U33255 ( .A(n33058), .B(n27543), .Z(n25348) );
  XOR U33256 ( .A(n28739), .B(n33059), .Z(n27543) );
  XOR U33257 ( .A(n32302), .B(n33060), .Z(n26994) );
  XOR U33258 ( .A(n33061), .B(n31598), .Z(n26993) );
  XNOR U33259 ( .A(n33064), .B(n27555), .Z(n24826) );
  XOR U33260 ( .A(n33065), .B(n32531), .Z(n27555) );
  NOR U33261 ( .A(n26623), .B(n26622), .Z(n33064) );
  XOR U33262 ( .A(n31669), .B(n33066), .Z(n26622) );
  XOR U33263 ( .A(n33067), .B(n33068), .Z(n26623) );
  XOR U33264 ( .A(n26239), .B(n33069), .Z(n33056) );
  XNOR U33265 ( .A(n27538), .B(n24985), .Z(n33069) );
  XNOR U33266 ( .A(n33070), .B(n27546), .Z(n24985) );
  XOR U33267 ( .A(n33071), .B(n30267), .Z(n27546) );
  IV U33268 ( .A(n32452), .Z(n30267) );
  XOR U33269 ( .A(n33072), .B(n33043), .Z(n32452) );
  XNOR U33270 ( .A(n33073), .B(n33074), .Z(n33043) );
  XNOR U33271 ( .A(n33075), .B(n33076), .Z(n33074) );
  XOR U33272 ( .A(n31571), .B(n33077), .Z(n33073) );
  XOR U33273 ( .A(n32748), .B(n33078), .Z(n33077) );
  XNOR U33274 ( .A(n33079), .B(n33080), .Z(n32748) );
  ANDN U33275 ( .B(n33081), .A(n33082), .Z(n33079) );
  XNOR U33276 ( .A(n33083), .B(n33084), .Z(n31571) );
  ANDN U33277 ( .B(n33085), .A(n33086), .Z(n33083) );
  ANDN U33278 ( .B(n29249), .A(n27547), .Z(n33070) );
  XOR U33279 ( .A(n29965), .B(n33087), .Z(n27547) );
  IV U33280 ( .A(n31357), .Z(n29249) );
  XOR U33281 ( .A(n31455), .B(n33088), .Z(n31357) );
  XNOR U33282 ( .A(n33089), .B(n27559), .Z(n27538) );
  XNOR U33283 ( .A(n32160), .B(n33090), .Z(n27559) );
  NOR U33284 ( .A(n31352), .B(n27558), .Z(n33089) );
  XOR U33285 ( .A(n33091), .B(n32511), .Z(n27558) );
  XOR U33286 ( .A(n32308), .B(n33092), .Z(n31352) );
  XNOR U33287 ( .A(n33093), .B(n27552), .Z(n26239) );
  XOR U33288 ( .A(n33094), .B(n32182), .Z(n27552) );
  ANDN U33289 ( .B(n31371), .A(n27551), .Z(n33093) );
  XOR U33290 ( .A(n33095), .B(n33096), .Z(n27582) );
  XNOR U33291 ( .A(n24850), .B(n22503), .Z(n33096) );
  XNOR U33292 ( .A(n33097), .B(n28036), .Z(n22503) );
  ANDN U33293 ( .B(n28037), .A(n29821), .Z(n33097) );
  XNOR U33294 ( .A(n29047), .B(n33098), .Z(n29821) );
  XNOR U33295 ( .A(n32422), .B(n31657), .Z(n28037) );
  XNOR U33296 ( .A(n33099), .B(n32545), .Z(n31657) );
  XNOR U33297 ( .A(n33100), .B(n33101), .Z(n32545) );
  XOR U33298 ( .A(n33102), .B(n29306), .Z(n33101) );
  XOR U33299 ( .A(n33103), .B(n33104), .Z(n29306) );
  NOR U33300 ( .A(n33105), .B(n33106), .Z(n33103) );
  XOR U33301 ( .A(n33107), .B(n33108), .Z(n33100) );
  XOR U33302 ( .A(n32253), .B(n31354), .Z(n33108) );
  XNOR U33303 ( .A(n33109), .B(n33110), .Z(n31354) );
  XNOR U33304 ( .A(n33113), .B(n33114), .Z(n32253) );
  XNOR U33305 ( .A(n33117), .B(n33118), .Z(n32422) );
  NOR U33306 ( .A(n33119), .B(n33120), .Z(n33117) );
  XOR U33307 ( .A(n33121), .B(n28863), .Z(n24850) );
  AND U33308 ( .A(n29825), .B(n28864), .Z(n33121) );
  XNOR U33309 ( .A(n33122), .B(n31440), .Z(n28864) );
  XOR U33310 ( .A(n28982), .B(n33123), .Z(n29825) );
  XNOR U33311 ( .A(n27056), .B(n33124), .Z(n33095) );
  XNOR U33312 ( .A(n25655), .B(n23340), .Z(n33124) );
  XNOR U33313 ( .A(n33125), .B(n33126), .Z(n23340) );
  ANDN U33314 ( .B(n29831), .A(n29832), .Z(n33125) );
  XOR U33315 ( .A(n31020), .B(n33127), .Z(n29832) );
  XNOR U33316 ( .A(n33128), .B(n27572), .Z(n25655) );
  ANDN U33317 ( .B(n27573), .A(n29829), .Z(n33128) );
  XNOR U33318 ( .A(n33129), .B(n30784), .Z(n29829) );
  XNOR U33319 ( .A(n33130), .B(n27947), .Z(n27573) );
  XNOR U33320 ( .A(n33131), .B(n27566), .Z(n27056) );
  ANDN U33321 ( .B(n29837), .A(n27565), .Z(n33131) );
  IV U33322 ( .A(n29835), .Z(n27565) );
  XOR U33323 ( .A(n33132), .B(n31314), .Z(n29835) );
  XNOR U33324 ( .A(n33133), .B(n29919), .Z(n29837) );
  IV U33325 ( .A(n27942), .Z(n29919) );
  XNOR U33326 ( .A(n33134), .B(n27551), .Z(n26538) );
  XOR U33327 ( .A(n27657), .B(n33135), .Z(n27551) );
  NOR U33328 ( .A(n31371), .B(n28970), .Z(n33134) );
  XOR U33329 ( .A(n33136), .B(n27939), .Z(n28970) );
  IV U33330 ( .A(n33137), .Z(n27939) );
  XNOR U33331 ( .A(n33138), .B(n30375), .Z(n31371) );
  XOR U33332 ( .A(n33139), .B(n33140), .Z(n23805) );
  XNOR U33333 ( .A(n19562), .B(n17532), .Z(n33140) );
  XOR U33334 ( .A(n33141), .B(n23228), .Z(n17532) );
  XNOR U33335 ( .A(n30710), .B(n23577), .Z(n23228) );
  XOR U33336 ( .A(n31731), .B(n27958), .Z(n23577) );
  XOR U33337 ( .A(n33142), .B(n33143), .Z(n27958) );
  XNOR U33338 ( .A(n25964), .B(n23327), .Z(n33143) );
  XNOR U33339 ( .A(n33144), .B(n28634), .Z(n23327) );
  XNOR U33340 ( .A(n33145), .B(n30381), .Z(n28634) );
  IV U33341 ( .A(n28793), .Z(n30381) );
  XOR U33342 ( .A(n33146), .B(n33147), .Z(n28793) );
  ANDN U33343 ( .B(n28635), .A(n30715), .Z(n33144) );
  XOR U33344 ( .A(n30148), .B(n33148), .Z(n30715) );
  XNOR U33345 ( .A(n28421), .B(n33149), .Z(n28635) );
  XNOR U33346 ( .A(n33150), .B(n31729), .Z(n25964) );
  XOR U33347 ( .A(n33151), .B(n31035), .Z(n31729) );
  XOR U33348 ( .A(n32987), .B(n33152), .Z(n31035) );
  XNOR U33349 ( .A(n33153), .B(n33154), .Z(n32987) );
  XNOR U33350 ( .A(n29925), .B(n32279), .Z(n33154) );
  XNOR U33351 ( .A(n33155), .B(n33156), .Z(n32279) );
  NOR U33352 ( .A(n33157), .B(n33158), .Z(n33155) );
  XNOR U33353 ( .A(n33159), .B(n33160), .Z(n29925) );
  ANDN U33354 ( .B(n33161), .A(n33162), .Z(n33159) );
  XNOR U33355 ( .A(n29958), .B(n33163), .Z(n33153) );
  XOR U33356 ( .A(n31837), .B(n33164), .Z(n33163) );
  XOR U33357 ( .A(n33165), .B(n33166), .Z(n31837) );
  ANDN U33358 ( .B(n33167), .A(n33168), .Z(n33165) );
  XNOR U33359 ( .A(n33169), .B(n33170), .Z(n29958) );
  NOR U33360 ( .A(n33171), .B(n33172), .Z(n33169) );
  ANDN U33361 ( .B(n30705), .A(n30703), .Z(n33150) );
  XOR U33362 ( .A(n33173), .B(n33137), .Z(n30703) );
  XOR U33363 ( .A(n33174), .B(n33175), .Z(n33137) );
  XOR U33364 ( .A(n33176), .B(n32402), .Z(n30705) );
  XOR U33365 ( .A(n24551), .B(n33177), .Z(n33142) );
  XNOR U33366 ( .A(n24448), .B(n26289), .Z(n33177) );
  XNOR U33367 ( .A(n33178), .B(n28639), .Z(n26289) );
  XNOR U33368 ( .A(n33179), .B(n29946), .Z(n28639) );
  NOR U33369 ( .A(n30712), .B(n28638), .Z(n33178) );
  XOR U33370 ( .A(n33182), .B(n32011), .Z(n28638) );
  XOR U33371 ( .A(n33183), .B(n31547), .Z(n30712) );
  XNOR U33372 ( .A(n33184), .B(n31903), .Z(n24448) );
  IV U33373 ( .A(n28643), .Z(n31903) );
  XNOR U33374 ( .A(n33185), .B(n32804), .Z(n28643) );
  ANDN U33375 ( .B(n32901), .A(n28642), .Z(n33184) );
  XNOR U33376 ( .A(n33186), .B(n28630), .Z(n24551) );
  XOR U33377 ( .A(n30961), .B(n33187), .Z(n28630) );
  NOR U33378 ( .A(n30707), .B(n28629), .Z(n33186) );
  XOR U33379 ( .A(n28747), .B(n33188), .Z(n28629) );
  XNOR U33380 ( .A(n33189), .B(n30535), .Z(n30707) );
  XOR U33381 ( .A(n33190), .B(n33191), .Z(n31731) );
  XNOR U33382 ( .A(n24786), .B(n24594), .Z(n33191) );
  XOR U33383 ( .A(n33192), .B(n27220), .Z(n24594) );
  XOR U33384 ( .A(n33193), .B(n30215), .Z(n27220) );
  NOR U33385 ( .A(n32070), .B(n32071), .Z(n33192) );
  XOR U33386 ( .A(n33194), .B(n32804), .Z(n32070) );
  XOR U33387 ( .A(n33195), .B(n27224), .Z(n24786) );
  XOR U33388 ( .A(n33196), .B(n30752), .Z(n27224) );
  NOR U33389 ( .A(n32068), .B(n27223), .Z(n33195) );
  XOR U33390 ( .A(n32538), .B(n33197), .Z(n27223) );
  XNOR U33391 ( .A(n33198), .B(n33199), .Z(n32538) );
  XOR U33392 ( .A(n26039), .B(n33200), .Z(n33190) );
  XOR U33393 ( .A(n27203), .B(n21720), .Z(n33200) );
  XNOR U33394 ( .A(n33201), .B(n27209), .Z(n21720) );
  ANDN U33395 ( .B(n27210), .A(n32074), .Z(n33201) );
  XOR U33396 ( .A(n33202), .B(n32139), .Z(n27210) );
  XNOR U33397 ( .A(n33203), .B(n29909), .Z(n27203) );
  XOR U33398 ( .A(n31810), .B(n33204), .Z(n29909) );
  ANDN U33399 ( .B(n29910), .A(n32077), .Z(n33203) );
  XOR U33400 ( .A(n33205), .B(n31680), .Z(n29910) );
  XNOR U33401 ( .A(n33206), .B(n27213), .Z(n26039) );
  XNOR U33402 ( .A(n28747), .B(n33207), .Z(n27213) );
  NOR U33403 ( .A(n32079), .B(n32080), .Z(n33206) );
  XOR U33404 ( .A(n33208), .B(n29934), .Z(n32079) );
  IV U33405 ( .A(n29741), .Z(n29934) );
  XNOR U33406 ( .A(n33209), .B(n33152), .Z(n29741) );
  XNOR U33407 ( .A(n33210), .B(n33211), .Z(n33152) );
  XOR U33408 ( .A(n33212), .B(n33213), .Z(n33211) );
  XOR U33409 ( .A(n33214), .B(n33215), .Z(n33210) );
  XNOR U33410 ( .A(n33216), .B(n33217), .Z(n33215) );
  XNOR U33411 ( .A(n33218), .B(n28642), .Z(n30710) );
  XNOR U33412 ( .A(n33219), .B(n30014), .Z(n28642) );
  XNOR U33413 ( .A(n33220), .B(n33221), .Z(n30014) );
  NOR U33414 ( .A(n32903), .B(n32901), .Z(n33218) );
  XOR U33415 ( .A(n32274), .B(n33222), .Z(n32901) );
  XOR U33416 ( .A(n33223), .B(n31584), .Z(n32903) );
  ANDN U33417 ( .B(n25141), .A(n25926), .Z(n33141) );
  IV U33418 ( .A(n23229), .Z(n25926) );
  XOR U33419 ( .A(n23714), .B(n26680), .Z(n23229) );
  XOR U33420 ( .A(n33224), .B(n31921), .Z(n26680) );
  ANDN U33421 ( .B(n27720), .A(n33225), .Z(n33224) );
  XNOR U33422 ( .A(n33212), .B(n33226), .Z(n27720) );
  XNOR U33423 ( .A(n33227), .B(n33228), .Z(n33212) );
  NOR U33424 ( .A(n33229), .B(n33230), .Z(n33227) );
  XNOR U33425 ( .A(n31644), .B(n30386), .Z(n23714) );
  XOR U33426 ( .A(n33231), .B(n33232), .Z(n30386) );
  XOR U33427 ( .A(n27200), .B(n25790), .Z(n33232) );
  XOR U33428 ( .A(n33233), .B(n29038), .Z(n25790) );
  XOR U33429 ( .A(n30200), .B(n33234), .Z(n29038) );
  ANDN U33430 ( .B(n29039), .A(n31767), .Z(n33233) );
  IV U33431 ( .A(n29461), .Z(n31767) );
  XOR U33432 ( .A(n33235), .B(n29713), .Z(n29461) );
  XOR U33433 ( .A(n33236), .B(n31223), .Z(n29039) );
  XNOR U33434 ( .A(n33237), .B(n28341), .Z(n27200) );
  XNOR U33435 ( .A(n30066), .B(n33238), .Z(n28341) );
  ANDN U33436 ( .B(n28342), .A(n30384), .Z(n33237) );
  XOR U33437 ( .A(n33239), .B(n31376), .Z(n30384) );
  XOR U33438 ( .A(n33240), .B(n28796), .Z(n28342) );
  XNOR U33439 ( .A(n25277), .B(n33241), .Z(n33231) );
  XOR U33440 ( .A(n24711), .B(n26636), .Z(n33241) );
  XNOR U33441 ( .A(n33242), .B(n28354), .Z(n26636) );
  XOR U33442 ( .A(n29064), .B(n33243), .Z(n28354) );
  IV U33443 ( .A(n29300), .Z(n29064) );
  XOR U33444 ( .A(n33099), .B(n33244), .Z(n29300) );
  XOR U33445 ( .A(n33245), .B(n33246), .Z(n33099) );
  XNOR U33446 ( .A(n30269), .B(n30070), .Z(n33246) );
  XNOR U33447 ( .A(n33247), .B(n33248), .Z(n30070) );
  NOR U33448 ( .A(n32432), .B(n32431), .Z(n33247) );
  XNOR U33449 ( .A(n33249), .B(n33250), .Z(n30269) );
  AND U33450 ( .A(n33119), .B(n33118), .Z(n33249) );
  XOR U33451 ( .A(n32910), .B(n33251), .Z(n33245) );
  XNOR U33452 ( .A(n32686), .B(n32938), .Z(n33251) );
  XNOR U33453 ( .A(n33252), .B(n33253), .Z(n32938) );
  NOR U33454 ( .A(n32858), .B(n32856), .Z(n33252) );
  XNOR U33455 ( .A(n33254), .B(n33255), .Z(n32686) );
  AND U33456 ( .A(n32426), .B(n32424), .Z(n33254) );
  XOR U33457 ( .A(n33256), .B(n33257), .Z(n32910) );
  ANDN U33458 ( .B(n32639), .A(n32637), .Z(n33256) );
  AND U33459 ( .A(n28355), .B(n29453), .Z(n33242) );
  XNOR U33460 ( .A(n28790), .B(n33258), .Z(n29453) );
  XOR U33461 ( .A(n33259), .B(n33260), .Z(n28355) );
  XNOR U33462 ( .A(n33261), .B(n28351), .Z(n24711) );
  XOR U33463 ( .A(n31238), .B(n33262), .Z(n28351) );
  NOR U33464 ( .A(n30019), .B(n28350), .Z(n33261) );
  XOR U33465 ( .A(n33263), .B(n29922), .Z(n28350) );
  XNOR U33466 ( .A(n32990), .B(n33264), .Z(n30019) );
  IV U33467 ( .A(n33265), .Z(n32990) );
  XNOR U33468 ( .A(n33266), .B(n28346), .Z(n25277) );
  XOR U33469 ( .A(n32101), .B(n33267), .Z(n28346) );
  NOR U33470 ( .A(n28347), .B(n29458), .Z(n33266) );
  XOR U33471 ( .A(n31810), .B(n33268), .Z(n29458) );
  XOR U33472 ( .A(n33269), .B(n29299), .Z(n28347) );
  IV U33473 ( .A(n30300), .Z(n29299) );
  XNOR U33474 ( .A(n32678), .B(n33270), .Z(n30300) );
  XOR U33475 ( .A(n33271), .B(n33272), .Z(n32678) );
  XOR U33476 ( .A(n33132), .B(n31313), .Z(n33272) );
  XOR U33477 ( .A(n33273), .B(n33274), .Z(n31313) );
  NOR U33478 ( .A(n33275), .B(n33276), .Z(n33273) );
  XNOR U33479 ( .A(n33277), .B(n33278), .Z(n33132) );
  ANDN U33480 ( .B(n33279), .A(n33280), .Z(n33277) );
  XOR U33481 ( .A(n33281), .B(n33282), .Z(n33271) );
  XOR U33482 ( .A(n32818), .B(n32485), .Z(n33282) );
  XNOR U33483 ( .A(n33283), .B(n33284), .Z(n32485) );
  NOR U33484 ( .A(n33285), .B(n33286), .Z(n33283) );
  XNOR U33485 ( .A(n33287), .B(n33288), .Z(n32818) );
  ANDN U33486 ( .B(n33289), .A(n33290), .Z(n33287) );
  XOR U33487 ( .A(n33291), .B(n33292), .Z(n31644) );
  XNOR U33488 ( .A(n25169), .B(n25866), .Z(n33292) );
  XOR U33489 ( .A(n33293), .B(n29855), .Z(n25866) );
  XOR U33490 ( .A(n28428), .B(n33294), .Z(n29855) );
  IV U33491 ( .A(n33295), .Z(n28428) );
  ANDN U33492 ( .B(n26684), .A(n26682), .Z(n33293) );
  IV U33493 ( .A(n29856), .Z(n26682) );
  XNOR U33494 ( .A(n28762), .B(n33296), .Z(n29856) );
  XOR U33495 ( .A(n33297), .B(n33298), .Z(n28762) );
  IV U33496 ( .A(n27715), .Z(n26684) );
  XOR U33497 ( .A(n33299), .B(n31233), .Z(n27715) );
  XOR U33498 ( .A(n33300), .B(n28333), .Z(n25169) );
  XOR U33499 ( .A(n33301), .B(n30219), .Z(n28333) );
  NOR U33500 ( .A(n26677), .B(n26676), .Z(n33300) );
  XOR U33501 ( .A(n33302), .B(n33303), .Z(n26676) );
  XOR U33502 ( .A(n33304), .B(n32032), .Z(n26677) );
  IV U33503 ( .A(n29734), .Z(n32032) );
  XOR U33504 ( .A(n28324), .B(n33305), .Z(n33291) );
  XNOR U33505 ( .A(n24407), .B(n26581), .Z(n33305) );
  XNOR U33506 ( .A(n33306), .B(n28329), .Z(n26581) );
  XOR U33507 ( .A(n31238), .B(n33307), .Z(n28329) );
  XOR U33508 ( .A(n32930), .B(n33308), .Z(n31238) );
  XOR U33509 ( .A(n33309), .B(n33310), .Z(n32930) );
  XNOR U33510 ( .A(n31554), .B(n33311), .Z(n33310) );
  XOR U33511 ( .A(n33312), .B(n33313), .Z(n31554) );
  XNOR U33512 ( .A(n33316), .B(n33317), .Z(n33309) );
  XNOR U33513 ( .A(n32165), .B(n33318), .Z(n33317) );
  XNOR U33514 ( .A(n33319), .B(n33320), .Z(n32165) );
  ANDN U33515 ( .B(n33321), .A(n33322), .Z(n33319) );
  ANDN U33516 ( .B(n26686), .A(n26688), .Z(n33306) );
  XNOR U33517 ( .A(n33323), .B(n32583), .Z(n26688) );
  XNOR U33518 ( .A(n33324), .B(n32053), .Z(n26686) );
  XNOR U33519 ( .A(n33325), .B(n31920), .Z(n24407) );
  XNOR U33520 ( .A(n33326), .B(n30215), .Z(n31920) );
  XNOR U33521 ( .A(n28995), .B(n33327), .Z(n31921) );
  IV U33522 ( .A(n27718), .Z(n33225) );
  XNOR U33523 ( .A(n33330), .B(n29032), .Z(n27718) );
  XNOR U33524 ( .A(n33331), .B(n32535), .Z(n29032) );
  XNOR U33525 ( .A(n33332), .B(n33333), .Z(n32535) );
  XOR U33526 ( .A(n31308), .B(n30656), .Z(n33333) );
  XOR U33527 ( .A(n33334), .B(n33335), .Z(n30656) );
  ANDN U33528 ( .B(n33336), .A(n33337), .Z(n33334) );
  XNOR U33529 ( .A(n33338), .B(n33339), .Z(n31308) );
  AND U33530 ( .A(n33340), .B(n33341), .Z(n33338) );
  XOR U33531 ( .A(n30228), .B(n33342), .Z(n33332) );
  XNOR U33532 ( .A(n32183), .B(n31889), .Z(n33342) );
  XNOR U33533 ( .A(n33343), .B(n33344), .Z(n31889) );
  ANDN U33534 ( .B(n33345), .A(n33346), .Z(n33343) );
  XOR U33535 ( .A(n33347), .B(n33348), .Z(n32183) );
  NOR U33536 ( .A(n33349), .B(n33350), .Z(n33347) );
  XNOR U33537 ( .A(n33351), .B(n33352), .Z(n30228) );
  NOR U33538 ( .A(n33353), .B(n33354), .Z(n33351) );
  XNOR U33539 ( .A(n33355), .B(n28335), .Z(n28324) );
  XNOR U33540 ( .A(n32622), .B(n33356), .Z(n28335) );
  ANDN U33541 ( .B(n27232), .A(n27230), .Z(n33355) );
  XNOR U33542 ( .A(n33357), .B(n30230), .Z(n27230) );
  XOR U33543 ( .A(n33358), .B(n33359), .Z(n27232) );
  XOR U33544 ( .A(n31508), .B(n25224), .Z(n25141) );
  IV U33545 ( .A(n25109), .Z(n25224) );
  XOR U33546 ( .A(n33360), .B(n33361), .Z(n30725) );
  XOR U33547 ( .A(n25485), .B(n25064), .Z(n33361) );
  XNOR U33548 ( .A(n33362), .B(n30457), .Z(n25064) );
  AND U33549 ( .A(n31511), .B(n31510), .Z(n33362) );
  XNOR U33550 ( .A(n29968), .B(n33366), .Z(n31510) );
  IV U33551 ( .A(n30248), .Z(n29968) );
  XOR U33552 ( .A(n33369), .B(n30639), .Z(n25485) );
  XOR U33553 ( .A(n33265), .B(n33370), .Z(n30639) );
  ANDN U33554 ( .B(n31514), .A(n33371), .Z(n33369) );
  XOR U33555 ( .A(n33372), .B(n30039), .Z(n31514) );
  XNOR U33556 ( .A(n32322), .B(n33373), .Z(n33360) );
  XNOR U33557 ( .A(n24824), .B(n27737), .Z(n33373) );
  XNOR U33558 ( .A(n33374), .B(n32327), .Z(n27737) );
  IV U33559 ( .A(n30443), .Z(n32327) );
  XOR U33560 ( .A(n33375), .B(n32205), .Z(n30443) );
  XOR U33561 ( .A(n33376), .B(n33377), .Z(n32205) );
  ANDN U33562 ( .B(n33378), .A(n32326), .Z(n33374) );
  XOR U33563 ( .A(n33380), .B(n30743), .Z(n30447) );
  AND U33564 ( .A(n31503), .B(n31502), .Z(n33379) );
  XOR U33565 ( .A(n33381), .B(n33382), .Z(n31502) );
  XOR U33566 ( .A(n33383), .B(n30453), .Z(n32322) );
  XOR U33567 ( .A(n33384), .B(n27947), .Z(n30453) );
  ANDN U33568 ( .B(n31505), .A(n31506), .Z(n33383) );
  XNOR U33569 ( .A(n33385), .B(n30784), .Z(n31505) );
  XOR U33570 ( .A(n33387), .B(n33388), .Z(n32742) );
  XNOR U33571 ( .A(n33389), .B(n28797), .Z(n33388) );
  XNOR U33572 ( .A(n33390), .B(n33391), .Z(n28797) );
  NOR U33573 ( .A(n33392), .B(n33393), .Z(n33390) );
  XOR U33574 ( .A(n30504), .B(n33394), .Z(n33387) );
  XOR U33575 ( .A(n33395), .B(n31978), .Z(n33394) );
  XNOR U33576 ( .A(n33396), .B(n33397), .Z(n31978) );
  ANDN U33577 ( .B(n33398), .A(n33399), .Z(n33396) );
  XNOR U33578 ( .A(n33400), .B(n33401), .Z(n30504) );
  NOR U33579 ( .A(n33402), .B(n33403), .Z(n33400) );
  XOR U33580 ( .A(n33404), .B(n33405), .Z(n28159) );
  XOR U33581 ( .A(n27953), .B(n24479), .Z(n33405) );
  XNOR U33582 ( .A(n33406), .B(n30477), .Z(n24479) );
  XNOR U33583 ( .A(n31190), .B(n33407), .Z(n30477) );
  AND U33584 ( .A(n30091), .B(n30093), .Z(n33406) );
  XOR U33585 ( .A(n33408), .B(n32625), .Z(n30093) );
  XOR U33586 ( .A(n33409), .B(n33053), .Z(n30091) );
  IV U33587 ( .A(n31348), .Z(n33053) );
  XOR U33588 ( .A(n33410), .B(n30463), .Z(n27953) );
  XNOR U33589 ( .A(n33411), .B(n28814), .Z(n30463) );
  ANDN U33590 ( .B(n30095), .A(n30096), .Z(n33410) );
  XOR U33591 ( .A(n33413), .B(n31539), .Z(n30095) );
  XOR U33592 ( .A(n24752), .B(n33414), .Z(n33404) );
  XOR U33593 ( .A(n24075), .B(n22830), .Z(n33414) );
  XNOR U33594 ( .A(n33415), .B(n30469), .Z(n22830) );
  XOR U33595 ( .A(n32662), .B(n30517), .Z(n30469) );
  XNOR U33596 ( .A(n33416), .B(n33417), .Z(n32662) );
  ANDN U33597 ( .B(n33418), .A(n33419), .Z(n33416) );
  ANDN U33598 ( .B(n30084), .A(n30082), .Z(n33415) );
  XOR U33599 ( .A(n32109), .B(n33420), .Z(n30082) );
  IV U33600 ( .A(n32806), .Z(n32109) );
  XOR U33601 ( .A(n33422), .B(n33423), .Z(n32931) );
  XOR U33602 ( .A(n31999), .B(n29074), .Z(n33423) );
  XOR U33603 ( .A(n33424), .B(n33425), .Z(n29074) );
  NOR U33604 ( .A(n33426), .B(n33427), .Z(n33424) );
  XNOR U33605 ( .A(n33428), .B(n33429), .Z(n31999) );
  ANDN U33606 ( .B(n33430), .A(n33431), .Z(n33428) );
  XOR U33607 ( .A(n32479), .B(n33432), .Z(n33422) );
  XOR U33608 ( .A(n33433), .B(n32036), .Z(n33432) );
  XNOR U33609 ( .A(n33434), .B(n33435), .Z(n32036) );
  ANDN U33610 ( .B(n33436), .A(n33437), .Z(n33434) );
  XNOR U33611 ( .A(n33438), .B(n33439), .Z(n32479) );
  ANDN U33612 ( .B(n33440), .A(n33441), .Z(n33438) );
  XNOR U33613 ( .A(n30903), .B(n33442), .Z(n30084) );
  XNOR U33614 ( .A(n33443), .B(n30473), .Z(n24075) );
  XOR U33615 ( .A(n32232), .B(n33444), .Z(n30473) );
  IV U33616 ( .A(n32571), .Z(n32232) );
  ANDN U33617 ( .B(n30086), .A(n30088), .Z(n33443) );
  XOR U33618 ( .A(n33446), .B(n33447), .Z(n30066) );
  XNOR U33619 ( .A(n33448), .B(n31434), .Z(n30086) );
  XNOR U33620 ( .A(n33451), .B(n30465), .Z(n24752) );
  XOR U33621 ( .A(n33452), .B(n30175), .Z(n30465) );
  IV U33622 ( .A(n31887), .Z(n30175) );
  XNOR U33623 ( .A(n33453), .B(n33454), .Z(n31887) );
  AND U33624 ( .A(n30101), .B(n30099), .Z(n33451) );
  XNOR U33625 ( .A(n33455), .B(n33456), .Z(n30099) );
  XOR U33626 ( .A(n33311), .B(n32166), .Z(n30101) );
  XNOR U33627 ( .A(n33457), .B(n33458), .Z(n33311) );
  ANDN U33628 ( .B(n33459), .A(n33460), .Z(n33457) );
  XOR U33629 ( .A(n33461), .B(n32326), .Z(n31508) );
  XOR U33630 ( .A(n32389), .B(n33462), .Z(n32326) );
  IV U33631 ( .A(n32480), .Z(n32389) );
  XOR U33632 ( .A(n33463), .B(n33464), .Z(n32480) );
  NOR U33633 ( .A(n30441), .B(n33378), .Z(n33461) );
  XNOR U33634 ( .A(n33465), .B(n20803), .Z(n19562) );
  XOR U33635 ( .A(n23066), .B(n27987), .Z(n20803) );
  XNOR U33636 ( .A(n33466), .B(n31498), .Z(n27987) );
  ANDN U33637 ( .B(n32784), .A(n32785), .Z(n33466) );
  IV U33638 ( .A(n26283), .Z(n23066) );
  XNOR U33639 ( .A(n31075), .B(n30640), .Z(n26283) );
  XOR U33640 ( .A(n33467), .B(n33468), .Z(n30640) );
  XNOR U33641 ( .A(n27096), .B(n24756), .Z(n33468) );
  XNOR U33642 ( .A(n33469), .B(n31503), .Z(n24756) );
  XOR U33643 ( .A(n30536), .B(n33470), .Z(n31503) );
  ANDN U33644 ( .B(n30445), .A(n30446), .Z(n33469) );
  XNOR U33645 ( .A(n33471), .B(n33359), .Z(n30446) );
  XOR U33646 ( .A(n31005), .B(n33472), .Z(n30445) );
  XOR U33647 ( .A(n33473), .B(n31506), .Z(n27096) );
  XNOR U33648 ( .A(n33474), .B(n30210), .Z(n31506) );
  ANDN U33649 ( .B(n30451), .A(n30452), .Z(n33473) );
  XOR U33650 ( .A(n33475), .B(n32887), .Z(n30452) );
  IV U33651 ( .A(n32064), .Z(n32887) );
  XOR U33652 ( .A(n31570), .B(n33078), .Z(n30451) );
  XNOR U33653 ( .A(n33478), .B(n33479), .Z(n33078) );
  NOR U33654 ( .A(n33480), .B(n33481), .Z(n33478) );
  XNOR U33655 ( .A(n28541), .B(n33482), .Z(n33467) );
  XOR U33656 ( .A(n23736), .B(n25155), .Z(n33482) );
  XNOR U33657 ( .A(n33483), .B(n31515), .Z(n25155) );
  IV U33658 ( .A(n33371), .Z(n31515) );
  XOR U33659 ( .A(n33484), .B(n32498), .Z(n33371) );
  XNOR U33660 ( .A(n33485), .B(n28473), .Z(n30637) );
  IV U33661 ( .A(n30125), .Z(n28473) );
  XOR U33662 ( .A(n33488), .B(n31068), .Z(n30638) );
  XNOR U33663 ( .A(n33491), .B(n33378), .Z(n23736) );
  XNOR U33664 ( .A(n33492), .B(n28825), .Z(n33378) );
  XOR U33665 ( .A(n33494), .B(n33495), .Z(n32970) );
  XOR U33666 ( .A(n30270), .B(n32238), .Z(n33495) );
  XNOR U33667 ( .A(n33496), .B(n33497), .Z(n32238) );
  ANDN U33668 ( .B(n32661), .A(n33498), .Z(n33496) );
  XNOR U33669 ( .A(n33499), .B(n32656), .Z(n30270) );
  ANDN U33670 ( .B(n32657), .A(n33500), .Z(n33499) );
  XNOR U33671 ( .A(n30901), .B(n33501), .Z(n33494) );
  XNOR U33672 ( .A(n29056), .B(n28749), .Z(n33501) );
  XOR U33673 ( .A(n33502), .B(n33503), .Z(n28749) );
  ANDN U33674 ( .B(n33504), .A(n33505), .Z(n33502) );
  XNOR U33675 ( .A(n33506), .B(n32674), .Z(n29056) );
  ANDN U33676 ( .B(n32673), .A(n33507), .Z(n33506) );
  XNOR U33677 ( .A(n33508), .B(n33419), .Z(n30901) );
  ANDN U33678 ( .B(n33509), .A(n33418), .Z(n33508) );
  ANDN U33679 ( .B(n30441), .A(n30442), .Z(n33491) );
  XNOR U33680 ( .A(n33510), .B(n30539), .Z(n30442) );
  XNOR U33681 ( .A(n33511), .B(n30764), .Z(n30441) );
  XNOR U33682 ( .A(n33514), .B(n31511), .Z(n28541) );
  XOR U33683 ( .A(n33515), .B(n31219), .Z(n31511) );
  ANDN U33684 ( .B(n30456), .A(n31512), .Z(n33514) );
  XNOR U33685 ( .A(n33516), .B(n30371), .Z(n31512) );
  XOR U33686 ( .A(n33517), .B(n32829), .Z(n30456) );
  XOR U33687 ( .A(n33518), .B(n33519), .Z(n31075) );
  XNOR U33688 ( .A(n25254), .B(n25349), .Z(n33519) );
  XOR U33689 ( .A(n33520), .B(n31497), .Z(n25349) );
  ANDN U33690 ( .B(n31498), .A(n32784), .Z(n33520) );
  XOR U33691 ( .A(n29943), .B(n33521), .Z(n32784) );
  XOR U33692 ( .A(n33522), .B(n31178), .Z(n31498) );
  XOR U33693 ( .A(n33523), .B(n31483), .Z(n25254) );
  ANDN U33694 ( .B(n28000), .A(n27999), .Z(n33523) );
  XNOR U33695 ( .A(n32368), .B(n33524), .Z(n27999) );
  XNOR U33696 ( .A(n33525), .B(n32456), .Z(n28000) );
  XNOR U33697 ( .A(n31478), .B(n33526), .Z(n33518) );
  XNOR U33698 ( .A(n26474), .B(n27235), .Z(n33526) );
  XOR U33699 ( .A(n33527), .B(n33528), .Z(n27235) );
  NOR U33700 ( .A(n27995), .B(n27996), .Z(n33527) );
  XNOR U33701 ( .A(n29528), .B(n33529), .Z(n27996) );
  XOR U33702 ( .A(n33530), .B(n33531), .Z(n27995) );
  XNOR U33703 ( .A(n33532), .B(n31486), .Z(n26474) );
  ANDN U33704 ( .B(n31487), .A(n32776), .Z(n33532) );
  IV U33705 ( .A(n31917), .Z(n32776) );
  XNOR U33706 ( .A(n33533), .B(n31448), .Z(n31917) );
  XNOR U33707 ( .A(n31618), .B(n33534), .Z(n31487) );
  XOR U33708 ( .A(n33535), .B(n31491), .Z(n31478) );
  NOR U33709 ( .A(n27991), .B(n27992), .Z(n33535) );
  XOR U33710 ( .A(n31666), .B(n33536), .Z(n27992) );
  XNOR U33711 ( .A(n33537), .B(n30507), .Z(n27991) );
  XNOR U33712 ( .A(n23831), .B(n31720), .Z(n25135) );
  XNOR U33713 ( .A(n33540), .B(n32075), .Z(n31720) );
  ANDN U33714 ( .B(n27208), .A(n27209), .Z(n33540) );
  XOR U33715 ( .A(n33541), .B(n32972), .Z(n27209) );
  XNOR U33716 ( .A(n27848), .B(n28714), .Z(n23831) );
  XNOR U33717 ( .A(n33542), .B(n33543), .Z(n28714) );
  XOR U33718 ( .A(n32048), .B(n25768), .Z(n33543) );
  XOR U33719 ( .A(n33544), .B(n32077), .Z(n25768) );
  XOR U33720 ( .A(n33318), .B(n32166), .Z(n32077) );
  XNOR U33721 ( .A(n33545), .B(n33546), .Z(n33318) );
  ANDN U33722 ( .B(n33547), .A(n33548), .Z(n33545) );
  ANDN U33723 ( .B(n31726), .A(n31725), .Z(n33544) );
  XOR U33724 ( .A(n33549), .B(n28425), .Z(n31725) );
  IV U33725 ( .A(n33550), .Z(n28425) );
  IV U33726 ( .A(n29908), .Z(n31726) );
  XOR U33727 ( .A(n33551), .B(n33552), .Z(n29908) );
  XNOR U33728 ( .A(n33553), .B(n32080), .Z(n32048) );
  XOR U33729 ( .A(n33554), .B(n32644), .Z(n32080) );
  ANDN U33730 ( .B(n31719), .A(n27212), .Z(n33553) );
  XNOR U33731 ( .A(n33555), .B(n32583), .Z(n27212) );
  XNOR U33732 ( .A(n33556), .B(n27937), .Z(n31719) );
  XNOR U33733 ( .A(n26222), .B(n33557), .Z(n33542) );
  XNOR U33734 ( .A(n24883), .B(n24030), .Z(n33557) );
  XNOR U33735 ( .A(n33558), .B(n32071), .Z(n24030) );
  XOR U33736 ( .A(n33559), .B(n27944), .Z(n32071) );
  IV U33737 ( .A(n30219), .Z(n27944) );
  XOR U33738 ( .A(n33367), .B(n33476), .Z(n30219) );
  XNOR U33739 ( .A(n33560), .B(n33561), .Z(n33476) );
  XNOR U33740 ( .A(n32792), .B(n32912), .Z(n33561) );
  XOR U33741 ( .A(n33562), .B(n33563), .Z(n32912) );
  ANDN U33742 ( .B(n33564), .A(n33565), .Z(n33562) );
  XOR U33743 ( .A(n33566), .B(n33567), .Z(n32792) );
  AND U33744 ( .A(n33568), .B(n33569), .Z(n33566) );
  XOR U33745 ( .A(n32688), .B(n33570), .Z(n33560) );
  XNOR U33746 ( .A(n32584), .B(n32922), .Z(n33570) );
  XNOR U33747 ( .A(n33571), .B(n33572), .Z(n32922) );
  AND U33748 ( .A(n33573), .B(n33574), .Z(n33571) );
  XOR U33749 ( .A(n33575), .B(n33576), .Z(n32584) );
  ANDN U33750 ( .B(n33577), .A(n33578), .Z(n33575) );
  XNOR U33751 ( .A(n33579), .B(n33580), .Z(n32688) );
  AND U33752 ( .A(n33581), .B(n33582), .Z(n33579) );
  XOR U33753 ( .A(n33583), .B(n33584), .Z(n33367) );
  XNOR U33754 ( .A(n31115), .B(n33585), .Z(n33584) );
  XNOR U33755 ( .A(n33586), .B(n33587), .Z(n31115) );
  ANDN U33756 ( .B(n33588), .A(n33589), .Z(n33586) );
  XOR U33757 ( .A(n33590), .B(n33591), .Z(n33583) );
  XNOR U33758 ( .A(n33592), .B(n30696), .Z(n33591) );
  XNOR U33759 ( .A(n33593), .B(n33594), .Z(n30696) );
  NOR U33760 ( .A(n33595), .B(n33596), .Z(n33593) );
  AND U33761 ( .A(n27218), .B(n31717), .Z(n33558) );
  XOR U33762 ( .A(n33597), .B(n31535), .Z(n31717) );
  IV U33763 ( .A(n32015), .Z(n31535) );
  XNOR U33764 ( .A(n33598), .B(n33599), .Z(n32015) );
  XOR U33765 ( .A(n33600), .B(n32891), .Z(n27218) );
  XNOR U33766 ( .A(n33601), .B(n32074), .Z(n24883) );
  XOR U33767 ( .A(n29930), .B(n33602), .Z(n32074) );
  XNOR U33768 ( .A(n33603), .B(n33604), .Z(n29930) );
  XOR U33769 ( .A(n28803), .B(n33605), .Z(n27208) );
  XNOR U33770 ( .A(n29324), .B(n33606), .Z(n32075) );
  XOR U33771 ( .A(n33607), .B(n32068), .Z(n26222) );
  XOR U33772 ( .A(n33608), .B(n31687), .Z(n32068) );
  ANDN U33773 ( .B(n31723), .A(n27222), .Z(n33607) );
  XNOR U33774 ( .A(n33609), .B(n30535), .Z(n27222) );
  XOR U33775 ( .A(n33463), .B(n33610), .Z(n30535) );
  XOR U33776 ( .A(n33611), .B(n33612), .Z(n33463) );
  XOR U33777 ( .A(n31099), .B(n33613), .Z(n33612) );
  XNOR U33778 ( .A(n33614), .B(n33615), .Z(n31099) );
  AND U33779 ( .A(n33616), .B(n33617), .Z(n33614) );
  XNOR U33780 ( .A(n31153), .B(n33618), .Z(n33611) );
  XOR U33781 ( .A(n32457), .B(n33619), .Z(n33618) );
  XOR U33782 ( .A(n33620), .B(n33621), .Z(n32457) );
  ANDN U33783 ( .B(n33622), .A(n33623), .Z(n33620) );
  XNOR U33784 ( .A(n33624), .B(n33625), .Z(n31153) );
  ANDN U33785 ( .B(n33626), .A(n33627), .Z(n33624) );
  XOR U33786 ( .A(n32117), .B(n33628), .Z(n31723) );
  XOR U33787 ( .A(n33629), .B(n33630), .Z(n27848) );
  XOR U33788 ( .A(n24660), .B(n24236), .Z(n33630) );
  XOR U33789 ( .A(n33631), .B(n31747), .Z(n24236) );
  XNOR U33790 ( .A(n33632), .B(n32175), .Z(n31747) );
  XNOR U33791 ( .A(n33633), .B(n33634), .Z(n32175) );
  NOR U33792 ( .A(n32056), .B(n29905), .Z(n33631) );
  XNOR U33793 ( .A(n33635), .B(n32248), .Z(n29905) );
  XNOR U33794 ( .A(n33636), .B(n28739), .Z(n32056) );
  XNOR U33795 ( .A(n33637), .B(n31740), .Z(n24660) );
  XNOR U33796 ( .A(n32101), .B(n33638), .Z(n31740) );
  NOR U33797 ( .A(n30054), .B(n29891), .Z(n33637) );
  XOR U33798 ( .A(n30911), .B(n33639), .Z(n29891) );
  XOR U33799 ( .A(n33640), .B(n30586), .Z(n30054) );
  IV U33800 ( .A(n30211), .Z(n30586) );
  XOR U33801 ( .A(n33641), .B(n33642), .Z(n30211) );
  XOR U33802 ( .A(n27069), .B(n33643), .Z(n33629) );
  XOR U33803 ( .A(n25088), .B(n26562), .Z(n33643) );
  XNOR U33804 ( .A(n33644), .B(n31744), .Z(n26562) );
  XNOR U33805 ( .A(n33645), .B(n30748), .Z(n31744) );
  ANDN U33806 ( .B(n29887), .A(n29888), .Z(n33644) );
  XOR U33807 ( .A(n33646), .B(n32117), .Z(n29888) );
  IV U33808 ( .A(n31394), .Z(n32117) );
  XOR U33809 ( .A(n33647), .B(n33368), .Z(n31394) );
  XNOR U33810 ( .A(n33648), .B(n33649), .Z(n33368) );
  XNOR U33811 ( .A(n27948), .B(n29322), .Z(n33649) );
  XNOR U33812 ( .A(n33650), .B(n33651), .Z(n29322) );
  XNOR U33813 ( .A(n33654), .B(n33655), .Z(n27948) );
  ANDN U33814 ( .B(n33656), .A(n33657), .Z(n33654) );
  XOR U33815 ( .A(n32095), .B(n33658), .Z(n33648) );
  XOR U33816 ( .A(n31675), .B(n33659), .Z(n33658) );
  XNOR U33817 ( .A(n33660), .B(n33661), .Z(n31675) );
  XNOR U33818 ( .A(n33664), .B(n33665), .Z(n32095) );
  NOR U33819 ( .A(n33666), .B(n33667), .Z(n33664) );
  XOR U33820 ( .A(n31005), .B(n33668), .Z(n29887) );
  IV U33821 ( .A(n31955), .Z(n31005) );
  XNOR U33822 ( .A(n33669), .B(n33670), .Z(n31955) );
  XOR U33823 ( .A(n33671), .B(n31736), .Z(n25088) );
  XOR U33824 ( .A(n33672), .B(n32743), .Z(n31736) );
  NOR U33825 ( .A(n29897), .B(n29896), .Z(n33671) );
  XNOR U33826 ( .A(n33673), .B(n31754), .Z(n29896) );
  IV U33827 ( .A(n30822), .Z(n31754) );
  XOR U33828 ( .A(n33674), .B(n28803), .Z(n29897) );
  XNOR U33829 ( .A(n32544), .B(n33675), .Z(n28803) );
  XOR U33830 ( .A(n33676), .B(n33677), .Z(n32544) );
  XNOR U33831 ( .A(n32311), .B(n33678), .Z(n33677) );
  XNOR U33832 ( .A(n33679), .B(n33680), .Z(n32311) );
  ANDN U33833 ( .B(n33681), .A(n33682), .Z(n33679) );
  XOR U33834 ( .A(n30499), .B(n33683), .Z(n33676) );
  XOR U33835 ( .A(n32578), .B(n31021), .Z(n33683) );
  XOR U33836 ( .A(n33684), .B(n33685), .Z(n31021) );
  AND U33837 ( .A(n33686), .B(n33687), .Z(n33684) );
  XNOR U33838 ( .A(n33688), .B(n33689), .Z(n32578) );
  ANDN U33839 ( .B(n33690), .A(n33691), .Z(n33688) );
  XOR U33840 ( .A(n33692), .B(n33693), .Z(n30499) );
  XNOR U33841 ( .A(n33696), .B(n31751), .Z(n27069) );
  XOR U33842 ( .A(n33697), .B(n31810), .Z(n31751) );
  IV U33843 ( .A(n33698), .Z(n31810) );
  NOR U33844 ( .A(n29902), .B(n29900), .Z(n33696) );
  XNOR U33845 ( .A(n33699), .B(n32235), .Z(n29900) );
  XNOR U33846 ( .A(n31026), .B(n33700), .Z(n29902) );
  XOR U33847 ( .A(n33701), .B(n33702), .Z(n31026) );
  XOR U33848 ( .A(n24423), .B(n31609), .Z(n23225) );
  XNOR U33849 ( .A(n33703), .B(n32772), .Z(n31609) );
  ANDN U33850 ( .B(n31088), .A(n30836), .Z(n33703) );
  XNOR U33851 ( .A(n30961), .B(n33704), .Z(n30836) );
  XNOR U33852 ( .A(n30319), .B(n30724), .Z(n24423) );
  XNOR U33853 ( .A(n33705), .B(n33706), .Z(n30724) );
  XOR U33854 ( .A(n26705), .B(n25265), .Z(n33706) );
  XOR U33855 ( .A(n33707), .B(n27997), .Z(n25265) );
  XOR U33856 ( .A(n33708), .B(n32602), .Z(n27997) );
  XOR U33857 ( .A(n33709), .B(n33710), .Z(n32602) );
  ANDN U33858 ( .B(n31494), .A(n31493), .Z(n33707) );
  IV U33859 ( .A(n32782), .Z(n31493) );
  XOR U33860 ( .A(n33711), .B(n33382), .Z(n32782) );
  IV U33861 ( .A(n33528), .Z(n31494) );
  XNOR U33862 ( .A(n31405), .B(n33712), .Z(n33528) );
  XOR U33863 ( .A(n33713), .B(n33714), .Z(n31405) );
  XNOR U33864 ( .A(n33715), .B(n31916), .Z(n26705) );
  XOR U33865 ( .A(n33716), .B(n30215), .Z(n31916) );
  ANDN U33866 ( .B(n31486), .A(n31485), .Z(n33715) );
  XNOR U33867 ( .A(n33719), .B(n27947), .Z(n31485) );
  XOR U33868 ( .A(n33720), .B(n33721), .Z(n31486) );
  XNOR U33869 ( .A(n23613), .B(n33722), .Z(n33705) );
  XOR U33870 ( .A(n22230), .B(n30932), .Z(n33722) );
  XOR U33871 ( .A(n33723), .B(n28001), .Z(n30932) );
  XOR U33872 ( .A(n33585), .B(n31116), .Z(n28001) );
  XOR U33873 ( .A(n33724), .B(n33725), .Z(n33585) );
  NOR U33874 ( .A(n33726), .B(n33727), .Z(n33724) );
  ANDN U33875 ( .B(n31482), .A(n31483), .Z(n33723) );
  XNOR U33876 ( .A(n33728), .B(n28462), .Z(n31483) );
  XOR U33877 ( .A(n33729), .B(n30990), .Z(n31482) );
  IV U33878 ( .A(n31250), .Z(n30990) );
  XOR U33879 ( .A(n33730), .B(n33731), .Z(n31250) );
  XOR U33880 ( .A(n33732), .B(n27993), .Z(n22230) );
  IV U33881 ( .A(n32778), .Z(n27993) );
  XOR U33882 ( .A(n33733), .B(n30559), .Z(n32778) );
  ANDN U33883 ( .B(n31490), .A(n31491), .Z(n33732) );
  XOR U33884 ( .A(n31364), .B(n33734), .Z(n31491) );
  IV U33885 ( .A(n31613), .Z(n31364) );
  XOR U33886 ( .A(n33735), .B(n33736), .Z(n31613) );
  XOR U33887 ( .A(n33737), .B(n33550), .Z(n31490) );
  XOR U33888 ( .A(n33738), .B(n32785), .Z(n23613) );
  XOR U33889 ( .A(n33739), .B(n30039), .Z(n32785) );
  NOR U33890 ( .A(n32786), .B(n31497), .Z(n33738) );
  XNOR U33891 ( .A(n30247), .B(n33740), .Z(n31497) );
  XOR U33892 ( .A(n31455), .B(n33741), .Z(n32786) );
  IV U33893 ( .A(n32768), .Z(n31455) );
  XOR U33894 ( .A(n33701), .B(n33742), .Z(n32768) );
  XOR U33895 ( .A(n33743), .B(n33744), .Z(n33701) );
  XNOR U33896 ( .A(n32014), .B(n33597), .Z(n33744) );
  XOR U33897 ( .A(n33745), .B(n33746), .Z(n33597) );
  ANDN U33898 ( .B(n33747), .A(n33748), .Z(n33745) );
  XNOR U33899 ( .A(n33749), .B(n33750), .Z(n32014) );
  NOR U33900 ( .A(n33751), .B(n33752), .Z(n33749) );
  XOR U33901 ( .A(n32004), .B(n33753), .Z(n33743) );
  XOR U33902 ( .A(n31534), .B(n32734), .Z(n33753) );
  XNOR U33903 ( .A(n33754), .B(n33755), .Z(n32734) );
  ANDN U33904 ( .B(n33756), .A(n33757), .Z(n33754) );
  XNOR U33905 ( .A(n33758), .B(n33759), .Z(n31534) );
  NOR U33906 ( .A(n33760), .B(n33761), .Z(n33758) );
  XNOR U33907 ( .A(n33762), .B(n33763), .Z(n32004) );
  ANDN U33908 ( .B(n33764), .A(n33765), .Z(n33762) );
  XOR U33909 ( .A(n33766), .B(n33767), .Z(n30319) );
  XNOR U33910 ( .A(n28781), .B(n27882), .Z(n33767) );
  XOR U33911 ( .A(n33768), .B(n30833), .Z(n27882) );
  XOR U33912 ( .A(n32705), .B(n33769), .Z(n30833) );
  NOR U33913 ( .A(n32769), .B(n31081), .Z(n33768) );
  XNOR U33914 ( .A(n30148), .B(n33770), .Z(n31081) );
  XNOR U33915 ( .A(n33771), .B(n33772), .Z(n30148) );
  IV U33916 ( .A(n31611), .Z(n32769) );
  XOR U33917 ( .A(n31459), .B(n33773), .Z(n31611) );
  XNOR U33918 ( .A(n33774), .B(n30837), .Z(n28781) );
  XOR U33919 ( .A(n33775), .B(n32306), .Z(n30837) );
  IV U33920 ( .A(n31840), .Z(n32306) );
  NOR U33921 ( .A(n32772), .B(n31088), .Z(n33774) );
  XNOR U33922 ( .A(n33776), .B(n30531), .Z(n31088) );
  XOR U33923 ( .A(n33777), .B(n33539), .Z(n30531) );
  XOR U33924 ( .A(n33778), .B(n33779), .Z(n33539) );
  XNOR U33925 ( .A(n29066), .B(n31212), .Z(n33779) );
  XNOR U33926 ( .A(n33780), .B(n33781), .Z(n31212) );
  NOR U33927 ( .A(n33782), .B(n33783), .Z(n33780) );
  XNOR U33928 ( .A(n33784), .B(n33393), .Z(n29066) );
  ANDN U33929 ( .B(n33785), .A(n33786), .Z(n33784) );
  XOR U33930 ( .A(n32350), .B(n33787), .Z(n33778) );
  XOR U33931 ( .A(n29971), .B(n32863), .Z(n33787) );
  XNOR U33932 ( .A(n33788), .B(n33402), .Z(n32863) );
  NOR U33933 ( .A(n33789), .B(n33790), .Z(n33788) );
  XOR U33934 ( .A(n33791), .B(n33792), .Z(n29971) );
  NOR U33935 ( .A(n33793), .B(n33794), .Z(n33791) );
  XNOR U33936 ( .A(n33795), .B(n33399), .Z(n32350) );
  NOR U33937 ( .A(n33796), .B(n33797), .Z(n33795) );
  XOR U33938 ( .A(n33798), .B(n31698), .Z(n32772) );
  XOR U33939 ( .A(n26452), .B(n33799), .Z(n33766) );
  XOR U33940 ( .A(n32756), .B(n26090), .Z(n33799) );
  XNOR U33941 ( .A(n33800), .B(n30841), .Z(n26090) );
  XNOR U33942 ( .A(n33801), .B(n29161), .Z(n30841) );
  IV U33943 ( .A(n30541), .Z(n29161) );
  XNOR U33944 ( .A(n33802), .B(n33633), .Z(n30541) );
  XOR U33945 ( .A(n33803), .B(n33804), .Z(n33633) );
  XNOR U33946 ( .A(n33805), .B(n33806), .Z(n33804) );
  XOR U33947 ( .A(n28768), .B(n33807), .Z(n33803) );
  XOR U33948 ( .A(n33808), .B(n32215), .Z(n33807) );
  XNOR U33949 ( .A(n33809), .B(n33286), .Z(n32215) );
  NOR U33950 ( .A(n33810), .B(n33811), .Z(n33809) );
  XNOR U33951 ( .A(n33812), .B(n33813), .Z(n28768) );
  ANDN U33952 ( .B(n33814), .A(n33815), .Z(n33812) );
  ANDN U33953 ( .B(n31079), .A(n31616), .Z(n33800) );
  XOR U33954 ( .A(n33816), .B(n30239), .Z(n31616) );
  XNOR U33955 ( .A(n33817), .B(n32044), .Z(n31079) );
  XNOR U33956 ( .A(n33818), .B(n30846), .Z(n32756) );
  XOR U33957 ( .A(n33819), .B(n33820), .Z(n30846) );
  ANDN U33958 ( .B(n31620), .A(n31090), .Z(n33818) );
  XOR U33959 ( .A(n32368), .B(n33821), .Z(n31090) );
  IV U33960 ( .A(n32743), .Z(n32368) );
  XOR U33961 ( .A(n33822), .B(n33823), .Z(n32743) );
  XNOR U33962 ( .A(n30644), .B(n33824), .Z(n31620) );
  XNOR U33963 ( .A(n33825), .B(n31092), .Z(n26452) );
  XOR U33964 ( .A(n33551), .B(n33826), .Z(n31092) );
  NOR U33965 ( .A(n31624), .B(n31084), .Z(n33825) );
  XOR U33966 ( .A(n33827), .B(n33828), .Z(n31084) );
  XOR U33967 ( .A(n33829), .B(n31542), .Z(n31624) );
  XNOR U33968 ( .A(n17582), .B(n33830), .Z(n33139) );
  XNOR U33969 ( .A(n19141), .B(n19024), .Z(n33830) );
  XNOR U33970 ( .A(n33831), .B(n20807), .Z(n19024) );
  XOR U33971 ( .A(n26568), .B(n27562), .Z(n20807) );
  XOR U33972 ( .A(n33832), .B(n30630), .Z(n27562) );
  ANDN U33973 ( .B(n33126), .A(n29831), .Z(n33832) );
  XOR U33974 ( .A(n33833), .B(n33834), .Z(n29831) );
  XNOR U33975 ( .A(n28479), .B(n26409), .Z(n26568) );
  XNOR U33976 ( .A(n33835), .B(n33836), .Z(n26409) );
  XNOR U33977 ( .A(n24463), .B(n25063), .Z(n33836) );
  XOR U33978 ( .A(n33837), .B(n29836), .Z(n25063) );
  XOR U33979 ( .A(n32359), .B(n33838), .Z(n29836) );
  ANDN U33980 ( .B(n27566), .A(n27564), .Z(n33837) );
  XOR U33981 ( .A(n33839), .B(n29071), .Z(n27564) );
  XOR U33982 ( .A(n33840), .B(n30928), .Z(n27566) );
  XOR U33983 ( .A(n33841), .B(n29828), .Z(n24463) );
  XNOR U33984 ( .A(n33217), .B(n33842), .Z(n29828) );
  XNOR U33985 ( .A(n33843), .B(n33844), .Z(n33217) );
  NOR U33986 ( .A(n33845), .B(n33846), .Z(n33843) );
  NOR U33987 ( .A(n27572), .B(n27571), .Z(n33841) );
  XOR U33988 ( .A(n33820), .B(n33847), .Z(n27571) );
  IV U33989 ( .A(n28811), .Z(n33820) );
  XNOR U33990 ( .A(n31054), .B(n33848), .Z(n27572) );
  XOR U33991 ( .A(n30607), .B(n33849), .Z(n33835) );
  XOR U33992 ( .A(n27357), .B(n22891), .Z(n33849) );
  XOR U33993 ( .A(n33850), .B(n29824), .Z(n22891) );
  XNOR U33994 ( .A(n33853), .B(n33854), .Z(n32386) );
  XOR U33995 ( .A(n33492), .B(n32173), .Z(n33854) );
  XOR U33996 ( .A(n33855), .B(n33856), .Z(n32173) );
  AND U33997 ( .A(n33857), .B(n33858), .Z(n33855) );
  XOR U33998 ( .A(n33859), .B(n33860), .Z(n33492) );
  XNOR U33999 ( .A(n30003), .B(n33863), .Z(n33853) );
  XNOR U34000 ( .A(n30172), .B(n28824), .Z(n33863) );
  XOR U34001 ( .A(n33864), .B(n33865), .Z(n28824) );
  XNOR U34002 ( .A(n33868), .B(n33869), .Z(n30172) );
  ANDN U34003 ( .B(n33870), .A(n33871), .Z(n33868) );
  XOR U34004 ( .A(n33872), .B(n33873), .Z(n30003) );
  ANDN U34005 ( .B(n33874), .A(n33875), .Z(n33872) );
  NOR U34006 ( .A(n28863), .B(n28862), .Z(n33850) );
  XNOR U34007 ( .A(n32160), .B(n33876), .Z(n28862) );
  IV U34008 ( .A(n32268), .Z(n32160) );
  XNOR U34009 ( .A(n33877), .B(n33878), .Z(n32268) );
  XOR U34010 ( .A(n33879), .B(n32829), .Z(n28863) );
  IV U34011 ( .A(n33721), .Z(n32829) );
  XOR U34012 ( .A(n33880), .B(n33881), .Z(n33721) );
  XNOR U34013 ( .A(n33882), .B(n29822), .Z(n27357) );
  XOR U34014 ( .A(n33883), .B(n30687), .Z(n29822) );
  XOR U34015 ( .A(n32755), .B(n33884), .Z(n30687) );
  XNOR U34016 ( .A(n33885), .B(n33886), .Z(n32755) );
  XNOR U34017 ( .A(n33887), .B(n32873), .Z(n33886) );
  XNOR U34018 ( .A(n33888), .B(n33889), .Z(n32873) );
  AND U34019 ( .A(n33890), .B(n33891), .Z(n33888) );
  XNOR U34020 ( .A(n31561), .B(n33892), .Z(n33885) );
  XNOR U34021 ( .A(n30864), .B(n33893), .Z(n33892) );
  XNOR U34022 ( .A(n33894), .B(n33895), .Z(n30864) );
  AND U34023 ( .A(n33896), .B(n33897), .Z(n33894) );
  XOR U34024 ( .A(n33898), .B(n33899), .Z(n31561) );
  ANDN U34025 ( .B(n33900), .A(n33901), .Z(n33898) );
  ANDN U34026 ( .B(n28036), .A(n28035), .Z(n33882) );
  XNOR U34027 ( .A(n33902), .B(n31148), .Z(n28035) );
  XOR U34028 ( .A(n33903), .B(n32531), .Z(n28036) );
  XNOR U34029 ( .A(n33904), .B(n29833), .Z(n30607) );
  XOR U34030 ( .A(n33905), .B(n32511), .Z(n29833) );
  XNOR U34031 ( .A(n33906), .B(n33907), .Z(n32511) );
  NOR U34032 ( .A(n33126), .B(n30630), .Z(n33904) );
  XNOR U34033 ( .A(n33908), .B(n33828), .Z(n30630) );
  XOR U34034 ( .A(n30869), .B(n33909), .Z(n33126) );
  IV U34035 ( .A(n29938), .Z(n30869) );
  XOR U34036 ( .A(n32385), .B(n33910), .Z(n29938) );
  XOR U34037 ( .A(n33911), .B(n33912), .Z(n32385) );
  XNOR U34038 ( .A(n32114), .B(n31367), .Z(n33912) );
  XOR U34039 ( .A(n33913), .B(n33504), .Z(n31367) );
  ANDN U34040 ( .B(n33505), .A(n33914), .Z(n33913) );
  XOR U34041 ( .A(n33915), .B(n32673), .Z(n32114) );
  XNOR U34042 ( .A(n33916), .B(n33917), .Z(n32673) );
  ANDN U34043 ( .B(n33507), .A(n33918), .Z(n33915) );
  XNOR U34044 ( .A(n32558), .B(n33919), .Z(n33911) );
  XNOR U34045 ( .A(n31263), .B(n32968), .Z(n33919) );
  XOR U34046 ( .A(n33920), .B(n32661), .Z(n32968) );
  XNOR U34047 ( .A(n33921), .B(n33922), .Z(n32661) );
  ANDN U34048 ( .B(n33923), .A(n33924), .Z(n33920) );
  XNOR U34049 ( .A(n33925), .B(n33418), .Z(n31263) );
  XOR U34050 ( .A(n33926), .B(n33927), .Z(n33418) );
  ANDN U34051 ( .B(n33928), .A(n33509), .Z(n33925) );
  XOR U34052 ( .A(n33929), .B(n32657), .Z(n32558) );
  XNOR U34053 ( .A(n33930), .B(n33931), .Z(n32657) );
  ANDN U34054 ( .B(n33500), .A(n33932), .Z(n33929) );
  XNOR U34055 ( .A(n33933), .B(n33934), .Z(n28479) );
  XOR U34056 ( .A(n24830), .B(n27050), .Z(n33934) );
  XNOR U34057 ( .A(n33935), .B(n29816), .Z(n27050) );
  XOR U34058 ( .A(n33214), .B(n33842), .Z(n29816) );
  IV U34059 ( .A(n33226), .Z(n33842) );
  XNOR U34060 ( .A(n33936), .B(n33937), .Z(n33214) );
  NOR U34061 ( .A(n30680), .B(n30621), .Z(n33935) );
  XNOR U34062 ( .A(n28790), .B(n33940), .Z(n30621) );
  IV U34063 ( .A(n33941), .Z(n28790) );
  XOR U34064 ( .A(n33942), .B(n33943), .Z(n30680) );
  XNOR U34065 ( .A(n33944), .B(n29813), .Z(n24830) );
  XOR U34066 ( .A(n33945), .B(n30743), .Z(n29813) );
  AND U34067 ( .A(n30623), .B(n30685), .Z(n33944) );
  XOR U34068 ( .A(n33947), .B(n31346), .Z(n30623) );
  XOR U34069 ( .A(n23581), .B(n33948), .Z(n33933) );
  XNOR U34070 ( .A(n24917), .B(n26977), .Z(n33948) );
  XOR U34071 ( .A(n33949), .B(n29802), .Z(n26977) );
  XOR U34072 ( .A(n30493), .B(n33950), .Z(n29802) );
  NOR U34073 ( .A(n30689), .B(n30616), .Z(n33949) );
  XOR U34074 ( .A(n33951), .B(n33952), .Z(n30616) );
  XOR U34075 ( .A(n33953), .B(n31233), .Z(n30689) );
  IV U34076 ( .A(n29262), .Z(n31233) );
  XNOR U34077 ( .A(n33954), .B(n33955), .Z(n29262) );
  XNOR U34078 ( .A(n33956), .B(n29807), .Z(n24917) );
  XNOR U34079 ( .A(n33957), .B(n31579), .Z(n29807) );
  ANDN U34080 ( .B(n30619), .A(n31144), .Z(n33956) );
  XOR U34081 ( .A(n33958), .B(n28821), .Z(n31144) );
  XOR U34082 ( .A(n33959), .B(n30651), .Z(n30619) );
  IV U34083 ( .A(n33359), .Z(n30651) );
  XNOR U34084 ( .A(n33962), .B(n30612), .Z(n23581) );
  XNOR U34085 ( .A(n30231), .B(n33963), .Z(n30612) );
  XOR U34086 ( .A(n33964), .B(n32239), .Z(n30231) );
  XOR U34087 ( .A(n33965), .B(n33966), .Z(n32239) );
  XNOR U34088 ( .A(n33967), .B(n33133), .Z(n33966) );
  XNOR U34089 ( .A(n33968), .B(n33969), .Z(n33133) );
  XOR U34090 ( .A(n27941), .B(n33972), .Z(n33965) );
  XNOR U34091 ( .A(n31581), .B(n29918), .Z(n33972) );
  XNOR U34092 ( .A(n33973), .B(n33974), .Z(n29918) );
  XOR U34093 ( .A(n33977), .B(n33978), .Z(n31581) );
  XNOR U34094 ( .A(n33981), .B(n33982), .Z(n27941) );
  ANDN U34095 ( .B(n33983), .A(n33984), .Z(n33981) );
  ANDN U34096 ( .B(n30693), .A(n31146), .Z(n33962) );
  XOR U34097 ( .A(n32101), .B(n33985), .Z(n31146) );
  XOR U34098 ( .A(n33619), .B(n31100), .Z(n30693) );
  IV U34099 ( .A(n31154), .Z(n31100) );
  XOR U34100 ( .A(n33986), .B(n33987), .Z(n33619) );
  ANDN U34101 ( .B(n23233), .A(n25126), .Z(n33831) );
  XOR U34102 ( .A(n25068), .B(n29385), .Z(n25126) );
  XNOR U34103 ( .A(n33990), .B(n30604), .Z(n29385) );
  NOR U34104 ( .A(n31024), .B(n29975), .Z(n33990) );
  XNOR U34105 ( .A(n31190), .B(n33991), .Z(n29975) );
  XOR U34106 ( .A(n33992), .B(n33993), .Z(n31190) );
  IV U34107 ( .A(n26924), .Z(n25068) );
  XOR U34108 ( .A(n31521), .B(n29656), .Z(n26924) );
  XOR U34109 ( .A(n33994), .B(n33995), .Z(n29656) );
  XOR U34110 ( .A(n27679), .B(n25718), .Z(n33995) );
  XOR U34111 ( .A(n33996), .B(n27322), .Z(n25718) );
  XNOR U34112 ( .A(n33997), .B(n30210), .Z(n27322) );
  IV U34113 ( .A(n30923), .Z(n30210) );
  XOR U34114 ( .A(n33998), .B(n33999), .Z(n30923) );
  ANDN U34115 ( .B(n29379), .A(n29378), .Z(n33996) );
  XOR U34116 ( .A(n34000), .B(n31348), .Z(n29378) );
  XNOR U34117 ( .A(n34001), .B(n34002), .Z(n33493) );
  XOR U34118 ( .A(n31138), .B(n31913), .Z(n34002) );
  XOR U34119 ( .A(n34003), .B(n34004), .Z(n31913) );
  ANDN U34120 ( .B(n33873), .A(n34005), .Z(n34003) );
  XNOR U34121 ( .A(n34006), .B(n34007), .Z(n31138) );
  ANDN U34122 ( .B(n33856), .A(n33858), .Z(n34006) );
  XOR U34123 ( .A(n32650), .B(n34008), .Z(n34001) );
  XNOR U34124 ( .A(n32206), .B(n31800), .Z(n34008) );
  XNOR U34125 ( .A(n34009), .B(n34010), .Z(n31800) );
  ANDN U34126 ( .B(n33869), .A(n33870), .Z(n34009) );
  XOR U34127 ( .A(n34011), .B(n34012), .Z(n32206) );
  ANDN U34128 ( .B(n33860), .A(n33862), .Z(n34011) );
  XOR U34129 ( .A(n34013), .B(n34014), .Z(n32650) );
  ANDN U34130 ( .B(n33865), .A(n33867), .Z(n34013) );
  XOR U34131 ( .A(n34016), .B(n32196), .Z(n29379) );
  XNOR U34132 ( .A(n34017), .B(n27917), .Z(n27679) );
  XOR U34133 ( .A(n32362), .B(n34018), .Z(n27917) );
  NOR U34134 ( .A(n29381), .B(n29382), .Z(n34017) );
  XOR U34135 ( .A(n34019), .B(n29734), .Z(n29382) );
  XNOR U34136 ( .A(n34021), .B(n34022), .Z(n33823) );
  XNOR U34137 ( .A(n34023), .B(n31288), .Z(n34022) );
  XNOR U34138 ( .A(n34024), .B(n34025), .Z(n31288) );
  NOR U34139 ( .A(n34026), .B(n34027), .Z(n34024) );
  XOR U34140 ( .A(n32217), .B(n34028), .Z(n34021) );
  XOR U34141 ( .A(n31686), .B(n33608), .Z(n34028) );
  XNOR U34142 ( .A(n34029), .B(n34030), .Z(n33608) );
  ANDN U34143 ( .B(n34031), .A(n34032), .Z(n34029) );
  XNOR U34144 ( .A(n34033), .B(n34034), .Z(n31686) );
  ANDN U34145 ( .B(n34035), .A(n34036), .Z(n34033) );
  XNOR U34146 ( .A(n34037), .B(n34038), .Z(n32217) );
  NOR U34147 ( .A(n34039), .B(n34040), .Z(n34037) );
  XOR U34148 ( .A(n34041), .B(n30197), .Z(n29381) );
  XOR U34149 ( .A(n34042), .B(n32257), .Z(n30197) );
  XNOR U34150 ( .A(n34043), .B(n34044), .Z(n32257) );
  XNOR U34151 ( .A(n31338), .B(n32614), .Z(n34044) );
  XNOR U34152 ( .A(n34045), .B(n34046), .Z(n32614) );
  ANDN U34153 ( .B(n34047), .A(n34048), .Z(n34045) );
  XNOR U34154 ( .A(n34049), .B(n34050), .Z(n31338) );
  ANDN U34155 ( .B(n34051), .A(n34052), .Z(n34049) );
  XNOR U34156 ( .A(n34053), .B(n34054), .Z(n34043) );
  XNOR U34157 ( .A(n31621), .B(n31638), .Z(n34054) );
  XNOR U34158 ( .A(n34055), .B(n34056), .Z(n31638) );
  ANDN U34159 ( .B(n34057), .A(n34058), .Z(n34055) );
  XNOR U34160 ( .A(n34059), .B(n34060), .Z(n31621) );
  ANDN U34161 ( .B(n34061), .A(n34062), .Z(n34059) );
  XNOR U34162 ( .A(n22520), .B(n34063), .Z(n33994) );
  XNOR U34163 ( .A(n23070), .B(n22984), .Z(n34063) );
  XOR U34164 ( .A(n34064), .B(n27318), .Z(n22984) );
  XNOR U34165 ( .A(n34065), .B(n30217), .Z(n27318) );
  IV U34166 ( .A(n31794), .Z(n30217) );
  XNOR U34167 ( .A(n34066), .B(n33731), .Z(n31794) );
  XNOR U34168 ( .A(n34067), .B(n34068), .Z(n33731) );
  XNOR U34169 ( .A(n29098), .B(n34069), .Z(n34068) );
  XNOR U34170 ( .A(n34070), .B(n34071), .Z(n29098) );
  NOR U34171 ( .A(n34072), .B(n34073), .Z(n34070) );
  XOR U34172 ( .A(n32494), .B(n34074), .Z(n34067) );
  XOR U34173 ( .A(n32375), .B(n31390), .Z(n34074) );
  XNOR U34174 ( .A(n34075), .B(n34076), .Z(n31390) );
  ANDN U34175 ( .B(n34077), .A(n34078), .Z(n34075) );
  XNOR U34176 ( .A(n34079), .B(n34080), .Z(n32375) );
  NOR U34177 ( .A(n34081), .B(n34082), .Z(n34079) );
  XNOR U34178 ( .A(n34083), .B(n34084), .Z(n32494) );
  NOR U34179 ( .A(n34085), .B(n34086), .Z(n34083) );
  XNOR U34180 ( .A(n34087), .B(n32044), .Z(n30599) );
  XNOR U34181 ( .A(n34088), .B(n33490), .Z(n32044) );
  XNOR U34182 ( .A(n34089), .B(n34090), .Z(n33490) );
  XNOR U34183 ( .A(n32293), .B(n29179), .Z(n34090) );
  XNOR U34184 ( .A(n34091), .B(n34092), .Z(n29179) );
  ANDN U34185 ( .B(n34093), .A(n34084), .Z(n34091) );
  XNOR U34186 ( .A(n34094), .B(n34095), .Z(n32293) );
  XOR U34187 ( .A(n33307), .B(n34097), .Z(n34089) );
  XOR U34188 ( .A(n33262), .B(n31239), .Z(n34097) );
  XNOR U34189 ( .A(n34098), .B(n34099), .Z(n31239) );
  ANDN U34190 ( .B(n34100), .A(n34071), .Z(n34098) );
  XNOR U34191 ( .A(n34101), .B(n34102), .Z(n33262) );
  ANDN U34192 ( .B(n34103), .A(n34080), .Z(n34101) );
  IV U34193 ( .A(n34104), .Z(n34080) );
  XNOR U34194 ( .A(n34105), .B(n34106), .Z(n33307) );
  NOR U34195 ( .A(n34107), .B(n34108), .Z(n34105) );
  XOR U34196 ( .A(n34109), .B(n33382), .Z(n30801) );
  XNOR U34197 ( .A(n34110), .B(n29977), .Z(n23070) );
  XOR U34198 ( .A(n34111), .B(n30170), .Z(n29977) );
  IV U34199 ( .A(n29747), .Z(n30170) );
  ANDN U34200 ( .B(n31024), .A(n30604), .Z(n34110) );
  XOR U34201 ( .A(n34114), .B(n30039), .Z(n30604) );
  IV U34202 ( .A(n34115), .Z(n30039) );
  XOR U34203 ( .A(n34116), .B(n31071), .Z(n31024) );
  XNOR U34204 ( .A(n32461), .B(n34117), .Z(n31071) );
  XOR U34205 ( .A(n34118), .B(n34119), .Z(n32461) );
  XNOR U34206 ( .A(n34120), .B(n33302), .Z(n34119) );
  XNOR U34207 ( .A(n34121), .B(n34122), .Z(n33302) );
  ANDN U34208 ( .B(n34123), .A(n34124), .Z(n34121) );
  XNOR U34209 ( .A(n34125), .B(n34126), .Z(n34118) );
  XOR U34210 ( .A(n30164), .B(n34127), .Z(n34126) );
  XNOR U34211 ( .A(n34128), .B(n34129), .Z(n30164) );
  ANDN U34212 ( .B(n34130), .A(n34131), .Z(n34128) );
  XNOR U34213 ( .A(n34132), .B(n27327), .Z(n22520) );
  XOR U34214 ( .A(n34133), .B(n32993), .Z(n27327) );
  XOR U34215 ( .A(n34134), .B(n28744), .Z(n29387) );
  XOR U34216 ( .A(n34135), .B(n34136), .Z(n28744) );
  XOR U34217 ( .A(n34137), .B(n29050), .Z(n29388) );
  XOR U34218 ( .A(n33489), .B(n34138), .Z(n29050) );
  XOR U34219 ( .A(n34139), .B(n34140), .Z(n33489) );
  XNOR U34220 ( .A(n32024), .B(n31273), .Z(n34140) );
  XNOR U34221 ( .A(n34141), .B(n34142), .Z(n31273) );
  NOR U34222 ( .A(n34143), .B(n34144), .Z(n34141) );
  XNOR U34223 ( .A(n34145), .B(n33315), .Z(n32024) );
  ANDN U34224 ( .B(n34146), .A(n33314), .Z(n34145) );
  XOR U34225 ( .A(n32283), .B(n34147), .Z(n34139) );
  XOR U34226 ( .A(n30861), .B(n32929), .Z(n34147) );
  XNOR U34227 ( .A(n34148), .B(n33321), .Z(n32929) );
  XNOR U34228 ( .A(n34150), .B(n33459), .Z(n30861) );
  IV U34229 ( .A(n34151), .Z(n33459) );
  XNOR U34230 ( .A(n34153), .B(n33547), .Z(n32283) );
  ANDN U34231 ( .B(n33548), .A(n34154), .Z(n34153) );
  XOR U34232 ( .A(n34155), .B(n34156), .Z(n31521) );
  XNOR U34233 ( .A(n25783), .B(n25763), .Z(n34156) );
  XOR U34234 ( .A(n34157), .B(n27685), .Z(n25763) );
  XOR U34235 ( .A(n34158), .B(n32139), .Z(n27685) );
  XOR U34236 ( .A(n33613), .B(n31154), .Z(n27684) );
  XOR U34237 ( .A(n34161), .B(n34162), .Z(n33613) );
  ANDN U34238 ( .B(n34163), .A(n34164), .Z(n34161) );
  XNOR U34239 ( .A(n34165), .B(n31369), .Z(n30373) );
  XOR U34240 ( .A(n34166), .B(n34167), .Z(n31369) );
  XNOR U34241 ( .A(n34168), .B(n27698), .Z(n25783) );
  XOR U34242 ( .A(n33433), .B(n32000), .Z(n27698) );
  IV U34243 ( .A(n29075), .Z(n32000) );
  XNOR U34244 ( .A(n34169), .B(n34170), .Z(n29075) );
  XNOR U34245 ( .A(n34171), .B(n34172), .Z(n33433) );
  NOR U34246 ( .A(n34173), .B(n34174), .Z(n34171) );
  ANDN U34247 ( .B(n27699), .A(n30363), .Z(n34168) );
  XOR U34248 ( .A(n30781), .B(n34175), .Z(n30363) );
  XNOR U34249 ( .A(n34176), .B(n34177), .Z(n30781) );
  XOR U34250 ( .A(n33678), .B(n31022), .Z(n27699) );
  IV U34251 ( .A(n30500), .Z(n31022) );
  XNOR U34252 ( .A(n34180), .B(n34181), .Z(n33678) );
  NOR U34253 ( .A(n34182), .B(n34183), .Z(n34180) );
  XOR U34254 ( .A(n25672), .B(n34184), .Z(n34155) );
  XOR U34255 ( .A(n26701), .B(n26574), .Z(n34184) );
  XNOR U34256 ( .A(n34185), .B(n27694), .Z(n26574) );
  XOR U34257 ( .A(n31566), .B(n34186), .Z(n27694) );
  ANDN U34258 ( .B(n27695), .A(n30368), .Z(n34185) );
  XOR U34259 ( .A(n34187), .B(n29922), .Z(n30368) );
  XNOR U34260 ( .A(n34188), .B(n34189), .Z(n33880) );
  XNOR U34261 ( .A(n30251), .B(n32061), .Z(n34189) );
  XOR U34262 ( .A(n34190), .B(n34191), .Z(n32061) );
  ANDN U34263 ( .B(n34192), .A(n34193), .Z(n34190) );
  XOR U34264 ( .A(n34194), .B(n34195), .Z(n30251) );
  XNOR U34265 ( .A(n31029), .B(n34198), .Z(n34188) );
  XOR U34266 ( .A(n32500), .B(n32221), .Z(n34198) );
  XNOR U34267 ( .A(n34199), .B(n34200), .Z(n32221) );
  NOR U34268 ( .A(n34201), .B(n34202), .Z(n34199) );
  XNOR U34269 ( .A(n34203), .B(n34204), .Z(n32500) );
  ANDN U34270 ( .B(n34205), .A(n34206), .Z(n34203) );
  XNOR U34271 ( .A(n34207), .B(n34208), .Z(n31029) );
  NOR U34272 ( .A(n34209), .B(n34210), .Z(n34207) );
  XNOR U34273 ( .A(n30247), .B(n34212), .Z(n27695) );
  XNOR U34274 ( .A(n34215), .B(n28119), .Z(n26701) );
  XNOR U34275 ( .A(n34216), .B(n30539), .Z(n28119) );
  AND U34276 ( .A(n31188), .B(n28127), .Z(n34215) );
  XNOR U34277 ( .A(n34217), .B(n32053), .Z(n28127) );
  XNOR U34278 ( .A(n34218), .B(n31820), .Z(n31188) );
  IV U34279 ( .A(n33531), .Z(n31820) );
  XNOR U34280 ( .A(n34219), .B(n27688), .Z(n25672) );
  XNOR U34281 ( .A(n30120), .B(n34220), .Z(n27688) );
  IV U34282 ( .A(n30200), .Z(n30120) );
  XOR U34283 ( .A(n34221), .B(n34222), .Z(n30200) );
  ANDN U34284 ( .B(n27689), .A(n30377), .Z(n34219) );
  XOR U34285 ( .A(n31020), .B(n34223), .Z(n30377) );
  IV U34286 ( .A(n30493), .Z(n31020) );
  XOR U34287 ( .A(n31240), .B(n34226), .Z(n27689) );
  XOR U34288 ( .A(n33180), .B(n34227), .Z(n31240) );
  XNOR U34289 ( .A(n34228), .B(n34229), .Z(n33180) );
  XNOR U34290 ( .A(n34230), .B(n31563), .Z(n34229) );
  XOR U34291 ( .A(n34231), .B(n34232), .Z(n31563) );
  NOR U34292 ( .A(n34233), .B(n34234), .Z(n34231) );
  XNOR U34293 ( .A(n32666), .B(n34235), .Z(n34228) );
  XOR U34294 ( .A(n32694), .B(n31339), .Z(n34235) );
  XNOR U34295 ( .A(n34236), .B(n34237), .Z(n31339) );
  XOR U34296 ( .A(n34240), .B(n34241), .Z(n32694) );
  XOR U34297 ( .A(n34244), .B(n34245), .Z(n32666) );
  ANDN U34298 ( .B(n34246), .A(n34247), .Z(n34244) );
  XOR U34299 ( .A(n25057), .B(n30162), .Z(n23233) );
  XOR U34300 ( .A(n34248), .B(n29987), .Z(n30162) );
  XNOR U34301 ( .A(n31459), .B(n34249), .Z(n29550) );
  IV U34302 ( .A(n31951), .Z(n31459) );
  XOR U34303 ( .A(n33220), .B(n34250), .Z(n31951) );
  XOR U34304 ( .A(n34251), .B(n34252), .Z(n33220) );
  XOR U34305 ( .A(n32628), .B(n34253), .Z(n34252) );
  XNOR U34306 ( .A(n34254), .B(n33623), .Z(n32628) );
  ANDN U34307 ( .B(n34255), .A(n34256), .Z(n34254) );
  XOR U34308 ( .A(n32854), .B(n34257), .Z(n34251) );
  XNOR U34309 ( .A(n32265), .B(n33035), .Z(n34257) );
  XOR U34310 ( .A(n34258), .B(n33627), .Z(n33035) );
  ANDN U34311 ( .B(n34259), .A(n34260), .Z(n34258) );
  XNOR U34312 ( .A(n34261), .B(n33616), .Z(n32265) );
  ANDN U34313 ( .B(n34262), .A(n34263), .Z(n34261) );
  XNOR U34314 ( .A(n34264), .B(n33989), .Z(n32854) );
  ANDN U34315 ( .B(n34265), .A(n34266), .Z(n34264) );
  XNOR U34316 ( .A(n26576), .B(n26014), .Z(n25057) );
  XNOR U34317 ( .A(n34267), .B(n34268), .Z(n26014) );
  XOR U34318 ( .A(n21224), .B(n24253), .Z(n34268) );
  XOR U34319 ( .A(n34269), .B(n27148), .Z(n24253) );
  XOR U34320 ( .A(n29315), .B(n34270), .Z(n27148) );
  XOR U34321 ( .A(n34271), .B(n31185), .Z(n29404) );
  IV U34322 ( .A(n30223), .Z(n31185) );
  XNOR U34323 ( .A(n34272), .B(n32865), .Z(n30223) );
  XNOR U34324 ( .A(n34273), .B(n34274), .Z(n32865) );
  XOR U34325 ( .A(n31152), .B(n34275), .Z(n34274) );
  XNOR U34326 ( .A(n34276), .B(n34277), .Z(n31152) );
  AND U34327 ( .A(n34278), .B(n34279), .Z(n34276) );
  XOR U34328 ( .A(n30558), .B(n34280), .Z(n34273) );
  XOR U34329 ( .A(n33733), .B(n30930), .Z(n34280) );
  XNOR U34330 ( .A(n34281), .B(n34282), .Z(n30930) );
  ANDN U34331 ( .B(n34283), .A(n34284), .Z(n34281) );
  XNOR U34332 ( .A(n34285), .B(n34286), .Z(n33733) );
  AND U34333 ( .A(n34287), .B(n34288), .Z(n34285) );
  XNOR U34334 ( .A(n34289), .B(n34290), .Z(n30558) );
  ANDN U34335 ( .B(n34291), .A(n34292), .Z(n34289) );
  XOR U34336 ( .A(n34293), .B(n31549), .Z(n28667) );
  XOR U34337 ( .A(n33634), .B(n34294), .Z(n31549) );
  XOR U34338 ( .A(n34295), .B(n34296), .Z(n33634) );
  XOR U34339 ( .A(n31368), .B(n32487), .Z(n34296) );
  XOR U34340 ( .A(n34297), .B(n34298), .Z(n32487) );
  NOR U34341 ( .A(n34299), .B(n34300), .Z(n34297) );
  XNOR U34342 ( .A(n34301), .B(n34302), .Z(n31368) );
  NOR U34343 ( .A(n34303), .B(n34304), .Z(n34301) );
  XOR U34344 ( .A(n28722), .B(n34305), .Z(n34295) );
  XOR U34345 ( .A(n32125), .B(n34165), .Z(n34305) );
  XNOR U34346 ( .A(n34306), .B(n34307), .Z(n34165) );
  ANDN U34347 ( .B(n34308), .A(n34309), .Z(n34306) );
  XNOR U34348 ( .A(n34310), .B(n34311), .Z(n32125) );
  ANDN U34349 ( .B(n34312), .A(n34313), .Z(n34310) );
  XNOR U34350 ( .A(n34314), .B(n34315), .Z(n28722) );
  NOR U34351 ( .A(n34316), .B(n34317), .Z(n34314) );
  XOR U34352 ( .A(n34318), .B(n27157), .Z(n21224) );
  XOR U34353 ( .A(n34319), .B(n33382), .Z(n27157) );
  IV U34354 ( .A(n34320), .Z(n33382) );
  XOR U34355 ( .A(n34321), .B(n31448), .Z(n29399) );
  XNOR U34356 ( .A(n29959), .B(n33164), .Z(n28660) );
  XNOR U34357 ( .A(n34322), .B(n34323), .Z(n33164) );
  NOR U34358 ( .A(n34324), .B(n34325), .Z(n34322) );
  XOR U34359 ( .A(n34117), .B(n34326), .Z(n29959) );
  XOR U34360 ( .A(n34327), .B(n34328), .Z(n34117) );
  XNOR U34361 ( .A(n30279), .B(n32918), .Z(n34328) );
  XNOR U34362 ( .A(n34329), .B(n34330), .Z(n32918) );
  ANDN U34363 ( .B(n34331), .A(n34332), .Z(n34329) );
  XNOR U34364 ( .A(n34333), .B(n34334), .Z(n30279) );
  ANDN U34365 ( .B(n34335), .A(n34336), .Z(n34333) );
  XOR U34366 ( .A(n30224), .B(n34337), .Z(n34327) );
  XOR U34367 ( .A(n29947), .B(n32959), .Z(n34337) );
  XOR U34368 ( .A(n34338), .B(n34339), .Z(n32959) );
  ANDN U34369 ( .B(n34340), .A(n34341), .Z(n34338) );
  XOR U34370 ( .A(n34342), .B(n34343), .Z(n29947) );
  ANDN U34371 ( .B(n34344), .A(n34345), .Z(n34342) );
  XNOR U34372 ( .A(n34346), .B(n34347), .Z(n30224) );
  ANDN U34373 ( .B(n34348), .A(n34349), .Z(n34346) );
  XOR U34374 ( .A(n27727), .B(n34350), .Z(n34267) );
  XNOR U34375 ( .A(n25933), .B(n25719), .Z(n34350) );
  XOR U34376 ( .A(n34351), .B(n27153), .Z(n25719) );
  XOR U34377 ( .A(n30144), .B(n34352), .Z(n27153) );
  ANDN U34378 ( .B(n29394), .A(n29395), .Z(n34351) );
  IV U34379 ( .A(n28664), .Z(n29395) );
  XOR U34380 ( .A(n34353), .B(n30275), .Z(n28664) );
  XNOR U34381 ( .A(n31947), .B(n34354), .Z(n29394) );
  IV U34382 ( .A(n30501), .Z(n31947) );
  XOR U34383 ( .A(n34355), .B(n27160), .Z(n25933) );
  XNOR U34384 ( .A(n34356), .B(n32402), .Z(n27160) );
  ANDN U34385 ( .B(n28658), .A(n29407), .Z(n34355) );
  IV U34386 ( .A(n30011), .Z(n29407) );
  XNOR U34387 ( .A(n34357), .B(n29916), .Z(n30011) );
  XNOR U34388 ( .A(n34358), .B(n34359), .Z(n29916) );
  XNOR U34389 ( .A(n33455), .B(n34360), .Z(n28658) );
  XNOR U34390 ( .A(n34361), .B(n28674), .Z(n27727) );
  XNOR U34391 ( .A(n32034), .B(n34362), .Z(n28674) );
  ANDN U34392 ( .B(n28669), .A(n29411), .Z(n34361) );
  XOR U34393 ( .A(n32665), .B(n30517), .Z(n29411) );
  XNOR U34394 ( .A(n34365), .B(n34366), .Z(n32665) );
  NOR U34395 ( .A(n33504), .B(n33503), .Z(n34365) );
  XOR U34396 ( .A(n34367), .B(n34368), .Z(n33504) );
  XOR U34397 ( .A(n34369), .B(n27929), .Z(n28669) );
  XOR U34398 ( .A(n34370), .B(n34371), .Z(n26576) );
  XNOR U34399 ( .A(n24373), .B(n26876), .Z(n34371) );
  XNOR U34400 ( .A(n34372), .B(n29992), .Z(n26876) );
  IV U34401 ( .A(n29543), .Z(n29992) );
  XOR U34402 ( .A(n30903), .B(n34373), .Z(n29543) );
  XNOR U34403 ( .A(n33878), .B(n34374), .Z(n30903) );
  XOR U34404 ( .A(n34375), .B(n34376), .Z(n33878) );
  XNOR U34405 ( .A(n28436), .B(n34377), .Z(n34376) );
  XNOR U34406 ( .A(n34378), .B(n34379), .Z(n28436) );
  AND U34407 ( .A(n34380), .B(n34381), .Z(n34378) );
  XNOR U34408 ( .A(n30563), .B(n34382), .Z(n34375) );
  XOR U34409 ( .A(n32377), .B(n34383), .Z(n34382) );
  XOR U34410 ( .A(n34384), .B(n34385), .Z(n32377) );
  ANDN U34411 ( .B(n34386), .A(n34387), .Z(n34384) );
  XOR U34412 ( .A(n34388), .B(n34389), .Z(n30563) );
  ANDN U34413 ( .B(n34390), .A(n34391), .Z(n34388) );
  ANDN U34414 ( .B(n29993), .A(n30127), .Z(n34372) );
  XNOR U34415 ( .A(n29047), .B(n34392), .Z(n30127) );
  XOR U34416 ( .A(n34393), .B(n32053), .Z(n29993) );
  XNOR U34417 ( .A(n34394), .B(n29538), .Z(n24373) );
  IV U34418 ( .A(n29996), .Z(n29538) );
  XNOR U34419 ( .A(n30306), .B(n34395), .Z(n29996) );
  NOR U34420 ( .A(n30119), .B(n29995), .Z(n34394) );
  XNOR U34421 ( .A(n29528), .B(n34396), .Z(n29995) );
  XOR U34422 ( .A(n34399), .B(n33009), .Z(n30119) );
  XOR U34423 ( .A(n29980), .B(n34400), .Z(n34370) );
  XOR U34424 ( .A(n24938), .B(n28724), .Z(n34400) );
  XOR U34425 ( .A(n34401), .B(n29547), .Z(n28724) );
  XOR U34426 ( .A(n34402), .B(n28897), .Z(n29547) );
  XNOR U34427 ( .A(n33884), .B(n34403), .Z(n28897) );
  XNOR U34428 ( .A(n34404), .B(n34405), .Z(n33884) );
  XOR U34429 ( .A(n31155), .B(n27938), .Z(n34405) );
  XOR U34430 ( .A(n34406), .B(n34407), .Z(n27938) );
  ANDN U34431 ( .B(n34408), .A(n34389), .Z(n34406) );
  XNOR U34432 ( .A(n34409), .B(n34410), .Z(n31155) );
  NOR U34433 ( .A(n34411), .B(n34412), .Z(n34409) );
  XOR U34434 ( .A(n33136), .B(n34413), .Z(n34404) );
  XOR U34435 ( .A(n33173), .B(n32839), .Z(n34413) );
  XNOR U34436 ( .A(n34414), .B(n34415), .Z(n32839) );
  XNOR U34437 ( .A(n34417), .B(n34418), .Z(n33173) );
  ANDN U34438 ( .B(n34419), .A(n34420), .Z(n34417) );
  XOR U34439 ( .A(n34421), .B(n34422), .Z(n33136) );
  NOR U34440 ( .A(n34423), .B(n34379), .Z(n34421) );
  ANDN U34441 ( .B(n29984), .A(n30123), .Z(n34401) );
  XOR U34442 ( .A(n34424), .B(n31322), .Z(n30123) );
  XNOR U34443 ( .A(n30644), .B(n34425), .Z(n29984) );
  XNOR U34444 ( .A(n34426), .B(n29556), .Z(n24938) );
  XOR U34445 ( .A(n34427), .B(n27929), .Z(n29556) );
  IV U34446 ( .A(n28875), .Z(n27929) );
  XNOR U34447 ( .A(n34428), .B(n34429), .Z(n28875) );
  ANDN U34448 ( .B(n29990), .A(n30110), .Z(n34426) );
  IV U34449 ( .A(n30168), .Z(n30110) );
  XOR U34450 ( .A(n28739), .B(n34430), .Z(n30168) );
  XNOR U34451 ( .A(n34431), .B(n34432), .Z(n28739) );
  XOR U34452 ( .A(n33590), .B(n31116), .Z(n29990) );
  XNOR U34453 ( .A(n34433), .B(n34434), .Z(n33590) );
  ANDN U34454 ( .B(n34435), .A(n34436), .Z(n34433) );
  XNOR U34455 ( .A(n34437), .B(n29552), .Z(n29980) );
  IV U34456 ( .A(n29986), .Z(n29552) );
  XNOR U34457 ( .A(n34438), .B(n31127), .Z(n29986) );
  ANDN U34458 ( .B(n29987), .A(n30114), .Z(n34437) );
  XOR U34459 ( .A(n31618), .B(n34439), .Z(n30114) );
  XNOR U34460 ( .A(n34440), .B(n31880), .Z(n29987) );
  XNOR U34461 ( .A(n34441), .B(n20811), .Z(n19141) );
  XOR U34462 ( .A(n21603), .B(n29700), .Z(n20811) );
  XNOR U34463 ( .A(n34442), .B(n29691), .Z(n29700) );
  ANDN U34464 ( .B(n32635), .A(n29687), .Z(n34442) );
  XOR U34465 ( .A(n30946), .B(n34443), .Z(n29687) );
  XOR U34466 ( .A(n33772), .B(n34159), .Z(n30946) );
  XNOR U34467 ( .A(n34444), .B(n34445), .Z(n34159) );
  XNOR U34468 ( .A(n31811), .B(n34446), .Z(n34445) );
  XNOR U34469 ( .A(n34447), .B(n34448), .Z(n31811) );
  NOR U34470 ( .A(n34449), .B(n34450), .Z(n34447) );
  XOR U34471 ( .A(n33204), .B(n34451), .Z(n34444) );
  XOR U34472 ( .A(n33697), .B(n33268), .Z(n34451) );
  XNOR U34473 ( .A(n34452), .B(n34453), .Z(n33268) );
  NOR U34474 ( .A(n34454), .B(n34455), .Z(n34452) );
  XNOR U34475 ( .A(n34456), .B(n34457), .Z(n33697) );
  NOR U34476 ( .A(n34458), .B(n34459), .Z(n34456) );
  XNOR U34477 ( .A(n34460), .B(n34461), .Z(n33204) );
  ANDN U34478 ( .B(n34462), .A(n34463), .Z(n34460) );
  XNOR U34479 ( .A(n34464), .B(n34465), .Z(n33772) );
  XNOR U34480 ( .A(n33470), .B(n30537), .Z(n34465) );
  XNOR U34481 ( .A(n34466), .B(n34467), .Z(n30537) );
  XNOR U34482 ( .A(n34470), .B(n34471), .Z(n33470) );
  ANDN U34483 ( .B(n34472), .A(n34473), .Z(n34470) );
  XNOR U34484 ( .A(n34474), .B(n34475), .Z(n34464) );
  XOR U34485 ( .A(n32141), .B(n34476), .Z(n34475) );
  XOR U34486 ( .A(n34477), .B(n34478), .Z(n32141) );
  NOR U34487 ( .A(n34479), .B(n34480), .Z(n34477) );
  XOR U34488 ( .A(n25887), .B(n26694), .Z(n21603) );
  XNOR U34489 ( .A(n34481), .B(n34482), .Z(n26694) );
  XOR U34490 ( .A(n23565), .B(n24774), .Z(n34482) );
  XNOR U34491 ( .A(n34483), .B(n29689), .Z(n24774) );
  XOR U34492 ( .A(n34484), .B(n31858), .Z(n29689) );
  IV U34493 ( .A(n32248), .Z(n31858) );
  XNOR U34494 ( .A(n34485), .B(n33709), .Z(n32248) );
  XOR U34495 ( .A(n34486), .B(n34487), .Z(n33709) );
  XOR U34496 ( .A(n30216), .B(n31402), .Z(n34487) );
  XNOR U34497 ( .A(n34488), .B(n34489), .Z(n31402) );
  ANDN U34498 ( .B(n34490), .A(n34106), .Z(n34488) );
  XOR U34499 ( .A(n34491), .B(n34078), .Z(n30216) );
  NOR U34500 ( .A(n34077), .B(n34095), .Z(n34491) );
  IV U34501 ( .A(n34492), .Z(n34077) );
  XNOR U34502 ( .A(n34065), .B(n34493), .Z(n34486) );
  XNOR U34503 ( .A(n31793), .B(n32252), .Z(n34493) );
  XOR U34504 ( .A(n34494), .B(n34495), .Z(n32252) );
  ANDN U34505 ( .B(n34073), .A(n34099), .Z(n34494) );
  XNOR U34506 ( .A(n34496), .B(n34497), .Z(n31793) );
  ANDN U34507 ( .B(n34086), .A(n34092), .Z(n34496) );
  XNOR U34508 ( .A(n34498), .B(n34082), .Z(n34065) );
  ANDN U34509 ( .B(n34081), .A(n34102), .Z(n34498) );
  ANDN U34510 ( .B(n29691), .A(n32635), .Z(n34483) );
  XNOR U34511 ( .A(n34499), .B(n28821), .Z(n32635) );
  XNOR U34512 ( .A(n29965), .B(n34500), .Z(n29691) );
  XOR U34513 ( .A(n34501), .B(n28317), .Z(n23565) );
  XOR U34514 ( .A(n34502), .B(n32956), .Z(n28317) );
  IV U34515 ( .A(n31148), .Z(n32956) );
  XNOR U34516 ( .A(n34504), .B(n34505), .Z(n32618) );
  XOR U34517 ( .A(n34506), .B(n31577), .Z(n34505) );
  XOR U34518 ( .A(n34507), .B(n34508), .Z(n31577) );
  ANDN U34519 ( .B(n34509), .A(n34510), .Z(n34507) );
  XOR U34520 ( .A(n30767), .B(n34511), .Z(n34504) );
  XOR U34521 ( .A(n32198), .B(n31559), .Z(n34511) );
  XNOR U34522 ( .A(n34512), .B(n34513), .Z(n31559) );
  ANDN U34523 ( .B(n34514), .A(n34515), .Z(n34512) );
  XOR U34524 ( .A(n34516), .B(n34517), .Z(n32198) );
  ANDN U34525 ( .B(n34518), .A(n34519), .Z(n34516) );
  XNOR U34526 ( .A(n34520), .B(n34521), .Z(n30767) );
  ANDN U34527 ( .B(n34522), .A(n34523), .Z(n34520) );
  ANDN U34528 ( .B(n28318), .A(n29704), .Z(n34501) );
  XOR U34529 ( .A(n34524), .B(n31636), .Z(n29704) );
  IV U34530 ( .A(n29329), .Z(n31636) );
  XOR U34531 ( .A(n34525), .B(n34526), .Z(n29329) );
  XNOR U34532 ( .A(n34527), .B(n32011), .Z(n28318) );
  IV U34533 ( .A(n31680), .Z(n32011) );
  XOR U34534 ( .A(n34528), .B(n34529), .Z(n31680) );
  XOR U34535 ( .A(n28301), .B(n34530), .Z(n34481) );
  XOR U34536 ( .A(n24312), .B(n26127), .Z(n34530) );
  XNOR U34537 ( .A(n34531), .B(n28311), .Z(n26127) );
  XNOR U34538 ( .A(n32203), .B(n34532), .Z(n28311) );
  XOR U34539 ( .A(n28811), .B(n34533), .Z(n28312) );
  XOR U34540 ( .A(n34534), .B(n34535), .Z(n29702) );
  XOR U34541 ( .A(n34536), .B(n28308), .Z(n24312) );
  XNOR U34542 ( .A(n34537), .B(n32053), .Z(n28308) );
  XNOR U34543 ( .A(n34538), .B(n34539), .Z(n33604) );
  XNOR U34544 ( .A(n28766), .B(n31244), .Z(n34539) );
  XNOR U34545 ( .A(n34540), .B(n34124), .Z(n31244) );
  NOR U34546 ( .A(n34541), .B(n34542), .Z(n34540) );
  XNOR U34547 ( .A(n34543), .B(n34544), .Z(n28766) );
  ANDN U34548 ( .B(n34545), .A(n34546), .Z(n34543) );
  XOR U34549 ( .A(n30735), .B(n34547), .Z(n34538) );
  XOR U34550 ( .A(n32711), .B(n32675), .Z(n34547) );
  XNOR U34551 ( .A(n34548), .B(n34131), .Z(n32675) );
  NOR U34552 ( .A(n34549), .B(n34550), .Z(n34548) );
  XNOR U34553 ( .A(n34551), .B(n34552), .Z(n32711) );
  NOR U34554 ( .A(n34553), .B(n34554), .Z(n34551) );
  XNOR U34555 ( .A(n34555), .B(n34556), .Z(n30735) );
  NOR U34556 ( .A(n34557), .B(n34558), .Z(n34555) );
  XOR U34557 ( .A(n34559), .B(n34560), .Z(n32373) );
  XNOR U34558 ( .A(n34561), .B(n29750), .Z(n34560) );
  XNOR U34559 ( .A(n34562), .B(n34345), .Z(n29750) );
  XOR U34560 ( .A(n32407), .B(n34565), .Z(n34559) );
  XOR U34561 ( .A(n29518), .B(n31168), .Z(n34565) );
  XNOR U34562 ( .A(n34566), .B(n34341), .Z(n31168) );
  NOR U34563 ( .A(n34567), .B(n34568), .Z(n34566) );
  XNOR U34564 ( .A(n34569), .B(n34349), .Z(n29518) );
  NOR U34565 ( .A(n34570), .B(n34571), .Z(n34569) );
  XNOR U34566 ( .A(n34572), .B(n34336), .Z(n32407) );
  ANDN U34567 ( .B(n34573), .A(n34574), .Z(n34572) );
  XOR U34568 ( .A(n32470), .B(n28890), .Z(n28307) );
  XNOR U34569 ( .A(n33907), .B(n34575), .Z(n28890) );
  XOR U34570 ( .A(n34576), .B(n34577), .Z(n33907) );
  XNOR U34571 ( .A(n30777), .B(n30574), .Z(n34577) );
  XNOR U34572 ( .A(n34578), .B(n34579), .Z(n30574) );
  ANDN U34573 ( .B(n34580), .A(n34581), .Z(n34578) );
  XNOR U34574 ( .A(n34582), .B(n34583), .Z(n30777) );
  AND U34575 ( .A(n34584), .B(n34585), .Z(n34582) );
  XNOR U34576 ( .A(n31063), .B(n34586), .Z(n34576) );
  XNOR U34577 ( .A(n32378), .B(n31842), .Z(n34586) );
  ANDN U34578 ( .B(n34589), .A(n34590), .Z(n34587) );
  ANDN U34579 ( .B(n34593), .A(n34594), .Z(n34591) );
  XOR U34580 ( .A(n34595), .B(n34596), .Z(n31063) );
  AND U34581 ( .A(n34597), .B(n34598), .Z(n34595) );
  XNOR U34582 ( .A(n34599), .B(n34600), .Z(n32470) );
  NOR U34583 ( .A(n34601), .B(n34602), .Z(n34599) );
  XOR U34584 ( .A(n34603), .B(n34604), .Z(n32642) );
  XOR U34585 ( .A(n34605), .B(n28322), .Z(n28301) );
  XOR U34586 ( .A(n34606), .B(n32804), .Z(n28322) );
  ANDN U34587 ( .B(n29698), .A(n28321), .Z(n34605) );
  XOR U34588 ( .A(n34607), .B(n33031), .Z(n28321) );
  XOR U34589 ( .A(n32926), .B(n34608), .Z(n29698) );
  IV U34590 ( .A(n31738), .Z(n32926) );
  XOR U34591 ( .A(n34609), .B(n34610), .Z(n25887) );
  XOR U34592 ( .A(n25184), .B(n32127), .Z(n34610) );
  XNOR U34593 ( .A(n34611), .B(n29670), .Z(n32127) );
  XOR U34594 ( .A(n30149), .B(n34612), .Z(n29670) );
  XNOR U34595 ( .A(n33964), .B(n33308), .Z(n30149) );
  XNOR U34596 ( .A(n34613), .B(n34614), .Z(n33308) );
  XNOR U34597 ( .A(n32601), .B(n30789), .Z(n34614) );
  XOR U34598 ( .A(n34615), .B(n34081), .Z(n30789) );
  XOR U34599 ( .A(n34616), .B(n34617), .Z(n34081) );
  ANDN U34600 ( .B(n34102), .A(n34103), .Z(n34615) );
  XOR U34601 ( .A(n34618), .B(n34619), .Z(n34102) );
  XOR U34602 ( .A(n34620), .B(n34490), .Z(n32601) );
  ANDN U34603 ( .B(n34106), .A(n34621), .Z(n34620) );
  XOR U34604 ( .A(n34622), .B(n34623), .Z(n34106) );
  XNOR U34605 ( .A(n31208), .B(n34624), .Z(n34613) );
  XOR U34606 ( .A(n32843), .B(n33708), .Z(n34624) );
  XNOR U34607 ( .A(n34625), .B(n34086), .Z(n33708) );
  XOR U34608 ( .A(n34626), .B(n34627), .Z(n34086) );
  ANDN U34609 ( .B(n34092), .A(n34093), .Z(n34625) );
  XOR U34610 ( .A(n34628), .B(n34629), .Z(n34092) );
  XNOR U34611 ( .A(n34630), .B(n34073), .Z(n32843) );
  XOR U34612 ( .A(n34631), .B(n34632), .Z(n34073) );
  ANDN U34613 ( .B(n34099), .A(n34100), .Z(n34630) );
  XNOR U34614 ( .A(n34633), .B(n34634), .Z(n34099) );
  XOR U34615 ( .A(n34635), .B(n34492), .Z(n31208) );
  XOR U34616 ( .A(n34636), .B(n34637), .Z(n34492) );
  ANDN U34617 ( .B(n34095), .A(n34096), .Z(n34635) );
  XNOR U34618 ( .A(n34638), .B(n34639), .Z(n34095) );
  XOR U34619 ( .A(n34640), .B(n34641), .Z(n33964) );
  XNOR U34620 ( .A(n34484), .B(n32399), .Z(n34641) );
  XOR U34621 ( .A(n34642), .B(n34643), .Z(n32399) );
  ANDN U34622 ( .B(n34644), .A(n34645), .Z(n34642) );
  XOR U34623 ( .A(n34646), .B(n34647), .Z(n34484) );
  ANDN U34624 ( .B(n34648), .A(n34649), .Z(n34646) );
  XOR U34625 ( .A(n32247), .B(n34650), .Z(n34640) );
  XOR U34626 ( .A(n31857), .B(n33635), .Z(n34650) );
  XNOR U34627 ( .A(n34651), .B(n34652), .Z(n33635) );
  XNOR U34628 ( .A(n34655), .B(n34656), .Z(n31857) );
  ANDN U34629 ( .B(n34657), .A(n34658), .Z(n34655) );
  XNOR U34630 ( .A(n34659), .B(n34660), .Z(n32247) );
  ANDN U34631 ( .B(n29600), .A(n29598), .Z(n34611) );
  XOR U34632 ( .A(n31411), .B(n34663), .Z(n29598) );
  XNOR U34633 ( .A(n34664), .B(n31738), .Z(n29600) );
  XOR U34634 ( .A(n34665), .B(n34666), .Z(n31738) );
  XNOR U34635 ( .A(n34667), .B(n32150), .Z(n25184) );
  IV U34636 ( .A(n31379), .Z(n32150) );
  XNOR U34637 ( .A(n32274), .B(n34668), .Z(n31379) );
  XNOR U34638 ( .A(n34669), .B(n33961), .Z(n32274) );
  XNOR U34639 ( .A(n34670), .B(n34671), .Z(n33961) );
  XOR U34640 ( .A(n34672), .B(n30259), .Z(n34671) );
  XNOR U34641 ( .A(n34673), .B(n34674), .Z(n30259) );
  NOR U34642 ( .A(n34675), .B(n34676), .Z(n34673) );
  XNOR U34643 ( .A(n34677), .B(n34678), .Z(n34670) );
  XNOR U34644 ( .A(n30302), .B(n31970), .Z(n34678) );
  XNOR U34645 ( .A(n34679), .B(n34680), .Z(n31970) );
  ANDN U34646 ( .B(n34681), .A(n34682), .Z(n34679) );
  XOR U34647 ( .A(n34683), .B(n34684), .Z(n30302) );
  NOR U34648 ( .A(n34685), .B(n34686), .Z(n34683) );
  ANDN U34649 ( .B(n29611), .A(n29613), .Z(n34667) );
  XOR U34650 ( .A(n34687), .B(n30116), .Z(n29613) );
  IV U34651 ( .A(n34688), .Z(n30116) );
  XOR U34652 ( .A(n34689), .B(n31448), .Z(n29611) );
  XNOR U34653 ( .A(n34690), .B(n33610), .Z(n31448) );
  XNOR U34654 ( .A(n34691), .B(n34692), .Z(n33610) );
  XNOR U34655 ( .A(n32590), .B(n34443), .Z(n34692) );
  XNOR U34656 ( .A(n34693), .B(n34463), .Z(n34443) );
  NOR U34657 ( .A(n34694), .B(n34462), .Z(n34693) );
  XNOR U34658 ( .A(n34695), .B(n34455), .Z(n32590) );
  ANDN U34659 ( .B(n34454), .A(n34696), .Z(n34695) );
  XNOR U34660 ( .A(n33001), .B(n34697), .Z(n34691) );
  XOR U34661 ( .A(n32964), .B(n30947), .Z(n34697) );
  XNOR U34662 ( .A(n34698), .B(n34699), .Z(n30947) );
  ANDN U34663 ( .B(n34700), .A(n34701), .Z(n34698) );
  XNOR U34664 ( .A(n34702), .B(n34450), .Z(n32964) );
  ANDN U34665 ( .B(n34449), .A(n34703), .Z(n34702) );
  XNOR U34666 ( .A(n34704), .B(n34459), .Z(n33001) );
  NOR U34667 ( .A(n34705), .B(n34706), .Z(n34704) );
  XOR U34668 ( .A(n30803), .B(n34707), .Z(n34609) );
  XNOR U34669 ( .A(n24454), .B(n26919), .Z(n34707) );
  XOR U34670 ( .A(n34708), .B(n29674), .Z(n26919) );
  XOR U34671 ( .A(n34709), .B(n33009), .Z(n29674) );
  IV U34672 ( .A(n29171), .Z(n33009) );
  XOR U34673 ( .A(n34272), .B(n34015), .Z(n29171) );
  XNOR U34674 ( .A(n34710), .B(n34711), .Z(n34015) );
  XNOR U34675 ( .A(n32580), .B(n30289), .Z(n34711) );
  XOR U34676 ( .A(n34712), .B(n34713), .Z(n30289) );
  AND U34677 ( .A(n34714), .B(n34715), .Z(n34712) );
  XOR U34678 ( .A(n34716), .B(n34717), .Z(n32580) );
  AND U34679 ( .A(n34718), .B(n34719), .Z(n34716) );
  XNOR U34680 ( .A(n32805), .B(n34720), .Z(n34710) );
  XOR U34681 ( .A(n28894), .B(n34721), .Z(n34720) );
  XNOR U34682 ( .A(n34722), .B(n34723), .Z(n28894) );
  ANDN U34683 ( .B(n34724), .A(n34725), .Z(n34722) );
  XOR U34684 ( .A(n34726), .B(n34727), .Z(n32805) );
  ANDN U34685 ( .B(n34728), .A(n34729), .Z(n34726) );
  XOR U34686 ( .A(n34730), .B(n34731), .Z(n34272) );
  XNOR U34687 ( .A(n33816), .B(n30238), .Z(n34731) );
  XOR U34688 ( .A(n34732), .B(n34733), .Z(n30238) );
  ANDN U34689 ( .B(n34734), .A(n34735), .Z(n34732) );
  XOR U34690 ( .A(n34736), .B(n34737), .Z(n33816) );
  ANDN U34691 ( .B(n34738), .A(n34739), .Z(n34736) );
  XOR U34692 ( .A(n34740), .B(n34741), .Z(n34730) );
  XOR U34693 ( .A(n34742), .B(n32224), .Z(n34741) );
  XNOR U34694 ( .A(n34743), .B(n34744), .Z(n32224) );
  NOR U34695 ( .A(n34745), .B(n34746), .Z(n34743) );
  XOR U34696 ( .A(n34747), .B(n32975), .Z(n29615) );
  XOR U34697 ( .A(n34748), .B(n33718), .Z(n32975) );
  XOR U34698 ( .A(n34749), .B(n34750), .Z(n33718) );
  XNOR U34699 ( .A(n32233), .B(n33444), .Z(n34750) );
  XOR U34700 ( .A(n34751), .B(n34752), .Z(n33444) );
  XOR U34701 ( .A(n34755), .B(n34756), .Z(n32233) );
  NOR U34702 ( .A(n34757), .B(n34758), .Z(n34755) );
  XNOR U34703 ( .A(n34759), .B(n34760), .Z(n34749) );
  XOR U34704 ( .A(n32709), .B(n32572), .Z(n34760) );
  XOR U34705 ( .A(n34761), .B(n34762), .Z(n32572) );
  ANDN U34706 ( .B(n34763), .A(n34764), .Z(n34761) );
  XNOR U34707 ( .A(n34765), .B(n34766), .Z(n32709) );
  ANDN U34708 ( .B(n34767), .A(n34768), .Z(n34765) );
  XOR U34709 ( .A(n33941), .B(n34769), .Z(n29617) );
  XNOR U34710 ( .A(n34770), .B(n34294), .Z(n33941) );
  XNOR U34711 ( .A(n34771), .B(n34772), .Z(n34294) );
  XNOR U34712 ( .A(n34392), .B(n34773), .Z(n34772) );
  XNOR U34713 ( .A(n34774), .B(n34775), .Z(n34392) );
  XOR U34714 ( .A(n33098), .B(n34777), .Z(n34771) );
  XOR U34715 ( .A(n32706), .B(n29048), .Z(n34777) );
  XNOR U34716 ( .A(n34778), .B(n34779), .Z(n29048) );
  ANDN U34717 ( .B(n34181), .A(n34780), .Z(n34778) );
  XNOR U34718 ( .A(n34781), .B(n34782), .Z(n32706) );
  NOR U34719 ( .A(n33685), .B(n34783), .Z(n34781) );
  XOR U34720 ( .A(n34784), .B(n34785), .Z(n33098) );
  ANDN U34721 ( .B(n33689), .A(n34786), .Z(n34784) );
  XNOR U34722 ( .A(n34787), .B(n29662), .Z(n24454) );
  XOR U34723 ( .A(n32595), .B(n34788), .Z(n29662) );
  XOR U34724 ( .A(n34789), .B(n34790), .Z(n32595) );
  XOR U34725 ( .A(n34791), .B(n29965), .Z(n29609) );
  XNOR U34726 ( .A(n34792), .B(n34793), .Z(n29965) );
  XOR U34727 ( .A(n34794), .B(n32196), .Z(n29607) );
  XOR U34728 ( .A(n34795), .B(n34796), .Z(n32196) );
  XNOR U34729 ( .A(n34797), .B(n29665), .Z(n30803) );
  XNOR U34730 ( .A(n30306), .B(n34798), .Z(n29665) );
  XNOR U34731 ( .A(n34799), .B(n33364), .Z(n30306) );
  XNOR U34732 ( .A(n34800), .B(n34801), .Z(n33364) );
  XNOR U34733 ( .A(n31353), .B(n32533), .Z(n34801) );
  XOR U34734 ( .A(n34802), .B(n33350), .Z(n32533) );
  ANDN U34735 ( .B(n34803), .A(n34804), .Z(n34802) );
  XOR U34736 ( .A(n34805), .B(n33354), .Z(n31353) );
  ANDN U34737 ( .B(n33353), .A(n34806), .Z(n34805) );
  XOR U34738 ( .A(n30772), .B(n34807), .Z(n34800) );
  XOR U34739 ( .A(n32023), .B(n30077), .Z(n34807) );
  XNOR U34740 ( .A(n34808), .B(n33336), .Z(n30077) );
  ANDN U34741 ( .B(n33337), .A(n34809), .Z(n34808) );
  XNOR U34742 ( .A(n34810), .B(n33341), .Z(n32023) );
  NOR U34743 ( .A(n33340), .B(n34811), .Z(n34810) );
  XOR U34744 ( .A(n34812), .B(n33346), .Z(n30772) );
  ANDN U34745 ( .B(n34813), .A(n33345), .Z(n34812) );
  NOR U34746 ( .A(n29602), .B(n29603), .Z(n34797) );
  XNOR U34747 ( .A(n34814), .B(n34815), .Z(n29603) );
  XOR U34748 ( .A(n34816), .B(n30544), .Z(n29602) );
  IV U34749 ( .A(n34604), .Z(n30544) );
  XNOR U34750 ( .A(n34817), .B(n34818), .Z(n33955) );
  XOR U34751 ( .A(n32043), .B(n32226), .Z(n34818) );
  XNOR U34752 ( .A(n34819), .B(n34654), .Z(n32226) );
  AND U34753 ( .A(n34820), .B(n34821), .Z(n34819) );
  XNOR U34754 ( .A(n34822), .B(n34661), .Z(n32043) );
  AND U34755 ( .A(n34823), .B(n34824), .Z(n34822) );
  XOR U34756 ( .A(n34087), .B(n34825), .Z(n34817) );
  XNOR U34757 ( .A(n32847), .B(n33817), .Z(n34825) );
  XNOR U34758 ( .A(n34826), .B(n34658), .Z(n33817) );
  AND U34759 ( .A(n34827), .B(n34828), .Z(n34826) );
  XOR U34760 ( .A(n34829), .B(n34645), .Z(n32847) );
  IV U34761 ( .A(n34830), .Z(n34645) );
  ANDN U34762 ( .B(n34831), .A(n34832), .Z(n34829) );
  XOR U34763 ( .A(n34833), .B(n34648), .Z(n34087) );
  ANDN U34764 ( .B(n34834), .A(n34835), .Z(n34833) );
  XOR U34765 ( .A(n34836), .B(n34837), .Z(n33910) );
  XNOR U34766 ( .A(n34158), .B(n34838), .Z(n34837) );
  XNOR U34767 ( .A(n34839), .B(n33970), .Z(n34158) );
  ANDN U34768 ( .B(n34840), .A(n34841), .Z(n34839) );
  XNOR U34769 ( .A(n32693), .B(n34842), .Z(n34836) );
  XOR U34770 ( .A(n32138), .B(n33202), .Z(n34842) );
  XNOR U34771 ( .A(n34843), .B(n33984), .Z(n33202) );
  NOR U34772 ( .A(n34844), .B(n34845), .Z(n34843) );
  XNOR U34773 ( .A(n33976), .B(n34846), .Z(n32138) );
  XOR U34774 ( .A(n4620), .B(n34847), .Z(n34846) );
  NANDN U34775 ( .A(n34848), .B(n34849), .Z(n34847) );
  ANDN U34776 ( .B(n31711), .A(rc_i[0]), .Z(n4620) );
  XNOR U34777 ( .A(n34850), .B(n33979), .Z(n32693) );
  ANDN U34778 ( .B(n34851), .A(n34852), .Z(n34850) );
  ANDN U34779 ( .B(n25921), .A(n25920), .Z(n34441) );
  XNOR U34780 ( .A(n28241), .B(n22820), .Z(n25920) );
  XNOR U34781 ( .A(n34853), .B(n34854), .Z(n29156) );
  XOR U34782 ( .A(n25161), .B(n26044), .Z(n34854) );
  XOR U34783 ( .A(n34855), .B(n26808), .Z(n26044) );
  XNOR U34784 ( .A(n30144), .B(n34856), .Z(n26808) );
  IV U34785 ( .A(n31411), .Z(n30144) );
  XNOR U34786 ( .A(n34857), .B(n33072), .Z(n31411) );
  XOR U34787 ( .A(n34858), .B(n34859), .Z(n33072) );
  XOR U34788 ( .A(n34396), .B(n33529), .Z(n34859) );
  XNOR U34789 ( .A(n34860), .B(n34861), .Z(n33529) );
  ANDN U34790 ( .B(n34862), .A(n34863), .Z(n34860) );
  XOR U34791 ( .A(n34864), .B(n34865), .Z(n34396) );
  ANDN U34792 ( .B(n34866), .A(n34727), .Z(n34864) );
  IV U34793 ( .A(n34867), .Z(n34727) );
  XOR U34794 ( .A(n30788), .B(n34868), .Z(n34858) );
  XNOR U34795 ( .A(n31838), .B(n29529), .Z(n34868) );
  XNOR U34796 ( .A(n34869), .B(n34870), .Z(n29529) );
  ANDN U34797 ( .B(n34713), .A(n34871), .Z(n34869) );
  XNOR U34798 ( .A(n34872), .B(n34873), .Z(n31838) );
  ANDN U34799 ( .B(n34717), .A(n34874), .Z(n34872) );
  XNOR U34800 ( .A(n34875), .B(n34876), .Z(n30788) );
  ANDN U34801 ( .B(n34877), .A(n34878), .Z(n34875) );
  ANDN U34802 ( .B(n26809), .A(n28151), .Z(n34855) );
  XOR U34803 ( .A(n32250), .B(n34879), .Z(n28151) );
  IV U34804 ( .A(n31844), .Z(n32250) );
  XNOR U34805 ( .A(n34880), .B(n33298), .Z(n31844) );
  XNOR U34806 ( .A(n34881), .B(n34882), .Z(n33298) );
  XOR U34807 ( .A(n28472), .B(n33485), .Z(n34882) );
  XOR U34808 ( .A(n34883), .B(n34884), .Z(n33485) );
  ANDN U34809 ( .B(n34885), .A(n34886), .Z(n34883) );
  XNOR U34810 ( .A(n34887), .B(n34888), .Z(n28472) );
  ANDN U34811 ( .B(n34889), .A(n33665), .Z(n34887) );
  XOR U34812 ( .A(n30007), .B(n34890), .Z(n34881) );
  XNOR U34813 ( .A(n30124), .B(n31175), .Z(n34890) );
  XNOR U34814 ( .A(n34891), .B(n34892), .Z(n31175) );
  NOR U34815 ( .A(n34893), .B(n33655), .Z(n34891) );
  XNOR U34816 ( .A(n34894), .B(n34895), .Z(n30124) );
  ANDN U34817 ( .B(n34896), .A(n33661), .Z(n34894) );
  XNOR U34818 ( .A(n34897), .B(n34898), .Z(n30007) );
  ANDN U34819 ( .B(n34899), .A(n33651), .Z(n34897) );
  XNOR U34820 ( .A(n34125), .B(n33303), .Z(n26809) );
  XNOR U34821 ( .A(n34900), .B(n34901), .Z(n34125) );
  ANDN U34822 ( .B(n34902), .A(n34552), .Z(n34900) );
  XNOR U34823 ( .A(n34903), .B(n32408), .Z(n25161) );
  XNOR U34824 ( .A(n34904), .B(n33531), .Z(n32408) );
  XOR U34825 ( .A(n32679), .B(n33221), .Z(n33531) );
  XNOR U34826 ( .A(n34905), .B(n34906), .Z(n33221) );
  XNOR U34827 ( .A(n34223), .B(n33950), .Z(n34906) );
  XOR U34828 ( .A(n34907), .B(n34908), .Z(n33950) );
  ANDN U34829 ( .B(n34909), .A(n34910), .Z(n34907) );
  XNOR U34830 ( .A(n34911), .B(n34912), .Z(n34223) );
  ANDN U34831 ( .B(n34913), .A(n34914), .Z(n34911) );
  XOR U34832 ( .A(n33127), .B(n34915), .Z(n34905) );
  XOR U34833 ( .A(n31019), .B(n30494), .Z(n34915) );
  XNOR U34834 ( .A(n34916), .B(n34917), .Z(n30494) );
  NOR U34835 ( .A(n34918), .B(n34919), .Z(n34916) );
  XNOR U34836 ( .A(n34920), .B(n34921), .Z(n31019) );
  NOR U34837 ( .A(n34922), .B(n34923), .Z(n34920) );
  XNOR U34838 ( .A(n34924), .B(n34925), .Z(n33127) );
  NOR U34839 ( .A(n34926), .B(n34927), .Z(n34924) );
  XOR U34840 ( .A(n34928), .B(n34929), .Z(n32679) );
  XNOR U34841 ( .A(n28468), .B(n34930), .Z(n34929) );
  XNOR U34842 ( .A(n34931), .B(n34932), .Z(n28468) );
  NOR U34843 ( .A(n34933), .B(n34934), .Z(n34931) );
  XOR U34844 ( .A(n32884), .B(n34935), .Z(n34928) );
  XOR U34845 ( .A(n32525), .B(n30792), .Z(n34935) );
  XNOR U34846 ( .A(n34936), .B(n34937), .Z(n30792) );
  ANDN U34847 ( .B(n34938), .A(n34939), .Z(n34936) );
  XNOR U34848 ( .A(n34940), .B(n34941), .Z(n32525) );
  XNOR U34849 ( .A(n34944), .B(n34945), .Z(n32884) );
  ANDN U34850 ( .B(n34946), .A(n34947), .Z(n34944) );
  ANDN U34851 ( .B(n28239), .A(n28139), .Z(n34903) );
  XOR U34852 ( .A(n34948), .B(n30956), .Z(n28139) );
  XNOR U34853 ( .A(n34949), .B(n34950), .Z(n30956) );
  XOR U34854 ( .A(n34951), .B(n31253), .Z(n28239) );
  IV U34855 ( .A(n34952), .Z(n31253) );
  XNOR U34856 ( .A(n25175), .B(n34953), .Z(n34853) );
  XOR U34857 ( .A(n26117), .B(n24234), .Z(n34953) );
  XNOR U34858 ( .A(n34954), .B(n26801), .Z(n24234) );
  XOR U34859 ( .A(n34955), .B(n31547), .Z(n26801) );
  XOR U34860 ( .A(n34957), .B(n34958), .Z(n33447) );
  XOR U34861 ( .A(n31668), .B(n30523), .Z(n34958) );
  XNOR U34862 ( .A(n34959), .B(n34960), .Z(n30523) );
  ANDN U34863 ( .B(n34961), .A(n34962), .Z(n34959) );
  XNOR U34864 ( .A(n34963), .B(n34964), .Z(n31668) );
  AND U34865 ( .A(n34680), .B(n34965), .Z(n34963) );
  XNOR U34866 ( .A(n33515), .B(n34966), .Z(n34957) );
  XNOR U34867 ( .A(n31218), .B(n34967), .Z(n34966) );
  XNOR U34868 ( .A(n34968), .B(n34969), .Z(n31218) );
  ANDN U34869 ( .B(n34674), .A(n34970), .Z(n34968) );
  XOR U34870 ( .A(n34971), .B(n34972), .Z(n33515) );
  ANDN U34871 ( .B(n34973), .A(n34974), .Z(n34971) );
  XNOR U34872 ( .A(n34975), .B(n31519), .Z(n26117) );
  XNOR U34873 ( .A(n31960), .B(n34976), .Z(n31519) );
  NOR U34874 ( .A(n29446), .B(n28147), .Z(n34975) );
  XOR U34875 ( .A(n34977), .B(n33834), .Z(n28147) );
  IV U34876 ( .A(n32583), .Z(n33834) );
  XOR U34877 ( .A(n34978), .B(n34374), .Z(n32583) );
  XNOR U34878 ( .A(n34979), .B(n34980), .Z(n34374) );
  XOR U34879 ( .A(n31049), .B(n29285), .Z(n34980) );
  XNOR U34880 ( .A(n34981), .B(n34982), .Z(n29285) );
  ANDN U34881 ( .B(n34983), .A(n34984), .Z(n34981) );
  XNOR U34882 ( .A(n34985), .B(n34986), .Z(n31049) );
  ANDN U34883 ( .B(n34987), .A(n34988), .Z(n34985) );
  XNOR U34884 ( .A(n34989), .B(n34990), .Z(n34979) );
  XOR U34885 ( .A(n32897), .B(n34991), .Z(n34990) );
  XNOR U34886 ( .A(n34992), .B(n33900), .Z(n32897) );
  ANDN U34887 ( .B(n34993), .A(n34994), .Z(n34992) );
  IV U34888 ( .A(n31520), .Z(n29446) );
  XNOR U34889 ( .A(n31570), .B(n33075), .Z(n31520) );
  XNOR U34890 ( .A(n34995), .B(n34996), .Z(n33075) );
  ANDN U34891 ( .B(n34997), .A(n34733), .Z(n34995) );
  XNOR U34892 ( .A(n34998), .B(n28729), .Z(n25175) );
  XNOR U34893 ( .A(n34999), .B(n31322), .Z(n28729) );
  XNOR U34894 ( .A(n30528), .B(n35000), .Z(n28154) );
  XNOR U34895 ( .A(n29324), .B(n35001), .Z(n28244) );
  XNOR U34896 ( .A(n35002), .B(n35003), .Z(n33062) );
  XNOR U34897 ( .A(n29966), .B(n32319), .Z(n35003) );
  XNOR U34898 ( .A(n35004), .B(n35005), .Z(n32319) );
  NOR U34899 ( .A(n35006), .B(n35007), .Z(n35004) );
  XNOR U34900 ( .A(n35008), .B(n35009), .Z(n29966) );
  NOR U34901 ( .A(n35010), .B(n35011), .Z(n35008) );
  XOR U34902 ( .A(n33087), .B(n35012), .Z(n35002) );
  XOR U34903 ( .A(n34791), .B(n34500), .Z(n35012) );
  XNOR U34904 ( .A(n35013), .B(n35014), .Z(n34500) );
  ANDN U34905 ( .B(n35015), .A(n35016), .Z(n35013) );
  XNOR U34906 ( .A(n35017), .B(n35018), .Z(n34791) );
  ANDN U34907 ( .B(n35019), .A(n35020), .Z(n35017) );
  XOR U34908 ( .A(n35021), .B(n35022), .Z(n33087) );
  ANDN U34909 ( .B(n35023), .A(n35024), .Z(n35021) );
  XNOR U34910 ( .A(n35025), .B(n35026), .Z(n34403) );
  XNOR U34911 ( .A(n33510), .B(n34216), .Z(n35026) );
  XOR U34912 ( .A(n35027), .B(n35028), .Z(n34216) );
  ANDN U34913 ( .B(n35029), .A(n35030), .Z(n35027) );
  XNOR U34914 ( .A(n35031), .B(n35032), .Z(n33510) );
  ANDN U34915 ( .B(n35033), .A(n35034), .Z(n35031) );
  XOR U34916 ( .A(n32336), .B(n35035), .Z(n35025) );
  XOR U34917 ( .A(n30538), .B(n35036), .Z(n35035) );
  XNOR U34918 ( .A(n35037), .B(n35038), .Z(n30538) );
  NOR U34919 ( .A(n35039), .B(n35040), .Z(n35037) );
  XOR U34920 ( .A(n35041), .B(n35042), .Z(n32336) );
  XNOR U34921 ( .A(n35045), .B(n35046), .Z(n26588) );
  XOR U34922 ( .A(n28366), .B(n27641), .Z(n35046) );
  XOR U34923 ( .A(n35047), .B(n28397), .Z(n27641) );
  XNOR U34924 ( .A(n35048), .B(n29284), .Z(n28397) );
  IV U34925 ( .A(n31698), .Z(n29284) );
  XNOR U34926 ( .A(n35049), .B(n32550), .Z(n31698) );
  XOR U34927 ( .A(n35050), .B(n35051), .Z(n32550) );
  XNOR U34928 ( .A(n30221), .B(n34524), .Z(n35051) );
  XNOR U34929 ( .A(n35052), .B(n35053), .Z(n34524) );
  ANDN U34930 ( .B(n35054), .A(n35055), .Z(n35052) );
  XNOR U34931 ( .A(n35056), .B(n35057), .Z(n30221) );
  ANDN U34932 ( .B(n35058), .A(n35059), .Z(n35056) );
  XOR U34933 ( .A(n31635), .B(n35060), .Z(n35050) );
  XNOR U34934 ( .A(n29328), .B(n32850), .Z(n35060) );
  XOR U34935 ( .A(n35061), .B(n35062), .Z(n32850) );
  XOR U34936 ( .A(n35065), .B(n35066), .Z(n29328) );
  ANDN U34937 ( .B(n35067), .A(n35068), .Z(n35065) );
  AND U34938 ( .A(n35071), .B(n35072), .Z(n35069) );
  ANDN U34939 ( .B(n27509), .A(n27507), .Z(n35047) );
  XNOR U34940 ( .A(n33316), .B(n32166), .Z(n27507) );
  IV U34941 ( .A(n31555), .Z(n32166) );
  XNOR U34942 ( .A(n34170), .B(n33710), .Z(n31555) );
  XNOR U34943 ( .A(n35073), .B(n35074), .Z(n33710) );
  XNOR U34944 ( .A(n31603), .B(n34976), .Z(n35074) );
  XNOR U34945 ( .A(n35075), .B(n35076), .Z(n34976) );
  ANDN U34946 ( .B(n33320), .A(n33321), .Z(n35075) );
  XOR U34947 ( .A(n35077), .B(n35078), .Z(n33321) );
  XNOR U34948 ( .A(n35079), .B(n35080), .Z(n31603) );
  NOR U34949 ( .A(n33315), .B(n33313), .Z(n35079) );
  XNOR U34950 ( .A(n35081), .B(n35082), .Z(n33315) );
  XOR U34951 ( .A(n31360), .B(n35083), .Z(n35073) );
  XOR U34952 ( .A(n31959), .B(n35084), .Z(n35083) );
  XOR U34953 ( .A(n35085), .B(n35086), .Z(n31959) );
  ANDN U34954 ( .B(n34151), .A(n35087), .Z(n35085) );
  XOR U34955 ( .A(n35088), .B(n35089), .Z(n34151) );
  XNOR U34956 ( .A(n35090), .B(n35091), .Z(n31360) );
  NOR U34957 ( .A(n33546), .B(n33547), .Z(n35090) );
  XNOR U34958 ( .A(n35092), .B(n35093), .Z(n33547) );
  XNOR U34959 ( .A(n35094), .B(n35095), .Z(n34170) );
  XNOR U34960 ( .A(n32859), .B(n35096), .Z(n35095) );
  XOR U34961 ( .A(n35097), .B(n35098), .Z(n32859) );
  ANDN U34962 ( .B(n33435), .A(n33436), .Z(n35097) );
  XOR U34963 ( .A(n30962), .B(n35099), .Z(n35094) );
  XNOR U34964 ( .A(n33704), .B(n33187), .Z(n35099) );
  XOR U34965 ( .A(n35100), .B(n35101), .Z(n33187) );
  XNOR U34966 ( .A(n35102), .B(n35103), .Z(n33704) );
  ANDN U34967 ( .B(n33425), .A(n35104), .Z(n35102) );
  XNOR U34968 ( .A(n35105), .B(n35106), .Z(n30962) );
  XNOR U34969 ( .A(n35107), .B(n35108), .Z(n33316) );
  AND U34970 ( .A(n34143), .B(n34142), .Z(n35107) );
  XOR U34971 ( .A(n30491), .B(n35109), .Z(n27509) );
  XNOR U34972 ( .A(n35110), .B(n28384), .Z(n28366) );
  XOR U34973 ( .A(n32101), .B(n35111), .Z(n28384) );
  XOR U34974 ( .A(n35112), .B(n35113), .Z(n32754) );
  XNOR U34975 ( .A(n35114), .B(n32721), .Z(n35113) );
  XNOR U34976 ( .A(n35115), .B(n34057), .Z(n32721) );
  AND U34977 ( .A(n35116), .B(n35117), .Z(n35115) );
  XNOR U34978 ( .A(n33223), .B(n35118), .Z(n35112) );
  XOR U34979 ( .A(n31583), .B(n35119), .Z(n35118) );
  XNOR U34980 ( .A(n35120), .B(n35121), .Z(n31583) );
  ANDN U34981 ( .B(n35122), .A(n35123), .Z(n35120) );
  XNOR U34982 ( .A(n35124), .B(n34051), .Z(n33223) );
  ANDN U34983 ( .B(n35125), .A(n35126), .Z(n35124) );
  XNOR U34984 ( .A(n35127), .B(n35128), .Z(n33742) );
  XOR U34985 ( .A(n31252), .B(n34951), .Z(n35128) );
  XOR U34986 ( .A(n35129), .B(n35130), .Z(n34951) );
  ANDN U34987 ( .B(n35131), .A(n35132), .Z(n35129) );
  XNOR U34988 ( .A(n35133), .B(n35134), .Z(n31252) );
  NOR U34989 ( .A(n35135), .B(n35136), .Z(n35133) );
  XOR U34990 ( .A(n32613), .B(n35137), .Z(n35127) );
  XOR U34991 ( .A(n32888), .B(n35138), .Z(n35137) );
  XNOR U34992 ( .A(n35139), .B(n35140), .Z(n32888) );
  XNOR U34993 ( .A(n35143), .B(n35144), .Z(n32613) );
  ANDN U34994 ( .B(n35145), .A(n35146), .Z(n35143) );
  ANDN U34995 ( .B(n27494), .A(n29509), .Z(n35110) );
  IV U34996 ( .A(n27496), .Z(n29509) );
  XOR U34997 ( .A(n33698), .B(n34446), .Z(n27496) );
  XNOR U34998 ( .A(n35147), .B(n35148), .Z(n34446) );
  ANDN U34999 ( .B(n34701), .A(n34699), .Z(n35147) );
  XOR U35000 ( .A(n34135), .B(n35149), .Z(n33698) );
  XOR U35001 ( .A(n35150), .B(n35151), .Z(n34135) );
  XNOR U35002 ( .A(n32414), .B(n31877), .Z(n35151) );
  XOR U35003 ( .A(n35152), .B(n35153), .Z(n31877) );
  AND U35004 ( .A(n34461), .B(n34463), .Z(n35152) );
  XOR U35005 ( .A(n35154), .B(n35155), .Z(n34463) );
  XOR U35006 ( .A(n35156), .B(n35157), .Z(n32414) );
  AND U35007 ( .A(n34448), .B(n34450), .Z(n35156) );
  XOR U35008 ( .A(n35158), .B(n35159), .Z(n34450) );
  XOR U35009 ( .A(n35160), .B(n35161), .Z(n35150) );
  XNOR U35010 ( .A(n32483), .B(n29174), .Z(n35161) );
  XOR U35011 ( .A(n35162), .B(n35163), .Z(n29174) );
  AND U35012 ( .A(n34453), .B(n34455), .Z(n35162) );
  XOR U35013 ( .A(n35164), .B(n35165), .Z(n34455) );
  XNOR U35014 ( .A(n35166), .B(n35167), .Z(n32483) );
  AND U35015 ( .A(n34459), .B(n34457), .Z(n35166) );
  XOR U35016 ( .A(n35168), .B(n35082), .Z(n34459) );
  XOR U35017 ( .A(n35169), .B(n31322), .Z(n27494) );
  XNOR U35018 ( .A(n35170), .B(n35171), .Z(n34690) );
  XOR U35019 ( .A(n31526), .B(n32532), .Z(n35171) );
  XNOR U35020 ( .A(n35172), .B(n35173), .Z(n32532) );
  XNOR U35021 ( .A(n35176), .B(n34473), .Z(n31526) );
  NOR U35022 ( .A(n34472), .B(n35177), .Z(n35176) );
  XNOR U35023 ( .A(n33148), .B(n35178), .Z(n35170) );
  XOR U35024 ( .A(n30147), .B(n33770), .Z(n35178) );
  XNOR U35025 ( .A(n35179), .B(n34468), .Z(n33770) );
  ANDN U35026 ( .B(n35180), .A(n34469), .Z(n35179) );
  XNOR U35027 ( .A(n35181), .B(n35182), .Z(n30147) );
  ANDN U35028 ( .B(n35183), .A(n35184), .Z(n35181) );
  XNOR U35029 ( .A(n35185), .B(n34479), .Z(n33148) );
  ANDN U35030 ( .B(n34480), .A(n35186), .Z(n35185) );
  XOR U35031 ( .A(n25022), .B(n35188), .Z(n35045) );
  XOR U35032 ( .A(n27336), .B(n26279), .Z(n35188) );
  XNOR U35033 ( .A(n35189), .B(n28394), .Z(n26279) );
  XOR U35034 ( .A(n35191), .B(n33329), .Z(n29045) );
  XOR U35035 ( .A(n35192), .B(n35193), .Z(n33329) );
  XOR U35036 ( .A(n31953), .B(n30553), .Z(n35193) );
  XOR U35037 ( .A(n35194), .B(n35195), .Z(n30553) );
  NOR U35038 ( .A(n35196), .B(n35197), .Z(n35194) );
  XNOR U35039 ( .A(n35198), .B(n35199), .Z(n31953) );
  NOR U35040 ( .A(n35200), .B(n35201), .Z(n35198) );
  XOR U35041 ( .A(n35202), .B(n35203), .Z(n35192) );
  XOR U35042 ( .A(n31979), .B(n32988), .Z(n35203) );
  XNOR U35043 ( .A(n35204), .B(n35205), .Z(n32988) );
  ANDN U35044 ( .B(n35206), .A(n35207), .Z(n35204) );
  XNOR U35045 ( .A(n35208), .B(n35209), .Z(n31979) );
  NOR U35046 ( .A(n35210), .B(n35211), .Z(n35208) );
  AND U35047 ( .A(n27499), .B(n27500), .Z(n35189) );
  XNOR U35048 ( .A(n28807), .B(n35212), .Z(n27500) );
  XOR U35049 ( .A(n33102), .B(n31355), .Z(n27499) );
  XOR U35050 ( .A(n35213), .B(n35214), .Z(n33102) );
  ANDN U35051 ( .B(n35215), .A(n35216), .Z(n35213) );
  XOR U35052 ( .A(n35217), .B(n28387), .Z(n27336) );
  XOR U35053 ( .A(n28435), .B(n34383), .Z(n28387) );
  XNOR U35054 ( .A(n35218), .B(n34411), .Z(n34383) );
  IV U35055 ( .A(n30562), .Z(n28435) );
  ANDN U35056 ( .B(n27492), .A(n27490), .Z(n35217) );
  XNOR U35057 ( .A(n34127), .B(n30165), .Z(n27490) );
  XNOR U35058 ( .A(n35221), .B(n35222), .Z(n34127) );
  ANDN U35059 ( .B(n35223), .A(n34544), .Z(n35221) );
  XOR U35060 ( .A(n33805), .B(n32216), .Z(n27492) );
  XNOR U35061 ( .A(n35224), .B(n33280), .Z(n33805) );
  NOR U35062 ( .A(n35225), .B(n35226), .Z(n35224) );
  XNOR U35063 ( .A(n35227), .B(n28391), .Z(n25022) );
  XOR U35064 ( .A(n35138), .B(n34952), .Z(n28391) );
  XOR U35065 ( .A(n33599), .B(n35228), .Z(n34952) );
  XOR U35066 ( .A(n35229), .B(n35230), .Z(n33599) );
  XOR U35067 ( .A(n32828), .B(n33517), .Z(n35230) );
  XNOR U35068 ( .A(n35231), .B(n35232), .Z(n33517) );
  AND U35069 ( .A(n33750), .B(n33752), .Z(n35231) );
  XOR U35070 ( .A(n35233), .B(n35234), .Z(n32828) );
  ANDN U35071 ( .B(n33760), .A(n35235), .Z(n35233) );
  XNOR U35072 ( .A(n33720), .B(n35236), .Z(n35229) );
  XOR U35073 ( .A(n33879), .B(n33002), .Z(n35236) );
  XNOR U35074 ( .A(n35237), .B(n35238), .Z(n33002) );
  NOR U35075 ( .A(n33746), .B(n33747), .Z(n35237) );
  XOR U35076 ( .A(n35239), .B(n35240), .Z(n33879) );
  ANDN U35077 ( .B(n33765), .A(n35241), .Z(n35239) );
  XOR U35078 ( .A(n35242), .B(n35243), .Z(n33720) );
  ANDN U35079 ( .B(n33755), .A(n33756), .Z(n35242) );
  XOR U35080 ( .A(n35244), .B(n35245), .Z(n35138) );
  NOR U35081 ( .A(n35246), .B(n35247), .Z(n35244) );
  ANDN U35082 ( .B(n27505), .A(n27503), .Z(n35227) );
  XOR U35083 ( .A(n35248), .B(n31663), .Z(n27503) );
  IV U35084 ( .A(n28802), .Z(n31663) );
  XOR U35085 ( .A(n35249), .B(n34956), .Z(n28802) );
  XNOR U35086 ( .A(n35250), .B(n35251), .Z(n34956) );
  XNOR U35087 ( .A(n34608), .B(n33014), .Z(n35251) );
  XNOR U35088 ( .A(n35252), .B(n35253), .Z(n33014) );
  ANDN U35089 ( .B(n35254), .A(n35255), .Z(n35252) );
  XNOR U35090 ( .A(n35256), .B(n35257), .Z(n34608) );
  ANDN U35091 ( .B(n35258), .A(n35259), .Z(n35256) );
  XOR U35092 ( .A(n32927), .B(n35260), .Z(n35250) );
  XOR U35093 ( .A(n34664), .B(n31739), .Z(n35260) );
  XNOR U35094 ( .A(n35261), .B(n35262), .Z(n31739) );
  NOR U35095 ( .A(n35263), .B(n35264), .Z(n35261) );
  XOR U35096 ( .A(n35265), .B(n35266), .Z(n34664) );
  ANDN U35097 ( .B(n35267), .A(n35268), .Z(n35265) );
  XNOR U35098 ( .A(n35269), .B(n35270), .Z(n32927) );
  ANDN U35099 ( .B(n35271), .A(n35272), .Z(n35269) );
  XOR U35100 ( .A(n33592), .B(n31116), .Z(n27505) );
  XNOR U35101 ( .A(n35273), .B(n35274), .Z(n32924) );
  XOR U35102 ( .A(n31965), .B(n33296), .Z(n35274) );
  XNOR U35103 ( .A(n35275), .B(n35276), .Z(n33296) );
  ANDN U35104 ( .B(n33596), .A(n35277), .Z(n35275) );
  XNOR U35105 ( .A(n35278), .B(n35279), .Z(n31965) );
  ANDN U35106 ( .B(n33726), .A(n33725), .Z(n35278) );
  XNOR U35107 ( .A(n31743), .B(n35280), .Z(n35273) );
  XOR U35108 ( .A(n31946), .B(n28763), .Z(n35280) );
  XOR U35109 ( .A(n35281), .B(n35282), .Z(n28763) );
  ANDN U35110 ( .B(n34434), .A(n34435), .Z(n35281) );
  XOR U35111 ( .A(n35283), .B(n35284), .Z(n31946) );
  ANDN U35112 ( .B(n33587), .A(n33588), .Z(n35283) );
  XNOR U35113 ( .A(n35285), .B(n35286), .Z(n31743) );
  ANDN U35114 ( .B(n35287), .A(n35288), .Z(n35285) );
  XOR U35115 ( .A(n35290), .B(n35287), .Z(n33592) );
  ANDN U35116 ( .B(n35288), .A(n35291), .Z(n35290) );
  XNOR U35117 ( .A(n35292), .B(n26802), .Z(n28241) );
  XNOR U35118 ( .A(n34838), .B(n32139), .Z(n26802) );
  XOR U35119 ( .A(n32969), .B(n34088), .Z(n32139) );
  XNOR U35120 ( .A(n35293), .B(n35294), .Z(n34088) );
  XNOR U35121 ( .A(n30150), .B(n34612), .Z(n35294) );
  XNOR U35122 ( .A(n35295), .B(n34644), .Z(n34612) );
  ANDN U35123 ( .B(n34832), .A(n34830), .Z(n35295) );
  XOR U35124 ( .A(n35296), .B(n35297), .Z(n34830) );
  XNOR U35125 ( .A(n35298), .B(n35299), .Z(n30150) );
  NOR U35126 ( .A(n34834), .B(n34648), .Z(n35298) );
  XNOR U35127 ( .A(n35300), .B(n35301), .Z(n34648) );
  XOR U35128 ( .A(n32134), .B(n35302), .Z(n35293) );
  XOR U35129 ( .A(n32732), .B(n32724), .Z(n35302) );
  XNOR U35130 ( .A(n35303), .B(n34657), .Z(n32724) );
  ANDN U35131 ( .B(n34658), .A(n34827), .Z(n35303) );
  XNOR U35132 ( .A(n35304), .B(n35305), .Z(n34658) );
  XNOR U35133 ( .A(n35306), .B(n34653), .Z(n32732) );
  NOR U35134 ( .A(n34654), .B(n34820), .Z(n35306) );
  XNOR U35135 ( .A(n35307), .B(n35308), .Z(n34654) );
  XNOR U35136 ( .A(n35309), .B(n34662), .Z(n32134) );
  ANDN U35137 ( .B(n34661), .A(n34824), .Z(n35309) );
  XNOR U35138 ( .A(n35310), .B(n35311), .Z(n34661) );
  XOR U35139 ( .A(n35312), .B(n35313), .Z(n32969) );
  XNOR U35140 ( .A(n33963), .B(n31227), .Z(n35313) );
  XNOR U35141 ( .A(n35314), .B(n33975), .Z(n31227) );
  ANDN U35142 ( .B(n34848), .A(n33976), .Z(n35314) );
  XOR U35143 ( .A(n35315), .B(n35316), .Z(n33976) );
  IV U35144 ( .A(n35317), .Z(n34848) );
  XNOR U35145 ( .A(n35318), .B(n33983), .Z(n33963) );
  XOR U35146 ( .A(n35319), .B(n35320), .Z(n33984) );
  XOR U35147 ( .A(n32495), .B(n35321), .Z(n35312) );
  XOR U35148 ( .A(n31625), .B(n30232), .Z(n35321) );
  XNOR U35149 ( .A(n35322), .B(n33971), .Z(n30232) );
  ANDN U35150 ( .B(n34841), .A(n33970), .Z(n35322) );
  XNOR U35151 ( .A(n35323), .B(n35324), .Z(n33970) );
  XNOR U35152 ( .A(n35325), .B(n35326), .Z(n31625) );
  NOR U35153 ( .A(n35327), .B(n35328), .Z(n35325) );
  XNOR U35154 ( .A(n35329), .B(n33980), .Z(n32495) );
  NOR U35155 ( .A(n34851), .B(n33979), .Z(n35329) );
  XOR U35156 ( .A(n35330), .B(n35331), .Z(n33979) );
  XNOR U35157 ( .A(n35332), .B(n35327), .Z(n34838) );
  ANDN U35158 ( .B(n35328), .A(n35333), .Z(n35332) );
  ANDN U35159 ( .B(n28144), .A(n28143), .Z(n35292) );
  XOR U35160 ( .A(n35334), .B(n29053), .Z(n28143) );
  IV U35161 ( .A(n29024), .Z(n29053) );
  XNOR U35162 ( .A(n33146), .B(n35335), .Z(n29024) );
  XOR U35163 ( .A(n35336), .B(n35337), .Z(n33146) );
  XOR U35164 ( .A(n31456), .B(n33741), .Z(n35337) );
  XNOR U35165 ( .A(n35338), .B(n35131), .Z(n33741) );
  ANDN U35166 ( .B(n35339), .A(n35340), .Z(n35338) );
  XNOR U35167 ( .A(n35341), .B(n35135), .Z(n31456) );
  ANDN U35168 ( .B(n35136), .A(n35342), .Z(n35341) );
  XNOR U35169 ( .A(n33088), .B(n35343), .Z(n35336) );
  XOR U35170 ( .A(n32767), .B(n33016), .Z(n35343) );
  XOR U35171 ( .A(n35344), .B(n35142), .Z(n33016) );
  ANDN U35172 ( .B(n35345), .A(n35141), .Z(n35344) );
  IV U35173 ( .A(n35346), .Z(n35141) );
  XNOR U35174 ( .A(n35347), .B(n35246), .Z(n32767) );
  ANDN U35175 ( .B(n35247), .A(n35348), .Z(n35347) );
  XNOR U35176 ( .A(n35349), .B(n35146), .Z(n33088) );
  NOR U35177 ( .A(n35350), .B(n35145), .Z(n35349) );
  XNOR U35178 ( .A(n35351), .B(n30075), .Z(n28144) );
  IV U35179 ( .A(n31226), .Z(n30075) );
  XOR U35180 ( .A(n35352), .B(n35353), .Z(n31226) );
  IV U35181 ( .A(n25129), .Z(n25921) );
  XOR U35182 ( .A(n25289), .B(n28465), .Z(n25129) );
  XNOR U35183 ( .A(n35354), .B(n28751), .Z(n28465) );
  XOR U35184 ( .A(n33389), .B(n28798), .Z(n26606) );
  IV U35185 ( .A(n30505), .Z(n28798) );
  XNOR U35186 ( .A(n35355), .B(n35356), .Z(n33389) );
  IV U35187 ( .A(n26904), .Z(n25289) );
  XNOR U35188 ( .A(n35358), .B(n35359), .Z(n29502) );
  XOR U35189 ( .A(n24837), .B(n22991), .Z(n35359) );
  XOR U35190 ( .A(n35360), .B(n26604), .Z(n22991) );
  XOR U35191 ( .A(n35361), .B(n30375), .Z(n26604) );
  XNOR U35192 ( .A(n34857), .B(n34364), .Z(n30375) );
  XNOR U35193 ( .A(n35362), .B(n35363), .Z(n34364) );
  XOR U35194 ( .A(n32195), .B(n31163), .Z(n35363) );
  XOR U35195 ( .A(n35364), .B(n33918), .Z(n31163) );
  ANDN U35196 ( .B(n32674), .A(n32672), .Z(n35364) );
  XNOR U35197 ( .A(n35365), .B(n35366), .Z(n32674) );
  XOR U35198 ( .A(n35367), .B(n33928), .Z(n32195) );
  AND U35199 ( .A(n33419), .B(n33417), .Z(n35367) );
  XOR U35200 ( .A(n35368), .B(n35369), .Z(n33419) );
  XNOR U35201 ( .A(n32917), .B(n35370), .Z(n35362) );
  XOR U35202 ( .A(n34016), .B(n34794), .Z(n35370) );
  XNOR U35203 ( .A(n35371), .B(n33923), .Z(n34794) );
  ANDN U35204 ( .B(n32659), .A(n32660), .Z(n35371) );
  IV U35205 ( .A(n33497), .Z(n32660) );
  XOR U35206 ( .A(n35372), .B(n35373), .Z(n33497) );
  XNOR U35207 ( .A(n35374), .B(n33914), .Z(n34016) );
  AND U35208 ( .A(n33503), .B(n34366), .Z(n35374) );
  XNOR U35209 ( .A(n35375), .B(n35376), .Z(n33503) );
  XOR U35210 ( .A(n35377), .B(n33932), .Z(n32917) );
  ANDN U35211 ( .B(n32655), .A(n32656), .Z(n35377) );
  XOR U35212 ( .A(n35378), .B(n35379), .Z(n32656) );
  XOR U35213 ( .A(n35380), .B(n35381), .Z(n34857) );
  XNOR U35214 ( .A(n32799), .B(n32312), .Z(n35381) );
  XOR U35215 ( .A(n35382), .B(n33871), .Z(n32312) );
  ANDN U35216 ( .B(n35383), .A(n35384), .Z(n35382) );
  XNOR U35217 ( .A(n35385), .B(n33857), .Z(n32799) );
  ANDN U35218 ( .B(n35386), .A(n35387), .Z(n35385) );
  XNOR U35219 ( .A(n35388), .B(n35389), .Z(n35380) );
  XOR U35220 ( .A(n29019), .B(n33046), .Z(n35389) );
  XNOR U35221 ( .A(n35390), .B(n33866), .Z(n33046) );
  XNOR U35222 ( .A(n35392), .B(n33861), .Z(n29019) );
  ANDN U35223 ( .B(n34012), .A(n35393), .Z(n35392) );
  ANDN U35224 ( .B(n28737), .A(n28475), .Z(n35360) );
  XOR U35225 ( .A(n35397), .B(n30027), .Z(n28737) );
  IV U35226 ( .A(n30662), .Z(n30027) );
  XNOR U35227 ( .A(n35398), .B(n26594), .Z(n24837) );
  XOR U35228 ( .A(n35399), .B(n29271), .Z(n26594) );
  XNOR U35229 ( .A(n33702), .B(n34177), .Z(n29271) );
  XNOR U35230 ( .A(n35400), .B(n35401), .Z(n34177) );
  XOR U35231 ( .A(n35402), .B(n31648), .Z(n35401) );
  XNOR U35232 ( .A(n35403), .B(n35404), .Z(n31648) );
  NOR U35233 ( .A(n35405), .B(n35406), .Z(n35403) );
  XNOR U35234 ( .A(n31166), .B(n35407), .Z(n35400) );
  XNOR U35235 ( .A(n28884), .B(n30647), .Z(n35407) );
  XNOR U35236 ( .A(n35408), .B(n35409), .Z(n30647) );
  ANDN U35237 ( .B(n35410), .A(n35411), .Z(n35408) );
  XNOR U35238 ( .A(n35412), .B(n35413), .Z(n28884) );
  ANDN U35239 ( .B(n35414), .A(n35415), .Z(n35412) );
  XOR U35240 ( .A(n35416), .B(n35417), .Z(n31166) );
  ANDN U35241 ( .B(n35418), .A(n35419), .Z(n35416) );
  XOR U35242 ( .A(n35420), .B(n35421), .Z(n33702) );
  XNOR U35243 ( .A(n35109), .B(n30492), .Z(n35421) );
  XNOR U35244 ( .A(n35422), .B(n34202), .Z(n30492) );
  ANDN U35245 ( .B(n35423), .A(n35424), .Z(n35422) );
  XNOR U35246 ( .A(n35425), .B(n34206), .Z(n35109) );
  ANDN U35247 ( .B(n35426), .A(n35427), .Z(n35425) );
  XOR U35248 ( .A(n32541), .B(n35428), .Z(n35420) );
  XOR U35249 ( .A(n32762), .B(n35429), .Z(n35428) );
  XNOR U35250 ( .A(n35430), .B(n34209), .Z(n32762) );
  ANDN U35251 ( .B(n35431), .A(n35432), .Z(n35430) );
  XOR U35252 ( .A(n35433), .B(n34193), .Z(n32541) );
  ANDN U35253 ( .B(n35434), .A(n35435), .Z(n35433) );
  ANDN U35254 ( .B(n28370), .A(n28467), .Z(n35398) );
  XOR U35255 ( .A(n30865), .B(n33887), .Z(n28467) );
  XNOR U35256 ( .A(n35436), .B(n35437), .Z(n33887) );
  XNOR U35257 ( .A(n30501), .B(n35439), .Z(n28370) );
  XNOR U35258 ( .A(n33603), .B(n32617), .Z(n30501) );
  XNOR U35259 ( .A(n35440), .B(n35441), .Z(n32617) );
  XOR U35260 ( .A(n35442), .B(n35443), .Z(n35441) );
  XOR U35261 ( .A(n30942), .B(n35444), .Z(n35440) );
  XOR U35262 ( .A(n31821), .B(n32944), .Z(n35444) );
  XNOR U35263 ( .A(n35445), .B(n35446), .Z(n32944) );
  NOR U35264 ( .A(n35447), .B(n34579), .Z(n35445) );
  XNOR U35265 ( .A(n35448), .B(n35449), .Z(n31821) );
  ANDN U35266 ( .B(n35450), .A(n34583), .Z(n35448) );
  IV U35267 ( .A(n35451), .Z(n34583) );
  XNOR U35268 ( .A(n35452), .B(n35453), .Z(n30942) );
  ANDN U35269 ( .B(n34592), .A(n35454), .Z(n35452) );
  XOR U35270 ( .A(n35455), .B(n35456), .Z(n33603) );
  XNOR U35271 ( .A(n32181), .B(n33094), .Z(n35456) );
  XOR U35272 ( .A(n35457), .B(n32473), .Z(n33094) );
  XNOR U35273 ( .A(n35460), .B(n32478), .Z(n32181) );
  XOR U35274 ( .A(n35463), .B(n35464), .Z(n35455) );
  XOR U35275 ( .A(n31864), .B(n32320), .Z(n35464) );
  XNOR U35276 ( .A(n35465), .B(n32467), .Z(n32320) );
  NOR U35277 ( .A(n35466), .B(n35467), .Z(n35465) );
  XNOR U35278 ( .A(n35468), .B(n34601), .Z(n31864) );
  NOR U35279 ( .A(n35469), .B(n35470), .Z(n35468) );
  XNOR U35280 ( .A(n27103), .B(n35471), .Z(n35358) );
  XOR U35281 ( .A(n24592), .B(n28730), .Z(n35471) );
  XOR U35282 ( .A(n35472), .B(n26608), .Z(n28730) );
  XNOR U35283 ( .A(n35473), .B(n31772), .Z(n26608) );
  ANDN U35284 ( .B(n28751), .A(n28376), .Z(n35472) );
  XNOR U35285 ( .A(n29047), .B(n34773), .Z(n28376) );
  XNOR U35286 ( .A(n35474), .B(n35475), .Z(n34773) );
  ANDN U35287 ( .B(n33693), .A(n35476), .Z(n35474) );
  XOR U35288 ( .A(n34528), .B(n34166), .Z(n29047) );
  XOR U35289 ( .A(n35477), .B(n35478), .Z(n34166) );
  XOR U35290 ( .A(n29298), .B(n32710), .Z(n35478) );
  XOR U35291 ( .A(n35479), .B(n35480), .Z(n32710) );
  ANDN U35292 ( .B(n34307), .A(n34308), .Z(n35479) );
  XNOR U35293 ( .A(n35481), .B(n35482), .Z(n29298) );
  AND U35294 ( .A(n34300), .B(n34298), .Z(n35481) );
  XNOR U35295 ( .A(n30299), .B(n35483), .Z(n35477) );
  XOR U35296 ( .A(n33269), .B(n31328), .Z(n35483) );
  XOR U35297 ( .A(n35484), .B(n35485), .Z(n31328) );
  AND U35298 ( .A(n34317), .B(n34315), .Z(n35484) );
  XNOR U35299 ( .A(n35486), .B(n35487), .Z(n33269) );
  AND U35300 ( .A(n34304), .B(n34302), .Z(n35486) );
  XOR U35301 ( .A(n35488), .B(n35489), .Z(n30299) );
  AND U35302 ( .A(n34313), .B(n34311), .Z(n35488) );
  XOR U35303 ( .A(n35490), .B(n35491), .Z(n34528) );
  XNOR U35304 ( .A(n30670), .B(n35492), .Z(n35491) );
  XNOR U35305 ( .A(n35493), .B(n33682), .Z(n30670) );
  ANDN U35306 ( .B(n34775), .A(n34776), .Z(n35493) );
  XNOR U35307 ( .A(n32281), .B(n35494), .Z(n35490) );
  XOR U35308 ( .A(n32809), .B(n32017), .Z(n35494) );
  XOR U35309 ( .A(n35495), .B(n33687), .Z(n32017) );
  AND U35310 ( .A(n34782), .B(n34783), .Z(n35495) );
  XNOR U35311 ( .A(n35496), .B(n34182), .Z(n32809) );
  XOR U35312 ( .A(n35497), .B(n33694), .Z(n32281) );
  ANDN U35313 ( .B(n35475), .A(n35498), .Z(n35497) );
  XOR U35314 ( .A(n35499), .B(n28881), .Z(n28751) );
  XNOR U35315 ( .A(n35500), .B(n35501), .Z(n28881) );
  XNOR U35316 ( .A(n35502), .B(n27063), .Z(n24592) );
  XNOR U35317 ( .A(n30562), .B(n34377), .Z(n27063) );
  XOR U35318 ( .A(n35503), .B(n34419), .Z(n34377) );
  ANDN U35319 ( .B(n35504), .A(n35505), .Z(n35503) );
  XOR U35320 ( .A(n32948), .B(n35506), .Z(n30562) );
  XOR U35321 ( .A(n35507), .B(n35508), .Z(n32948) );
  XOR U35322 ( .A(n30740), .B(n33883), .Z(n35508) );
  XNOR U35323 ( .A(n35509), .B(n34420), .Z(n33883) );
  ANDN U35324 ( .B(n35505), .A(n34419), .Z(n35509) );
  XNOR U35325 ( .A(n35510), .B(n35511), .Z(n34419) );
  IV U35326 ( .A(n35512), .Z(n35505) );
  XNOR U35327 ( .A(n35513), .B(n35514), .Z(n30740) );
  ANDN U35328 ( .B(n34379), .A(n34380), .Z(n35513) );
  XOR U35329 ( .A(n35515), .B(n35516), .Z(n34379) );
  XOR U35330 ( .A(n30953), .B(n35517), .Z(n35507) );
  XNOR U35331 ( .A(n32282), .B(n30686), .Z(n35517) );
  XNOR U35332 ( .A(n35518), .B(n34412), .Z(n30686) );
  ANDN U35333 ( .B(n34411), .A(n35219), .Z(n35518) );
  XNOR U35334 ( .A(n35519), .B(n35520), .Z(n34411) );
  XNOR U35335 ( .A(n35521), .B(n34416), .Z(n32282) );
  NOR U35336 ( .A(n34386), .B(n34385), .Z(n35521) );
  XNOR U35337 ( .A(n35522), .B(n35523), .Z(n34385) );
  XNOR U35338 ( .A(n35524), .B(n34408), .Z(n30953) );
  ANDN U35339 ( .B(n34389), .A(n34390), .Z(n35524) );
  XOR U35340 ( .A(n35525), .B(n35526), .Z(n34389) );
  ANDN U35341 ( .B(n28460), .A(n28463), .Z(n35502) );
  XNOR U35342 ( .A(n35527), .B(n29717), .Z(n28463) );
  XOR U35343 ( .A(n32894), .B(n33512), .Z(n29717) );
  XNOR U35344 ( .A(n35528), .B(n35529), .Z(n33512) );
  XOR U35345 ( .A(n31439), .B(n32394), .Z(n35529) );
  XOR U35346 ( .A(n35530), .B(n34174), .Z(n32394) );
  XNOR U35347 ( .A(n35532), .B(n33427), .Z(n31439) );
  ANDN U35348 ( .B(n35533), .A(n35103), .Z(n35532) );
  XOR U35349 ( .A(n35534), .B(n35535), .Z(n35528) );
  XNOR U35350 ( .A(n33122), .B(n31572), .Z(n35535) );
  XNOR U35351 ( .A(n35536), .B(n33437), .Z(n31572) );
  ANDN U35352 ( .B(n35098), .A(n35537), .Z(n35536) );
  XNOR U35353 ( .A(n35538), .B(n33431), .Z(n33122) );
  NOR U35354 ( .A(n35106), .B(n35539), .Z(n35538) );
  XNOR U35355 ( .A(n35540), .B(n35541), .Z(n32894) );
  XOR U35356 ( .A(n32592), .B(n35542), .Z(n35541) );
  XNOR U35357 ( .A(n35543), .B(n35544), .Z(n32592) );
  ANDN U35358 ( .B(n35545), .A(n35546), .Z(n35543) );
  XOR U35359 ( .A(n28424), .B(n35547), .Z(n35540) );
  XOR U35360 ( .A(n33737), .B(n33549), .Z(n35547) );
  XNOR U35361 ( .A(n35548), .B(n35549), .Z(n33549) );
  ANDN U35362 ( .B(n35550), .A(n35551), .Z(n35548) );
  XNOR U35363 ( .A(n35552), .B(n35553), .Z(n33737) );
  ANDN U35364 ( .B(n35554), .A(n35555), .Z(n35552) );
  XNOR U35365 ( .A(n35556), .B(n35557), .Z(n28424) );
  ANDN U35366 ( .B(n35558), .A(n35559), .Z(n35556) );
  XOR U35367 ( .A(n31666), .B(n35560), .Z(n28460) );
  XOR U35368 ( .A(n33328), .B(n35561), .Z(n31666) );
  XOR U35369 ( .A(n35562), .B(n35563), .Z(n33328) );
  XNOR U35370 ( .A(n29961), .B(n35564), .Z(n35563) );
  XNOR U35371 ( .A(n35565), .B(n35566), .Z(n29961) );
  ANDN U35372 ( .B(n35066), .A(n35567), .Z(n35565) );
  XOR U35373 ( .A(n32791), .B(n35568), .Z(n35562) );
  XOR U35374 ( .A(n32690), .B(n35569), .Z(n35568) );
  XNOR U35375 ( .A(n35570), .B(n35571), .Z(n32690) );
  ANDN U35376 ( .B(n35062), .A(n35572), .Z(n35570) );
  XNOR U35377 ( .A(n35573), .B(n35574), .Z(n32791) );
  NOR U35378 ( .A(n35575), .B(n35057), .Z(n35573) );
  XOR U35379 ( .A(n35576), .B(n26597), .Z(n27103) );
  XNOR U35380 ( .A(n32376), .B(n34069), .Z(n26597) );
  XNOR U35381 ( .A(n35577), .B(n34108), .Z(n34069) );
  NOR U35382 ( .A(n34490), .B(n34489), .Z(n35577) );
  XNOR U35383 ( .A(n35578), .B(n35579), .Z(n34490) );
  XOR U35384 ( .A(n33954), .B(n33513), .Z(n32376) );
  XOR U35385 ( .A(n35580), .B(n35581), .Z(n33513) );
  XOR U35386 ( .A(n30282), .B(n32241), .Z(n35581) );
  XNOR U35387 ( .A(n35582), .B(n33460), .Z(n32241) );
  XNOR U35388 ( .A(n35583), .B(n35584), .Z(n33460) );
  ANDN U35389 ( .B(n35086), .A(n34152), .Z(n35582) );
  XOR U35390 ( .A(n35585), .B(n33548), .Z(n30282) );
  XNOR U35391 ( .A(n35586), .B(n35587), .Z(n33548) );
  ANDN U35392 ( .B(n34154), .A(n35091), .Z(n35585) );
  IV U35393 ( .A(n35588), .Z(n35091) );
  XNOR U35394 ( .A(n31207), .B(n35589), .Z(n35580) );
  XOR U35395 ( .A(n34137), .B(n29049), .Z(n35589) );
  XOR U35396 ( .A(n35590), .B(n33314), .Z(n29049) );
  NOR U35397 ( .A(n35080), .B(n34146), .Z(n35590) );
  IV U35398 ( .A(n35592), .Z(n35080) );
  XNOR U35399 ( .A(n35593), .B(n33322), .Z(n34137) );
  XNOR U35400 ( .A(n35594), .B(n35595), .Z(n33322) );
  NOR U35401 ( .A(n34149), .B(n35076), .Z(n35593) );
  XNOR U35402 ( .A(n35596), .B(n34143), .Z(n31207) );
  XOR U35403 ( .A(n35597), .B(n35598), .Z(n34143) );
  ANDN U35404 ( .B(n34144), .A(n35599), .Z(n35596) );
  XOR U35405 ( .A(n35600), .B(n35601), .Z(n33954) );
  XOR U35406 ( .A(n33488), .B(n31067), .Z(n35601) );
  XOR U35407 ( .A(n35602), .B(n34100), .Z(n31067) );
  ANDN U35408 ( .B(n34071), .A(n34495), .Z(n35602) );
  IV U35409 ( .A(n34072), .Z(n34495) );
  XOR U35410 ( .A(n35605), .B(n35606), .Z(n34072) );
  XNOR U35411 ( .A(n35378), .B(n35607), .Z(n34071) );
  XNOR U35412 ( .A(n35608), .B(n34621), .Z(n33488) );
  IV U35413 ( .A(n34107), .Z(n34621) );
  XNOR U35414 ( .A(n35609), .B(n35093), .Z(n34107) );
  AND U35415 ( .A(n34108), .B(n34489), .Z(n35608) );
  XOR U35416 ( .A(n35610), .B(n35611), .Z(n34489) );
  XNOR U35417 ( .A(n35612), .B(n35613), .Z(n34108) );
  XOR U35418 ( .A(n32436), .B(n35614), .Z(n35600) );
  XNOR U35419 ( .A(n31824), .B(n32909), .Z(n35614) );
  XOR U35420 ( .A(n35615), .B(n34096), .Z(n32909) );
  XOR U35421 ( .A(n35616), .B(n35617), .Z(n34096) );
  ANDN U35422 ( .B(n34078), .A(n34076), .Z(n35615) );
  XNOR U35423 ( .A(n35618), .B(n35619), .Z(n34076) );
  XOR U35424 ( .A(n35620), .B(n35621), .Z(n34078) );
  XNOR U35425 ( .A(n35622), .B(n34093), .Z(n31824) );
  XNOR U35426 ( .A(n35583), .B(n35623), .Z(n34093) );
  ANDN U35427 ( .B(n34084), .A(n34497), .Z(n35622) );
  IV U35428 ( .A(n34085), .Z(n34497) );
  XOR U35429 ( .A(n35624), .B(n35625), .Z(n34085) );
  XNOR U35430 ( .A(n35626), .B(n35627), .Z(n34084) );
  XNOR U35431 ( .A(n35628), .B(n34103), .Z(n32436) );
  XNOR U35432 ( .A(n35629), .B(n35630), .Z(n34103) );
  ANDN U35433 ( .B(n34082), .A(n34104), .Z(n35628) );
  XOR U35434 ( .A(n35631), .B(n35632), .Z(n34104) );
  XOR U35435 ( .A(n35633), .B(n35634), .Z(n34082) );
  AND U35436 ( .A(n28372), .B(n28471), .Z(n35576) );
  XNOR U35437 ( .A(n35635), .B(n31454), .Z(n28471) );
  XNOR U35438 ( .A(n33199), .B(n32502), .Z(n31454) );
  XNOR U35439 ( .A(n35636), .B(n35637), .Z(n32502) );
  XNOR U35440 ( .A(n35638), .B(n33412), .Z(n35637) );
  XOR U35441 ( .A(n35639), .B(n35640), .Z(n33412) );
  NOR U35442 ( .A(n34197), .B(n34195), .Z(n35639) );
  XOR U35443 ( .A(n33380), .B(n35641), .Z(n35636) );
  XOR U35444 ( .A(n33945), .B(n30742), .Z(n35641) );
  XNOR U35445 ( .A(n35642), .B(n35435), .Z(n30742) );
  NOR U35446 ( .A(n34192), .B(n34191), .Z(n35642) );
  XNOR U35447 ( .A(n35643), .B(n35424), .Z(n33945) );
  ANDN U35448 ( .B(n34201), .A(n34200), .Z(n35643) );
  XNOR U35449 ( .A(n35644), .B(n35432), .Z(n33380) );
  ANDN U35450 ( .B(n34210), .A(n34208), .Z(n35644) );
  XNOR U35451 ( .A(n35645), .B(n35646), .Z(n33199) );
  XNOR U35452 ( .A(n31631), .B(n35647), .Z(n35646) );
  XNOR U35453 ( .A(n35648), .B(n33757), .Z(n31631) );
  NOR U35454 ( .A(n35649), .B(n35243), .Z(n35648) );
  XNOR U35455 ( .A(n32437), .B(n35650), .Z(n35645) );
  XNOR U35456 ( .A(n35651), .B(n35652), .Z(n35650) );
  XNOR U35457 ( .A(n35653), .B(n33761), .Z(n32437) );
  NOR U35458 ( .A(n35234), .B(n35654), .Z(n35653) );
  XOR U35459 ( .A(n35655), .B(n28796), .Z(n28372) );
  IV U35460 ( .A(n31595), .Z(n28796) );
  XOR U35461 ( .A(n35656), .B(n35657), .Z(n31595) );
  XNOR U35462 ( .A(n35658), .B(n35659), .Z(n26980) );
  XNOR U35463 ( .A(n23557), .B(n28358), .Z(n35659) );
  XNOR U35464 ( .A(n35660), .B(n30325), .Z(n28358) );
  XNOR U35465 ( .A(n35661), .B(n31772), .Z(n30325) );
  XNOR U35466 ( .A(n35662), .B(n35663), .Z(n32211) );
  XOR U35467 ( .A(n32684), .B(n33905), .Z(n35663) );
  XNOR U35468 ( .A(n35664), .B(n34580), .Z(n33905) );
  XOR U35469 ( .A(n35665), .B(n34593), .Z(n32684) );
  ANDN U35470 ( .B(n34594), .A(n35453), .Z(n35665) );
  XOR U35471 ( .A(n33091), .B(n35666), .Z(n35662) );
  XNOR U35472 ( .A(n32510), .B(n33044), .Z(n35666) );
  XNOR U35473 ( .A(n35667), .B(n34584), .Z(n33044) );
  NOR U35474 ( .A(n34585), .B(n35449), .Z(n35667) );
  XOR U35475 ( .A(n35668), .B(n34590), .Z(n32510) );
  IV U35476 ( .A(n35669), .Z(n34590) );
  ANDN U35477 ( .B(n35670), .A(n34589), .Z(n35668) );
  XNOR U35478 ( .A(n35671), .B(n34597), .Z(n33091) );
  NOR U35479 ( .A(n34598), .B(n35672), .Z(n35671) );
  XNOR U35480 ( .A(n35673), .B(n35674), .Z(n34227) );
  XNOR U35481 ( .A(n33023), .B(n35675), .Z(n35674) );
  XNOR U35482 ( .A(n35676), .B(n35677), .Z(n33023) );
  XOR U35483 ( .A(n28422), .B(n35679), .Z(n35673) );
  XNOR U35484 ( .A(n32736), .B(n33149), .Z(n35679) );
  XNOR U35485 ( .A(n35680), .B(n35681), .Z(n33149) );
  NOR U35486 ( .A(n34508), .B(n35682), .Z(n35680) );
  XNOR U35487 ( .A(n35683), .B(n35684), .Z(n32736) );
  NOR U35488 ( .A(n34521), .B(n35685), .Z(n35683) );
  XNOR U35489 ( .A(n35686), .B(n35687), .Z(n28422) );
  NOR U35490 ( .A(n35688), .B(n35689), .Z(n35686) );
  NOR U35491 ( .A(n27404), .B(n30850), .Z(n35660) );
  XOR U35492 ( .A(n28831), .B(n35690), .Z(n30850) );
  IV U35493 ( .A(n32622), .Z(n28831) );
  XOR U35494 ( .A(n35691), .B(n34160), .Z(n32622) );
  XNOR U35495 ( .A(n35692), .B(n35693), .Z(n34160) );
  XNOR U35496 ( .A(n31874), .B(n32343), .Z(n35693) );
  NOR U35497 ( .A(n33626), .B(n33625), .Z(n35694) );
  XNOR U35498 ( .A(n35695), .B(n34256), .Z(n31874) );
  NOR U35499 ( .A(n33622), .B(n33621), .Z(n35695) );
  XOR U35500 ( .A(n34134), .B(n35696), .Z(n35692) );
  XOR U35501 ( .A(n32106), .B(n28743), .Z(n35696) );
  XNOR U35502 ( .A(n35697), .B(n35698), .Z(n28743) );
  ANDN U35503 ( .B(n33988), .A(n33987), .Z(n35697) );
  XNOR U35504 ( .A(n35699), .B(n35700), .Z(n32106) );
  NOR U35505 ( .A(n34163), .B(n34162), .Z(n35699) );
  XNOR U35506 ( .A(n35701), .B(n34263), .Z(n34134) );
  NOR U35507 ( .A(n33617), .B(n33615), .Z(n35701) );
  XNOR U35508 ( .A(n31700), .B(n35702), .Z(n27404) );
  XNOR U35509 ( .A(n35703), .B(n30335), .Z(n23557) );
  XNOR U35510 ( .A(n34677), .B(n30303), .Z(n30335) );
  XNOR U35511 ( .A(n35704), .B(n34961), .Z(n34677) );
  NOR U35512 ( .A(n35705), .B(n35706), .Z(n35704) );
  NOR U35513 ( .A(n30859), .B(n30826), .Z(n35703) );
  XOR U35514 ( .A(n35707), .B(n29315), .Z(n30826) );
  IV U35515 ( .A(n32359), .Z(n29315) );
  XNOR U35516 ( .A(n35708), .B(n35709), .Z(n32359) );
  XOR U35517 ( .A(n35710), .B(n33455), .Z(n30859) );
  IV U35518 ( .A(n30528), .Z(n33455) );
  XNOR U35519 ( .A(n35711), .B(n33647), .Z(n30528) );
  XNOR U35520 ( .A(n35712), .B(n35713), .Z(n33647) );
  XOR U35521 ( .A(n35714), .B(n31782), .Z(n35713) );
  XOR U35522 ( .A(n35715), .B(n35716), .Z(n31782) );
  ANDN U35523 ( .B(n35717), .A(n35718), .Z(n35715) );
  XNOR U35524 ( .A(n32609), .B(n35719), .Z(n35712) );
  XNOR U35525 ( .A(n31833), .B(n35720), .Z(n35719) );
  XOR U35526 ( .A(n35721), .B(n35722), .Z(n31833) );
  ANDN U35527 ( .B(n35723), .A(n35724), .Z(n35721) );
  XNOR U35528 ( .A(n35725), .B(n35726), .Z(n32609) );
  XOR U35529 ( .A(n26383), .B(n35729), .Z(n35658) );
  XOR U35530 ( .A(n24980), .B(n31606), .Z(n35729) );
  XNOR U35531 ( .A(n35730), .B(n30323), .Z(n31606) );
  XNOR U35532 ( .A(n28747), .B(n35731), .Z(n30323) );
  XOR U35533 ( .A(n35732), .B(n32528), .Z(n28747) );
  XNOR U35534 ( .A(n35733), .B(n35734), .Z(n32528) );
  XOR U35535 ( .A(n33525), .B(n35735), .Z(n35734) );
  XNOR U35536 ( .A(n35736), .B(n35737), .Z(n33525) );
  ANDN U35537 ( .B(n35738), .A(n35739), .Z(n35736) );
  XOR U35538 ( .A(n32455), .B(n35740), .Z(n35733) );
  XOR U35539 ( .A(n35741), .B(n35742), .Z(n35740) );
  XNOR U35540 ( .A(n35743), .B(n35744), .Z(n32455) );
  ANDN U35541 ( .B(n35745), .A(n35746), .Z(n35743) );
  ANDN U35542 ( .B(n30867), .A(n27399), .Z(n35730) );
  XOR U35543 ( .A(n35747), .B(n30674), .Z(n27399) );
  XOR U35544 ( .A(n35748), .B(n32362), .Z(n30867) );
  XNOR U35545 ( .A(n35749), .B(n30331), .Z(n24980) );
  XNOR U35546 ( .A(n32034), .B(n35750), .Z(n30331) );
  IV U35547 ( .A(n33942), .Z(n32034) );
  XNOR U35548 ( .A(n35752), .B(n35753), .Z(n33675) );
  XOR U35549 ( .A(n32439), .B(n35754), .Z(n35753) );
  XOR U35550 ( .A(n35755), .B(n34303), .Z(n32439) );
  ANDN U35551 ( .B(n35487), .A(n35756), .Z(n35755) );
  XOR U35552 ( .A(n30958), .B(n35757), .Z(n35752) );
  XOR U35553 ( .A(n32121), .B(n31997), .Z(n35757) );
  XNOR U35554 ( .A(n35758), .B(n34309), .Z(n31997) );
  ANDN U35555 ( .B(n35759), .A(n35480), .Z(n35758) );
  XNOR U35556 ( .A(n35760), .B(n34299), .Z(n32121) );
  ANDN U35557 ( .B(n35761), .A(n35482), .Z(n35760) );
  XNOR U35558 ( .A(n35762), .B(n34316), .Z(n30958) );
  NOR U35559 ( .A(n35485), .B(n35763), .Z(n35762) );
  NOR U35560 ( .A(n27535), .B(n30854), .Z(n35749) );
  XNOR U35561 ( .A(n35764), .B(n32008), .Z(n30854) );
  XOR U35562 ( .A(n29072), .B(n35765), .Z(n27535) );
  IV U35563 ( .A(n32038), .Z(n29072) );
  XNOR U35564 ( .A(n34795), .B(n33730), .Z(n32038) );
  XNOR U35565 ( .A(n35766), .B(n35767), .Z(n33730) );
  XNOR U35566 ( .A(n29261), .B(n32547), .Z(n35767) );
  XOR U35567 ( .A(n35769), .B(n35770), .Z(n34832) );
  NOR U35568 ( .A(n34831), .B(n34643), .Z(n35768) );
  XNOR U35569 ( .A(n35771), .B(n34834), .Z(n29261) );
  XNOR U35570 ( .A(n35772), .B(n35773), .Z(n34834) );
  NOR U35571 ( .A(n35774), .B(n34647), .Z(n35771) );
  XOR U35572 ( .A(n31232), .B(n35775), .Z(n35766) );
  XOR U35573 ( .A(n33299), .B(n33953), .Z(n35775) );
  XNOR U35574 ( .A(n35776), .B(n34827), .Z(n33953) );
  XOR U35575 ( .A(n35777), .B(n35778), .Z(n34827) );
  NOR U35576 ( .A(n34656), .B(n34828), .Z(n35776) );
  XNOR U35577 ( .A(n35779), .B(n34820), .Z(n33299) );
  XNOR U35578 ( .A(n35780), .B(n35606), .Z(n34820) );
  NOR U35579 ( .A(n34652), .B(n34821), .Z(n35779) );
  XNOR U35580 ( .A(n35781), .B(n34824), .Z(n31232) );
  XNOR U35581 ( .A(n35782), .B(n35783), .Z(n34824) );
  NOR U35582 ( .A(n34660), .B(n34823), .Z(n35781) );
  XOR U35583 ( .A(n35784), .B(n35785), .Z(n34795) );
  XOR U35584 ( .A(n31703), .B(n34603), .Z(n35785) );
  XOR U35585 ( .A(n35786), .B(n35328), .Z(n34603) );
  XOR U35586 ( .A(n35787), .B(n35788), .Z(n35328) );
  ANDN U35587 ( .B(n35333), .A(n35789), .Z(n35786) );
  XNOR U35588 ( .A(n35790), .B(n34851), .Z(n31703) );
  XNOR U35589 ( .A(n35791), .B(n35792), .Z(n34851) );
  ANDN U35590 ( .B(n34852), .A(n33978), .Z(n35790) );
  XOR U35591 ( .A(n31815), .B(n35793), .Z(n35784) );
  XOR U35592 ( .A(n30543), .B(n34816), .Z(n35793) );
  XNOR U35593 ( .A(n35794), .B(n35317), .Z(n34816) );
  XOR U35594 ( .A(n35795), .B(n35796), .Z(n35317) );
  NOR U35595 ( .A(n33974), .B(n34849), .Z(n35794) );
  XOR U35596 ( .A(n35797), .B(n34841), .Z(n30543) );
  XNOR U35597 ( .A(n35798), .B(n35799), .Z(n34841) );
  NOR U35598 ( .A(n33969), .B(n34840), .Z(n35797) );
  XOR U35599 ( .A(n35800), .B(n34844), .Z(n31815) );
  XNOR U35600 ( .A(n35510), .B(n35801), .Z(n34844) );
  ANDN U35601 ( .B(n34845), .A(n33982), .Z(n35800) );
  XNOR U35602 ( .A(n35802), .B(n30329), .Z(n26383) );
  XNOR U35603 ( .A(n31669), .B(n35803), .Z(n30329) );
  IV U35604 ( .A(n32365), .Z(n31669) );
  XNOR U35605 ( .A(n32841), .B(n33421), .Z(n32365) );
  XNOR U35606 ( .A(n35804), .B(n35805), .Z(n33421) );
  XNOR U35607 ( .A(n35806), .B(n28735), .Z(n35805) );
  XNOR U35608 ( .A(n35807), .B(n35808), .Z(n28735) );
  NOR U35609 ( .A(n35809), .B(n35549), .Z(n35807) );
  XNOR U35610 ( .A(n30496), .B(n35810), .Z(n35804) );
  XOR U35611 ( .A(n33947), .B(n31345), .Z(n35810) );
  XOR U35612 ( .A(n35811), .B(n35812), .Z(n31345) );
  NOR U35613 ( .A(n35544), .B(n35813), .Z(n35811) );
  IV U35614 ( .A(n35814), .Z(n35544) );
  XNOR U35615 ( .A(n35815), .B(n35816), .Z(n33947) );
  NOR U35616 ( .A(n35817), .B(n35557), .Z(n35815) );
  XNOR U35617 ( .A(n35818), .B(n35819), .Z(n30496) );
  NOR U35618 ( .A(n35820), .B(n35821), .Z(n35818) );
  XOR U35619 ( .A(n35822), .B(n35823), .Z(n32841) );
  XNOR U35620 ( .A(n33475), .B(n32827), .Z(n35823) );
  XNOR U35621 ( .A(n35824), .B(n35825), .Z(n32827) );
  ANDN U35622 ( .B(n35826), .A(n35827), .Z(n35824) );
  XNOR U35623 ( .A(n35828), .B(n35829), .Z(n33475) );
  NOR U35624 ( .A(n35830), .B(n35831), .Z(n35828) );
  XOR U35625 ( .A(n32063), .B(n35832), .Z(n35822) );
  XNOR U35626 ( .A(n32886), .B(n33054), .Z(n35832) );
  XNOR U35627 ( .A(n35833), .B(n35834), .Z(n33054) );
  ANDN U35628 ( .B(n35835), .A(n35836), .Z(n35833) );
  XOR U35629 ( .A(n35837), .B(n35838), .Z(n32886) );
  NOR U35630 ( .A(n35839), .B(n35840), .Z(n35837) );
  XNOR U35631 ( .A(n35841), .B(n35842), .Z(n32063) );
  NOR U35632 ( .A(n35843), .B(n35844), .Z(n35841) );
  NOR U35633 ( .A(n27393), .B(n30863), .Z(n35802) );
  XNOR U35634 ( .A(n33265), .B(n35845), .Z(n30863) );
  XOR U35635 ( .A(n33551), .B(n35846), .Z(n27393) );
  IV U35636 ( .A(n30911), .Z(n33551) );
  XOR U35637 ( .A(n32087), .B(n35847), .Z(n30911) );
  XOR U35638 ( .A(n35848), .B(n35849), .Z(n32087) );
  XOR U35639 ( .A(n33484), .B(n32997), .Z(n35849) );
  XNOR U35640 ( .A(n35850), .B(n35851), .Z(n32997) );
  ANDN U35641 ( .B(n35852), .A(n35853), .Z(n35850) );
  XNOR U35642 ( .A(n35854), .B(n34031), .Z(n33484) );
  ANDN U35643 ( .B(n35855), .A(n35856), .Z(n35854) );
  XNOR U35644 ( .A(n32497), .B(n35857), .Z(n35848) );
  XNOR U35645 ( .A(n29532), .B(n35858), .Z(n35857) );
  XOR U35646 ( .A(n35859), .B(n35860), .Z(n29532) );
  NOR U35647 ( .A(n35861), .B(n35862), .Z(n35859) );
  XOR U35648 ( .A(n35863), .B(n34039), .Z(n32497) );
  NOR U35649 ( .A(n35864), .B(n35865), .Z(n35863) );
  XOR U35650 ( .A(n35866), .B(n20797), .Z(n17582) );
  XNOR U35651 ( .A(n27862), .B(n24835), .Z(n20797) );
  XNOR U35652 ( .A(n26271), .B(n28779), .Z(n24835) );
  XNOR U35653 ( .A(n35867), .B(n35868), .Z(n28779) );
  XOR U35654 ( .A(n27725), .B(n26508), .Z(n35868) );
  XNOR U35655 ( .A(n35869), .B(n27762), .Z(n26508) );
  XOR U35656 ( .A(n35870), .B(n32006), .Z(n27762) );
  XOR U35657 ( .A(n33453), .B(n35871), .Z(n32006) );
  XOR U35658 ( .A(n35872), .B(n35873), .Z(n33453) );
  XNOR U35659 ( .A(n35874), .B(n32600), .Z(n35873) );
  XNOR U35660 ( .A(n35875), .B(n35876), .Z(n32600) );
  AND U35661 ( .A(n35877), .B(n35878), .Z(n35875) );
  XOR U35662 ( .A(n33092), .B(n35879), .Z(n35872) );
  XOR U35663 ( .A(n35880), .B(n32309), .Z(n35879) );
  XNOR U35664 ( .A(n35881), .B(n35882), .Z(n32309) );
  ANDN U35665 ( .B(n35883), .A(n35884), .Z(n35881) );
  XNOR U35666 ( .A(n35885), .B(n35886), .Z(n33092) );
  AND U35667 ( .A(n35887), .B(n35888), .Z(n35885) );
  AND U35668 ( .A(n27763), .B(n35889), .Z(n35869) );
  XOR U35669 ( .A(n35890), .B(n30192), .Z(n27725) );
  XOR U35670 ( .A(n28807), .B(n35891), .Z(n30192) );
  AND U35671 ( .A(n27857), .B(n27855), .Z(n35890) );
  XOR U35672 ( .A(n31840), .B(n35892), .Z(n27855) );
  XOR U35673 ( .A(n35708), .B(n35893), .Z(n31840) );
  XOR U35674 ( .A(n35894), .B(n35895), .Z(n35708) );
  XNOR U35675 ( .A(n32234), .B(n28876), .Z(n35895) );
  XOR U35676 ( .A(n35896), .B(n35897), .Z(n28876) );
  AND U35677 ( .A(n35898), .B(n35899), .Z(n35896) );
  XOR U35678 ( .A(n35900), .B(n35901), .Z(n32234) );
  AND U35679 ( .A(n35902), .B(n35903), .Z(n35900) );
  XOR U35680 ( .A(n28758), .B(n35904), .Z(n35894) );
  XOR U35681 ( .A(n35905), .B(n33699), .Z(n35904) );
  XOR U35682 ( .A(n35906), .B(n35907), .Z(n33699) );
  XNOR U35683 ( .A(n35910), .B(n35911), .Z(n28758) );
  XNOR U35684 ( .A(n25007), .B(n35914), .Z(n35867) );
  XNOR U35685 ( .A(n27738), .B(n26550), .Z(n35914) );
  XOR U35686 ( .A(n35915), .B(n31419), .Z(n26550) );
  IV U35687 ( .A(n27768), .Z(n31419) );
  XOR U35688 ( .A(n35647), .B(n35916), .Z(n27768) );
  XOR U35689 ( .A(n35917), .B(n33764), .Z(n35647) );
  ANDN U35690 ( .B(n35918), .A(n35240), .Z(n35917) );
  NOR U35691 ( .A(n27868), .B(n27767), .Z(n35915) );
  XOR U35692 ( .A(n35919), .B(n30928), .Z(n27767) );
  XOR U35693 ( .A(n35920), .B(n35921), .Z(n30928) );
  XOR U35694 ( .A(n35922), .B(n27771), .Z(n27738) );
  XOR U35695 ( .A(n35534), .B(n32395), .Z(n27771) );
  IV U35696 ( .A(n31440), .Z(n32395) );
  XNOR U35697 ( .A(n35923), .B(n35924), .Z(n34138) );
  XNOR U35698 ( .A(n33420), .B(n32807), .Z(n35924) );
  XNOR U35699 ( .A(n35925), .B(n33436), .Z(n32807) );
  XNOR U35700 ( .A(n35926), .B(n35927), .Z(n33436) );
  XOR U35701 ( .A(n35928), .B(n35929), .Z(n33437) );
  XNOR U35702 ( .A(n35930), .B(n34173), .Z(n33420) );
  XOR U35703 ( .A(n35931), .B(n35932), .Z(n34173) );
  ANDN U35704 ( .B(n34174), .A(n35531), .Z(n35930) );
  XOR U35705 ( .A(n35933), .B(n35934), .Z(n34174) );
  XOR U35706 ( .A(n32646), .B(n35935), .Z(n35923) );
  XNOR U35707 ( .A(n32110), .B(n32507), .Z(n35935) );
  XNOR U35708 ( .A(n35936), .B(n33430), .Z(n32507) );
  XNOR U35709 ( .A(n35937), .B(n35938), .Z(n33430) );
  AND U35710 ( .A(n33431), .B(n35539), .Z(n35936) );
  XOR U35711 ( .A(n35939), .B(n35940), .Z(n33431) );
  XNOR U35712 ( .A(n35941), .B(n33426), .Z(n32110) );
  IV U35713 ( .A(n35104), .Z(n33426) );
  ANDN U35714 ( .B(n33427), .A(n35533), .Z(n35941) );
  XNOR U35715 ( .A(n35944), .B(n35945), .Z(n33427) );
  XOR U35716 ( .A(n35946), .B(n33441), .Z(n32646) );
  ANDN U35717 ( .B(n35947), .A(n33440), .Z(n35946) );
  IV U35718 ( .A(n35948), .Z(n33440) );
  XNOR U35719 ( .A(n35950), .B(n35948), .Z(n35534) );
  XOR U35720 ( .A(n35951), .B(n35952), .Z(n35948) );
  NOR U35721 ( .A(n35953), .B(n35947), .Z(n35950) );
  XOR U35722 ( .A(n35954), .B(n30583), .Z(n27772) );
  XOR U35723 ( .A(n35955), .B(n27775), .Z(n25007) );
  XOR U35724 ( .A(n32747), .B(n35956), .Z(n27775) );
  XOR U35725 ( .A(n32419), .B(n35957), .Z(n32747) );
  XOR U35726 ( .A(n35958), .B(n35959), .Z(n32419) );
  XNOR U35727 ( .A(n29400), .B(n30550), .Z(n35959) );
  XNOR U35728 ( .A(n35960), .B(n35216), .Z(n30550) );
  NOR U35729 ( .A(n35961), .B(n35215), .Z(n35960) );
  XOR U35730 ( .A(n35962), .B(n35963), .Z(n29400) );
  ANDN U35731 ( .B(n33106), .A(n35964), .Z(n35962) );
  XNOR U35732 ( .A(n32543), .B(n35965), .Z(n35958) );
  XOR U35733 ( .A(n30111), .B(n31041), .Z(n35965) );
  XOR U35734 ( .A(n35966), .B(n33112), .Z(n31041) );
  NOR U35735 ( .A(n33111), .B(n35967), .Z(n35966) );
  XOR U35736 ( .A(n35968), .B(n33116), .Z(n30111) );
  NOR U35737 ( .A(n35969), .B(n33115), .Z(n35968) );
  XNOR U35738 ( .A(n35970), .B(n35971), .Z(n32543) );
  ANDN U35739 ( .B(n35972), .A(n35973), .Z(n35970) );
  ANDN U35740 ( .B(n27860), .A(n27859), .Z(n35955) );
  IV U35741 ( .A(n27776), .Z(n27859) );
  XOR U35742 ( .A(n34120), .B(n30165), .Z(n27776) );
  IV U35743 ( .A(n33303), .Z(n30165) );
  XNOR U35744 ( .A(n35974), .B(n35975), .Z(n32961) );
  XNOR U35745 ( .A(n35976), .B(n32301), .Z(n35975) );
  XOR U35746 ( .A(n35977), .B(n34554), .Z(n32301) );
  NOR U35747 ( .A(n34902), .B(n34901), .Z(n35977) );
  XOR U35748 ( .A(n31567), .B(n35978), .Z(n35974) );
  XOR U35749 ( .A(n32212), .B(n34186), .Z(n35978) );
  XNOR U35750 ( .A(n35979), .B(n34550), .Z(n34186) );
  NOR U35751 ( .A(n34130), .B(n34129), .Z(n35979) );
  XNOR U35752 ( .A(n35980), .B(n34558), .Z(n32212) );
  NOR U35753 ( .A(n35981), .B(n35982), .Z(n35980) );
  XNOR U35754 ( .A(n35983), .B(n34542), .Z(n31567) );
  NOR U35755 ( .A(n34123), .B(n34122), .Z(n35983) );
  XOR U35756 ( .A(n35984), .B(n35985), .Z(n34575) );
  XOR U35757 ( .A(n31780), .B(n30513), .Z(n35985) );
  XNOR U35758 ( .A(n35986), .B(n35987), .Z(n30513) );
  ANDN U35759 ( .B(n32880), .A(n32878), .Z(n35986) );
  XNOR U35760 ( .A(n35988), .B(n35467), .Z(n31780) );
  AND U35761 ( .A(n32466), .B(n32468), .Z(n35988) );
  XOR U35762 ( .A(n32277), .B(n35989), .Z(n35984) );
  XOR U35763 ( .A(n35990), .B(n31317), .Z(n35989) );
  XNOR U35764 ( .A(n35991), .B(n35458), .Z(n31317) );
  AND U35765 ( .A(n32472), .B(n32474), .Z(n35991) );
  XNOR U35766 ( .A(n35992), .B(n35461), .Z(n32277) );
  AND U35767 ( .A(n32477), .B(n32476), .Z(n35992) );
  XOR U35768 ( .A(n35993), .B(n35994), .Z(n34120) );
  ANDN U35769 ( .B(n35982), .A(n34556), .Z(n35993) );
  XOR U35770 ( .A(n35995), .B(n35996), .Z(n26271) );
  XOR U35771 ( .A(n25509), .B(n25592), .Z(n35996) );
  XOR U35772 ( .A(n35997), .B(n27750), .Z(n25592) );
  XOR U35773 ( .A(n35998), .B(n31542), .Z(n27750) );
  AND U35774 ( .A(n26435), .B(n26433), .Z(n35997) );
  XNOR U35775 ( .A(n30674), .B(n35999), .Z(n26433) );
  IV U35776 ( .A(n27657), .Z(n30674) );
  XNOR U35777 ( .A(n36000), .B(n32893), .Z(n27657) );
  XNOR U35778 ( .A(n36001), .B(n36002), .Z(n32893) );
  XNOR U35779 ( .A(n32913), .B(n32557), .Z(n36002) );
  XNOR U35780 ( .A(n36003), .B(n35827), .Z(n32557) );
  ANDN U35781 ( .B(n36004), .A(n36005), .Z(n36003) );
  XNOR U35782 ( .A(n36006), .B(n35839), .Z(n32913) );
  ANDN U35783 ( .B(n36007), .A(n36008), .Z(n36006) );
  XOR U35784 ( .A(n32263), .B(n36009), .Z(n36001) );
  XOR U35785 ( .A(n31653), .B(n32552), .Z(n36009) );
  XNOR U35786 ( .A(n36010), .B(n35831), .Z(n32552) );
  NOR U35787 ( .A(n36011), .B(n36012), .Z(n36010) );
  XNOR U35788 ( .A(n36013), .B(n35844), .Z(n31653) );
  NOR U35789 ( .A(n36014), .B(n36015), .Z(n36013) );
  XNOR U35790 ( .A(n36016), .B(n35836), .Z(n32263) );
  ANDN U35791 ( .B(n36017), .A(n36018), .Z(n36016) );
  XNOR U35792 ( .A(n36019), .B(n36020), .Z(n35675) );
  XNOR U35793 ( .A(n33906), .B(n36022), .Z(n28421) );
  XOR U35794 ( .A(n36023), .B(n36024), .Z(n33906) );
  XNOR U35795 ( .A(n36025), .B(n36026), .Z(n36024) );
  XNOR U35796 ( .A(n32704), .B(n36027), .Z(n36023) );
  XNOR U35797 ( .A(n30855), .B(n33769), .Z(n36027) );
  XNOR U35798 ( .A(n36028), .B(n34523), .Z(n33769) );
  IV U35799 ( .A(n36029), .Z(n34523) );
  AND U35800 ( .A(n35685), .B(n35684), .Z(n36028) );
  XOR U35801 ( .A(n36030), .B(n36031), .Z(n30855) );
  AND U35802 ( .A(n35682), .B(n35681), .Z(n36030) );
  XOR U35803 ( .A(n36032), .B(n34519), .Z(n32704) );
  ANDN U35804 ( .B(n35677), .A(n35678), .Z(n36032) );
  XNOR U35805 ( .A(n36033), .B(n30189), .Z(n25509) );
  XOR U35806 ( .A(n33806), .B(n28769), .Z(n30189) );
  XNOR U35807 ( .A(n36034), .B(n33290), .Z(n33806) );
  ANDN U35808 ( .B(n26428), .A(n26429), .Z(n36033) );
  XNOR U35809 ( .A(n36037), .B(n31467), .Z(n26429) );
  XOR U35810 ( .A(n31659), .B(n36038), .Z(n26428) );
  XOR U35811 ( .A(n26244), .B(n36039), .Z(n35995) );
  XOR U35812 ( .A(n26197), .B(n25381), .Z(n36039) );
  XOR U35813 ( .A(n36040), .B(n27743), .Z(n25381) );
  XOR U35814 ( .A(n33216), .B(n33226), .Z(n27743) );
  XNOR U35815 ( .A(n36041), .B(n36042), .Z(n33216) );
  NOR U35816 ( .A(n36043), .B(n36044), .Z(n36041) );
  ANDN U35817 ( .B(n26437), .A(n26438), .Z(n36040) );
  XOR U35818 ( .A(n36045), .B(n31223), .Z(n26438) );
  IV U35819 ( .A(n33068), .Z(n31223) );
  XNOR U35820 ( .A(n34428), .B(n33999), .Z(n33068) );
  XNOR U35821 ( .A(n36046), .B(n36047), .Z(n33999) );
  XNOR U35822 ( .A(n33712), .B(n32089), .Z(n36047) );
  XNOR U35823 ( .A(n36048), .B(n36049), .Z(n32089) );
  NOR U35824 ( .A(n36050), .B(n36051), .Z(n36048) );
  XNOR U35825 ( .A(n36052), .B(n36053), .Z(n33712) );
  NOR U35826 ( .A(n36054), .B(n36055), .Z(n36052) );
  XOR U35827 ( .A(n31576), .B(n36056), .Z(n36046) );
  XOR U35828 ( .A(n31990), .B(n31406), .Z(n36056) );
  XNOR U35829 ( .A(n36057), .B(n36058), .Z(n31406) );
  ANDN U35830 ( .B(n36059), .A(n36060), .Z(n36057) );
  XNOR U35831 ( .A(n36061), .B(n36062), .Z(n31990) );
  ANDN U35832 ( .B(n36063), .A(n36064), .Z(n36061) );
  XOR U35833 ( .A(n36065), .B(n36066), .Z(n31576) );
  ANDN U35834 ( .B(n36067), .A(n36068), .Z(n36065) );
  XOR U35835 ( .A(n36069), .B(n36070), .Z(n34428) );
  XNOR U35836 ( .A(n36037), .B(n32981), .Z(n36070) );
  XNOR U35837 ( .A(n36071), .B(n36072), .Z(n32981) );
  ANDN U35838 ( .B(n36073), .A(n36074), .Z(n36071) );
  XNOR U35839 ( .A(n36075), .B(n36076), .Z(n36037) );
  ANDN U35840 ( .B(n36077), .A(n36078), .Z(n36075) );
  XNOR U35841 ( .A(n31466), .B(n36079), .Z(n36069) );
  XOR U35842 ( .A(n36080), .B(n32996), .Z(n36079) );
  XOR U35843 ( .A(n36081), .B(n36082), .Z(n32996) );
  ANDN U35844 ( .B(n36083), .A(n36084), .Z(n36081) );
  XOR U35845 ( .A(n36085), .B(n36086), .Z(n31466) );
  ANDN U35846 ( .B(n36087), .A(n36088), .Z(n36085) );
  XNOR U35847 ( .A(n32571), .B(n34759), .Z(n26437) );
  XOR U35848 ( .A(n36089), .B(n36090), .Z(n34759) );
  ANDN U35849 ( .B(n36091), .A(n36092), .Z(n36089) );
  XNOR U35850 ( .A(n36093), .B(n36094), .Z(n35732) );
  XNOR U35851 ( .A(n31956), .B(n32016), .Z(n36094) );
  XNOR U35852 ( .A(n36095), .B(n36096), .Z(n32016) );
  NOR U35853 ( .A(n36097), .B(n36098), .Z(n36095) );
  XNOR U35854 ( .A(n36099), .B(n36100), .Z(n31956) );
  XNOR U35855 ( .A(n33472), .B(n36103), .Z(n36093) );
  XOR U35856 ( .A(n33668), .B(n31006), .Z(n36103) );
  XNOR U35857 ( .A(n36104), .B(n36105), .Z(n31006) );
  ANDN U35858 ( .B(n36106), .A(n36107), .Z(n36104) );
  XNOR U35859 ( .A(n36108), .B(n36109), .Z(n33668) );
  ANDN U35860 ( .B(n36110), .A(n36111), .Z(n36108) );
  XOR U35861 ( .A(n36112), .B(n36113), .Z(n33472) );
  ANDN U35862 ( .B(n36114), .A(n36115), .Z(n36112) );
  XOR U35863 ( .A(n36117), .B(n30187), .Z(n26197) );
  IV U35864 ( .A(n27753), .Z(n30187) );
  XOR U35865 ( .A(n34967), .B(n31219), .Z(n27753) );
  IV U35866 ( .A(n30524), .Z(n31219) );
  XNOR U35867 ( .A(n36118), .B(n36119), .Z(n34666) );
  XOR U35868 ( .A(n32314), .B(n33541), .Z(n36119) );
  ANDN U35869 ( .B(n34964), .A(n34965), .Z(n36120) );
  XNOR U35870 ( .A(n36121), .B(n34676), .Z(n32314) );
  XOR U35871 ( .A(n32971), .B(n36122), .Z(n36118) );
  XOR U35872 ( .A(n32398), .B(n36123), .Z(n36122) );
  XNOR U35873 ( .A(n36124), .B(n34686), .Z(n32398) );
  ANDN U35874 ( .B(n36125), .A(n36126), .Z(n36124) );
  XNOR U35875 ( .A(n36127), .B(n35706), .Z(n32971) );
  ANDN U35876 ( .B(n34962), .A(n34960), .Z(n36127) );
  XOR U35877 ( .A(n36128), .B(n36129), .Z(n35893) );
  XNOR U35878 ( .A(n32434), .B(n29712), .Z(n36129) );
  XNOR U35879 ( .A(n36130), .B(n36131), .Z(n29712) );
  NOR U35880 ( .A(n36132), .B(n36133), .Z(n36130) );
  XNOR U35881 ( .A(n36134), .B(n36135), .Z(n32434) );
  ANDN U35882 ( .B(n36136), .A(n36137), .Z(n36134) );
  XNOR U35883 ( .A(n36138), .B(n36139), .Z(n36128) );
  XOR U35884 ( .A(n33235), .B(n31673), .Z(n36139) );
  XNOR U35885 ( .A(n36140), .B(n36141), .Z(n31673) );
  ANDN U35886 ( .B(n36142), .A(n36143), .Z(n36140) );
  XOR U35887 ( .A(n36144), .B(n36145), .Z(n33235) );
  ANDN U35888 ( .B(n36146), .A(n36147), .Z(n36144) );
  XOR U35889 ( .A(n36148), .B(n36125), .Z(n34967) );
  ANDN U35890 ( .B(n36126), .A(n34684), .Z(n36148) );
  ANDN U35891 ( .B(n26441), .A(n26442), .Z(n36117) );
  XOR U35892 ( .A(n35564), .B(n32691), .Z(n26442) );
  XNOR U35893 ( .A(n36149), .B(n36150), .Z(n35564) );
  ANDN U35894 ( .B(n35070), .A(n36151), .Z(n36149) );
  XOR U35895 ( .A(n36152), .B(n29927), .Z(n26441) );
  XNOR U35896 ( .A(n36153), .B(n27756), .Z(n26244) );
  XNOR U35897 ( .A(n27661), .B(n36154), .Z(n27756) );
  IV U35898 ( .A(n32008), .Z(n27661) );
  XNOR U35899 ( .A(n33777), .B(n36155), .Z(n32008) );
  XOR U35900 ( .A(n36156), .B(n36157), .Z(n33777) );
  XOR U35901 ( .A(n32208), .B(n31184), .Z(n36157) );
  XOR U35902 ( .A(n36158), .B(n34291), .Z(n31184) );
  NOR U35903 ( .A(n36159), .B(n36160), .Z(n36158) );
  XOR U35904 ( .A(n36161), .B(n36162), .Z(n32208) );
  NOR U35905 ( .A(n36163), .B(n36164), .Z(n36161) );
  XOR U35906 ( .A(n34271), .B(n36165), .Z(n36156) );
  XNOR U35907 ( .A(n32294), .B(n30222), .Z(n36165) );
  XOR U35908 ( .A(n36166), .B(n34284), .Z(n30222) );
  NOR U35909 ( .A(n34283), .B(n36167), .Z(n36166) );
  XNOR U35910 ( .A(n36168), .B(n34279), .Z(n32294) );
  NOR U35911 ( .A(n34278), .B(n36169), .Z(n36168) );
  XNOR U35912 ( .A(n36170), .B(n34287), .Z(n34271) );
  NOR U35913 ( .A(n34288), .B(n36171), .Z(n36170) );
  AND U35914 ( .A(n26424), .B(n26425), .Z(n36153) );
  XNOR U35915 ( .A(n31618), .B(n36172), .Z(n26425) );
  XOR U35916 ( .A(n36173), .B(n36174), .Z(n31618) );
  XNOR U35917 ( .A(n36175), .B(n31471), .Z(n26424) );
  IV U35918 ( .A(n32191), .Z(n31471) );
  XNOR U35919 ( .A(n36176), .B(n27763), .Z(n27862) );
  XNOR U35920 ( .A(n36177), .B(n31579), .Z(n27763) );
  NOR U35921 ( .A(n36178), .B(n35889), .Z(n36176) );
  XOR U35922 ( .A(n28199), .B(n22943), .Z(n23238) );
  XNOR U35923 ( .A(n26511), .B(n27362), .Z(n22943) );
  XNOR U35924 ( .A(n36179), .B(n36180), .Z(n27362) );
  XOR U35925 ( .A(n25539), .B(n24574), .Z(n36180) );
  XNOR U35926 ( .A(n36181), .B(n27603), .Z(n24574) );
  XNOR U35927 ( .A(n36182), .B(n31178), .Z(n27603) );
  XNOR U35928 ( .A(n36183), .B(n32914), .Z(n31178) );
  XOR U35929 ( .A(n36184), .B(n36185), .Z(n32914) );
  XNOR U35930 ( .A(n36186), .B(n33827), .Z(n36185) );
  XNOR U35931 ( .A(n36187), .B(n33574), .Z(n33827) );
  XNOR U35932 ( .A(n36190), .B(n36191), .Z(n36184) );
  XOR U35933 ( .A(n32410), .B(n33908), .Z(n36191) );
  XNOR U35934 ( .A(n36192), .B(n33569), .Z(n33908) );
  NOR U35935 ( .A(n36193), .B(n36194), .Z(n36192) );
  XNOR U35936 ( .A(n36195), .B(n33582), .Z(n32410) );
  ANDN U35937 ( .B(n36196), .A(n36197), .Z(n36195) );
  XOR U35938 ( .A(n33659), .B(n31676), .Z(n27604) );
  IV U35939 ( .A(n27949), .Z(n31676) );
  XNOR U35940 ( .A(n36198), .B(n36199), .Z(n35289) );
  XOR U35941 ( .A(n32251), .B(n32345), .Z(n36199) );
  XNOR U35942 ( .A(n36200), .B(n34899), .Z(n32345) );
  ANDN U35943 ( .B(n33651), .A(n33653), .Z(n36200) );
  XOR U35944 ( .A(n36201), .B(n36202), .Z(n33651) );
  XOR U35945 ( .A(n36203), .B(n34885), .Z(n32251) );
  AND U35946 ( .A(n34886), .B(n36204), .Z(n36203) );
  XNOR U35947 ( .A(n33037), .B(n36205), .Z(n36198) );
  XNOR U35948 ( .A(n31845), .B(n34879), .Z(n36205) );
  XOR U35949 ( .A(n36206), .B(n34893), .Z(n34879) );
  ANDN U35950 ( .B(n33655), .A(n33656), .Z(n36206) );
  IV U35951 ( .A(n36207), .Z(n33656) );
  XNOR U35952 ( .A(n36208), .B(n36209), .Z(n33655) );
  XOR U35953 ( .A(n36210), .B(n34896), .Z(n31845) );
  ANDN U35954 ( .B(n33661), .A(n33663), .Z(n36210) );
  XOR U35955 ( .A(n36213), .B(n34889), .Z(n33037) );
  AND U35956 ( .A(n33665), .B(n33667), .Z(n36213) );
  XOR U35957 ( .A(n36214), .B(n36215), .Z(n33665) );
  XNOR U35958 ( .A(n36217), .B(n34886), .Z(n33659) );
  XOR U35959 ( .A(n36218), .B(n36219), .Z(n34886) );
  NOR U35960 ( .A(n36220), .B(n36204), .Z(n36217) );
  XNOR U35961 ( .A(n36221), .B(n27607), .Z(n25539) );
  XOR U35962 ( .A(n35905), .B(n32235), .Z(n27607) );
  XOR U35963 ( .A(n36222), .B(n34113), .Z(n32235) );
  XNOR U35964 ( .A(n36223), .B(n36224), .Z(n34113) );
  XOR U35965 ( .A(n31141), .B(n31291), .Z(n36224) );
  XNOR U35966 ( .A(n36225), .B(n33796), .Z(n31291) );
  IV U35967 ( .A(n36226), .Z(n33796) );
  ANDN U35968 ( .B(n33797), .A(n33397), .Z(n36225) );
  XNOR U35969 ( .A(n36227), .B(n33785), .Z(n31141) );
  ANDN U35970 ( .B(n33786), .A(n33391), .Z(n36227) );
  XNOR U35971 ( .A(n31242), .B(n36228), .Z(n36223) );
  XNOR U35972 ( .A(n33776), .B(n30530), .Z(n36228) );
  XNOR U35973 ( .A(n36229), .B(n33794), .Z(n30530) );
  ANDN U35974 ( .B(n33793), .A(n35356), .Z(n36229) );
  XOR U35975 ( .A(n36230), .B(n36231), .Z(n33776) );
  ANDN U35976 ( .B(n33783), .A(n36232), .Z(n36230) );
  XNOR U35977 ( .A(n36233), .B(n33790), .Z(n31242) );
  ANDN U35978 ( .B(n33789), .A(n33401), .Z(n36233) );
  XNOR U35979 ( .A(n36234), .B(n36235), .Z(n35905) );
  ANDN U35980 ( .B(n36236), .A(n36237), .Z(n36234) );
  AND U35981 ( .A(n36238), .B(n27608), .Z(n36221) );
  XNOR U35982 ( .A(n25997), .B(n36239), .Z(n36179) );
  XOR U35983 ( .A(n24389), .B(n21600), .Z(n36239) );
  XOR U35984 ( .A(n36240), .B(n27595), .Z(n21600) );
  XOR U35985 ( .A(n36241), .B(n32191), .Z(n27595) );
  ANDN U35986 ( .B(n28203), .A(n28201), .Z(n36240) );
  IV U35987 ( .A(n27594), .Z(n28201) );
  XOR U35988 ( .A(n36242), .B(n32644), .Z(n27594) );
  IV U35989 ( .A(n31872), .Z(n32644) );
  XOR U35990 ( .A(n33735), .B(n36243), .Z(n31872) );
  XOR U35991 ( .A(n36244), .B(n36245), .Z(n33735) );
  XOR U35992 ( .A(n31925), .B(n28801), .Z(n36245) );
  XNOR U35993 ( .A(n36246), .B(n36247), .Z(n28801) );
  ANDN U35994 ( .B(n36248), .A(n36249), .Z(n36246) );
  XNOR U35995 ( .A(n36250), .B(n36251), .Z(n31925) );
  NOR U35996 ( .A(n36252), .B(n36253), .Z(n36250) );
  XNOR U35997 ( .A(n35248), .B(n36254), .Z(n36244) );
  XOR U35998 ( .A(n31074), .B(n31662), .Z(n36254) );
  XNOR U35999 ( .A(n36255), .B(n36256), .Z(n31662) );
  NOR U36000 ( .A(n36257), .B(n36258), .Z(n36255) );
  XNOR U36001 ( .A(n36259), .B(n36260), .Z(n31074) );
  NOR U36002 ( .A(n36261), .B(n36262), .Z(n36259) );
  XNOR U36003 ( .A(n36263), .B(n36264), .Z(n35248) );
  ANDN U36004 ( .B(n36265), .A(n36266), .Z(n36263) );
  XNOR U36005 ( .A(n36267), .B(n27600), .Z(n24389) );
  XOR U36006 ( .A(n34230), .B(n31340), .Z(n27600) );
  XOR U36007 ( .A(n36022), .B(n36268), .Z(n31340) );
  XOR U36008 ( .A(n36269), .B(n36270), .Z(n36022) );
  XNOR U36009 ( .A(n33061), .B(n32800), .Z(n36270) );
  XNOR U36010 ( .A(n36271), .B(n36272), .Z(n32800) );
  XNOR U36011 ( .A(n36273), .B(n36274), .Z(n33061) );
  ANDN U36012 ( .B(n34237), .A(n34239), .Z(n36273) );
  XOR U36013 ( .A(n31597), .B(n36275), .Z(n36269) );
  XOR U36014 ( .A(n32454), .B(n32237), .Z(n36275) );
  XNOR U36015 ( .A(n36276), .B(n36277), .Z(n32237) );
  NOR U36016 ( .A(n34242), .B(n34241), .Z(n36276) );
  XOR U36017 ( .A(n36278), .B(n36279), .Z(n32454) );
  AND U36018 ( .A(n34232), .B(n34234), .Z(n36278) );
  XNOR U36019 ( .A(n36280), .B(n36281), .Z(n31597) );
  ANDN U36020 ( .B(n36282), .A(n36283), .Z(n36280) );
  XNOR U36021 ( .A(n36284), .B(n36282), .Z(n34230) );
  XNOR U36022 ( .A(n31622), .B(n34053), .Z(n27599) );
  XNOR U36023 ( .A(n36286), .B(n36287), .Z(n34053) );
  AND U36024 ( .A(n36288), .B(n35121), .Z(n36286) );
  IV U36025 ( .A(n31337), .Z(n31622) );
  XNOR U36026 ( .A(n33198), .B(n34978), .Z(n31337) );
  XNOR U36027 ( .A(n36289), .B(n36290), .Z(n34978) );
  XNOR U36028 ( .A(n29052), .B(n29023), .Z(n36290) );
  XNOR U36029 ( .A(n36291), .B(n36292), .Z(n29023) );
  NOR U36030 ( .A(n34047), .B(n34046), .Z(n36291) );
  XOR U36031 ( .A(n36293), .B(n35122), .Z(n29052) );
  NOR U36032 ( .A(n36288), .B(n36287), .Z(n36293) );
  XOR U36033 ( .A(n35334), .B(n36294), .Z(n36289) );
  XNOR U36034 ( .A(n32872), .B(n31157), .Z(n36294) );
  XNOR U36035 ( .A(n36295), .B(n36296), .Z(n31157) );
  ANDN U36036 ( .B(n34060), .A(n34061), .Z(n36295) );
  XOR U36037 ( .A(n36297), .B(n35125), .Z(n32872) );
  ANDN U36038 ( .B(n34052), .A(n34050), .Z(n36297) );
  XOR U36039 ( .A(n36298), .B(n35116), .Z(n35334) );
  NOR U36040 ( .A(n36299), .B(n34056), .Z(n36298) );
  XOR U36041 ( .A(n36300), .B(n36301), .Z(n33198) );
  XNOR U36042 ( .A(n30380), .B(n28792), .Z(n36301) );
  XNOR U36043 ( .A(n36302), .B(n35132), .Z(n28792) );
  IV U36044 ( .A(n35340), .Z(n35132) );
  XOR U36045 ( .A(n36303), .B(n36304), .Z(n35340) );
  ANDN U36046 ( .B(n36305), .A(n35339), .Z(n36302) );
  XNOR U36047 ( .A(n36306), .B(n35136), .Z(n30380) );
  XOR U36048 ( .A(n36307), .B(n36308), .Z(n35136) );
  XOR U36049 ( .A(n32726), .B(n36310), .Z(n36300) );
  XOR U36050 ( .A(n30273), .B(n33145), .Z(n36310) );
  XNOR U36051 ( .A(n36311), .B(n35346), .Z(n33145) );
  XNOR U36052 ( .A(n36312), .B(n35630), .Z(n35346) );
  NOR U36053 ( .A(n36313), .B(n35345), .Z(n36311) );
  XOR U36054 ( .A(n36314), .B(n35145), .Z(n30273) );
  XNOR U36055 ( .A(n36315), .B(n36316), .Z(n35145) );
  ANDN U36056 ( .B(n35350), .A(n36317), .Z(n36314) );
  XNOR U36057 ( .A(n36318), .B(n35247), .Z(n32726) );
  XNOR U36058 ( .A(n36319), .B(n36320), .Z(n35247) );
  ANDN U36059 ( .B(n35348), .A(n36321), .Z(n36318) );
  XNOR U36060 ( .A(n36322), .B(n27590), .Z(n25997) );
  XOR U36061 ( .A(n36323), .B(n34688), .Z(n27590) );
  XNOR U36062 ( .A(n32372), .B(n36324), .Z(n34688) );
  XOR U36063 ( .A(n36325), .B(n36326), .Z(n32372) );
  XNOR U36064 ( .A(n32985), .B(n30207), .Z(n36326) );
  XNOR U36065 ( .A(n36327), .B(n33157), .Z(n30207) );
  ANDN U36066 ( .B(n33158), .A(n36328), .Z(n36327) );
  XNOR U36067 ( .A(n36329), .B(n34325), .Z(n32985) );
  ANDN U36068 ( .B(n34324), .A(n36330), .Z(n36329) );
  XOR U36069 ( .A(n31678), .B(n36331), .Z(n36325) );
  XOR U36070 ( .A(n31914), .B(n32957), .Z(n36331) );
  XOR U36071 ( .A(n36332), .B(n33161), .Z(n32957) );
  ANDN U36072 ( .B(n33162), .A(n36333), .Z(n36332) );
  XNOR U36073 ( .A(n36334), .B(n33172), .Z(n31914) );
  ANDN U36074 ( .B(n33171), .A(n36335), .Z(n36334) );
  XNOR U36075 ( .A(n36336), .B(n33167), .Z(n31678) );
  ANDN U36076 ( .B(n33168), .A(n36337), .Z(n36336) );
  XOR U36077 ( .A(n31943), .B(n36338), .Z(n27591) );
  XNOR U36078 ( .A(n36339), .B(n36340), .Z(n26511) );
  XOR U36079 ( .A(n26717), .B(n26029), .Z(n36340) );
  XOR U36080 ( .A(n36341), .B(n29841), .Z(n26029) );
  XNOR U36081 ( .A(n34253), .B(n33036), .Z(n29841) );
  IV U36082 ( .A(n32266), .Z(n33036) );
  XOR U36083 ( .A(n36342), .B(n34225), .Z(n32266) );
  XNOR U36084 ( .A(n36343), .B(n36344), .Z(n34225) );
  XNOR U36085 ( .A(n32416), .B(n33609), .Z(n36344) );
  XOR U36086 ( .A(n36345), .B(n34163), .Z(n33609) );
  XOR U36087 ( .A(n36346), .B(n36347), .Z(n34163) );
  ANDN U36088 ( .B(n34164), .A(n36348), .Z(n36345) );
  XOR U36089 ( .A(n36349), .B(n33617), .Z(n32416) );
  XOR U36090 ( .A(n36350), .B(n36351), .Z(n33617) );
  NOR U36091 ( .A(n33616), .B(n34262), .Z(n36349) );
  XNOR U36092 ( .A(n36352), .B(n36353), .Z(n33616) );
  XOR U36093 ( .A(n30534), .B(n36354), .Z(n36343) );
  XNOR U36094 ( .A(n31935), .B(n33189), .Z(n36354) );
  XOR U36095 ( .A(n36355), .B(n33622), .Z(n33189) );
  XOR U36096 ( .A(n36356), .B(n36357), .Z(n33622) );
  ANDN U36097 ( .B(n33623), .A(n34255), .Z(n36355) );
  XOR U36098 ( .A(n36358), .B(n36359), .Z(n33623) );
  XNOR U36099 ( .A(n36360), .B(n33988), .Z(n31935) );
  XOR U36100 ( .A(n36361), .B(n36362), .Z(n33988) );
  XOR U36101 ( .A(n36363), .B(n36364), .Z(n33989) );
  XNOR U36102 ( .A(n36365), .B(n33626), .Z(n30534) );
  XNOR U36103 ( .A(n36366), .B(n36367), .Z(n33626) );
  XOR U36104 ( .A(n36368), .B(n36369), .Z(n33627) );
  XOR U36105 ( .A(n36370), .B(n34164), .Z(n34253) );
  XNOR U36106 ( .A(n35378), .B(n36371), .Z(n34164) );
  ANDN U36107 ( .B(n36348), .A(n35700), .Z(n36370) );
  XOR U36108 ( .A(n31570), .B(n33076), .Z(n28191) );
  XNOR U36109 ( .A(n36372), .B(n36373), .Z(n33076) );
  NOR U36110 ( .A(n36374), .B(n34744), .Z(n36372) );
  XNOR U36111 ( .A(n36375), .B(n34398), .Z(n31570) );
  XNOR U36112 ( .A(n36376), .B(n36377), .Z(n34398) );
  XOR U36113 ( .A(n31989), .B(n33851), .Z(n36377) );
  XOR U36114 ( .A(n36378), .B(n34718), .Z(n33851) );
  ANDN U36115 ( .B(n34874), .A(n34873), .Z(n36378) );
  IV U36116 ( .A(n36379), .Z(n34874) );
  XOR U36117 ( .A(n36380), .B(n34725), .Z(n31989) );
  ANDN U36118 ( .B(n34861), .A(n34862), .Z(n36380) );
  XOR U36119 ( .A(n28835), .B(n36381), .Z(n36376) );
  XOR U36120 ( .A(n32716), .B(n32509), .Z(n36381) );
  XNOR U36121 ( .A(n36382), .B(n34728), .Z(n32509) );
  ANDN U36122 ( .B(n34865), .A(n34866), .Z(n36382) );
  XNOR U36123 ( .A(n36383), .B(n34714), .Z(n32716) );
  ANDN U36124 ( .B(n34871), .A(n34870), .Z(n36383) );
  XNOR U36125 ( .A(n36384), .B(n36385), .Z(n28835) );
  ANDN U36126 ( .B(n34876), .A(n34877), .Z(n36384) );
  XOR U36127 ( .A(n35542), .B(n33550), .Z(n28193) );
  XOR U36128 ( .A(n32915), .B(n35949), .Z(n33550) );
  XNOR U36129 ( .A(n36386), .B(n36387), .Z(n35949) );
  XNOR U36130 ( .A(n32681), .B(n33066), .Z(n36387) );
  XNOR U36131 ( .A(n36388), .B(n35813), .Z(n33066) );
  NOR U36132 ( .A(n35814), .B(n35545), .Z(n36388) );
  XOR U36133 ( .A(n36389), .B(n36390), .Z(n35814) );
  XNOR U36134 ( .A(n36391), .B(n35809), .Z(n32681) );
  ANDN U36135 ( .B(n35549), .A(n35550), .Z(n36391) );
  XOR U36136 ( .A(n36392), .B(n36393), .Z(n35549) );
  XNOR U36137 ( .A(n35803), .B(n36394), .Z(n36386) );
  XOR U36138 ( .A(n32366), .B(n31670), .Z(n36394) );
  XNOR U36139 ( .A(n36395), .B(n36396), .Z(n31670) );
  ANDN U36140 ( .B(n35553), .A(n35554), .Z(n36395) );
  XNOR U36141 ( .A(n36397), .B(n35817), .Z(n32366) );
  ANDN U36142 ( .B(n35557), .A(n35558), .Z(n36397) );
  XOR U36143 ( .A(n36398), .B(n36369), .Z(n35557) );
  XNOR U36144 ( .A(n36399), .B(n35820), .Z(n35803) );
  ANDN U36145 ( .B(n35821), .A(n36400), .Z(n36399) );
  XNOR U36146 ( .A(n36401), .B(n36402), .Z(n32915) );
  XOR U36147 ( .A(n32596), .B(n31893), .Z(n36402) );
  XNOR U36148 ( .A(n36403), .B(n36404), .Z(n31893) );
  XOR U36149 ( .A(n36405), .B(n36406), .Z(n35836) );
  XOR U36150 ( .A(n36407), .B(n35826), .Z(n32596) );
  ANDN U36151 ( .B(n35827), .A(n36004), .Z(n36407) );
  XNOR U36152 ( .A(n36408), .B(n36409), .Z(n35827) );
  XNOR U36153 ( .A(n32188), .B(n36410), .Z(n36401) );
  XOR U36154 ( .A(n32840), .B(n32516), .Z(n36410) );
  XNOR U36155 ( .A(n36411), .B(n35843), .Z(n32516) );
  AND U36156 ( .A(n36015), .B(n35844), .Z(n36411) );
  XOR U36157 ( .A(n36412), .B(n36413), .Z(n35844) );
  XNOR U36158 ( .A(n36414), .B(n35830), .Z(n32840) );
  ANDN U36159 ( .B(n35831), .A(n36415), .Z(n36414) );
  XNOR U36160 ( .A(n36416), .B(n36417), .Z(n35831) );
  XNOR U36161 ( .A(n36418), .B(n35840), .Z(n32188) );
  XOR U36162 ( .A(n36419), .B(n36420), .Z(n35839) );
  XOR U36163 ( .A(n36421), .B(n35821), .Z(n35542) );
  XNOR U36164 ( .A(n36422), .B(n36423), .Z(n35821) );
  ANDN U36165 ( .B(n36400), .A(n36424), .Z(n36421) );
  XNOR U36166 ( .A(n36425), .B(n26300), .Z(n26717) );
  XOR U36167 ( .A(n36426), .B(n28462), .Z(n26300) );
  ANDN U36168 ( .B(n28196), .A(n28195), .Z(n36425) );
  XOR U36169 ( .A(n36427), .B(n31539), .Z(n28195) );
  XOR U36170 ( .A(n35463), .B(n31865), .Z(n28196) );
  IV U36171 ( .A(n32182), .Z(n31865) );
  XOR U36172 ( .A(n32713), .B(n36428), .Z(n32182) );
  XOR U36173 ( .A(n36429), .B(n36430), .Z(n32713) );
  XNOR U36174 ( .A(n31261), .B(n31266), .Z(n36430) );
  XNOR U36175 ( .A(n36431), .B(n32474), .Z(n31266) );
  XNOR U36176 ( .A(n36432), .B(n35632), .Z(n32474) );
  NOR U36177 ( .A(n35459), .B(n32473), .Z(n36431) );
  XOR U36178 ( .A(n36433), .B(n36434), .Z(n32473) );
  XNOR U36179 ( .A(n36435), .B(n32468), .Z(n31261) );
  XOR U36180 ( .A(n36436), .B(n36437), .Z(n32468) );
  AND U36181 ( .A(n32467), .B(n35466), .Z(n36435) );
  XOR U36182 ( .A(n36438), .B(n36439), .Z(n32467) );
  XNOR U36183 ( .A(n32209), .B(n36440), .Z(n36429) );
  XOR U36184 ( .A(n30257), .B(n31746), .Z(n36440) );
  XNOR U36185 ( .A(n36441), .B(n32477), .Z(n31746) );
  XOR U36186 ( .A(n36442), .B(n36443), .Z(n32477) );
  ANDN U36187 ( .B(n32478), .A(n35462), .Z(n36441) );
  XNOR U36188 ( .A(n36444), .B(n36445), .Z(n32478) );
  XNOR U36189 ( .A(n36446), .B(n34602), .Z(n30257) );
  AND U36190 ( .A(n34601), .B(n35470), .Z(n36446) );
  XOR U36191 ( .A(n36447), .B(n35952), .Z(n34601) );
  XNOR U36192 ( .A(n36448), .B(n32880), .Z(n32209) );
  XOR U36193 ( .A(n36449), .B(n36450), .Z(n32880) );
  ANDN U36194 ( .B(n32879), .A(n36451), .Z(n36448) );
  XNOR U36195 ( .A(n36452), .B(n32879), .Z(n35463) );
  XOR U36196 ( .A(n35769), .B(n36453), .Z(n32879) );
  XOR U36197 ( .A(n30157), .B(n36454), .Z(n36339) );
  XNOR U36198 ( .A(n29278), .B(n33010), .Z(n36454) );
  XOR U36199 ( .A(n36455), .B(n26310), .Z(n33010) );
  XOR U36200 ( .A(n35114), .B(n31584), .Z(n26310) );
  XOR U36201 ( .A(n36456), .B(n34062), .Z(n35114) );
  ANDN U36202 ( .B(n28183), .A(n28184), .Z(n36455) );
  XNOR U36203 ( .A(n31943), .B(n36458), .Z(n28184) );
  IV U36204 ( .A(n31785), .Z(n31943) );
  XNOR U36205 ( .A(n33992), .B(n34525), .Z(n31785) );
  XNOR U36206 ( .A(n36459), .B(n36460), .Z(n34525) );
  XNOR U36207 ( .A(n31332), .B(n36461), .Z(n36460) );
  XNOR U36208 ( .A(n36462), .B(n36463), .Z(n31332) );
  NOR U36209 ( .A(n36464), .B(n36465), .Z(n36462) );
  XOR U36210 ( .A(n31937), .B(n36466), .Z(n36459) );
  XOR U36211 ( .A(n31830), .B(n28878), .Z(n36466) );
  XOR U36212 ( .A(n36467), .B(n36468), .Z(n28878) );
  ANDN U36213 ( .B(n36469), .A(n36470), .Z(n36467) );
  ANDN U36214 ( .B(n36473), .A(n36474), .Z(n36471) );
  XNOR U36215 ( .A(n36475), .B(n36476), .Z(n31937) );
  NOR U36216 ( .A(n36477), .B(n36478), .Z(n36475) );
  XOR U36217 ( .A(n36479), .B(n36480), .Z(n33992) );
  XOR U36218 ( .A(n30750), .B(n36481), .Z(n36480) );
  XNOR U36219 ( .A(n36482), .B(n36483), .Z(n30750) );
  XOR U36220 ( .A(n32561), .B(n36485), .Z(n36479) );
  XNOR U36221 ( .A(n32149), .B(n30128), .Z(n36485) );
  XNOR U36222 ( .A(n36486), .B(n36487), .Z(n30128) );
  ANDN U36223 ( .B(n36488), .A(n36058), .Z(n36486) );
  IV U36224 ( .A(n36489), .Z(n36058) );
  XNOR U36225 ( .A(n36490), .B(n36491), .Z(n32149) );
  ANDN U36226 ( .B(n36492), .A(n36049), .Z(n36490) );
  XNOR U36227 ( .A(n36493), .B(n36494), .Z(n32561) );
  ANDN U36228 ( .B(n36495), .A(n36062), .Z(n36493) );
  XOR U36229 ( .A(n30198), .B(n36496), .Z(n28183) );
  XOR U36230 ( .A(n36497), .B(n26315), .Z(n29278) );
  XOR U36231 ( .A(n36498), .B(n31707), .Z(n26315) );
  XOR U36232 ( .A(n36499), .B(n36500), .Z(n31707) );
  NOR U36233 ( .A(n28189), .B(n28188), .Z(n36497) );
  XOR U36234 ( .A(n35858), .B(n32498), .Z(n28188) );
  XOR U36235 ( .A(n36501), .B(n33450), .Z(n32498) );
  XNOR U36236 ( .A(n36502), .B(n36503), .Z(n33450) );
  XNOR U36237 ( .A(n32369), .B(n33524), .Z(n36503) );
  XOR U36238 ( .A(n36504), .B(n34040), .Z(n33524) );
  ANDN U36239 ( .B(n34039), .A(n36505), .Z(n36504) );
  XOR U36240 ( .A(n36506), .B(n36507), .Z(n34039) );
  XOR U36241 ( .A(n36508), .B(n34027), .Z(n32369) );
  ANDN U36242 ( .B(n34026), .A(n36509), .Z(n36508) );
  XOR U36243 ( .A(n33821), .B(n36510), .Z(n36502) );
  XOR U36244 ( .A(n33672), .B(n32744), .Z(n36510) );
  XOR U36245 ( .A(n36511), .B(n34032), .Z(n32744) );
  NOR U36246 ( .A(n34031), .B(n35855), .Z(n36511) );
  XOR U36247 ( .A(n36512), .B(n36513), .Z(n34031) );
  XNOR U36248 ( .A(n36514), .B(n36515), .Z(n33672) );
  ANDN U36249 ( .B(n35851), .A(n35852), .Z(n36514) );
  XNOR U36250 ( .A(n36516), .B(n36517), .Z(n33821) );
  ANDN U36251 ( .B(n35861), .A(n34035), .Z(n36516) );
  IV U36252 ( .A(n35860), .Z(n34035) );
  XOR U36253 ( .A(n36518), .B(n36519), .Z(n35860) );
  XNOR U36254 ( .A(n36520), .B(n34026), .Z(n35858) );
  XNOR U36255 ( .A(n36521), .B(n36522), .Z(n34026) );
  ANDN U36256 ( .B(n36509), .A(n36523), .Z(n36520) );
  XOR U36257 ( .A(n36524), .B(n32875), .Z(n28189) );
  XNOR U36258 ( .A(n36525), .B(n33021), .Z(n30157) );
  IV U36259 ( .A(n26304), .Z(n33021) );
  XOR U36260 ( .A(n35735), .B(n32456), .Z(n26304) );
  XNOR U36261 ( .A(n36526), .B(n36527), .Z(n35735) );
  ANDN U36262 ( .B(n36528), .A(n36529), .Z(n36526) );
  ANDN U36263 ( .B(n28181), .A(n33020), .Z(n36525) );
  IV U36264 ( .A(n28180), .Z(n33020) );
  XOR U36265 ( .A(n34721), .B(n28895), .Z(n28180) );
  IV U36266 ( .A(n30290), .Z(n28895) );
  XOR U36267 ( .A(n32651), .B(n36530), .Z(n30290) );
  XNOR U36268 ( .A(n36531), .B(n36532), .Z(n32651) );
  XOR U36269 ( .A(n33138), .B(n31692), .Z(n36532) );
  XOR U36270 ( .A(n36533), .B(n35383), .Z(n31692) );
  NOR U36271 ( .A(n34010), .B(n33869), .Z(n36533) );
  XOR U36272 ( .A(n36534), .B(n36535), .Z(n33869) );
  IV U36273 ( .A(n35384), .Z(n34010) );
  XOR U36274 ( .A(n36536), .B(n36537), .Z(n35384) );
  XOR U36275 ( .A(n36538), .B(n36539), .Z(n33138) );
  NOR U36276 ( .A(n33873), .B(n34004), .Z(n36538) );
  XOR U36277 ( .A(n36540), .B(n36541), .Z(n33873) );
  XOR U36278 ( .A(n35361), .B(n36542), .Z(n36531) );
  XOR U36279 ( .A(n30374), .B(n32977), .Z(n36542) );
  XNOR U36280 ( .A(n36543), .B(n35391), .Z(n32977) );
  NOR U36281 ( .A(n33865), .B(n34014), .Z(n36543) );
  XOR U36282 ( .A(n36544), .B(n36545), .Z(n34014) );
  XOR U36283 ( .A(n36546), .B(n36547), .Z(n33865) );
  XNOR U36284 ( .A(n36548), .B(n36549), .Z(n30374) );
  NOR U36285 ( .A(n33860), .B(n34012), .Z(n36548) );
  XOR U36286 ( .A(n36550), .B(n36551), .Z(n34012) );
  XOR U36287 ( .A(n36356), .B(n36552), .Z(n33860) );
  XNOR U36288 ( .A(n36553), .B(n35386), .Z(n35361) );
  NOR U36289 ( .A(n34007), .B(n33856), .Z(n36553) );
  XNOR U36290 ( .A(n36554), .B(n36555), .Z(n33856) );
  IV U36291 ( .A(n35387), .Z(n34007) );
  XOR U36292 ( .A(n36556), .B(n36557), .Z(n35387) );
  XNOR U36293 ( .A(n36558), .B(n34878), .Z(n34721) );
  ANDN U36294 ( .B(n36559), .A(n36385), .Z(n36558) );
  XNOR U36295 ( .A(n36561), .B(n36562), .Z(n33960) );
  XOR U36296 ( .A(n30064), .B(n30010), .Z(n36562) );
  XNOR U36297 ( .A(n36563), .B(n35268), .Z(n30010) );
  IV U36298 ( .A(n36564), .Z(n35268) );
  AND U36299 ( .A(n36565), .B(n36566), .Z(n36563) );
  XOR U36300 ( .A(n36567), .B(n35272), .Z(n30064) );
  ANDN U36301 ( .B(n36568), .A(n36569), .Z(n36567) );
  XOR U36302 ( .A(n33521), .B(n36570), .Z(n36561) );
  XNOR U36303 ( .A(n36571), .B(n29944), .Z(n36570) );
  XOR U36304 ( .A(n36572), .B(n35259), .Z(n29944) );
  XNOR U36305 ( .A(n36575), .B(n35264), .Z(n33521) );
  AND U36306 ( .A(n36576), .B(n36577), .Z(n36575) );
  XNOR U36307 ( .A(n36578), .B(n36579), .Z(n35353) );
  XNOR U36308 ( .A(n32689), .B(n36242), .Z(n36579) );
  XNOR U36309 ( .A(n36580), .B(n36261), .Z(n36242) );
  AND U36310 ( .A(n36262), .B(n36581), .Z(n36580) );
  ANDN U36311 ( .B(n36583), .A(n36248), .Z(n36582) );
  XOR U36312 ( .A(n32643), .B(n36584), .Z(n36578) );
  XOR U36313 ( .A(n33554), .B(n31871), .Z(n36584) );
  XNOR U36314 ( .A(n36585), .B(n36257), .Z(n31871) );
  AND U36315 ( .A(n36258), .B(n36586), .Z(n36585) );
  XNOR U36316 ( .A(n36587), .B(n36253), .Z(n33554) );
  ANDN U36317 ( .B(n36252), .A(n36588), .Z(n36587) );
  XNOR U36318 ( .A(n36589), .B(n36265), .Z(n32643) );
  XNOR U36319 ( .A(n36591), .B(n27608), .Z(n28199) );
  XOR U36320 ( .A(n35442), .B(n31822), .Z(n27608) );
  IV U36321 ( .A(n30943), .Z(n31822) );
  XOR U36322 ( .A(n36592), .B(n35670), .Z(n35442) );
  ANDN U36323 ( .B(n36593), .A(n34588), .Z(n36592) );
  NOR U36324 ( .A(n36238), .B(n31284), .Z(n36591) );
  XOR U36325 ( .A(n25488), .B(n27654), .Z(n25138) );
  XNOR U36326 ( .A(n36594), .B(n31101), .Z(n27654) );
  ANDN U36327 ( .B(n26361), .A(n26362), .Z(n36594) );
  XOR U36328 ( .A(n36595), .B(n28462), .Z(n26362) );
  XNOR U36329 ( .A(n35352), .B(n32501), .Z(n28462) );
  XNOR U36330 ( .A(n36596), .B(n36597), .Z(n32501) );
  XNOR U36331 ( .A(n32450), .B(n31213), .Z(n36597) );
  XNOR U36332 ( .A(n36598), .B(n35406), .Z(n31213) );
  ANDN U36333 ( .B(n36599), .A(n36600), .Z(n36598) );
  XNOR U36334 ( .A(n36601), .B(n35411), .Z(n32450) );
  ANDN U36335 ( .B(n36602), .A(n36603), .Z(n36601) );
  XOR U36336 ( .A(n28983), .B(n36604), .Z(n36596) );
  XOR U36337 ( .A(n36605), .B(n33123), .Z(n36604) );
  XNOR U36338 ( .A(n36606), .B(n35415), .Z(n33123) );
  ANDN U36339 ( .B(n36607), .A(n36608), .Z(n36606) );
  XNOR U36340 ( .A(n36609), .B(n35419), .Z(n28983) );
  NOR U36341 ( .A(n36610), .B(n36611), .Z(n36609) );
  XOR U36342 ( .A(n36612), .B(n36613), .Z(n35352) );
  XOR U36343 ( .A(n32565), .B(n31365), .Z(n36613) );
  XNOR U36344 ( .A(n36614), .B(n36615), .Z(n31365) );
  ANDN U36345 ( .B(n36616), .A(n36617), .Z(n36614) );
  XOR U36346 ( .A(n36618), .B(n36619), .Z(n32565) );
  NOR U36347 ( .A(n36620), .B(n36621), .Z(n36618) );
  XNOR U36348 ( .A(n33734), .B(n36622), .Z(n36612) );
  XOR U36349 ( .A(n31612), .B(n32815), .Z(n36622) );
  XNOR U36350 ( .A(n36623), .B(n36624), .Z(n32815) );
  ANDN U36351 ( .B(n36625), .A(n36626), .Z(n36623) );
  XNOR U36352 ( .A(n36627), .B(n36628), .Z(n31612) );
  ANDN U36353 ( .B(n36629), .A(n36630), .Z(n36627) );
  XOR U36354 ( .A(n36631), .B(n36632), .Z(n33734) );
  ANDN U36355 ( .B(n36633), .A(n36634), .Z(n36631) );
  XOR U36356 ( .A(n30106), .B(n25103), .Z(n25488) );
  XOR U36357 ( .A(n36635), .B(n36636), .Z(n25103) );
  XOR U36358 ( .A(n25205), .B(n26765), .Z(n36636) );
  XOR U36359 ( .A(n36637), .B(n27132), .Z(n26765) );
  XOR U36360 ( .A(n35741), .B(n32456), .Z(n27132) );
  XNOR U36361 ( .A(n36638), .B(n36639), .Z(n35741) );
  NOR U36362 ( .A(n36640), .B(n36641), .Z(n36638) );
  ANDN U36363 ( .B(n31101), .A(n26361), .Z(n36637) );
  XOR U36364 ( .A(n36642), .B(n32993), .Z(n26361) );
  IV U36365 ( .A(n32891), .Z(n32993) );
  XOR U36366 ( .A(n34792), .B(n34503), .Z(n32891) );
  XNOR U36367 ( .A(n36643), .B(n36644), .Z(n34503) );
  XNOR U36368 ( .A(n34439), .B(n36172), .Z(n36644) );
  XNOR U36369 ( .A(n36645), .B(n34238), .Z(n36172) );
  ANDN U36370 ( .B(n36646), .A(n36274), .Z(n36645) );
  XNOR U36371 ( .A(n36647), .B(n36285), .Z(n34439) );
  ANDN U36372 ( .B(n36648), .A(n36281), .Z(n36647) );
  XNOR U36373 ( .A(n33534), .B(n36649), .Z(n36643) );
  XNOR U36374 ( .A(n31617), .B(n31791), .Z(n36649) );
  XNOR U36375 ( .A(n36650), .B(n34243), .Z(n31791) );
  ANDN U36376 ( .B(n36277), .A(n36651), .Z(n36650) );
  XOR U36377 ( .A(n36652), .B(n34233), .Z(n31617) );
  AND U36378 ( .A(n36279), .B(n36653), .Z(n36652) );
  XNOR U36379 ( .A(n36654), .B(n36655), .Z(n33534) );
  ANDN U36380 ( .B(n36656), .A(n36272), .Z(n36654) );
  XOR U36381 ( .A(n36657), .B(n36658), .Z(n34792) );
  XNOR U36382 ( .A(n33839), .B(n36659), .Z(n36658) );
  XNOR U36383 ( .A(n36660), .B(n36661), .Z(n33839) );
  ANDN U36384 ( .B(n35024), .A(n35022), .Z(n36660) );
  XNOR U36385 ( .A(n29275), .B(n36662), .Z(n36657) );
  XOR U36386 ( .A(n31305), .B(n29070), .Z(n36662) );
  XNOR U36387 ( .A(n36663), .B(n36664), .Z(n29070) );
  ANDN U36388 ( .B(n35014), .A(n35015), .Z(n36663) );
  XNOR U36389 ( .A(n36665), .B(n36666), .Z(n31305) );
  ANDN U36390 ( .B(n35005), .A(n36667), .Z(n36665) );
  XNOR U36391 ( .A(n36668), .B(n36669), .Z(n29275) );
  XOR U36392 ( .A(n36186), .B(n33828), .Z(n31101) );
  IV U36393 ( .A(n32411), .Z(n33828) );
  XOR U36394 ( .A(n36670), .B(n36671), .Z(n36186) );
  NOR U36395 ( .A(n36672), .B(n36673), .Z(n36670) );
  XOR U36396 ( .A(n36674), .B(n27138), .Z(n25205) );
  XOR U36397 ( .A(n34930), .B(n32885), .Z(n27138) );
  XOR U36398 ( .A(n34224), .B(n36675), .Z(n32885) );
  XNOR U36399 ( .A(n36676), .B(n36677), .Z(n34224) );
  XOR U36400 ( .A(n32481), .B(n33462), .Z(n36677) );
  XNOR U36401 ( .A(n36678), .B(n36679), .Z(n33462) );
  NOR U36402 ( .A(n34909), .B(n34908), .Z(n36678) );
  XOR U36403 ( .A(n36680), .B(n36681), .Z(n32481) );
  ANDN U36404 ( .B(n34914), .A(n36682), .Z(n36680) );
  XOR U36405 ( .A(n32390), .B(n36683), .Z(n36676) );
  XOR U36406 ( .A(n32735), .B(n32790), .Z(n36683) );
  XOR U36407 ( .A(n36684), .B(n36685), .Z(n32790) );
  XNOR U36408 ( .A(n36686), .B(n36687), .Z(n32735) );
  XNOR U36409 ( .A(n36688), .B(n36689), .Z(n32390) );
  AND U36410 ( .A(n34927), .B(n34925), .Z(n36688) );
  XNOR U36411 ( .A(n36690), .B(n36691), .Z(n34930) );
  ANDN U36412 ( .B(n36692), .A(n36693), .Z(n36690) );
  NOR U36413 ( .A(n28721), .B(n27665), .Z(n36674) );
  XOR U36414 ( .A(n36694), .B(n29927), .Z(n27665) );
  XNOR U36415 ( .A(n33377), .B(n32185), .Z(n29927) );
  XNOR U36416 ( .A(n36695), .B(n36696), .Z(n32185) );
  XNOR U36417 ( .A(n29301), .B(n31246), .Z(n36696) );
  XNOR U36418 ( .A(n36697), .B(n36698), .Z(n31246) );
  ANDN U36419 ( .B(n33354), .A(n36699), .Z(n36697) );
  XNOR U36420 ( .A(n36700), .B(n36701), .Z(n33354) );
  XNOR U36421 ( .A(n36702), .B(n36703), .Z(n29301) );
  NOR U36422 ( .A(n33335), .B(n33336), .Z(n36702) );
  XOR U36423 ( .A(n36704), .B(n36705), .Z(n33336) );
  XNOR U36424 ( .A(n29065), .B(n36706), .Z(n36695) );
  XNOR U36425 ( .A(n32725), .B(n33243), .Z(n36706) );
  XNOR U36426 ( .A(n36707), .B(n36708), .Z(n33243) );
  AND U36427 ( .A(n33346), .B(n33344), .Z(n36707) );
  XNOR U36428 ( .A(n36709), .B(n36710), .Z(n33346) );
  XOR U36429 ( .A(n36711), .B(n36712), .Z(n32725) );
  ANDN U36430 ( .B(n33339), .A(n33341), .Z(n36711) );
  XOR U36431 ( .A(n36713), .B(n36437), .Z(n33341) );
  XNOR U36432 ( .A(n36714), .B(n36715), .Z(n29065) );
  ANDN U36433 ( .B(n33350), .A(n33348), .Z(n36714) );
  XOR U36434 ( .A(n36716), .B(n36717), .Z(n33350) );
  XNOR U36435 ( .A(n36718), .B(n36719), .Z(n33377) );
  XNOR U36436 ( .A(n36720), .B(n33957), .Z(n36719) );
  XOR U36437 ( .A(n36721), .B(n36722), .Z(n33957) );
  XNOR U36438 ( .A(n36177), .B(n36725), .Z(n36718) );
  XOR U36439 ( .A(n34534), .B(n31578), .Z(n36725) );
  XOR U36440 ( .A(n36726), .B(n36727), .Z(n31578) );
  AND U36441 ( .A(n36728), .B(n36729), .Z(n36726) );
  XNOR U36442 ( .A(n36730), .B(n36731), .Z(n34534) );
  ANDN U36443 ( .B(n36732), .A(n36733), .Z(n36730) );
  XOR U36444 ( .A(n36734), .B(n36735), .Z(n36177) );
  AND U36445 ( .A(n36736), .B(n36737), .Z(n36734) );
  XNOR U36446 ( .A(n30198), .B(n36738), .Z(n28721) );
  XOR U36447 ( .A(n33209), .B(n36739), .Z(n30198) );
  XOR U36448 ( .A(n36740), .B(n36741), .Z(n33209) );
  XOR U36449 ( .A(n36427), .B(n31695), .Z(n36741) );
  XOR U36450 ( .A(n36742), .B(n36743), .Z(n31695) );
  NOR U36451 ( .A(n36744), .B(n36745), .Z(n36742) );
  XNOR U36452 ( .A(n36746), .B(n36747), .Z(n36427) );
  NOR U36453 ( .A(n36748), .B(n36749), .Z(n36746) );
  XOR U36454 ( .A(n31538), .B(n36750), .Z(n36740) );
  XOR U36455 ( .A(n36751), .B(n33413), .Z(n36750) );
  XNOR U36456 ( .A(n36752), .B(n36753), .Z(n33413) );
  NOR U36457 ( .A(n36754), .B(n36755), .Z(n36752) );
  XNOR U36458 ( .A(n36756), .B(n36757), .Z(n31538) );
  NOR U36459 ( .A(n36758), .B(n36759), .Z(n36756) );
  XOR U36460 ( .A(n30802), .B(n36760), .Z(n36635) );
  XNOR U36461 ( .A(n31093), .B(n25234), .Z(n36760) );
  XOR U36462 ( .A(n36761), .B(n31111), .Z(n25234) );
  IV U36463 ( .A(n27126), .Z(n31111) );
  XOR U36464 ( .A(n36762), .B(n33260), .Z(n27126) );
  IV U36465 ( .A(n31159), .Z(n33260) );
  XNOR U36466 ( .A(n36763), .B(n36764), .Z(n33049) );
  XNOR U36467 ( .A(n33324), .B(n34393), .Z(n36764) );
  XNOR U36468 ( .A(n36765), .B(n36766), .Z(n34393) );
  ANDN U36469 ( .B(n34334), .A(n34573), .Z(n36765) );
  XOR U36470 ( .A(n36767), .B(n34564), .Z(n33324) );
  ANDN U36471 ( .B(n34563), .A(n34343), .Z(n36767) );
  XOR U36472 ( .A(n34537), .B(n36768), .Z(n36763) );
  XNOR U36473 ( .A(n32052), .B(n34217), .Z(n36768) );
  XNOR U36474 ( .A(n36769), .B(n34568), .Z(n34217) );
  ANDN U36475 ( .B(n34567), .A(n34339), .Z(n36769) );
  XOR U36476 ( .A(n36770), .B(n34571), .Z(n32052) );
  NOR U36477 ( .A(n36771), .B(n34347), .Z(n36770) );
  XNOR U36478 ( .A(n36772), .B(n36773), .Z(n34537) );
  XNOR U36479 ( .A(n36775), .B(n36776), .Z(n36500) );
  XOR U36480 ( .A(n30278), .B(n31602), .Z(n36776) );
  XNOR U36481 ( .A(n36777), .B(n34324), .Z(n31602) );
  XNOR U36482 ( .A(n36778), .B(n36779), .Z(n34324) );
  XOR U36483 ( .A(n36781), .B(n33171), .Z(n30278) );
  XNOR U36484 ( .A(n36782), .B(n36783), .Z(n33171) );
  XNOR U36485 ( .A(n31256), .B(n36785), .Z(n36775) );
  XNOR U36486 ( .A(n32371), .B(n31798), .Z(n36785) );
  XOR U36487 ( .A(n36786), .B(n33168), .Z(n31798) );
  XNOR U36488 ( .A(n36787), .B(n35606), .Z(n33168) );
  XNOR U36489 ( .A(n36789), .B(n33158), .Z(n32371) );
  XNOR U36490 ( .A(n36790), .B(n35595), .Z(n33158) );
  XOR U36491 ( .A(n36792), .B(n33162), .Z(n31256) );
  XNOR U36492 ( .A(n36793), .B(n36794), .Z(n33162) );
  ANDN U36493 ( .B(n36333), .A(n36795), .Z(n36792) );
  XOR U36494 ( .A(n36796), .B(n27933), .Z(n27660) );
  XNOR U36495 ( .A(n36798), .B(n36799), .Z(n35847) );
  XNOR U36496 ( .A(n32354), .B(n32001), .Z(n36799) );
  XNOR U36497 ( .A(n36800), .B(n36801), .Z(n32001) );
  ANDN U36498 ( .B(n35744), .A(n36802), .Z(n36800) );
  XNOR U36499 ( .A(n36803), .B(n36804), .Z(n32354) );
  NOR U36500 ( .A(n36805), .B(n36806), .Z(n36803) );
  XOR U36501 ( .A(n32902), .B(n36807), .Z(n36798) );
  XOR U36502 ( .A(n31433), .B(n33448), .Z(n36807) );
  XNOR U36503 ( .A(n36808), .B(n36809), .Z(n33448) );
  NOR U36504 ( .A(n36810), .B(n36639), .Z(n36808) );
  XNOR U36505 ( .A(n36811), .B(n36812), .Z(n31433) );
  ANDN U36506 ( .B(n36813), .A(n36527), .Z(n36811) );
  IV U36507 ( .A(n36814), .Z(n36527) );
  XNOR U36508 ( .A(n36815), .B(n36816), .Z(n32902) );
  NOR U36509 ( .A(n36817), .B(n35737), .Z(n36815) );
  XOR U36510 ( .A(n31054), .B(n36818), .Z(n26355) );
  XNOR U36511 ( .A(n36819), .B(n27135), .Z(n31093) );
  IV U36512 ( .A(n31108), .Z(n27135) );
  XOR U36513 ( .A(n36820), .B(n28814), .Z(n31108) );
  IV U36514 ( .A(n31807), .Z(n28814) );
  XNOR U36515 ( .A(n34669), .B(n33538), .Z(n31807) );
  XNOR U36516 ( .A(n36821), .B(n36822), .Z(n33538) );
  XOR U36517 ( .A(n28808), .B(n35212), .Z(n36822) );
  XOR U36518 ( .A(n36823), .B(n36824), .Z(n35212) );
  ANDN U36519 ( .B(n36825), .A(n36235), .Z(n36823) );
  XNOR U36520 ( .A(n36826), .B(n36827), .Z(n28808) );
  AND U36521 ( .A(n35907), .B(n36828), .Z(n36826) );
  XOR U36522 ( .A(n35891), .B(n36829), .Z(n36821) );
  XOR U36523 ( .A(n36830), .B(n31661), .Z(n36829) );
  XOR U36524 ( .A(n36831), .B(n36832), .Z(n31661) );
  ANDN U36525 ( .B(n36833), .A(n35901), .Z(n36831) );
  XNOR U36526 ( .A(n36834), .B(n36835), .Z(n35891) );
  ANDN U36527 ( .B(n36836), .A(n35911), .Z(n36834) );
  XOR U36528 ( .A(n36837), .B(n36838), .Z(n34669) );
  XNOR U36529 ( .A(n29917), .B(n33059), .Z(n36838) );
  XNOR U36530 ( .A(n36839), .B(n36840), .Z(n33059) );
  NOR U36531 ( .A(n36131), .B(n36841), .Z(n36839) );
  XNOR U36532 ( .A(n36842), .B(n36843), .Z(n29917) );
  ANDN U36533 ( .B(n36844), .A(n36845), .Z(n36842) );
  XOR U36534 ( .A(n34430), .B(n36846), .Z(n36837) );
  XNOR U36535 ( .A(n33636), .B(n28740), .Z(n36846) );
  XOR U36536 ( .A(n36847), .B(n36848), .Z(n28740) );
  AND U36537 ( .A(n36145), .B(n36849), .Z(n36847) );
  XNOR U36538 ( .A(n36850), .B(n36851), .Z(n33636) );
  NOR U36539 ( .A(n36852), .B(n36141), .Z(n36850) );
  XOR U36540 ( .A(n36853), .B(n36854), .Z(n34430) );
  ANDN U36541 ( .B(n36855), .A(n36135), .Z(n36853) );
  IV U36542 ( .A(n36856), .Z(n36135) );
  ANDN U36543 ( .B(n26365), .A(n27656), .Z(n36819) );
  XNOR U36544 ( .A(n36857), .B(n28892), .Z(n27656) );
  XOR U36545 ( .A(n36858), .B(n33031), .Z(n26365) );
  IV U36546 ( .A(n31123), .Z(n33031) );
  XNOR U36547 ( .A(n36859), .B(n27129), .Z(n30802) );
  XOR U36548 ( .A(n34742), .B(n30239), .Z(n27129) );
  XNOR U36549 ( .A(n36860), .B(n33481), .Z(n34742) );
  ANDN U36550 ( .B(n36861), .A(n36862), .Z(n36860) );
  XOR U36551 ( .A(n35569), .B(n32691), .Z(n27650) );
  XNOR U36552 ( .A(n36864), .B(n36865), .Z(n34790) );
  XOR U36553 ( .A(n30922), .B(n33474), .Z(n36865) );
  XNOR U36554 ( .A(n36866), .B(n36867), .Z(n33474) );
  ANDN U36555 ( .B(n36476), .A(n36868), .Z(n36866) );
  XOR U36556 ( .A(n36869), .B(n36870), .Z(n30922) );
  XNOR U36557 ( .A(n31629), .B(n36872), .Z(n36864) );
  XOR U36558 ( .A(n33997), .B(n30209), .Z(n36872) );
  XNOR U36559 ( .A(n36873), .B(n36874), .Z(n30209) );
  ANDN U36560 ( .B(n36875), .A(n36468), .Z(n36873) );
  IV U36561 ( .A(n36876), .Z(n36468) );
  XOR U36562 ( .A(n36877), .B(n36878), .Z(n33997) );
  XOR U36563 ( .A(n36880), .B(n36881), .Z(n31629) );
  NOR U36564 ( .A(n36882), .B(n36883), .Z(n36880) );
  XNOR U36565 ( .A(n36884), .B(n36885), .Z(n35569) );
  ANDN U36566 ( .B(n35053), .A(n36886), .Z(n36884) );
  XOR U36567 ( .A(n36887), .B(n34320), .Z(n26946) );
  XNOR U36568 ( .A(n36888), .B(n36889), .Z(n36268) );
  XNOR U36569 ( .A(n32271), .B(n35001), .Z(n36889) );
  XOR U36570 ( .A(n36890), .B(n35006), .Z(n35001) );
  IV U36571 ( .A(n36667), .Z(n35006) );
  XNOR U36572 ( .A(n36891), .B(n36541), .Z(n36667) );
  ANDN U36573 ( .B(n35007), .A(n36892), .Z(n36890) );
  XNOR U36574 ( .A(n36893), .B(n35010), .Z(n32271) );
  XOR U36575 ( .A(n36894), .B(n36895), .Z(n35010) );
  ANDN U36576 ( .B(n35011), .A(n36896), .Z(n36893) );
  XNOR U36577 ( .A(n31160), .B(n36897), .Z(n36888) );
  XNOR U36578 ( .A(n29325), .B(n33606), .Z(n36897) );
  XNOR U36579 ( .A(n36898), .B(n35015), .Z(n33606) );
  XOR U36580 ( .A(n36899), .B(n36900), .Z(n35015) );
  ANDN U36581 ( .B(n35016), .A(n36901), .Z(n36898) );
  XNOR U36582 ( .A(n36902), .B(n35020), .Z(n29325) );
  IV U36583 ( .A(n36903), .Z(n35020) );
  ANDN U36584 ( .B(n36904), .A(n35019), .Z(n36902) );
  XNOR U36585 ( .A(n36905), .B(n35024), .Z(n31160) );
  XOR U36586 ( .A(n36906), .B(n36907), .Z(n35024) );
  ANDN U36587 ( .B(n36908), .A(n35023), .Z(n36905) );
  XOR U36588 ( .A(n36909), .B(n36910), .Z(n32949) );
  XOR U36589 ( .A(n28896), .B(n34402), .Z(n36910) );
  XOR U36590 ( .A(n36911), .B(n36912), .Z(n34402) );
  ANDN U36591 ( .B(n36913), .A(n36914), .Z(n36911) );
  XNOR U36592 ( .A(n36915), .B(n35029), .Z(n28896) );
  NOR U36593 ( .A(n36916), .B(n36917), .Z(n36915) );
  XNOR U36594 ( .A(n31475), .B(n36918), .Z(n36909) );
  XNOR U36595 ( .A(n32489), .B(n30036), .Z(n36918) );
  XNOR U36596 ( .A(n36919), .B(n36920), .Z(n30036) );
  NOR U36597 ( .A(n35033), .B(n36921), .Z(n36919) );
  XNOR U36598 ( .A(n36922), .B(n35043), .Z(n32489) );
  ANDN U36599 ( .B(n36923), .A(n35044), .Z(n36922) );
  XOR U36600 ( .A(n36924), .B(n36925), .Z(n31475) );
  ANDN U36601 ( .B(n35040), .A(n36926), .Z(n36924) );
  XNOR U36602 ( .A(n36927), .B(n36928), .Z(n30106) );
  XOR U36603 ( .A(n25073), .B(n26914), .Z(n36928) );
  XOR U36604 ( .A(n36929), .B(n28131), .Z(n26914) );
  XNOR U36605 ( .A(n35036), .B(n30539), .Z(n28131) );
  XNOR U36606 ( .A(n34793), .B(n33175), .Z(n30539) );
  XNOR U36607 ( .A(n36930), .B(n36931), .Z(n33175) );
  XNOR U36608 ( .A(n36932), .B(n29408), .Z(n36931) );
  XNOR U36609 ( .A(n36933), .B(n35220), .Z(n29408) );
  AND U36610 ( .A(n34410), .B(n34412), .Z(n36933) );
  XOR U36611 ( .A(n36934), .B(n36935), .Z(n34412) );
  XNOR U36612 ( .A(n32514), .B(n36936), .Z(n36930) );
  XOR U36613 ( .A(n31216), .B(n32100), .Z(n36936) );
  XNOR U36614 ( .A(n36937), .B(n34381), .Z(n32100) );
  ANDN U36615 ( .B(n34423), .A(n34422), .Z(n36937) );
  IV U36616 ( .A(n35514), .Z(n34423) );
  XOR U36617 ( .A(n36938), .B(n36939), .Z(n35514) );
  XNOR U36618 ( .A(n36940), .B(n34387), .Z(n31216) );
  ANDN U36619 ( .B(n34415), .A(n34416), .Z(n36940) );
  XOR U36620 ( .A(n36941), .B(n36942), .Z(n34416) );
  XOR U36621 ( .A(n36943), .B(n34391), .Z(n32514) );
  IV U36622 ( .A(n36944), .Z(n34391) );
  ANDN U36623 ( .B(n34407), .A(n34408), .Z(n36943) );
  XOR U36624 ( .A(n36945), .B(n36946), .Z(n34408) );
  XOR U36625 ( .A(n36947), .B(n36948), .Z(n34793) );
  XOR U36626 ( .A(n30955), .B(n32403), .Z(n36948) );
  XOR U36627 ( .A(n36949), .B(n36950), .Z(n32403) );
  ANDN U36628 ( .B(n35032), .A(n36920), .Z(n36949) );
  IV U36629 ( .A(n35034), .Z(n36920) );
  XNOR U36630 ( .A(n36951), .B(n35606), .Z(n35034) );
  XNOR U36631 ( .A(n36952), .B(n36953), .Z(n30955) );
  ANDN U36632 ( .B(n35038), .A(n36925), .Z(n36952) );
  IV U36633 ( .A(n35039), .Z(n36925) );
  XOR U36634 ( .A(n36954), .B(n36955), .Z(n35039) );
  XOR U36635 ( .A(n31262), .B(n36956), .Z(n36947) );
  XNOR U36636 ( .A(n32055), .B(n34948), .Z(n36956) );
  XNOR U36637 ( .A(n36957), .B(n36958), .Z(n34948) );
  ANDN U36638 ( .B(n36959), .A(n36912), .Z(n36957) );
  XOR U36639 ( .A(n36960), .B(n36961), .Z(n32055) );
  NOR U36640 ( .A(n35029), .B(n35028), .Z(n36960) );
  XNOR U36641 ( .A(n36962), .B(n36963), .Z(n35029) );
  XNOR U36642 ( .A(n36964), .B(n36965), .Z(n31262) );
  ANDN U36643 ( .B(n35043), .A(n35042), .Z(n36964) );
  XNOR U36644 ( .A(n36966), .B(n36967), .Z(n35043) );
  XNOR U36645 ( .A(n36968), .B(n36959), .Z(n35036) );
  ANDN U36646 ( .B(n36912), .A(n36913), .Z(n36968) );
  XOR U36647 ( .A(n36969), .B(n36970), .Z(n36912) );
  NOR U36648 ( .A(n31124), .B(n28283), .Z(n36929) );
  XOR U36649 ( .A(n33107), .B(n31355), .Z(n28283) );
  XOR U36650 ( .A(n34178), .B(n32940), .Z(n31355) );
  XNOR U36651 ( .A(n36971), .B(n36972), .Z(n32940) );
  XOR U36652 ( .A(n32591), .B(n33258), .Z(n36972) );
  XNOR U36653 ( .A(n36973), .B(n36974), .Z(n33258) );
  ANDN U36654 ( .B(n33110), .A(n33112), .Z(n36973) );
  XOR U36655 ( .A(n36975), .B(n36976), .Z(n33112) );
  XNOR U36656 ( .A(n36977), .B(n36978), .Z(n32591) );
  ANDN U36657 ( .B(n33114), .A(n33116), .Z(n36977) );
  XOR U36658 ( .A(n36979), .B(n36980), .Z(n33116) );
  XNOR U36659 ( .A(n33940), .B(n36981), .Z(n36971) );
  XNOR U36660 ( .A(n34769), .B(n28791), .Z(n36981) );
  XNOR U36661 ( .A(n36982), .B(n36983), .Z(n28791) );
  ANDN U36662 ( .B(n33104), .A(n35963), .Z(n36982) );
  IV U36663 ( .A(n33105), .Z(n35963) );
  XOR U36664 ( .A(n36550), .B(n36984), .Z(n33105) );
  XNOR U36665 ( .A(n36985), .B(n36986), .Z(n34769) );
  ANDN U36666 ( .B(n35216), .A(n35214), .Z(n36985) );
  XNOR U36667 ( .A(n36987), .B(n36988), .Z(n35216) );
  XNOR U36668 ( .A(n36989), .B(n36990), .Z(n33940) );
  XOR U36669 ( .A(n36992), .B(n36993), .Z(n34178) );
  XOR U36670 ( .A(n34293), .B(n29290), .Z(n36993) );
  XNOR U36671 ( .A(n36994), .B(n34783), .Z(n29290) );
  XNOR U36672 ( .A(n36995), .B(n36996), .Z(n34783) );
  ANDN U36673 ( .B(n33685), .A(n33686), .Z(n36994) );
  XNOR U36674 ( .A(n36997), .B(n35630), .Z(n33685) );
  XNOR U36675 ( .A(n36998), .B(n34780), .Z(n34293) );
  XNOR U36676 ( .A(n36999), .B(n37000), .Z(n34780) );
  ANDN U36677 ( .B(n34183), .A(n34181), .Z(n36998) );
  XOR U36678 ( .A(n37001), .B(n37002), .Z(n34181) );
  XOR U36679 ( .A(n31548), .B(n37003), .Z(n36992) );
  XOR U36680 ( .A(n31601), .B(n31934), .Z(n37003) );
  XNOR U36681 ( .A(n37004), .B(n34776), .Z(n31934) );
  XNOR U36682 ( .A(n37005), .B(n37006), .Z(n34776) );
  XOR U36683 ( .A(n37007), .B(n37008), .Z(n33680) );
  XNOR U36684 ( .A(n37009), .B(n34786), .Z(n31601) );
  NOR U36685 ( .A(n33690), .B(n33689), .Z(n37009) );
  XNOR U36686 ( .A(n37010), .B(n37011), .Z(n33689) );
  XNOR U36687 ( .A(n37012), .B(n35498), .Z(n31548) );
  IV U36688 ( .A(n35476), .Z(n35498) );
  XOR U36689 ( .A(n37013), .B(n37014), .Z(n35476) );
  NOR U36690 ( .A(n33695), .B(n33693), .Z(n37012) );
  XNOR U36691 ( .A(n37015), .B(n37016), .Z(n33693) );
  XNOR U36692 ( .A(n37017), .B(n36991), .Z(n33107) );
  NOR U36693 ( .A(n35972), .B(n35971), .Z(n37017) );
  XOR U36694 ( .A(n37018), .B(n37019), .Z(n35971) );
  XOR U36695 ( .A(n37020), .B(n27937), .Z(n31124) );
  XNOR U36696 ( .A(n33641), .B(n32960), .Z(n27937) );
  XOR U36697 ( .A(n37021), .B(n37022), .Z(n32960) );
  XNOR U36698 ( .A(n31214), .B(n30950), .Z(n37022) );
  XOR U36699 ( .A(n37023), .B(n34573), .Z(n30950) );
  XOR U36700 ( .A(n37024), .B(n37025), .Z(n34573) );
  NOR U36701 ( .A(n34334), .B(n34335), .Z(n37023) );
  XNOR U36702 ( .A(n37026), .B(n37027), .Z(n34334) );
  XNOR U36703 ( .A(n37028), .B(n34563), .Z(n31214) );
  XNOR U36704 ( .A(n37029), .B(n37030), .Z(n34563) );
  XOR U36705 ( .A(n37031), .B(n37032), .Z(n34343) );
  XOR U36706 ( .A(n33047), .B(n37033), .Z(n37021) );
  XOR U36707 ( .A(n29288), .B(n32171), .Z(n37033) );
  XNOR U36708 ( .A(n37034), .B(n34570), .Z(n32171) );
  IV U36709 ( .A(n36771), .Z(n34570) );
  XOR U36710 ( .A(n37035), .B(n37036), .Z(n36771) );
  ANDN U36711 ( .B(n34347), .A(n34348), .Z(n37034) );
  XOR U36712 ( .A(n37037), .B(n36406), .Z(n34347) );
  XNOR U36713 ( .A(n37038), .B(n34567), .Z(n29288) );
  XNOR U36714 ( .A(n37039), .B(n37040), .Z(n34567) );
  ANDN U36715 ( .B(n34339), .A(n34340), .Z(n37038) );
  XNOR U36716 ( .A(n37041), .B(n35320), .Z(n34339) );
  XNOR U36717 ( .A(n37042), .B(n36774), .Z(n33047) );
  NOR U36718 ( .A(n34331), .B(n34330), .Z(n37042) );
  XOR U36719 ( .A(n37043), .B(n37044), .Z(n34330) );
  XOR U36720 ( .A(n37045), .B(n37046), .Z(n33641) );
  XOR U36721 ( .A(n33259), .B(n32570), .Z(n37046) );
  XOR U36722 ( .A(n37047), .B(n36333), .Z(n32570) );
  XOR U36723 ( .A(n37048), .B(n35611), .Z(n36333) );
  XNOR U36724 ( .A(n37049), .B(n36335), .Z(n33259) );
  XNOR U36725 ( .A(n37050), .B(n37051), .Z(n36335) );
  NOR U36726 ( .A(n36784), .B(n33170), .Z(n37049) );
  XOR U36727 ( .A(n31179), .B(n37052), .Z(n37045) );
  XOR U36728 ( .A(n36762), .B(n31158), .Z(n37052) );
  XNOR U36729 ( .A(n37053), .B(n36328), .Z(n31158) );
  XOR U36730 ( .A(n37054), .B(n37055), .Z(n36328) );
  ANDN U36731 ( .B(n36791), .A(n33156), .Z(n37053) );
  XNOR U36732 ( .A(n37056), .B(n36337), .Z(n36762) );
  XOR U36733 ( .A(n37057), .B(n36939), .Z(n36337) );
  NOR U36734 ( .A(n37058), .B(n36788), .Z(n37056) );
  XNOR U36735 ( .A(n37059), .B(n36330), .Z(n31179) );
  XOR U36736 ( .A(n37060), .B(n37061), .Z(n36330) );
  NOR U36737 ( .A(n36780), .B(n34323), .Z(n37059) );
  XNOR U36738 ( .A(n31130), .B(n37062), .Z(n25073) );
  XOR U36739 ( .A(n37063), .B(n37064), .Z(n37062) );
  NANDN U36740 ( .A(rc_i[2]), .B(n11417), .Z(n37064) );
  ANDN U36741 ( .B(n28279), .A(n29517), .Z(n37063) );
  XOR U36742 ( .A(n34740), .B(n32225), .Z(n29517) );
  IV U36743 ( .A(n30239), .Z(n32225) );
  XOR U36744 ( .A(n37065), .B(n36530), .Z(n30239) );
  XNOR U36745 ( .A(n37066), .B(n37067), .Z(n36530) );
  XNOR U36746 ( .A(n34663), .B(n34352), .Z(n37067) );
  XNOR U36747 ( .A(n37068), .B(n34862), .Z(n34352) );
  XNOR U36748 ( .A(n37069), .B(n37070), .Z(n34862) );
  NOR U36749 ( .A(n34723), .B(n34724), .Z(n37068) );
  IV U36750 ( .A(n34863), .Z(n34723) );
  XNOR U36751 ( .A(n37071), .B(n37072), .Z(n34863) );
  XNOR U36752 ( .A(n37073), .B(n34877), .Z(n34663) );
  XOR U36753 ( .A(n37074), .B(n36364), .Z(n34877) );
  ANDN U36754 ( .B(n34878), .A(n36559), .Z(n37073) );
  XOR U36755 ( .A(n37075), .B(n37076), .Z(n34878) );
  XOR U36756 ( .A(n30145), .B(n37077), .Z(n37066) );
  XOR U36757 ( .A(n31412), .B(n34856), .Z(n37077) );
  XOR U36758 ( .A(n37078), .B(n34871), .Z(n34856) );
  XOR U36759 ( .A(n37079), .B(n35159), .Z(n34871) );
  NOR U36760 ( .A(n34715), .B(n34713), .Z(n37078) );
  XOR U36761 ( .A(n37080), .B(n37081), .Z(n34713) );
  XNOR U36762 ( .A(n37082), .B(n36379), .Z(n31412) );
  XOR U36763 ( .A(n37083), .B(n36219), .Z(n36379) );
  NOR U36764 ( .A(n34719), .B(n34717), .Z(n37082) );
  XOR U36765 ( .A(n37084), .B(n37085), .Z(n34717) );
  XNOR U36766 ( .A(n37086), .B(n34866), .Z(n30145) );
  XNOR U36767 ( .A(n35315), .B(n37087), .Z(n34866) );
  ANDN U36768 ( .B(n34729), .A(n34867), .Z(n37086) );
  XOR U36769 ( .A(n37088), .B(n37089), .Z(n34867) );
  IV U36770 ( .A(n37090), .Z(n34729) );
  XNOR U36771 ( .A(n37091), .B(n33086), .Z(n34740) );
  ANDN U36772 ( .B(n37092), .A(n37093), .Z(n37091) );
  XNOR U36773 ( .A(n37094), .B(n28821), .Z(n28279) );
  XOR U36774 ( .A(n36375), .B(n34112), .Z(n28821) );
  XNOR U36775 ( .A(n37095), .B(n37096), .Z(n34112) );
  XNOR U36776 ( .A(n27662), .B(n31969), .Z(n37096) );
  XNOR U36777 ( .A(n37097), .B(n34278), .Z(n31969) );
  XOR U36778 ( .A(n37098), .B(n37099), .Z(n34278) );
  ANDN U36779 ( .B(n36169), .A(n37100), .Z(n37097) );
  XOR U36780 ( .A(n37101), .B(n34292), .Z(n27662) );
  IV U36781 ( .A(n36159), .Z(n34292) );
  XOR U36782 ( .A(n37102), .B(n37103), .Z(n36159) );
  ANDN U36783 ( .B(n36160), .A(n37104), .Z(n37101) );
  XNOR U36784 ( .A(n36154), .B(n37105), .Z(n37095) );
  XOR U36785 ( .A(n35764), .B(n32009), .Z(n37105) );
  XNOR U36786 ( .A(n37106), .B(n36163), .Z(n32009) );
  ANDN U36787 ( .B(n36164), .A(n37107), .Z(n37106) );
  XNOR U36788 ( .A(n37108), .B(n34283), .Z(n35764) );
  XOR U36789 ( .A(n35089), .B(n37109), .Z(n34283) );
  IV U36790 ( .A(n37110), .Z(n35089) );
  ANDN U36791 ( .B(n36167), .A(n37111), .Z(n37108) );
  XNOR U36792 ( .A(n37112), .B(n34288), .Z(n36154) );
  XOR U36793 ( .A(n37113), .B(n37114), .Z(n34288) );
  AND U36794 ( .A(n37115), .B(n36171), .Z(n37112) );
  XOR U36795 ( .A(n37116), .B(n37117), .Z(n36375) );
  XNOR U36796 ( .A(n32836), .B(n31590), .Z(n37117) );
  XNOR U36797 ( .A(n37118), .B(n36861), .Z(n31590) );
  ANDN U36798 ( .B(n33480), .A(n33479), .Z(n37118) );
  ANDN U36799 ( .B(n34996), .A(n34997), .Z(n37119) );
  XOR U36800 ( .A(n31474), .B(n37120), .Z(n37116) );
  XOR U36801 ( .A(n30745), .B(n37121), .Z(n37120) );
  XOR U36802 ( .A(n37122), .B(n34739), .Z(n30745) );
  ANDN U36803 ( .B(n33082), .A(n33080), .Z(n37122) );
  NOR U36804 ( .A(n33084), .B(n33085), .Z(n37123) );
  IV U36805 ( .A(n27110), .Z(n31130) );
  XOR U36806 ( .A(n36720), .B(n34535), .Z(n27110) );
  IV U36807 ( .A(n31579), .Z(n34535) );
  XNOR U36808 ( .A(n37124), .B(n37125), .Z(n34213) );
  XNOR U36809 ( .A(n32291), .B(n37126), .Z(n37125) );
  XNOR U36810 ( .A(n37127), .B(n37128), .Z(n32291) );
  ANDN U36811 ( .B(n36735), .A(n36736), .Z(n37127) );
  XOR U36812 ( .A(n30796), .B(n37129), .Z(n37124) );
  XOR U36813 ( .A(n29094), .B(n30653), .Z(n37129) );
  XNOR U36814 ( .A(n37130), .B(n37131), .Z(n30653) );
  ANDN U36815 ( .B(n37132), .A(n37133), .Z(n37130) );
  XNOR U36816 ( .A(n37134), .B(n37135), .Z(n29094) );
  NOR U36817 ( .A(n37136), .B(n36732), .Z(n37134) );
  XNOR U36818 ( .A(n37137), .B(n37138), .Z(n30796) );
  ANDN U36819 ( .B(n36722), .A(n36724), .Z(n37137) );
  XNOR U36820 ( .A(n37139), .B(n37140), .Z(n33244) );
  XNOR U36821 ( .A(n37141), .B(n29318), .Z(n37140) );
  NOR U36822 ( .A(n33344), .B(n36708), .Z(n37142) );
  XOR U36823 ( .A(n37143), .B(n37144), .Z(n33344) );
  XOR U36824 ( .A(n37145), .B(n37146), .Z(n37139) );
  XOR U36825 ( .A(n36857), .B(n28891), .Z(n37146) );
  XOR U36826 ( .A(n37147), .B(n34803), .Z(n28891) );
  XOR U36827 ( .A(n37148), .B(n37149), .Z(n33348) );
  XNOR U36828 ( .A(n37150), .B(n34811), .Z(n36857) );
  NOR U36829 ( .A(n36712), .B(n33339), .Z(n37150) );
  XOR U36830 ( .A(n37151), .B(n37152), .Z(n33339) );
  XOR U36831 ( .A(n37133), .B(n37153), .Z(n36720) );
  XNOR U36832 ( .A(n11417), .B(n37154), .Z(n37153) );
  NANDN U36833 ( .A(n37132), .B(n37155), .Z(n37154) );
  XOR U36834 ( .A(n30158), .B(n37156), .Z(n36927) );
  XNOR U36835 ( .A(n25675), .B(n21215), .Z(n37156) );
  XOR U36836 ( .A(n37157), .B(n27121), .Z(n21215) );
  XOR U36837 ( .A(n37158), .B(n30748), .Z(n27121) );
  XNOR U36838 ( .A(n33877), .B(n33181), .Z(n30748) );
  XOR U36839 ( .A(n37159), .B(n37160), .Z(n33181) );
  XNOR U36840 ( .A(n34319), .B(n36887), .Z(n37160) );
  XNOR U36841 ( .A(n37161), .B(n35023), .Z(n36887) );
  XOR U36842 ( .A(n37162), .B(n36445), .Z(n35023) );
  IV U36843 ( .A(n37163), .Z(n36445) );
  ANDN U36844 ( .B(n36661), .A(n36908), .Z(n37161) );
  XOR U36845 ( .A(n37164), .B(n35011), .Z(n34319) );
  XNOR U36846 ( .A(n37165), .B(n37166), .Z(n35011) );
  ANDN U36847 ( .B(n36669), .A(n37167), .Z(n37164) );
  XNOR U36848 ( .A(n33381), .B(n37168), .Z(n37159) );
  XNOR U36849 ( .A(n34109), .B(n33711), .Z(n37168) );
  XOR U36850 ( .A(n37169), .B(n35007), .Z(n33711) );
  XOR U36851 ( .A(n37170), .B(n35617), .Z(n35007) );
  AND U36852 ( .A(n36666), .B(n36892), .Z(n37169) );
  XNOR U36853 ( .A(n37171), .B(n35016), .Z(n34109) );
  XNOR U36854 ( .A(n37172), .B(n37173), .Z(n35016) );
  AND U36855 ( .A(n36664), .B(n36901), .Z(n37171) );
  XNOR U36856 ( .A(n37175), .B(n37176), .Z(n35019) );
  NOR U36857 ( .A(n36904), .B(n37177), .Z(n37174) );
  IV U36858 ( .A(n37178), .Z(n36904) );
  XOR U36859 ( .A(n37179), .B(n37180), .Z(n33877) );
  XNOR U36860 ( .A(n30690), .B(n32568), .Z(n37180) );
  XNOR U36861 ( .A(n37181), .B(n35044), .Z(n32568) );
  XNOR U36862 ( .A(n37182), .B(n37183), .Z(n35044) );
  NOR U36863 ( .A(n36965), .B(n36923), .Z(n37181) );
  IV U36864 ( .A(n37184), .Z(n36965) );
  XOR U36865 ( .A(n37185), .B(n36913), .Z(n30690) );
  XNOR U36866 ( .A(n37186), .B(n37187), .Z(n36913) );
  ANDN U36867 ( .B(n36914), .A(n36958), .Z(n37185) );
  IV U36868 ( .A(n37188), .Z(n36958) );
  XNOR U36869 ( .A(n32298), .B(n37189), .Z(n37179) );
  XOR U36870 ( .A(n32947), .B(n32895), .Z(n37189) );
  XOR U36871 ( .A(n37190), .B(n36916), .Z(n32895) );
  IV U36872 ( .A(n35030), .Z(n36916) );
  XNOR U36873 ( .A(n37191), .B(n33927), .Z(n35030) );
  ANDN U36874 ( .B(n36917), .A(n36961), .Z(n37190) );
  IV U36875 ( .A(n37192), .Z(n36961) );
  XNOR U36876 ( .A(n37193), .B(n35033), .Z(n32947) );
  XOR U36877 ( .A(n37194), .B(n35373), .Z(n35033) );
  ANDN U36878 ( .B(n36921), .A(n36950), .Z(n37193) );
  XOR U36879 ( .A(n37195), .B(n35040), .Z(n32298) );
  XOR U36880 ( .A(n37196), .B(n37197), .Z(n35040) );
  ANDN U36881 ( .B(n36926), .A(n37198), .Z(n37195) );
  ANDN U36882 ( .B(n28276), .A(n29531), .Z(n37157) );
  XNOR U36883 ( .A(n33265), .B(n37199), .Z(n29531) );
  XNOR U36884 ( .A(n34176), .B(n35249), .Z(n33265) );
  XNOR U36885 ( .A(n37200), .B(n37201), .Z(n35249) );
  XOR U36886 ( .A(n33130), .B(n33719), .Z(n37201) );
  XOR U36887 ( .A(n37202), .B(n37203), .Z(n33719) );
  ANDN U36888 ( .B(n36249), .A(n36247), .Z(n37202) );
  XOR U36889 ( .A(n37204), .B(n37205), .Z(n36249) );
  XOR U36890 ( .A(n37206), .B(n37207), .Z(n33130) );
  ANDN U36891 ( .B(n36253), .A(n37208), .Z(n37206) );
  XNOR U36892 ( .A(n37209), .B(n37210), .Z(n36253) );
  XOR U36893 ( .A(n27946), .B(n37211), .Z(n37200) );
  XNOR U36894 ( .A(n37212), .B(n33384), .Z(n37211) );
  XNOR U36895 ( .A(n37213), .B(n37214), .Z(n33384) );
  ANDN U36896 ( .B(n36257), .A(n36256), .Z(n37213) );
  XNOR U36897 ( .A(n37215), .B(n37216), .Z(n36257) );
  XNOR U36898 ( .A(n37217), .B(n37218), .Z(n27946) );
  ANDN U36899 ( .B(n36264), .A(n36265), .Z(n37217) );
  XOR U36900 ( .A(n37219), .B(n37220), .Z(n36265) );
  XOR U36901 ( .A(n37221), .B(n37222), .Z(n34176) );
  XNOR U36902 ( .A(n30582), .B(n31882), .Z(n37222) );
  XNOR U36903 ( .A(n37223), .B(n37224), .Z(n31882) );
  NOR U36904 ( .A(n36632), .B(n37225), .Z(n37223) );
  XNOR U36905 ( .A(n37226), .B(n37227), .Z(n30582) );
  ANDN U36906 ( .B(n37228), .A(n36628), .Z(n37226) );
  XOR U36907 ( .A(n37229), .B(n37230), .Z(n37221) );
  XOR U36908 ( .A(n33946), .B(n35954), .Z(n37230) );
  XNOR U36909 ( .A(n37231), .B(n37232), .Z(n35954) );
  NOR U36910 ( .A(n37233), .B(n36615), .Z(n37231) );
  XNOR U36911 ( .A(n37234), .B(n37235), .Z(n33946) );
  ANDN U36912 ( .B(n37236), .A(n36624), .Z(n37234) );
  XOR U36913 ( .A(n35160), .B(n32415), .Z(n28276) );
  XOR U36914 ( .A(n37237), .B(n37238), .Z(n34748) );
  XOR U36915 ( .A(n31755), .B(n30823), .Z(n37238) );
  XNOR U36916 ( .A(n37239), .B(n35174), .Z(n30823) );
  ANDN U36917 ( .B(n37240), .A(n37241), .Z(n37239) );
  XNOR U36918 ( .A(n37242), .B(n35177), .Z(n31755) );
  ANDN U36919 ( .B(n37243), .A(n37244), .Z(n37242) );
  XOR U36920 ( .A(n37245), .B(n37246), .Z(n37237) );
  XOR U36921 ( .A(n33673), .B(n32752), .Z(n37246) );
  XOR U36922 ( .A(n37247), .B(n35184), .Z(n32752) );
  ANDN U36923 ( .B(n37248), .A(n37249), .Z(n37247) );
  XOR U36924 ( .A(n37250), .B(n35186), .Z(n33673) );
  ANDN U36925 ( .B(n37251), .A(n34478), .Z(n37250) );
  XNOR U36926 ( .A(n37252), .B(n37253), .Z(n34250) );
  XNOR U36927 ( .A(n37254), .B(n31701), .Z(n37253) );
  XNOR U36928 ( .A(n37255), .B(n37256), .Z(n31701) );
  NOR U36929 ( .A(n34448), .B(n35157), .Z(n37255) );
  XNOR U36930 ( .A(n37257), .B(n37258), .Z(n34448) );
  XNOR U36931 ( .A(n32943), .B(n37259), .Z(n37252) );
  XOR U36932 ( .A(n35702), .B(n30365), .Z(n37259) );
  XNOR U36933 ( .A(n37260), .B(n34700), .Z(n30365) );
  NOR U36934 ( .A(n37261), .B(n35148), .Z(n37260) );
  XOR U36935 ( .A(n37262), .B(n34696), .Z(n35702) );
  ANDN U36936 ( .B(n35163), .A(n34453), .Z(n37262) );
  XNOR U36937 ( .A(n37263), .B(n37264), .Z(n34453) );
  XOR U36938 ( .A(n37265), .B(n34694), .Z(n32943) );
  NOR U36939 ( .A(n34461), .B(n35153), .Z(n37265) );
  XOR U36940 ( .A(n37266), .B(n37267), .Z(n34461) );
  XNOR U36941 ( .A(n37268), .B(n37261), .Z(n35160) );
  AND U36942 ( .A(n34699), .B(n35148), .Z(n37268) );
  XOR U36943 ( .A(n37269), .B(n37270), .Z(n35148) );
  XOR U36944 ( .A(n37271), .B(n37272), .Z(n34699) );
  XNOR U36945 ( .A(n37273), .B(n28286), .Z(n25675) );
  XOR U36946 ( .A(n36481), .B(n30129), .Z(n28286) );
  XOR U36947 ( .A(n37274), .B(n37275), .Z(n33376) );
  XOR U36948 ( .A(n32484), .B(n31691), .Z(n37275) );
  XNOR U36949 ( .A(n37276), .B(n36088), .Z(n31691) );
  ANDN U36950 ( .B(n37277), .A(n37278), .Z(n37276) );
  XOR U36951 ( .A(n37279), .B(n36074), .Z(n32484) );
  XNOR U36952 ( .A(n33740), .B(n37282), .Z(n37274) );
  XOR U36953 ( .A(n30246), .B(n34212), .Z(n37282) );
  XNOR U36954 ( .A(n37283), .B(n37284), .Z(n34212) );
  XNOR U36955 ( .A(n37287), .B(n36084), .Z(n30246) );
  ANDN U36956 ( .B(n37288), .A(n37289), .Z(n37287) );
  XNOR U36957 ( .A(n37290), .B(n37291), .Z(n33740) );
  ANDN U36958 ( .B(n37292), .A(n37293), .Z(n37290) );
  XOR U36959 ( .A(n37295), .B(n37296), .Z(n36481) );
  NOR U36960 ( .A(n29513), .B(n30103), .Z(n37273) );
  XOR U36961 ( .A(n36190), .B(n32411), .Z(n30103) );
  XNOR U36962 ( .A(n37300), .B(n37301), .Z(n32842) );
  XOR U36963 ( .A(n30945), .B(n27943), .Z(n37301) );
  XOR U36964 ( .A(n37302), .B(n33568), .Z(n27943) );
  ANDN U36965 ( .B(n36193), .A(n33569), .Z(n37302) );
  XNOR U36966 ( .A(n37303), .B(n35320), .Z(n33569) );
  XNOR U36967 ( .A(n37304), .B(n33564), .Z(n30945) );
  ANDN U36968 ( .B(n33565), .A(n37305), .Z(n37304) );
  XOR U36969 ( .A(n33559), .B(n37306), .Z(n37300) );
  XOR U36970 ( .A(n33301), .B(n30218), .Z(n37306) );
  XNOR U36971 ( .A(n37307), .B(n33573), .Z(n30218) );
  NOR U36972 ( .A(n36189), .B(n33574), .Z(n37307) );
  XNOR U36973 ( .A(n37308), .B(n36907), .Z(n33574) );
  XNOR U36974 ( .A(n37309), .B(n37310), .Z(n33301) );
  ANDN U36975 ( .B(n36672), .A(n33577), .Z(n37309) );
  IV U36976 ( .A(n36671), .Z(n33577) );
  XOR U36977 ( .A(n37311), .B(n35526), .Z(n36671) );
  XNOR U36978 ( .A(n37312), .B(n33581), .Z(n33559) );
  NOR U36979 ( .A(n37313), .B(n33582), .Z(n37312) );
  XNOR U36980 ( .A(n37314), .B(n37315), .Z(n33582) );
  XOR U36981 ( .A(n37316), .B(n33565), .Z(n36190) );
  XOR U36982 ( .A(n37317), .B(n37318), .Z(n33565) );
  ANDN U36983 ( .B(n37305), .A(n37319), .Z(n37316) );
  XOR U36984 ( .A(n36123), .B(n32972), .Z(n29513) );
  XNOR U36985 ( .A(n37320), .B(n37321), .Z(n35657) );
  XNOR U36986 ( .A(n32275), .B(n34668), .Z(n37321) );
  XNOR U36987 ( .A(n37322), .B(n34675), .Z(n34668) );
  ANDN U36988 ( .B(n34676), .A(n34969), .Z(n37322) );
  XOR U36989 ( .A(n37323), .B(n37324), .Z(n34969) );
  XOR U36990 ( .A(n37325), .B(n37326), .Z(n34676) );
  XNOR U36991 ( .A(n37327), .B(n35705), .Z(n32275) );
  XOR U36992 ( .A(n37328), .B(n37329), .Z(n34960) );
  XNOR U36993 ( .A(n33004), .B(n37332), .Z(n37320) );
  XOR U36994 ( .A(n32370), .B(n33222), .Z(n37332) );
  XNOR U36995 ( .A(n37333), .B(n34682), .Z(n33222) );
  NOR U36996 ( .A(n34681), .B(n34964), .Z(n37333) );
  XNOR U36997 ( .A(n37334), .B(n36976), .Z(n34964) );
  XOR U36998 ( .A(n37071), .B(n37335), .Z(n34681) );
  XNOR U36999 ( .A(n37336), .B(n37337), .Z(n32370) );
  ANDN U37000 ( .B(n37338), .A(n34972), .Z(n37336) );
  XNOR U37001 ( .A(n37339), .B(n34685), .Z(n33004) );
  ANDN U37002 ( .B(n34686), .A(n36125), .Z(n37339) );
  XOR U37003 ( .A(n37340), .B(n36541), .Z(n36125) );
  XOR U37004 ( .A(n37341), .B(n35155), .Z(n34686) );
  XNOR U37005 ( .A(n37343), .B(n37338), .Z(n36123) );
  ANDN U37006 ( .B(n34972), .A(n34973), .Z(n37343) );
  XNOR U37007 ( .A(n37344), .B(n37345), .Z(n34972) );
  XNOR U37008 ( .A(n37346), .B(n27115), .Z(n30158) );
  XOR U37009 ( .A(n37141), .B(n28892), .Z(n27115) );
  XNOR U37010 ( .A(n37347), .B(n34809), .Z(n37141) );
  ANDN U37011 ( .B(n33335), .A(n36703), .Z(n37347) );
  XOR U37012 ( .A(n37348), .B(n37349), .Z(n33335) );
  NOR U37013 ( .A(n29523), .B(n29521), .Z(n37346) );
  XOR U37014 ( .A(n33281), .B(n32819), .Z(n29521) );
  IV U37015 ( .A(n31314), .Z(n32819) );
  XNOR U37016 ( .A(n35751), .B(n36675), .Z(n31314) );
  XNOR U37017 ( .A(n37350), .B(n37351), .Z(n36675) );
  XNOR U37018 ( .A(n37352), .B(n37353), .Z(n37351) );
  XNOR U37019 ( .A(n34532), .B(n37354), .Z(n37350) );
  XOR U37020 ( .A(n32202), .B(n29061), .Z(n37354) );
  XNOR U37021 ( .A(n37355), .B(n37356), .Z(n29061) );
  ANDN U37022 ( .B(n36691), .A(n36692), .Z(n37355) );
  XOR U37023 ( .A(n37357), .B(n37358), .Z(n32202) );
  ANDN U37024 ( .B(n34937), .A(n34938), .Z(n37357) );
  XNOR U37025 ( .A(n37359), .B(n37360), .Z(n34532) );
  ANDN U37026 ( .B(n34932), .A(n37361), .Z(n37359) );
  XNOR U37027 ( .A(n37362), .B(n37363), .Z(n35751) );
  XOR U37028 ( .A(n37364), .B(n32717), .Z(n37363) );
  XNOR U37029 ( .A(n37365), .B(n37366), .Z(n32717) );
  ANDN U37030 ( .B(n33274), .A(n37367), .Z(n37365) );
  XOR U37031 ( .A(n33060), .B(n37368), .Z(n37362) );
  XOR U37032 ( .A(n32751), .B(n32303), .Z(n37368) );
  XNOR U37033 ( .A(n37369), .B(n36036), .Z(n32303) );
  ANDN U37034 ( .B(n33288), .A(n33289), .Z(n37369) );
  XOR U37035 ( .A(n37370), .B(n33810), .Z(n32751) );
  ANDN U37036 ( .B(n33284), .A(n37371), .Z(n37370) );
  XNOR U37037 ( .A(n37372), .B(n33815), .Z(n33060) );
  ANDN U37038 ( .B(n37373), .A(n37374), .Z(n37372) );
  XNOR U37039 ( .A(n37375), .B(n37373), .Z(n33281) );
  NOR U37040 ( .A(n37376), .B(n33813), .Z(n37375) );
  XOR U37041 ( .A(n32705), .B(n36025), .Z(n29523) );
  XOR U37042 ( .A(n37377), .B(n37378), .Z(n36025) );
  AND U37043 ( .A(n35689), .B(n35687), .Z(n37377) );
  XNOR U37044 ( .A(n37379), .B(n23467), .Z(n25905) );
  XNOR U37045 ( .A(n32812), .B(n25410), .Z(n23467) );
  IV U37046 ( .A(n21382), .Z(n25410) );
  XOR U37047 ( .A(n26929), .B(n27923), .Z(n21382) );
  XNOR U37048 ( .A(n37380), .B(n37381), .Z(n27923) );
  XNOR U37049 ( .A(n21822), .B(n27236), .Z(n37381) );
  XNOR U37050 ( .A(n37382), .B(n27825), .Z(n27236) );
  XOR U37051 ( .A(n35402), .B(n31649), .Z(n27825) );
  IV U37052 ( .A(n28885), .Z(n31649) );
  XNOR U37053 ( .A(n37383), .B(n37384), .Z(n28885) );
  XNOR U37054 ( .A(n37385), .B(n37386), .Z(n35402) );
  ANDN U37055 ( .B(n37387), .A(n37388), .Z(n37385) );
  ANDN U37056 ( .B(n27529), .A(n27527), .Z(n37382) );
  XOR U37057 ( .A(n37389), .B(n31258), .Z(n27527) );
  IV U37058 ( .A(n31229), .Z(n31258) );
  XOR U37059 ( .A(n33449), .B(n35395), .Z(n31229) );
  XNOR U37060 ( .A(n37390), .B(n37391), .Z(n35395) );
  XOR U37061 ( .A(n33829), .B(n37392), .Z(n37391) );
  XNOR U37062 ( .A(n37393), .B(n36107), .Z(n33829) );
  ANDN U37063 ( .B(n37394), .A(n37395), .Z(n37393) );
  XOR U37064 ( .A(n31541), .B(n37396), .Z(n37390) );
  XOR U37065 ( .A(n35998), .B(n31298), .Z(n37396) );
  XNOR U37066 ( .A(n37397), .B(n36111), .Z(n31298) );
  ANDN U37067 ( .B(n37398), .A(n37399), .Z(n37397) );
  XNOR U37068 ( .A(n37400), .B(n36115), .Z(n35998) );
  ANDN U37069 ( .B(n37401), .A(n37402), .Z(n37400) );
  XNOR U37070 ( .A(n37403), .B(n36098), .Z(n31541) );
  ANDN U37071 ( .B(n37404), .A(n37405), .Z(n37403) );
  XOR U37072 ( .A(n37406), .B(n37407), .Z(n33449) );
  XOR U37073 ( .A(n32031), .B(n34019), .Z(n37407) );
  XOR U37074 ( .A(n37408), .B(n36641), .Z(n34019) );
  ANDN U37075 ( .B(n36810), .A(n37409), .Z(n37408) );
  XNOR U37076 ( .A(n37410), .B(n37411), .Z(n32031) );
  XOR U37077 ( .A(n33304), .B(n37412), .Z(n37406) );
  XOR U37078 ( .A(n29733), .B(n31129), .Z(n37412) );
  XNOR U37079 ( .A(n37413), .B(n36529), .Z(n31129) );
  ANDN U37080 ( .B(n36812), .A(n36813), .Z(n37413) );
  XOR U37081 ( .A(n37414), .B(n35738), .Z(n29733) );
  AND U37082 ( .A(n36816), .B(n36817), .Z(n37414) );
  XNOR U37083 ( .A(n37415), .B(n35746), .Z(n33304) );
  XOR U37084 ( .A(n33808), .B(n32216), .Z(n27529) );
  IV U37085 ( .A(n28769), .Z(n32216) );
  XOR U37086 ( .A(n35921), .B(n34167), .Z(n28769) );
  XNOR U37087 ( .A(n37416), .B(n37417), .Z(n34167) );
  XNOR U37088 ( .A(n28988), .B(n32677), .Z(n37417) );
  XNOR U37089 ( .A(n37418), .B(n33279), .Z(n32677) );
  AND U37090 ( .A(n35226), .B(n33280), .Z(n37418) );
  XNOR U37091 ( .A(n37419), .B(n37420), .Z(n33280) );
  XNOR U37092 ( .A(n37421), .B(n37376), .Z(n28988) );
  IV U37093 ( .A(n37374), .Z(n37376) );
  XNOR U37094 ( .A(n37422), .B(n35619), .Z(n37374) );
  ANDN U37095 ( .B(n33813), .A(n33814), .Z(n37421) );
  XNOR U37096 ( .A(n35933), .B(n37423), .Z(n33813) );
  XOR U37097 ( .A(n30033), .B(n37424), .Z(n37416) );
  XNOR U37098 ( .A(n31988), .B(n32244), .Z(n37424) );
  XNOR U37099 ( .A(n37425), .B(n33289), .Z(n32244) );
  XOR U37100 ( .A(n37426), .B(n37427), .Z(n33289) );
  ANDN U37101 ( .B(n33290), .A(n36035), .Z(n37425) );
  XOR U37102 ( .A(n37428), .B(n37429), .Z(n33290) );
  XNOR U37103 ( .A(n37430), .B(n33285), .Z(n31988) );
  IV U37104 ( .A(n37371), .Z(n33285) );
  XOR U37105 ( .A(n37431), .B(n37432), .Z(n37371) );
  AND U37106 ( .A(n33811), .B(n33286), .Z(n37430) );
  XNOR U37107 ( .A(n37433), .B(n37434), .Z(n33286) );
  XNOR U37108 ( .A(n37435), .B(n33275), .Z(n30033) );
  IV U37109 ( .A(n37367), .Z(n33275) );
  XOR U37110 ( .A(n37436), .B(n37437), .Z(n37367) );
  ANDN U37111 ( .B(n33276), .A(n37438), .Z(n37435) );
  XOR U37112 ( .A(n37439), .B(n37440), .Z(n35921) );
  XNOR U37113 ( .A(n34218), .B(n33530), .Z(n37440) );
  XOR U37114 ( .A(n37441), .B(n34946), .Z(n33530) );
  XOR U37115 ( .A(n37443), .B(n34938), .Z(n34218) );
  XOR U37116 ( .A(n37015), .B(n37444), .Z(n34938) );
  ANDN U37117 ( .B(n37445), .A(n37446), .Z(n37443) );
  XNOR U37118 ( .A(n31819), .B(n37447), .Z(n37439) );
  XOR U37119 ( .A(n32597), .B(n34904), .Z(n37447) );
  XOR U37120 ( .A(n37448), .B(n36692), .Z(n34904) );
  XOR U37121 ( .A(n37449), .B(n37450), .Z(n36692) );
  AND U37122 ( .A(n37451), .B(n36693), .Z(n37448) );
  XOR U37123 ( .A(n37452), .B(n34943), .Z(n32597) );
  ANDN U37124 ( .B(n34942), .A(n37453), .Z(n37452) );
  XOR U37125 ( .A(n37454), .B(n37361), .Z(n31819) );
  IV U37126 ( .A(n34933), .Z(n37361) );
  XNOR U37127 ( .A(n37455), .B(n37176), .Z(n34933) );
  ANDN U37128 ( .B(n34934), .A(n37456), .Z(n37454) );
  XNOR U37129 ( .A(n37457), .B(n33276), .Z(n33808) );
  XOR U37130 ( .A(n37458), .B(n37176), .Z(n33276) );
  NOR U37131 ( .A(n37459), .B(n37366), .Z(n37457) );
  XNOR U37132 ( .A(n37460), .B(n27815), .Z(n21822) );
  XOR U37133 ( .A(n32308), .B(n35874), .Z(n27815) );
  XNOR U37134 ( .A(n37461), .B(n37462), .Z(n35874) );
  ANDN U37135 ( .B(n37463), .A(n37464), .Z(n37461) );
  IV U37136 ( .A(n37465), .Z(n32308) );
  ANDN U37137 ( .B(n27952), .A(n27814), .Z(n37460) );
  XOR U37138 ( .A(n37126), .B(n30654), .Z(n27814) );
  IV U37139 ( .A(n29095), .Z(n30654) );
  XOR U37140 ( .A(n34429), .B(n37466), .Z(n29095) );
  XOR U37141 ( .A(n37467), .B(n37468), .Z(n34429) );
  XNOR U37142 ( .A(n29737), .B(n33363), .Z(n37468) );
  XNOR U37143 ( .A(n37469), .B(n37470), .Z(n33363) );
  XOR U37144 ( .A(n37471), .B(n37472), .Z(n37133) );
  XOR U37145 ( .A(n37473), .B(n37474), .Z(n29737) );
  ANDN U37146 ( .B(n37128), .A(n36735), .Z(n37473) );
  XOR U37147 ( .A(n37475), .B(n37055), .Z(n36735) );
  XNOR U37148 ( .A(n32448), .B(n37476), .Z(n37467) );
  XOR U37149 ( .A(n31846), .B(n32493), .Z(n37476) );
  XOR U37150 ( .A(n37477), .B(n37478), .Z(n32493) );
  ANDN U37151 ( .B(n37138), .A(n36722), .Z(n37477) );
  XOR U37152 ( .A(n37479), .B(n37480), .Z(n36722) );
  XOR U37153 ( .A(n37481), .B(n37482), .Z(n31846) );
  ANDN U37154 ( .B(n36727), .A(n37483), .Z(n37481) );
  XOR U37155 ( .A(n37484), .B(n37485), .Z(n32448) );
  ANDN U37156 ( .B(n37135), .A(n36731), .Z(n37484) );
  IV U37157 ( .A(n37136), .Z(n36731) );
  XOR U37158 ( .A(n37486), .B(n34368), .Z(n37136) );
  NOR U37159 ( .A(n36729), .B(n36727), .Z(n37487) );
  XOR U37160 ( .A(n35943), .B(n37488), .Z(n36727) );
  XNOR U37161 ( .A(n30364), .B(n37254), .Z(n27952) );
  XOR U37162 ( .A(n37489), .B(n34706), .Z(n37254) );
  ANDN U37163 ( .B(n35167), .A(n34457), .Z(n37489) );
  XOR U37164 ( .A(n37490), .B(n37491), .Z(n34457) );
  IV U37165 ( .A(n31700), .Z(n30364) );
  XNOR U37166 ( .A(n36342), .B(n37492), .Z(n31700) );
  XOR U37167 ( .A(n37493), .B(n37494), .Z(n36342) );
  XNOR U37168 ( .A(n33533), .B(n34321), .Z(n37494) );
  XNOR U37169 ( .A(n37495), .B(n34454), .Z(n34321) );
  XOR U37170 ( .A(n37496), .B(n37497), .Z(n34454) );
  XNOR U37171 ( .A(n37498), .B(n36955), .Z(n35163) );
  XOR U37172 ( .A(n37499), .B(n37500), .Z(n34696) );
  XOR U37173 ( .A(n37501), .B(n34701), .Z(n33533) );
  XOR U37174 ( .A(n37502), .B(n37187), .Z(n34701) );
  ANDN U37175 ( .B(n37261), .A(n34700), .Z(n37501) );
  XOR U37176 ( .A(n37503), .B(n37504), .Z(n34700) );
  XOR U37177 ( .A(n37148), .B(n37505), .Z(n37261) );
  XOR U37178 ( .A(n32795), .B(n37506), .Z(n37493) );
  XOR U37179 ( .A(n31447), .B(n34689), .Z(n37506) );
  XOR U37180 ( .A(n37507), .B(n34462), .Z(n34689) );
  XOR U37181 ( .A(n37508), .B(n37014), .Z(n34462) );
  XOR U37182 ( .A(n37509), .B(n37510), .Z(n34694) );
  XOR U37183 ( .A(n37511), .B(n37512), .Z(n35153) );
  XNOR U37184 ( .A(n37513), .B(n34458), .Z(n31447) );
  IV U37185 ( .A(n34705), .Z(n34458) );
  XOR U37186 ( .A(n37514), .B(n37515), .Z(n34705) );
  ANDN U37187 ( .B(n34706), .A(n35167), .Z(n37513) );
  XOR U37188 ( .A(n37516), .B(n37517), .Z(n35167) );
  XNOR U37189 ( .A(n37518), .B(n35519), .Z(n34706) );
  XNOR U37190 ( .A(n37519), .B(n34449), .Z(n32795) );
  XOR U37191 ( .A(n37520), .B(n37521), .Z(n34449) );
  ANDN U37192 ( .B(n35157), .A(n37256), .Z(n37519) );
  IV U37193 ( .A(n34703), .Z(n37256) );
  XOR U37194 ( .A(n37522), .B(n37523), .Z(n34703) );
  XNOR U37195 ( .A(n37524), .B(n37525), .Z(n35157) );
  XOR U37196 ( .A(n25962), .B(n37526), .Z(n37380) );
  XNOR U37197 ( .A(n25597), .B(n27797), .Z(n37526) );
  XNOR U37198 ( .A(n37527), .B(n32520), .Z(n27797) );
  XNOR U37199 ( .A(n35119), .B(n31584), .Z(n32520) );
  XNOR U37200 ( .A(n37528), .B(n37529), .Z(n35228) );
  XOR U37201 ( .A(n35397), .B(n37530), .Z(n37529) );
  XNOR U37202 ( .A(n37531), .B(n37532), .Z(n35397) );
  XNOR U37203 ( .A(n4687), .B(n37533), .Z(n37532) );
  NANDN U37204 ( .A(n35245), .B(n35246), .Z(n37533) );
  XOR U37205 ( .A(n37534), .B(n37535), .Z(n35246) );
  XNOR U37206 ( .A(n32822), .B(n37536), .Z(n37528) );
  XNOR U37207 ( .A(n30661), .B(n30026), .Z(n37536) );
  XOR U37208 ( .A(n37537), .B(n36305), .Z(n30026) );
  ANDN U37209 ( .B(n35130), .A(n35131), .Z(n37537) );
  XOR U37210 ( .A(n37538), .B(n35598), .Z(n35131) );
  XNOR U37211 ( .A(n37539), .B(n36309), .Z(n30661) );
  XOR U37212 ( .A(n37540), .B(n36717), .Z(n35135) );
  XOR U37213 ( .A(n37541), .B(n36313), .Z(n32822) );
  ANDN U37214 ( .B(n35140), .A(n35142), .Z(n37541) );
  XOR U37215 ( .A(n37542), .B(n37543), .Z(n35142) );
  XOR U37216 ( .A(n37545), .B(n34048), .Z(n35119) );
  IV U37217 ( .A(n37546), .Z(n34048) );
  ANDN U37218 ( .B(n37547), .A(n36292), .Z(n37545) );
  IV U37219 ( .A(n37548), .Z(n36292) );
  AND U37220 ( .A(n27521), .B(n27522), .Z(n37527) );
  XNOR U37221 ( .A(n31642), .B(n37549), .Z(n27522) );
  XOR U37222 ( .A(n34880), .B(n35049), .Z(n31642) );
  XOR U37223 ( .A(n37550), .B(n37551), .Z(n35049) );
  XOR U37224 ( .A(n36241), .B(n37552), .Z(n37551) );
  XNOR U37225 ( .A(n37553), .B(n37554), .Z(n36241) );
  XOR U37226 ( .A(n31470), .B(n37557), .Z(n37550) );
  XNOR U37227 ( .A(n32190), .B(n36175), .Z(n37557) );
  XOR U37228 ( .A(n37558), .B(n35211), .Z(n36175) );
  XNOR U37229 ( .A(n37561), .B(n35207), .Z(n32190) );
  ANDN U37230 ( .B(n37562), .A(n37563), .Z(n37561) );
  XNOR U37231 ( .A(n37564), .B(n35197), .Z(n31470) );
  ANDN U37232 ( .B(n37565), .A(n37566), .Z(n37564) );
  XOR U37233 ( .A(n37567), .B(n37568), .Z(n34880) );
  XOR U37234 ( .A(n33357), .B(n31251), .Z(n37568) );
  XOR U37235 ( .A(n37569), .B(n37570), .Z(n31251) );
  XNOR U37236 ( .A(n37572), .B(n37573), .Z(n33357) );
  ANDN U37237 ( .B(n37574), .A(n35716), .Z(n37572) );
  XOR U37238 ( .A(n37575), .B(n37576), .Z(n37567) );
  XNOR U37239 ( .A(n30229), .B(n33025), .Z(n37576) );
  XNOR U37240 ( .A(n37577), .B(n37578), .Z(n33025) );
  ANDN U37241 ( .B(n35722), .A(n37579), .Z(n37577) );
  XOR U37242 ( .A(n37580), .B(n37581), .Z(n30229) );
  NOR U37243 ( .A(n37582), .B(n37583), .Z(n37580) );
  XNOR U37244 ( .A(n35652), .B(n35916), .Z(n27521) );
  IV U37245 ( .A(n31632), .Z(n35916) );
  XOR U37246 ( .A(n37584), .B(n37585), .Z(n35652) );
  ANDN U37247 ( .B(n35238), .A(n37586), .Z(n37584) );
  XNOR U37248 ( .A(n37587), .B(n27822), .Z(n25597) );
  XNOR U37249 ( .A(n37588), .B(n31127), .Z(n27822) );
  XNOR U37250 ( .A(n37589), .B(n37590), .Z(n32534) );
  XOR U37251 ( .A(n32418), .B(n29397), .Z(n37590) );
  XNOR U37252 ( .A(n37591), .B(n32432), .Z(n29397) );
  XNOR U37253 ( .A(n37592), .B(n37593), .Z(n32432) );
  AND U37254 ( .A(n32433), .B(n37594), .Z(n37591) );
  XNOR U37255 ( .A(n37595), .B(n32639), .Z(n32418) );
  XNOR U37256 ( .A(n37596), .B(n36359), .Z(n32639) );
  ANDN U37257 ( .B(n37597), .A(n32638), .Z(n37595) );
  IV U37258 ( .A(n37598), .Z(n32638) );
  XNOR U37259 ( .A(n31104), .B(n37599), .Z(n37589) );
  XOR U37260 ( .A(n31408), .B(n32318), .Z(n37599) );
  XNOR U37261 ( .A(n37600), .B(n32426), .Z(n32318) );
  XOR U37262 ( .A(n37601), .B(n37602), .Z(n32426) );
  ANDN U37263 ( .B(n37603), .A(n32425), .Z(n37600) );
  IV U37264 ( .A(n37604), .Z(n32425) );
  XOR U37265 ( .A(n37605), .B(n32858), .Z(n31408) );
  XOR U37266 ( .A(n37606), .B(n35778), .Z(n32858) );
  NOR U37267 ( .A(n32857), .B(n37607), .Z(n37605) );
  XNOR U37268 ( .A(n37608), .B(n33119), .Z(n31104) );
  XOR U37269 ( .A(n37609), .B(n37610), .Z(n33119) );
  XNOR U37270 ( .A(n37612), .B(n37613), .Z(n34529) );
  XNOR U37271 ( .A(n29267), .B(n31031), .Z(n37613) );
  XOR U37272 ( .A(n37614), .B(n33115), .Z(n31031) );
  XNOR U37273 ( .A(n37615), .B(n36970), .Z(n33115) );
  ANDN U37274 ( .B(n35969), .A(n37616), .Z(n37614) );
  XNOR U37275 ( .A(n37617), .B(n35972), .Z(n29267) );
  XOR U37276 ( .A(n37479), .B(n37618), .Z(n35972) );
  ANDN U37277 ( .B(n36990), .A(n37619), .Z(n37617) );
  XOR U37278 ( .A(n35956), .B(n37620), .Z(n37612) );
  XOR U37279 ( .A(n32746), .B(n32835), .Z(n37620) );
  XOR U37280 ( .A(n37621), .B(n33111), .Z(n32835) );
  XNOR U37281 ( .A(n37622), .B(n36316), .Z(n33111) );
  IV U37282 ( .A(n37623), .Z(n36316) );
  AND U37283 ( .A(n35967), .B(n36974), .Z(n37621) );
  XNOR U37284 ( .A(n37624), .B(n33106), .Z(n32746) );
  XOR U37285 ( .A(n37625), .B(n37626), .Z(n33106) );
  ANDN U37286 ( .B(n35964), .A(n37627), .Z(n37624) );
  XOR U37287 ( .A(n37628), .B(n35215), .Z(n35956) );
  XOR U37288 ( .A(n37629), .B(n37630), .Z(n35215) );
  AND U37289 ( .A(n27519), .B(n27517), .Z(n37587) );
  XOR U37290 ( .A(n37631), .B(n33952), .Z(n27517) );
  IV U37291 ( .A(n31880), .Z(n33952) );
  XNOR U37292 ( .A(n35691), .B(n33802), .Z(n31880) );
  XNOR U37293 ( .A(n37632), .B(n37633), .Z(n33802) );
  XOR U37294 ( .A(n35919), .B(n30927), .Z(n37633) );
  XOR U37295 ( .A(n37634), .B(n34942), .Z(n30927) );
  XNOR U37296 ( .A(n37635), .B(n37636), .Z(n34942) );
  ANDN U37297 ( .B(n37453), .A(n37637), .Z(n37634) );
  XNOR U37298 ( .A(n37638), .B(n34934), .Z(n35919) );
  XNOR U37299 ( .A(n37639), .B(n37640), .Z(n34934) );
  XOR U37300 ( .A(n33840), .B(n37641), .Z(n37632) );
  XNOR U37301 ( .A(n31372), .B(n31016), .Z(n37641) );
  XOR U37302 ( .A(n37642), .B(n37446), .Z(n31016) );
  IV U37303 ( .A(n34939), .Z(n37446) );
  XOR U37304 ( .A(n37643), .B(n35619), .Z(n34939) );
  ANDN U37305 ( .B(n37358), .A(n37445), .Z(n37642) );
  XNOR U37306 ( .A(n37644), .B(n36693), .Z(n31372) );
  XNOR U37307 ( .A(n37645), .B(n37646), .Z(n36693) );
  NOR U37308 ( .A(n37356), .B(n37451), .Z(n37644) );
  XNOR U37309 ( .A(n37647), .B(n34947), .Z(n33840) );
  XOR U37310 ( .A(n35943), .B(n37648), .Z(n34947) );
  ANDN U37311 ( .B(n37649), .A(n37442), .Z(n37647) );
  IV U37312 ( .A(n37650), .Z(n37442) );
  XOR U37313 ( .A(n37651), .B(n37652), .Z(n35691) );
  XOR U37314 ( .A(n37653), .B(n36524), .Z(n37652) );
  XOR U37315 ( .A(n37654), .B(n34910), .Z(n36524) );
  ANDN U37316 ( .B(n37655), .A(n37656), .Z(n37654) );
  XOR U37317 ( .A(n31392), .B(n37657), .Z(n37651) );
  XOR U37318 ( .A(n30797), .B(n32874), .Z(n37657) );
  XNOR U37319 ( .A(n37658), .B(n34926), .Z(n32874) );
  NOR U37320 ( .A(n36689), .B(n37659), .Z(n37658) );
  XOR U37321 ( .A(n37660), .B(n34913), .Z(n30797) );
  NOR U37322 ( .A(n37661), .B(n36681), .Z(n37660) );
  XNOR U37323 ( .A(n37662), .B(n34919), .Z(n31392) );
  ANDN U37324 ( .B(n36687), .A(n37663), .Z(n37662) );
  XOR U37325 ( .A(n33967), .B(n27942), .Z(n27519) );
  XOR U37326 ( .A(n34485), .B(n34363), .Z(n27942) );
  XNOR U37327 ( .A(n37664), .B(n37665), .Z(n34363) );
  XNOR U37328 ( .A(n29073), .B(n32039), .Z(n37665) );
  XNOR U37329 ( .A(n37666), .B(n35333), .Z(n32039) );
  XOR U37330 ( .A(n36987), .B(n37667), .Z(n35333) );
  ANDN U37331 ( .B(n35789), .A(n35326), .Z(n37666) );
  IV U37332 ( .A(n37668), .Z(n35326) );
  XOR U37333 ( .A(n37669), .B(n34849), .Z(n29073) );
  ANDN U37334 ( .B(n33974), .A(n33975), .Z(n37669) );
  XNOR U37335 ( .A(n37671), .B(n36434), .Z(n33975) );
  XOR U37336 ( .A(n37672), .B(n37673), .Z(n33974) );
  XNOR U37337 ( .A(n32012), .B(n37674), .Z(n37664) );
  XNOR U37338 ( .A(n35765), .B(n32731), .Z(n37674) );
  XOR U37339 ( .A(n37675), .B(n34852), .Z(n32731) );
  XOR U37340 ( .A(n37676), .B(n35929), .Z(n34852) );
  ANDN U37341 ( .B(n33978), .A(n33980), .Z(n37675) );
  XOR U37342 ( .A(n37677), .B(n37678), .Z(n33980) );
  XOR U37343 ( .A(n37679), .B(n37680), .Z(n33978) );
  XOR U37344 ( .A(n37681), .B(n34840), .Z(n35765) );
  XNOR U37345 ( .A(n37682), .B(n37683), .Z(n34840) );
  ANDN U37346 ( .B(n33969), .A(n33971), .Z(n37681) );
  XOR U37347 ( .A(n37684), .B(n37685), .Z(n33971) );
  XOR U37348 ( .A(n37686), .B(n37687), .Z(n33969) );
  XOR U37349 ( .A(n37688), .B(n34845), .Z(n32012) );
  XNOR U37350 ( .A(n37689), .B(n35082), .Z(n34845) );
  ANDN U37351 ( .B(n33982), .A(n33983), .Z(n37688) );
  XOR U37352 ( .A(n37690), .B(n37691), .Z(n33983) );
  XOR U37353 ( .A(n37692), .B(n37197), .Z(n33982) );
  XOR U37354 ( .A(n37693), .B(n37694), .Z(n34485) );
  XNOR U37355 ( .A(n33729), .B(n31249), .Z(n37694) );
  XOR U37356 ( .A(n37695), .B(n34823), .Z(n31249) );
  XOR U37357 ( .A(n37102), .B(n37696), .Z(n34823) );
  IV U37358 ( .A(n37314), .Z(n37102) );
  ANDN U37359 ( .B(n34660), .A(n34662), .Z(n37695) );
  XOR U37360 ( .A(n37697), .B(n37197), .Z(n34662) );
  XNOR U37361 ( .A(n37698), .B(n37699), .Z(n34660) );
  XNOR U37362 ( .A(n37700), .B(n34831), .Z(n33729) );
  XNOR U37363 ( .A(n37701), .B(n35619), .Z(n34831) );
  ANDN U37364 ( .B(n34643), .A(n34644), .Z(n37700) );
  XNOR U37365 ( .A(n36513), .B(n37702), .Z(n34644) );
  XNOR U37366 ( .A(n37703), .B(n35630), .Z(n34643) );
  XOR U37367 ( .A(n31174), .B(n37704), .Z(n37693) );
  XOR U37368 ( .A(n31977), .B(n30989), .Z(n37704) );
  XOR U37369 ( .A(n37705), .B(n34835), .Z(n30989) );
  IV U37370 ( .A(n35774), .Z(n34835) );
  XOR U37371 ( .A(n37706), .B(n37707), .Z(n35774) );
  ANDN U37372 ( .B(n34647), .A(n35299), .Z(n37705) );
  IV U37373 ( .A(n34649), .Z(n35299) );
  XOR U37374 ( .A(n37708), .B(n36212), .Z(n34649) );
  XOR U37375 ( .A(n37709), .B(n37710), .Z(n34647) );
  XNOR U37376 ( .A(n37711), .B(n34828), .Z(n31977) );
  XOR U37377 ( .A(n37712), .B(n35611), .Z(n34828) );
  ANDN U37378 ( .B(n34656), .A(n34657), .Z(n37711) );
  XOR U37379 ( .A(n37713), .B(n37714), .Z(n34657) );
  XNOR U37380 ( .A(n37715), .B(n37716), .Z(n34656) );
  XOR U37381 ( .A(n37717), .B(n34821), .Z(n31174) );
  XOR U37382 ( .A(n37718), .B(n37719), .Z(n34821) );
  ANDN U37383 ( .B(n34652), .A(n34653), .Z(n37717) );
  XNOR U37384 ( .A(n37720), .B(n37721), .Z(n34653) );
  XNOR U37385 ( .A(n37722), .B(n35938), .Z(n34652) );
  XNOR U37386 ( .A(n37723), .B(n35789), .Z(n33967) );
  XNOR U37387 ( .A(n37724), .B(n37725), .Z(n35789) );
  ANDN U37388 ( .B(n35327), .A(n37668), .Z(n37723) );
  XOR U37389 ( .A(n37726), .B(n37727), .Z(n37668) );
  XOR U37390 ( .A(n37718), .B(n37728), .Z(n35327) );
  XNOR U37391 ( .A(n37729), .B(n27819), .Z(n25962) );
  XNOR U37392 ( .A(n35202), .B(n30554), .Z(n27819) );
  XNOR U37393 ( .A(n35711), .B(n36863), .Z(n30554) );
  XNOR U37394 ( .A(n37730), .B(n37731), .Z(n36863) );
  XNOR U37395 ( .A(n28429), .B(n37732), .Z(n37731) );
  XOR U37396 ( .A(n37733), .B(n35067), .Z(n28429) );
  ANDN U37397 ( .B(n35567), .A(n37734), .Z(n37733) );
  XOR U37398 ( .A(n37735), .B(n37736), .Z(n37730) );
  XOR U37399 ( .A(n31957), .B(n33294), .Z(n37736) );
  XNOR U37400 ( .A(n37737), .B(n35055), .Z(n33294) );
  ANDN U37401 ( .B(n36886), .A(n37738), .Z(n37737) );
  XOR U37402 ( .A(n37739), .B(n35072), .Z(n31957) );
  XOR U37403 ( .A(n37740), .B(n37741), .Z(n35711) );
  XOR U37404 ( .A(n30136), .B(n32685), .Z(n37741) );
  XNOR U37405 ( .A(n37742), .B(n37559), .Z(n32685) );
  ANDN U37406 ( .B(n35209), .A(n37743), .Z(n37742) );
  XOR U37407 ( .A(n37744), .B(n37566), .Z(n30136) );
  XNOR U37408 ( .A(n35499), .B(n37745), .Z(n37740) );
  XNOR U37409 ( .A(n28880), .B(n32868), .Z(n37745) );
  XOR U37410 ( .A(n37746), .B(n37563), .Z(n32868) );
  ANDN U37411 ( .B(n35205), .A(n35206), .Z(n37746) );
  XNOR U37412 ( .A(n37747), .B(n37555), .Z(n28880) );
  AND U37413 ( .A(n37748), .B(n37749), .Z(n37747) );
  XNOR U37414 ( .A(n37750), .B(n37751), .Z(n35499) );
  AND U37415 ( .A(n35200), .B(n35199), .Z(n37750) );
  XNOR U37416 ( .A(n37752), .B(n37748), .Z(n35202) );
  NOR U37417 ( .A(n37749), .B(n37554), .Z(n37752) );
  XOR U37418 ( .A(n34665), .B(n37753), .Z(n27947) );
  XOR U37419 ( .A(n37754), .B(n37755), .Z(n34665) );
  XNOR U37420 ( .A(n33240), .B(n31984), .Z(n37755) );
  XNOR U37421 ( .A(n37756), .B(n36573), .Z(n31984) );
  NOR U37422 ( .A(n35257), .B(n35258), .Z(n37756) );
  XNOR U37423 ( .A(n37757), .B(n36577), .Z(n33240) );
  ANDN U37424 ( .B(n35263), .A(n35262), .Z(n37757) );
  XOR U37425 ( .A(n35655), .B(n37758), .Z(n37754) );
  XOR U37426 ( .A(n31594), .B(n28795), .Z(n37758) );
  XOR U37427 ( .A(n37759), .B(n36569), .Z(n28795) );
  IV U37428 ( .A(n37760), .Z(n36569) );
  NOR U37429 ( .A(n35270), .B(n35271), .Z(n37759) );
  XNOR U37430 ( .A(n37761), .B(n37762), .Z(n31594) );
  ANDN U37431 ( .B(n35255), .A(n35253), .Z(n37761) );
  XOR U37432 ( .A(n37763), .B(n36566), .Z(n35655) );
  XOR U37433 ( .A(n37764), .B(n37765), .Z(n37212) );
  IV U37434 ( .A(n28565), .Z(n27533) );
  XOR U37435 ( .A(n37767), .B(n34815), .Z(n28565) );
  XOR U37436 ( .A(n37768), .B(n37769), .Z(n26929) );
  XNOR U37437 ( .A(n25511), .B(n24553), .Z(n37769) );
  XOR U37438 ( .A(n37770), .B(n27303), .Z(n24553) );
  XNOR U37439 ( .A(n33213), .B(n33226), .Z(n27303) );
  XNOR U37440 ( .A(n37772), .B(n37773), .Z(n34326) );
  XNOR U37441 ( .A(n27936), .B(n37020), .Z(n37773) );
  XOR U37442 ( .A(n37774), .B(n36791), .Z(n37020) );
  XOR U37443 ( .A(n37775), .B(n37776), .Z(n36791) );
  AND U37444 ( .A(n33156), .B(n33157), .Z(n37774) );
  XNOR U37445 ( .A(n37777), .B(n36308), .Z(n33157) );
  XNOR U37446 ( .A(n37778), .B(n37163), .Z(n33156) );
  XOR U37447 ( .A(n37779), .B(n36795), .Z(n27936) );
  XOR U37448 ( .A(n37449), .B(n37780), .Z(n36795) );
  ANDN U37449 ( .B(n33160), .A(n33161), .Z(n37779) );
  XOR U37450 ( .A(n36413), .B(n37781), .Z(n33161) );
  XNOR U37451 ( .A(n37782), .B(n37783), .Z(n33160) );
  XNOR U37452 ( .A(n32670), .B(n37784), .Z(n37772) );
  XOR U37453 ( .A(n33556), .B(n31013), .Z(n37784) );
  XNOR U37454 ( .A(n37785), .B(n36780), .Z(n31013) );
  XNOR U37455 ( .A(n37786), .B(n37787), .Z(n36780) );
  AND U37456 ( .A(n34325), .B(n34323), .Z(n37785) );
  XNOR U37457 ( .A(n37788), .B(n37789), .Z(n34323) );
  XOR U37458 ( .A(n37790), .B(n37791), .Z(n34325) );
  XNOR U37459 ( .A(n37792), .B(n36788), .Z(n33556) );
  XOR U37460 ( .A(n37793), .B(n35320), .Z(n36788) );
  NOR U37461 ( .A(n33166), .B(n33167), .Z(n37792) );
  XOR U37462 ( .A(n37794), .B(n37795), .Z(n33167) );
  IV U37463 ( .A(n37058), .Z(n33166) );
  XOR U37464 ( .A(n37796), .B(n37797), .Z(n37058) );
  XNOR U37465 ( .A(n37798), .B(n36784), .Z(n32670) );
  XOR U37466 ( .A(n37799), .B(n37800), .Z(n36784) );
  AND U37467 ( .A(n33172), .B(n33170), .Z(n37798) );
  XNOR U37468 ( .A(n37801), .B(n37802), .Z(n33170) );
  XNOR U37469 ( .A(n37803), .B(n37804), .Z(n33172) );
  XOR U37470 ( .A(n37805), .B(n37806), .Z(n33213) );
  ANDN U37471 ( .B(n37807), .A(n37808), .Z(n37805) );
  ANDN U37472 ( .B(n28560), .A(n32814), .Z(n37770) );
  XOR U37473 ( .A(n30536), .B(n34474), .Z(n32814) );
  XNOR U37474 ( .A(n37809), .B(n37248), .Z(n34474) );
  ANDN U37475 ( .B(n35182), .A(n35183), .Z(n37809) );
  IV U37476 ( .A(n32142), .Z(n30536) );
  XNOR U37477 ( .A(n37575), .B(n30230), .Z(n28560) );
  XNOR U37478 ( .A(n37810), .B(n33487), .Z(n30230) );
  XOR U37479 ( .A(n37811), .B(n37812), .Z(n33487) );
  XOR U37480 ( .A(n35190), .B(n29046), .Z(n37812) );
  XOR U37481 ( .A(n37813), .B(n35723), .Z(n29046) );
  ANDN U37482 ( .B(n37578), .A(n37814), .Z(n37813) );
  XNOR U37483 ( .A(n37815), .B(n35717), .Z(n35190) );
  ANDN U37484 ( .B(n37573), .A(n37574), .Z(n37815) );
  XOR U37485 ( .A(n30730), .B(n37816), .Z(n37811) );
  XOR U37486 ( .A(n31705), .B(n32186), .Z(n37816) );
  XNOR U37487 ( .A(n37817), .B(n37818), .Z(n32186) );
  AND U37488 ( .A(n37582), .B(n37581), .Z(n37817) );
  NOR U37489 ( .A(n37571), .B(n37570), .Z(n37819) );
  XNOR U37490 ( .A(n37820), .B(n37821), .Z(n30730) );
  ANDN U37491 ( .B(n37822), .A(n37823), .Z(n37820) );
  XNOR U37492 ( .A(n37824), .B(n37822), .Z(n37575) );
  ANDN U37493 ( .B(n37823), .A(n37825), .Z(n37824) );
  XNOR U37494 ( .A(n37826), .B(n27292), .Z(n25511) );
  XNOR U37495 ( .A(n37827), .B(n34815), .Z(n27292) );
  IV U37496 ( .A(n31001), .Z(n34815) );
  ANDN U37497 ( .B(n28549), .A(n32821), .Z(n37826) );
  XOR U37498 ( .A(n35388), .B(n32313), .Z(n32821) );
  IV U37499 ( .A(n29020), .Z(n32313) );
  XOR U37500 ( .A(n34397), .B(n34796), .Z(n29020) );
  XNOR U37501 ( .A(n37830), .B(n37831), .Z(n34796) );
  XOR U37502 ( .A(n33909), .B(n29939), .Z(n37831) );
  XNOR U37503 ( .A(n37832), .B(n33498), .Z(n29939) );
  IV U37504 ( .A(n33924), .Z(n33498) );
  XOR U37505 ( .A(n37833), .B(n37834), .Z(n33924) );
  NOR U37506 ( .A(n32659), .B(n33923), .Z(n37832) );
  XNOR U37507 ( .A(n37835), .B(n37437), .Z(n33923) );
  XNOR U37508 ( .A(n37836), .B(n37837), .Z(n32659) );
  XNOR U37509 ( .A(n37838), .B(n33500), .Z(n33909) );
  XOR U37510 ( .A(n37839), .B(n36557), .Z(n33500) );
  ANDN U37511 ( .B(n33932), .A(n32655), .Z(n37838) );
  XOR U37512 ( .A(n37840), .B(n37841), .Z(n32655) );
  XOR U37513 ( .A(n37842), .B(n34637), .Z(n33932) );
  XOR U37514 ( .A(n32444), .B(n37843), .Z(n37830) );
  XOR U37515 ( .A(n30868), .B(n31672), .Z(n37843) );
  XNOR U37516 ( .A(n37844), .B(n33505), .Z(n31672) );
  ANDN U37517 ( .B(n33914), .A(n34366), .Z(n37844) );
  XOR U37518 ( .A(n37846), .B(n36701), .Z(n34366) );
  XNOR U37519 ( .A(n37847), .B(n37848), .Z(n33914) );
  XNOR U37520 ( .A(n37849), .B(n33507), .Z(n30868) );
  XOR U37521 ( .A(n37850), .B(n35331), .Z(n33507) );
  IV U37522 ( .A(n37851), .Z(n35331) );
  AND U37523 ( .A(n32672), .B(n33918), .Z(n37849) );
  XOR U37524 ( .A(n37690), .B(n37852), .Z(n33918) );
  XOR U37525 ( .A(n37853), .B(n37854), .Z(n32672) );
  XOR U37526 ( .A(n37855), .B(n33509), .Z(n32444) );
  XOR U37527 ( .A(n37856), .B(n37857), .Z(n33509) );
  NOR U37528 ( .A(n33417), .B(n33928), .Z(n37855) );
  XOR U37529 ( .A(n37858), .B(n37859), .Z(n33928) );
  XNOR U37530 ( .A(n37860), .B(n37267), .Z(n33417) );
  XNOR U37531 ( .A(n37861), .B(n37862), .Z(n34397) );
  XNOR U37532 ( .A(n32259), .B(n32131), .Z(n37862) );
  XNOR U37533 ( .A(n37863), .B(n33867), .Z(n32131) );
  XOR U37534 ( .A(n37864), .B(n36967), .Z(n33867) );
  NOR U37535 ( .A(n35391), .B(n33866), .Z(n37863) );
  XOR U37536 ( .A(n37328), .B(n37865), .Z(n33866) );
  XNOR U37537 ( .A(n37866), .B(n35940), .Z(n35391) );
  XNOR U37538 ( .A(n37867), .B(n33858), .Z(n32259) );
  XNOR U37539 ( .A(n37868), .B(n37869), .Z(n33858) );
  NOR U37540 ( .A(n35386), .B(n33857), .Z(n37867) );
  XNOR U37541 ( .A(n37870), .B(n37871), .Z(n33857) );
  XOR U37542 ( .A(n37872), .B(n36996), .Z(n35386) );
  XNOR U37543 ( .A(n32384), .B(n37873), .Z(n37861) );
  XOR U37544 ( .A(n30518), .B(n30203), .Z(n37873) );
  XNOR U37545 ( .A(n37874), .B(n34005), .Z(n30203) );
  IV U37546 ( .A(n33875), .Z(n34005) );
  XOR U37547 ( .A(n37875), .B(n37876), .Z(n33875) );
  ANDN U37548 ( .B(n36539), .A(n33874), .Z(n37874) );
  XNOR U37549 ( .A(n37877), .B(n33862), .Z(n30518) );
  XOR U37550 ( .A(n34633), .B(n37878), .Z(n33862) );
  ANDN U37551 ( .B(n35393), .A(n33861), .Z(n37877) );
  XNOR U37552 ( .A(n37879), .B(n37880), .Z(n33861) );
  IV U37553 ( .A(n36549), .Z(n35393) );
  XNOR U37554 ( .A(n37881), .B(n37472), .Z(n36549) );
  XNOR U37555 ( .A(n37882), .B(n33870), .Z(n32384) );
  XNOR U37556 ( .A(n37883), .B(n37884), .Z(n33870) );
  ANDN U37557 ( .B(n33871), .A(n35383), .Z(n37882) );
  XNOR U37558 ( .A(n37885), .B(n37854), .Z(n35383) );
  IV U37559 ( .A(n37523), .Z(n37854) );
  XOR U37560 ( .A(n37886), .B(n37887), .Z(n33871) );
  XNOR U37561 ( .A(n37888), .B(n33874), .Z(n35388) );
  XOR U37562 ( .A(n37889), .B(n37837), .Z(n33874) );
  ANDN U37563 ( .B(n34004), .A(n36539), .Z(n37888) );
  XOR U37564 ( .A(n37890), .B(n37891), .Z(n36539) );
  XNOR U37565 ( .A(n37892), .B(n35301), .Z(n34004) );
  XNOR U37566 ( .A(n34989), .B(n29286), .Z(n28549) );
  XNOR U37567 ( .A(n37893), .B(n33890), .Z(n34989) );
  ANDN U37568 ( .B(n37894), .A(n37895), .Z(n37893) );
  XNOR U37569 ( .A(n25269), .B(n37896), .Z(n37768) );
  XNOR U37570 ( .A(n22898), .B(n25136), .Z(n37896) );
  XNOR U37571 ( .A(n37897), .B(n32122), .Z(n25136) );
  IV U37572 ( .A(n27299), .Z(n32122) );
  XOR U37573 ( .A(n37898), .B(n32625), .Z(n27299) );
  XNOR U37574 ( .A(n36000), .B(n33297), .Z(n32625) );
  XOR U37575 ( .A(n37899), .B(n37900), .Z(n33297) );
  XNOR U37576 ( .A(n37901), .B(n33194), .Z(n37900) );
  XOR U37577 ( .A(n37902), .B(n37903), .Z(n33194) );
  ANDN U37578 ( .B(n35282), .A(n34434), .Z(n37902) );
  XNOR U37579 ( .A(n36899), .B(n37904), .Z(n34434) );
  XNOR U37580 ( .A(n34606), .B(n37905), .Z(n37899) );
  XNOR U37581 ( .A(n32803), .B(n33185), .Z(n37905) );
  XNOR U37582 ( .A(n37906), .B(n37907), .Z(n33185) );
  ANDN U37583 ( .B(n33725), .A(n35279), .Z(n37906) );
  XNOR U37584 ( .A(n37908), .B(n37909), .Z(n33725) );
  XNOR U37585 ( .A(n37910), .B(n37911), .Z(n32803) );
  ANDN U37586 ( .B(n35284), .A(n33587), .Z(n37910) );
  XNOR U37587 ( .A(n37912), .B(n37913), .Z(n33587) );
  XNOR U37588 ( .A(n37914), .B(n37915), .Z(n34606) );
  NOR U37589 ( .A(n35286), .B(n35287), .Z(n37914) );
  XNOR U37590 ( .A(n35604), .B(n37916), .Z(n35287) );
  XOR U37591 ( .A(n37917), .B(n37918), .Z(n36000) );
  XNOR U37592 ( .A(n33522), .B(n36182), .Z(n37918) );
  XNOR U37593 ( .A(n37919), .B(n37313), .Z(n36182) );
  IV U37594 ( .A(n36197), .Z(n37313) );
  XOR U37595 ( .A(n36303), .B(n37920), .Z(n36197) );
  ANDN U37596 ( .B(n37921), .A(n33580), .Z(n37919) );
  XOR U37597 ( .A(n37922), .B(n37305), .Z(n33522) );
  XOR U37598 ( .A(n36356), .B(n37923), .Z(n37305) );
  NOR U37599 ( .A(n37924), .B(n33563), .Z(n37922) );
  XNOR U37600 ( .A(n31177), .B(n37925), .Z(n37917) );
  XOR U37601 ( .A(n31975), .B(n32157), .Z(n37925) );
  XOR U37602 ( .A(n37926), .B(n36189), .Z(n32157) );
  XOR U37603 ( .A(n37927), .B(n37928), .Z(n36189) );
  NOR U37604 ( .A(n33572), .B(n36188), .Z(n37926) );
  XNOR U37605 ( .A(n37929), .B(n36672), .Z(n31975) );
  XOR U37606 ( .A(n37930), .B(n37931), .Z(n36672) );
  AND U37607 ( .A(n33576), .B(n36673), .Z(n37929) );
  XNOR U37608 ( .A(n37932), .B(n36193), .Z(n31177) );
  ANDN U37609 ( .B(n36194), .A(n33567), .Z(n37932) );
  ANDN U37610 ( .B(n32123), .A(n28547), .Z(n37897) );
  XNOR U37611 ( .A(n37934), .B(n28573), .Z(n22898) );
  XOR U37612 ( .A(n37901), .B(n32804), .Z(n28573) );
  XOR U37613 ( .A(n36183), .B(n33486), .Z(n32804) );
  XNOR U37614 ( .A(n37935), .B(n37936), .Z(n33486) );
  XNOR U37615 ( .A(n32867), .B(n30254), .Z(n37936) );
  XNOR U37616 ( .A(n37937), .B(n36220), .Z(n30254) );
  ANDN U37617 ( .B(n34884), .A(n34885), .Z(n37937) );
  XOR U37618 ( .A(n37938), .B(n37939), .Z(n34885) );
  XNOR U37619 ( .A(n37940), .B(n33652), .Z(n32867) );
  ANDN U37620 ( .B(n34898), .A(n34899), .Z(n37940) );
  XNOR U37621 ( .A(n37941), .B(n35792), .Z(n34899) );
  XOR U37622 ( .A(n37942), .B(n37943), .Z(n37935) );
  XOR U37623 ( .A(n32355), .B(n31944), .Z(n37943) );
  XOR U37624 ( .A(n37944), .B(n33657), .Z(n31944) );
  XOR U37625 ( .A(n37945), .B(n35598), .Z(n34893) );
  XOR U37626 ( .A(n37946), .B(n33666), .Z(n32355) );
  ANDN U37627 ( .B(n34888), .A(n34889), .Z(n37946) );
  XOR U37628 ( .A(n37947), .B(n37948), .Z(n34889) );
  XOR U37629 ( .A(n37949), .B(n37950), .Z(n36183) );
  XNOR U37630 ( .A(n31461), .B(n29721), .Z(n37950) );
  XNOR U37631 ( .A(n37951), .B(n33589), .Z(n29721) );
  IV U37632 ( .A(n37952), .Z(n33589) );
  NOR U37633 ( .A(n37911), .B(n35284), .Z(n37951) );
  XOR U37634 ( .A(n37953), .B(n37954), .Z(n35284) );
  XNOR U37635 ( .A(n37955), .B(n35291), .Z(n31461) );
  XOR U37636 ( .A(n37956), .B(n36423), .Z(n35286) );
  XOR U37637 ( .A(n29940), .B(n37957), .Z(n37949) );
  XOR U37638 ( .A(n37958), .B(n32564), .Z(n37957) );
  XNOR U37639 ( .A(n33595), .B(n37959), .Z(n32564) );
  XNOR U37640 ( .A(n11417), .B(n37960), .Z(n37959) );
  OR U37641 ( .A(n37961), .B(n35276), .Z(n37960) );
  XNOR U37642 ( .A(n37962), .B(n34436), .Z(n29940) );
  ANDN U37643 ( .B(n37903), .A(n35282), .Z(n37962) );
  XOR U37644 ( .A(n37963), .B(n37964), .Z(n35282) );
  XNOR U37645 ( .A(n37965), .B(n37961), .Z(n37901) );
  ANDN U37646 ( .B(n35276), .A(n33594), .Z(n37965) );
  IV U37647 ( .A(n35277), .Z(n33594) );
  XOR U37648 ( .A(n37966), .B(n35938), .Z(n35277) );
  XOR U37649 ( .A(n37967), .B(n36939), .Z(n35276) );
  IV U37650 ( .A(n37968), .Z(n36939) );
  ANDN U37651 ( .B(n32107), .A(n32824), .Z(n37934) );
  XNOR U37652 ( .A(n37969), .B(n31376), .Z(n32824) );
  XNOR U37653 ( .A(n33822), .B(n36739), .Z(n31376) );
  XNOR U37654 ( .A(n37970), .B(n37971), .Z(n36739) );
  XOR U37655 ( .A(n32005), .B(n32499), .Z(n37971) );
  XOR U37656 ( .A(n37972), .B(n37973), .Z(n32499) );
  NOR U37657 ( .A(n37974), .B(n37975), .Z(n37972) );
  XNOR U37658 ( .A(n37976), .B(n37463), .Z(n32005) );
  ANDN U37659 ( .B(n37464), .A(n37977), .Z(n37976) );
  XOR U37660 ( .A(n35870), .B(n37978), .Z(n37970) );
  XOR U37661 ( .A(n29294), .B(n32801), .Z(n37978) );
  XNOR U37662 ( .A(n37979), .B(n35877), .Z(n32801) );
  NOR U37663 ( .A(n37980), .B(n35878), .Z(n37979) );
  XNOR U37664 ( .A(n37981), .B(n35883), .Z(n29294) );
  NOR U37665 ( .A(n37982), .B(n37983), .Z(n37981) );
  XNOR U37666 ( .A(n37984), .B(n35888), .Z(n35870) );
  NOR U37667 ( .A(n37985), .B(n35887), .Z(n37984) );
  XOR U37668 ( .A(n37986), .B(n37987), .Z(n33822) );
  XNOR U37669 ( .A(n30174), .B(n33452), .Z(n37987) );
  XNOR U37670 ( .A(n37988), .B(n37989), .Z(n33452) );
  NOR U37671 ( .A(n37990), .B(n37991), .Z(n37988) );
  XNOR U37672 ( .A(n37992), .B(n37993), .Z(n30174) );
  NOR U37673 ( .A(n37994), .B(n37995), .Z(n37992) );
  XOR U37674 ( .A(n33034), .B(n37996), .Z(n37986) );
  XOR U37675 ( .A(n31886), .B(n32967), .Z(n37996) );
  XNOR U37676 ( .A(n37997), .B(n37998), .Z(n32967) );
  ANDN U37677 ( .B(n37999), .A(n38000), .Z(n37997) );
  XNOR U37678 ( .A(n38001), .B(n38002), .Z(n31886) );
  NOR U37679 ( .A(n38003), .B(n38004), .Z(n38001) );
  XNOR U37680 ( .A(n38005), .B(n38006), .Z(n33034) );
  ANDN U37681 ( .B(n38007), .A(n38008), .Z(n38005) );
  XOR U37682 ( .A(n38009), .B(n31123), .Z(n32107) );
  XNOR U37683 ( .A(n33713), .B(n32551), .Z(n31123) );
  XNOR U37684 ( .A(n38010), .B(n38011), .Z(n32551) );
  XOR U37685 ( .A(n31786), .B(n36458), .Z(n38011) );
  XNOR U37686 ( .A(n38012), .B(n36464), .Z(n36458) );
  ANDN U37687 ( .B(n36465), .A(n36878), .Z(n38012) );
  XNOR U37688 ( .A(n38013), .B(n38014), .Z(n31786) );
  NOR U37689 ( .A(n36881), .B(n38015), .Z(n38013) );
  XOR U37690 ( .A(n36338), .B(n38016), .Z(n38010) );
  XOR U37691 ( .A(n31942), .B(n32882), .Z(n38016) );
  XOR U37692 ( .A(n38017), .B(n36477), .Z(n32882) );
  ANDN U37693 ( .B(n36478), .A(n36867), .Z(n38017) );
  XNOR U37694 ( .A(n38018), .B(n36474), .Z(n31942) );
  NOR U37695 ( .A(n36870), .B(n36473), .Z(n38018) );
  XNOR U37696 ( .A(n38019), .B(n36469), .Z(n36338) );
  AND U37697 ( .A(n36470), .B(n36874), .Z(n38019) );
  XOR U37698 ( .A(n38020), .B(n38021), .Z(n33713) );
  XNOR U37699 ( .A(n33407), .B(n31973), .Z(n38021) );
  XNOR U37700 ( .A(n38022), .B(n36492), .Z(n31973) );
  XOR U37701 ( .A(n38023), .B(n38024), .Z(n36049) );
  XNOR U37702 ( .A(n38025), .B(n36484), .Z(n33407) );
  NOR U37703 ( .A(n36067), .B(n36066), .Z(n38025) );
  XOR U37704 ( .A(n38026), .B(n38027), .Z(n36066) );
  XOR U37705 ( .A(n31191), .B(n38028), .Z(n38020) );
  XOR U37706 ( .A(n32760), .B(n33991), .Z(n38028) );
  XNOR U37707 ( .A(n38029), .B(n36488), .Z(n33991) );
  NOR U37708 ( .A(n36489), .B(n36059), .Z(n38029) );
  XOR U37709 ( .A(n38030), .B(n38031), .Z(n36489) );
  XNOR U37710 ( .A(n38032), .B(n37298), .Z(n32760) );
  ANDN U37711 ( .B(n36054), .A(n37297), .Z(n38032) );
  IV U37712 ( .A(n36053), .Z(n37297) );
  XOR U37713 ( .A(n38033), .B(n38034), .Z(n36053) );
  XNOR U37714 ( .A(n38035), .B(n36495), .Z(n31191) );
  XOR U37715 ( .A(n38036), .B(n38037), .Z(n36062) );
  XNOR U37716 ( .A(n38038), .B(n27288), .Z(n25269) );
  XOR U37717 ( .A(n30483), .B(n38039), .Z(n27288) );
  XOR U37718 ( .A(n38040), .B(n38041), .Z(n36499) );
  XOR U37719 ( .A(n30115), .B(n34687), .Z(n38041) );
  XNOR U37720 ( .A(n38042), .B(n33939), .Z(n34687) );
  ANDN U37721 ( .B(n38043), .A(n38044), .Z(n38042) );
  XNOR U37722 ( .A(n38045), .B(n33846), .Z(n30115) );
  ANDN U37723 ( .B(n38046), .A(n38047), .Z(n38045) );
  XOR U37724 ( .A(n30237), .B(n38048), .Z(n38040) );
  XNOR U37725 ( .A(n36323), .B(n32980), .Z(n38048) );
  XOR U37726 ( .A(n38049), .B(n37808), .Z(n32980) );
  ANDN U37727 ( .B(n38050), .A(n38051), .Z(n38049) );
  XNOR U37728 ( .A(n38052), .B(n33229), .Z(n36323) );
  AND U37729 ( .A(n38053), .B(n38054), .Z(n38052) );
  XNOR U37730 ( .A(n38055), .B(n36043), .Z(n30237) );
  ANDN U37731 ( .B(n38056), .A(n38057), .Z(n38055) );
  XNOR U37732 ( .A(n38058), .B(n38059), .Z(n34359) );
  XOR U37733 ( .A(n32530), .B(n32796), .Z(n38059) );
  XNOR U37734 ( .A(n38060), .B(n36749), .Z(n32796) );
  ANDN U37735 ( .B(n38061), .A(n38062), .Z(n38060) );
  XOR U37736 ( .A(n38063), .B(n36758), .Z(n32530) );
  ANDN U37737 ( .B(n38064), .A(n38065), .Z(n38063) );
  XOR U37738 ( .A(n33903), .B(n38066), .Z(n38058) );
  XOR U37739 ( .A(n38067), .B(n33065), .Z(n38066) );
  XNOR U37740 ( .A(n38068), .B(n38069), .Z(n33065) );
  ANDN U37741 ( .B(n38070), .A(n38071), .Z(n38068) );
  XNOR U37742 ( .A(n38072), .B(n36745), .Z(n33903) );
  NOR U37743 ( .A(n38073), .B(n38074), .Z(n38072) );
  ANDN U37744 ( .B(n32115), .A(n28556), .Z(n38038) );
  XOR U37745 ( .A(n37145), .B(n28892), .Z(n28556) );
  XOR U37746 ( .A(n32939), .B(n37466), .Z(n28892) );
  XNOR U37747 ( .A(n38075), .B(n38076), .Z(n37466) );
  XOR U37748 ( .A(n34798), .B(n34395), .Z(n38076) );
  XNOR U37749 ( .A(n38077), .B(n33337), .Z(n34395) );
  XNOR U37750 ( .A(n37857), .B(n38078), .Z(n33337) );
  AND U37751 ( .A(n36703), .B(n34809), .Z(n38077) );
  XNOR U37752 ( .A(n38079), .B(n38080), .Z(n34809) );
  XOR U37753 ( .A(n38081), .B(n38082), .Z(n36703) );
  XNOR U37754 ( .A(n38083), .B(n33340), .Z(n34798) );
  XOR U37755 ( .A(n38084), .B(n37687), .Z(n33340) );
  AND U37756 ( .A(n36712), .B(n34811), .Z(n38083) );
  XOR U37757 ( .A(n38085), .B(n37183), .Z(n34811) );
  XNOR U37758 ( .A(n30307), .B(n38087), .Z(n38075) );
  XNOR U37759 ( .A(n30485), .B(n31171), .Z(n38087) );
  XNOR U37760 ( .A(n38088), .B(n33345), .Z(n31171) );
  XOR U37761 ( .A(n38089), .B(n38090), .Z(n33345) );
  ANDN U37762 ( .B(n36708), .A(n34813), .Z(n38088) );
  XOR U37763 ( .A(n37868), .B(n38091), .Z(n34813) );
  XNOR U37764 ( .A(n38092), .B(n38093), .Z(n36708) );
  XNOR U37765 ( .A(n38094), .B(n33353), .Z(n30485) );
  XNOR U37766 ( .A(n38095), .B(n38096), .Z(n33353) );
  XNOR U37767 ( .A(n38097), .B(n34804), .Z(n30307) );
  IV U37768 ( .A(n33349), .Z(n34804) );
  XOR U37769 ( .A(n38098), .B(n37051), .Z(n33349) );
  ANDN U37770 ( .B(n36715), .A(n34803), .Z(n38097) );
  XNOR U37771 ( .A(n38099), .B(n38100), .Z(n34803) );
  XOR U37772 ( .A(n37503), .B(n38101), .Z(n36715) );
  XOR U37773 ( .A(n38102), .B(n38103), .Z(n32939) );
  XNOR U37774 ( .A(n32881), .B(n31587), .Z(n38103) );
  XOR U37775 ( .A(n38104), .B(n37611), .Z(n31587) );
  NOR U37776 ( .A(n33118), .B(n33250), .Z(n38104) );
  XOR U37777 ( .A(n35799), .B(n38105), .Z(n33118) );
  XOR U37778 ( .A(n38106), .B(n37603), .Z(n32881) );
  NOR U37779 ( .A(n33255), .B(n32424), .Z(n38106) );
  XOR U37780 ( .A(n37216), .B(n38107), .Z(n32424) );
  XOR U37781 ( .A(n30919), .B(n38108), .Z(n38102) );
  XOR U37782 ( .A(n32718), .B(n38109), .Z(n38108) );
  XOR U37783 ( .A(n38110), .B(n37594), .Z(n32718) );
  ANDN U37784 ( .B(n32431), .A(n33248), .Z(n38110) );
  XNOR U37785 ( .A(n38111), .B(n36393), .Z(n32431) );
  XNOR U37786 ( .A(n38112), .B(n37607), .Z(n30919) );
  XNOR U37787 ( .A(n38113), .B(n38114), .Z(n32856) );
  XNOR U37788 ( .A(n38115), .B(n34806), .Z(n37145) );
  XNOR U37789 ( .A(n38116), .B(n37909), .Z(n34806) );
  ANDN U37790 ( .B(n36699), .A(n36698), .Z(n38115) );
  XOR U37791 ( .A(n38117), .B(n38118), .Z(n36698) );
  IV U37792 ( .A(n33352), .Z(n36699) );
  XOR U37793 ( .A(n38119), .B(n38120), .Z(n33352) );
  XNOR U37794 ( .A(n36659), .B(n29071), .Z(n32115) );
  XNOR U37795 ( .A(n38121), .B(n38122), .Z(n34949) );
  XNOR U37796 ( .A(n32269), .B(n33090), .Z(n38122) );
  XNOR U37797 ( .A(n38123), .B(n36921), .Z(n33090) );
  XNOR U37798 ( .A(n38124), .B(n38125), .Z(n36921) );
  ANDN U37799 ( .B(n36950), .A(n35032), .Z(n38123) );
  XOR U37800 ( .A(n38126), .B(n38127), .Z(n35032) );
  XOR U37801 ( .A(n38128), .B(n37841), .Z(n36950) );
  XOR U37802 ( .A(n38129), .B(n36923), .Z(n32269) );
  XNOR U37803 ( .A(n38130), .B(n36347), .Z(n36923) );
  ANDN U37804 ( .B(n35042), .A(n37184), .Z(n38129) );
  XOR U37805 ( .A(n38131), .B(n38132), .Z(n37184) );
  XNOR U37806 ( .A(n38133), .B(n38134), .Z(n35042) );
  XOR U37807 ( .A(n33055), .B(n38135), .Z(n38121) );
  XOR U37808 ( .A(n32161), .B(n33876), .Z(n38135) );
  XNOR U37809 ( .A(n38136), .B(n36914), .Z(n33876) );
  XOR U37810 ( .A(n38137), .B(n37176), .Z(n36914) );
  NOR U37811 ( .A(n37188), .B(n36959), .Z(n38136) );
  XOR U37812 ( .A(n38138), .B(n37025), .Z(n36959) );
  XOR U37813 ( .A(n38139), .B(n37909), .Z(n37188) );
  XNOR U37814 ( .A(n38140), .B(n36917), .Z(n32161) );
  XNOR U37815 ( .A(n38141), .B(n37472), .Z(n36917) );
  ANDN U37816 ( .B(n35028), .A(n37192), .Z(n38140) );
  XOR U37817 ( .A(n38142), .B(n38143), .Z(n37192) );
  XOR U37818 ( .A(n37890), .B(n38144), .Z(n35028) );
  XNOR U37819 ( .A(n38145), .B(n36926), .Z(n33055) );
  XOR U37820 ( .A(n38146), .B(n38147), .Z(n36926) );
  NOR U37821 ( .A(n36953), .B(n35038), .Z(n38145) );
  XNOR U37822 ( .A(n38148), .B(n38149), .Z(n35038) );
  IV U37823 ( .A(n37198), .Z(n36953) );
  XOR U37824 ( .A(n38150), .B(n38151), .Z(n37198) );
  XNOR U37825 ( .A(n38152), .B(n38153), .Z(n36174) );
  XNOR U37826 ( .A(n33645), .B(n37158), .Z(n38153) );
  XOR U37827 ( .A(n38155), .B(n37027), .Z(n36908) );
  ANDN U37828 ( .B(n35022), .A(n36661), .Z(n38154) );
  XNOR U37829 ( .A(n38156), .B(n34623), .Z(n36661) );
  XOR U37830 ( .A(n38157), .B(n38158), .Z(n35022) );
  XNOR U37831 ( .A(n38159), .B(n36892), .Z(n33645) );
  XOR U37832 ( .A(n38160), .B(n38161), .Z(n36892) );
  NOR U37833 ( .A(n36666), .B(n35005), .Z(n38159) );
  XOR U37834 ( .A(n38162), .B(n38163), .Z(n35005) );
  XOR U37835 ( .A(n38164), .B(n35165), .Z(n36666) );
  IV U37836 ( .A(n36967), .Z(n35165) );
  XOR U37837 ( .A(n32607), .B(n38165), .Z(n38152) );
  XNOR U37838 ( .A(n31193), .B(n30747), .Z(n38165) );
  XNOR U37839 ( .A(n38166), .B(n36901), .Z(n30747) );
  XNOR U37840 ( .A(n38124), .B(n38167), .Z(n36901) );
  NOR U37841 ( .A(n36664), .B(n35014), .Z(n38166) );
  XNOR U37842 ( .A(n38168), .B(n38169), .Z(n35014) );
  XOR U37843 ( .A(n38170), .B(n38171), .Z(n36664) );
  XOR U37844 ( .A(n38172), .B(n37178), .Z(n31193) );
  XOR U37845 ( .A(n38173), .B(n38174), .Z(n37178) );
  ANDN U37846 ( .B(n37177), .A(n35018), .Z(n38172) );
  XNOR U37847 ( .A(n38175), .B(n36896), .Z(n32607) );
  IV U37848 ( .A(n37167), .Z(n36896) );
  XNOR U37849 ( .A(n38176), .B(n38177), .Z(n37167) );
  NOR U37850 ( .A(n36669), .B(n35009), .Z(n38175) );
  XOR U37851 ( .A(n36408), .B(n38178), .Z(n35009) );
  XOR U37852 ( .A(n38179), .B(n33931), .Z(n36669) );
  XOR U37853 ( .A(n38180), .B(n37177), .Z(n36659) );
  XNOR U37854 ( .A(n38181), .B(n38182), .Z(n37177) );
  ANDN U37855 ( .B(n35018), .A(n36903), .Z(n38180) );
  XOR U37856 ( .A(n38183), .B(n38184), .Z(n36903) );
  XOR U37857 ( .A(n38185), .B(n37797), .Z(n35018) );
  XNOR U37858 ( .A(n38186), .B(n32123), .Z(n32812) );
  XNOR U37859 ( .A(n30852), .B(n38187), .Z(n32123) );
  XOR U37860 ( .A(n38188), .B(n34211), .Z(n30852) );
  XOR U37861 ( .A(n38189), .B(n38190), .Z(n34211) );
  XNOR U37862 ( .A(n36426), .B(n33728), .Z(n38190) );
  XNOR U37863 ( .A(n38191), .B(n38192), .Z(n33728) );
  NOR U37864 ( .A(n36602), .B(n35409), .Z(n38191) );
  XNOR U37865 ( .A(n38193), .B(n36599), .Z(n36426) );
  AND U37866 ( .A(n36600), .B(n35404), .Z(n38193) );
  XNOR U37867 ( .A(n36595), .B(n38194), .Z(n38189) );
  XNOR U37868 ( .A(n28461), .B(n31932), .Z(n38194) );
  XOR U37869 ( .A(n38195), .B(n38196), .Z(n31932) );
  ANDN U37870 ( .B(n35413), .A(n36607), .Z(n38195) );
  XNOR U37871 ( .A(n38197), .B(n38198), .Z(n28461) );
  ANDN U37872 ( .B(n38199), .A(n37386), .Z(n38197) );
  XNOR U37873 ( .A(n38200), .B(n36611), .Z(n36595) );
  ANDN U37874 ( .B(n36610), .A(n35417), .Z(n38200) );
  ANDN U37875 ( .B(n28547), .A(n27297), .Z(n38186) );
  XOR U37876 ( .A(n38201), .B(n31268), .Z(n27297) );
  XOR U37877 ( .A(n33670), .B(n35187), .Z(n31268) );
  XNOR U37878 ( .A(n38202), .B(n38203), .Z(n35187) );
  XNOR U37879 ( .A(n34018), .B(n38204), .Z(n38203) );
  XNOR U37880 ( .A(n38205), .B(n38206), .Z(n34018) );
  NOR U37881 ( .A(n34762), .B(n38207), .Z(n38205) );
  XOR U37882 ( .A(n32363), .B(n38208), .Z(n38202) );
  XOR U37883 ( .A(n35748), .B(n38209), .Z(n38208) );
  XNOR U37884 ( .A(n38210), .B(n38211), .Z(n35748) );
  NOR U37885 ( .A(n34752), .B(n38212), .Z(n38210) );
  XNOR U37886 ( .A(n38213), .B(n38214), .Z(n32363) );
  NOR U37887 ( .A(n34756), .B(n38215), .Z(n38213) );
  XOR U37888 ( .A(n38216), .B(n38217), .Z(n33670) );
  XNOR U37889 ( .A(n31688), .B(n31802), .Z(n38217) );
  XOR U37890 ( .A(n38218), .B(n37401), .Z(n31802) );
  ANDN U37891 ( .B(n36113), .A(n36114), .Z(n38218) );
  XOR U37892 ( .A(n38219), .B(n37394), .Z(n31688) );
  NOR U37893 ( .A(n36106), .B(n36105), .Z(n38219) );
  XNOR U37894 ( .A(n27932), .B(n38220), .Z(n38216) );
  XNOR U37895 ( .A(n36796), .B(n29068), .Z(n38220) );
  XOR U37896 ( .A(n38221), .B(n37398), .Z(n29068) );
  NOR U37897 ( .A(n36109), .B(n36110), .Z(n38221) );
  XNOR U37898 ( .A(n38222), .B(n38223), .Z(n36796) );
  NOR U37899 ( .A(n36102), .B(n36100), .Z(n38222) );
  XNOR U37900 ( .A(n38224), .B(n37404), .Z(n27932) );
  ANDN U37901 ( .B(n36097), .A(n36096), .Z(n38224) );
  XOR U37902 ( .A(n35638), .B(n30743), .Z(n28547) );
  XOR U37903 ( .A(n38227), .B(n38228), .Z(n35638) );
  NOR U37904 ( .A(n34205), .B(n34204), .Z(n38227) );
  ANDN U37905 ( .B(n23680), .A(n23679), .Z(n37379) );
  XOR U37906 ( .A(n31436), .B(n23592), .Z(n23679) );
  XOR U37907 ( .A(n38229), .B(n38230), .Z(n26081) );
  XOR U37908 ( .A(n25500), .B(n24784), .Z(n38230) );
  XOR U37909 ( .A(n38231), .B(n27868), .Z(n24784) );
  XOR U37910 ( .A(n32362), .B(n38209), .Z(n27868) );
  XNOR U37911 ( .A(n38232), .B(n38233), .Z(n38209) );
  ANDN U37912 ( .B(n34766), .A(n38234), .Z(n38232) );
  XOR U37913 ( .A(n35443), .B(n30943), .Z(n27766) );
  XOR U37914 ( .A(n38235), .B(n36428), .Z(n30943) );
  XNOR U37915 ( .A(n38236), .B(n38237), .Z(n36428) );
  XOR U37916 ( .A(n31097), .B(n31771), .Z(n38237) );
  XNOR U37917 ( .A(n38238), .B(n34598), .Z(n31771) );
  XOR U37918 ( .A(n38239), .B(n36783), .Z(n34598) );
  ANDN U37919 ( .B(n35672), .A(n38240), .Z(n38238) );
  XNOR U37920 ( .A(n38241), .B(n34594), .Z(n31097) );
  XNOR U37921 ( .A(n38242), .B(n38243), .Z(n34594) );
  AND U37922 ( .A(n35453), .B(n35454), .Z(n38241) );
  XOR U37923 ( .A(n38244), .B(n37152), .Z(n35453) );
  XNOR U37924 ( .A(n35473), .B(n38245), .Z(n38236) );
  XOR U37925 ( .A(n30519), .B(n35661), .Z(n38245) );
  XNOR U37926 ( .A(n38246), .B(n34585), .Z(n35661) );
  XOR U37927 ( .A(n38247), .B(n38248), .Z(n34585) );
  ANDN U37928 ( .B(n35449), .A(n35450), .Z(n38246) );
  IV U37929 ( .A(n38249), .Z(n35450) );
  XOR U37930 ( .A(n38252), .B(n38253), .Z(n34589) );
  NOR U37931 ( .A(n35670), .B(n36593), .Z(n38251) );
  XNOR U37932 ( .A(n38254), .B(n38255), .Z(n35670) );
  XOR U37933 ( .A(n38256), .B(n34581), .Z(n35473) );
  XOR U37934 ( .A(n36941), .B(n38257), .Z(n34581) );
  AND U37935 ( .A(n35447), .B(n35446), .Z(n38256) );
  XNOR U37936 ( .A(n38258), .B(n37089), .Z(n35446) );
  XOR U37937 ( .A(n38259), .B(n35672), .Z(n35443) );
  XOR U37938 ( .A(n38260), .B(n38261), .Z(n35672) );
  XOR U37939 ( .A(n35806), .B(n28736), .Z(n27869) );
  IV U37940 ( .A(n31346), .Z(n28736) );
  XOR U37941 ( .A(n34169), .B(n33477), .Z(n31346) );
  XOR U37942 ( .A(n38262), .B(n38263), .Z(n33477) );
  XOR U37943 ( .A(n28812), .B(n38264), .Z(n38263) );
  XNOR U37944 ( .A(n38265), .B(n36012), .Z(n28812) );
  ANDN U37945 ( .B(n35830), .A(n35829), .Z(n38265) );
  IV U37946 ( .A(n38266), .Z(n35829) );
  XNOR U37947 ( .A(n38267), .B(n38268), .Z(n35830) );
  XOR U37948 ( .A(n33847), .B(n38269), .Z(n38262) );
  XNOR U37949 ( .A(n33819), .B(n34533), .Z(n38269) );
  XNOR U37950 ( .A(n38270), .B(n36014), .Z(n34533) );
  ANDN U37951 ( .B(n35843), .A(n35842), .Z(n38270) );
  XNOR U37952 ( .A(n38271), .B(n38272), .Z(n35843) );
  XNOR U37953 ( .A(n38273), .B(n36018), .Z(n33819) );
  ANDN U37954 ( .B(n35834), .A(n35835), .Z(n38273) );
  IV U37955 ( .A(n36404), .Z(n35835) );
  XOR U37956 ( .A(n38274), .B(n37848), .Z(n36404) );
  XNOR U37957 ( .A(n38275), .B(n36005), .Z(n33847) );
  ANDN U37958 ( .B(n35825), .A(n35826), .Z(n38275) );
  XOR U37959 ( .A(n38276), .B(n38277), .Z(n35826) );
  XOR U37960 ( .A(n38278), .B(n38279), .Z(n34169) );
  XOR U37961 ( .A(n31000), .B(n37827), .Z(n38279) );
  XNOR U37962 ( .A(n38280), .B(n38281), .Z(n37827) );
  ANDN U37963 ( .B(n35813), .A(n35812), .Z(n38280) );
  XOR U37964 ( .A(n38282), .B(n38283), .Z(n35813) );
  XNOR U37965 ( .A(n38284), .B(n35559), .Z(n31000) );
  ANDN U37966 ( .B(n35817), .A(n35816), .Z(n38284) );
  XNOR U37967 ( .A(n38285), .B(n38286), .Z(n35817) );
  XOR U37968 ( .A(n34814), .B(n38287), .Z(n38278) );
  XOR U37969 ( .A(n31702), .B(n37767), .Z(n38287) );
  XOR U37970 ( .A(n38288), .B(n35555), .Z(n37767) );
  ANDN U37971 ( .B(n36396), .A(n38289), .Z(n38288) );
  XOR U37972 ( .A(n38290), .B(n35551), .Z(n31702) );
  XNOR U37973 ( .A(n38291), .B(n38268), .Z(n35809) );
  IV U37974 ( .A(n36783), .Z(n38268) );
  XNOR U37975 ( .A(n38292), .B(n36424), .Z(n34814) );
  IV U37976 ( .A(n38293), .Z(n36424) );
  AND U37977 ( .A(n35819), .B(n35820), .Z(n38292) );
  XOR U37978 ( .A(n38294), .B(n38295), .Z(n35820) );
  NOR U37979 ( .A(n36396), .B(n35553), .Z(n38296) );
  XOR U37980 ( .A(n38297), .B(n38298), .Z(n35553) );
  XOR U37981 ( .A(n38299), .B(n35159), .Z(n36396) );
  XNOR U37982 ( .A(n38300), .B(n27860), .Z(n25500) );
  XNOR U37983 ( .A(n35754), .B(n30959), .Z(n27860) );
  XOR U37984 ( .A(n38301), .B(n38302), .Z(n34179) );
  XNOR U37985 ( .A(n32176), .B(n31983), .Z(n38302) );
  XNOR U37986 ( .A(n38303), .B(n34308), .Z(n31983) );
  XOR U37987 ( .A(n38304), .B(n38305), .Z(n34308) );
  XOR U37988 ( .A(n38306), .B(n38307), .Z(n34309) );
  XOR U37989 ( .A(n38308), .B(n34304), .Z(n32176) );
  XOR U37990 ( .A(n38309), .B(n35627), .Z(n34304) );
  AND U37991 ( .A(n35756), .B(n34303), .Z(n38308) );
  XNOR U37992 ( .A(n38310), .B(n35595), .Z(n34303) );
  XOR U37993 ( .A(n32270), .B(n38311), .Z(n38301) );
  XNOR U37994 ( .A(n33632), .B(n32364), .Z(n38311) );
  XOR U37995 ( .A(n38312), .B(n34317), .Z(n32364) );
  XOR U37996 ( .A(n38313), .B(n37727), .Z(n34317) );
  IV U37997 ( .A(n37710), .Z(n37727) );
  AND U37998 ( .A(n35763), .B(n34316), .Z(n38312) );
  XNOR U37999 ( .A(n38314), .B(n36439), .Z(n34316) );
  XNOR U38000 ( .A(n38315), .B(n34300), .Z(n33632) );
  XNOR U38001 ( .A(n38316), .B(n36545), .Z(n34300) );
  IV U38002 ( .A(n36955), .Z(n36545) );
  ANDN U38003 ( .B(n34299), .A(n35761), .Z(n38315) );
  XNOR U38004 ( .A(n38317), .B(n38318), .Z(n34299) );
  XOR U38005 ( .A(n38319), .B(n34313), .Z(n32270) );
  XOR U38006 ( .A(n38320), .B(n38321), .Z(n34313) );
  ANDN U38007 ( .B(n38322), .A(n34312), .Z(n38319) );
  XOR U38008 ( .A(n38324), .B(n34312), .Z(n35754) );
  XOR U38009 ( .A(n38325), .B(n38326), .Z(n34312) );
  NOR U38010 ( .A(n35489), .B(n38322), .Z(n38324) );
  ANDN U38011 ( .B(n27861), .A(n27774), .Z(n38300) );
  XOR U38012 ( .A(n38327), .B(n31444), .Z(n27774) );
  XOR U38013 ( .A(n34789), .B(n34214), .Z(n31444) );
  XOR U38014 ( .A(n38328), .B(n38329), .Z(n34214) );
  XOR U38015 ( .A(n28874), .B(n34427), .Z(n38329) );
  XOR U38016 ( .A(n38330), .B(n36077), .Z(n34427) );
  NOR U38017 ( .A(n37291), .B(n37292), .Z(n38330) );
  IV U38018 ( .A(n36078), .Z(n37291) );
  XOR U38019 ( .A(n38331), .B(n38332), .Z(n36078) );
  XNOR U38020 ( .A(n38333), .B(n36087), .Z(n28874) );
  ANDN U38021 ( .B(n36088), .A(n37277), .Z(n38333) );
  XNOR U38022 ( .A(n38334), .B(n35598), .Z(n36088) );
  XOR U38023 ( .A(n27928), .B(n38335), .Z(n38328) );
  XOR U38024 ( .A(n32287), .B(n34369), .Z(n38335) );
  XOR U38025 ( .A(n38336), .B(n38337), .Z(n34369) );
  NOR U38026 ( .A(n37286), .B(n37284), .Z(n38336) );
  XNOR U38027 ( .A(n38338), .B(n36083), .Z(n32287) );
  ANDN U38028 ( .B(n36084), .A(n37288), .Z(n38338) );
  XOR U38029 ( .A(n38339), .B(n38340), .Z(n36084) );
  XNOR U38030 ( .A(n38341), .B(n36073), .Z(n27928) );
  ANDN U38031 ( .B(n36074), .A(n37281), .Z(n38341) );
  XOR U38032 ( .A(n38342), .B(n38343), .Z(n36074) );
  XOR U38033 ( .A(n38344), .B(n38345), .Z(n34789) );
  XOR U38034 ( .A(n36045), .B(n33067), .Z(n38345) );
  XOR U38035 ( .A(n38346), .B(n36063), .Z(n33067) );
  XOR U38036 ( .A(n38347), .B(n38118), .Z(n36063) );
  XOR U38037 ( .A(n36054), .B(n38348), .Z(n36045) );
  XOR U38038 ( .A(n38349), .B(n38350), .Z(n38348) );
  NANDN U38039 ( .A(rc_i[0]), .B(n4549), .Z(n38350) );
  ANDN U38040 ( .B(n36055), .A(n37296), .Z(n38349) );
  XOR U38041 ( .A(n38351), .B(n38352), .Z(n36054) );
  XOR U38042 ( .A(n33236), .B(n38353), .Z(n38344) );
  XNOR U38043 ( .A(n32178), .B(n31222), .Z(n38353) );
  XNOR U38044 ( .A(n38354), .B(n36051), .Z(n31222) );
  XOR U38045 ( .A(n38355), .B(n35579), .Z(n36051) );
  XNOR U38046 ( .A(n38356), .B(n36059), .Z(n32178) );
  XOR U38047 ( .A(n38357), .B(n37081), .Z(n36059) );
  XNOR U38048 ( .A(n38358), .B(n36067), .Z(n33236) );
  XOR U38049 ( .A(n38359), .B(n38360), .Z(n36067) );
  AND U38050 ( .A(n36483), .B(n36068), .Z(n38358) );
  XOR U38051 ( .A(n34023), .B(n31687), .Z(n27861) );
  XNOR U38052 ( .A(n33454), .B(n32527), .Z(n31687) );
  XNOR U38053 ( .A(n38361), .B(n38362), .Z(n32527) );
  XNOR U38054 ( .A(n30121), .B(n34220), .Z(n38362) );
  XNOR U38055 ( .A(n38363), .B(n35862), .Z(n34220) );
  ANDN U38056 ( .B(n34034), .A(n36517), .Z(n38363) );
  IV U38057 ( .A(n34036), .Z(n36517) );
  XOR U38058 ( .A(n38364), .B(n35082), .Z(n34036) );
  XNOR U38059 ( .A(n38365), .B(n35853), .Z(n30121) );
  ANDN U38060 ( .B(n38366), .A(n36515), .Z(n38365) );
  XNOR U38061 ( .A(n32837), .B(n38367), .Z(n38361) );
  XOR U38062 ( .A(n33234), .B(n30201), .Z(n38367) );
  XNOR U38063 ( .A(n38368), .B(n35856), .Z(n30201) );
  ANDN U38064 ( .B(n34032), .A(n38369), .Z(n38368) );
  XNOR U38065 ( .A(n38370), .B(n37427), .Z(n34032) );
  XNOR U38066 ( .A(n38371), .B(n35865), .Z(n33234) );
  ANDN U38067 ( .B(n34040), .A(n38372), .Z(n38371) );
  XNOR U38068 ( .A(n38373), .B(n38374), .Z(n34040) );
  XOR U38069 ( .A(n38375), .B(n36523), .Z(n32837) );
  ANDN U38070 ( .B(n34027), .A(n38376), .Z(n38375) );
  XOR U38071 ( .A(n35304), .B(n38377), .Z(n34027) );
  XNOR U38072 ( .A(n38378), .B(n38379), .Z(n33454) );
  XNOR U38073 ( .A(n38380), .B(n33372), .Z(n38379) );
  XOR U38074 ( .A(n38381), .B(n38382), .Z(n33372) );
  AND U38075 ( .A(n38002), .B(n38004), .Z(n38381) );
  XOR U38076 ( .A(n34114), .B(n38383), .Z(n38378) );
  XOR U38077 ( .A(n30038), .B(n33739), .Z(n38383) );
  XOR U38078 ( .A(n38384), .B(n38385), .Z(n33739) );
  AND U38079 ( .A(n37993), .B(n37995), .Z(n38384) );
  ANDN U38080 ( .B(n38000), .A(n37998), .Z(n38386) );
  IV U38081 ( .A(n38388), .Z(n38000) );
  XNOR U38082 ( .A(n38389), .B(n38390), .Z(n34114) );
  XNOR U38083 ( .A(n38391), .B(n38366), .Z(n34023) );
  XNOR U38084 ( .A(n38392), .B(n37880), .Z(n35851) );
  XOR U38085 ( .A(n37069), .B(n38393), .Z(n36515) );
  XNOR U38086 ( .A(n26235), .B(n38394), .Z(n38229) );
  XNOR U38087 ( .A(n24246), .B(n26419), .Z(n38394) );
  XNOR U38088 ( .A(n38395), .B(n27857), .Z(n26419) );
  XOR U38089 ( .A(n38067), .B(n32531), .Z(n27857) );
  XNOR U38090 ( .A(n36324), .B(n38396), .Z(n32531) );
  XNOR U38091 ( .A(n38397), .B(n38398), .Z(n36324) );
  XNOR U38092 ( .A(n32170), .B(n33151), .Z(n38398) );
  XNOR U38093 ( .A(n38399), .B(n36044), .Z(n33151) );
  ANDN U38094 ( .B(n36043), .A(n38056), .Z(n38399) );
  XNOR U38095 ( .A(n38400), .B(n38401), .Z(n36043) );
  XNOR U38096 ( .A(n38402), .B(n33230), .Z(n32170) );
  ANDN U38097 ( .B(n33229), .A(n38053), .Z(n38402) );
  XNOR U38098 ( .A(n38403), .B(n37264), .Z(n33229) );
  XNOR U38099 ( .A(n27651), .B(n38404), .Z(n38397) );
  XOR U38100 ( .A(n31034), .B(n32567), .Z(n38404) );
  XOR U38101 ( .A(n38405), .B(n37807), .Z(n32567) );
  ANDN U38102 ( .B(n37808), .A(n38050), .Z(n38405) );
  XOR U38103 ( .A(n38406), .B(n36701), .Z(n37808) );
  XNOR U38104 ( .A(n38407), .B(n33845), .Z(n31034) );
  ANDN U38105 ( .B(n33846), .A(n38046), .Z(n38407) );
  XNOR U38106 ( .A(n38408), .B(n37776), .Z(n33846) );
  XNOR U38107 ( .A(n38409), .B(n33938), .Z(n27651) );
  NOR U38108 ( .A(n33939), .B(n38043), .Z(n38409) );
  XOR U38109 ( .A(n38410), .B(n38411), .Z(n33939) );
  XNOR U38110 ( .A(n38412), .B(n36755), .Z(n38067) );
  ANDN U38111 ( .B(n38413), .A(n38414), .Z(n38412) );
  NOR U38112 ( .A(n27856), .B(n30191), .Z(n38395) );
  XOR U38113 ( .A(n36461), .B(n28879), .Z(n30191) );
  XOR U38114 ( .A(n35561), .B(n37294), .Z(n28879) );
  XOR U38115 ( .A(n38415), .B(n38416), .Z(n37294) );
  XNOR U38116 ( .A(n31443), .B(n38327), .Z(n38416) );
  XOR U38117 ( .A(n38417), .B(n36055), .Z(n38327) );
  XNOR U38118 ( .A(n38418), .B(n38419), .Z(n36055) );
  ANDN U38119 ( .B(n37296), .A(n37298), .Z(n38417) );
  XNOR U38120 ( .A(n38124), .B(n38420), .Z(n37298) );
  XNOR U38121 ( .A(n38421), .B(n38422), .Z(n37296) );
  XOR U38122 ( .A(n38423), .B(n36060), .Z(n31443) );
  XOR U38123 ( .A(n38424), .B(n38151), .Z(n36060) );
  NOR U38124 ( .A(n36488), .B(n36487), .Z(n38423) );
  XNOR U38125 ( .A(n38425), .B(n38426), .Z(n36487) );
  XNOR U38126 ( .A(n38427), .B(n36976), .Z(n36488) );
  XNOR U38127 ( .A(n33019), .B(n38428), .Z(n38415) );
  XNOR U38128 ( .A(n32619), .B(n33032), .Z(n38428) );
  XOR U38129 ( .A(n38429), .B(n36064), .Z(n33032) );
  XNOR U38130 ( .A(n38430), .B(n37272), .Z(n36064) );
  ANDN U38131 ( .B(n36494), .A(n36495), .Z(n38429) );
  XNOR U38132 ( .A(n38431), .B(n38432), .Z(n36495) );
  XNOR U38133 ( .A(n37857), .B(n38433), .Z(n36494) );
  IV U38134 ( .A(n36941), .Z(n37857) );
  XNOR U38135 ( .A(n38434), .B(n38435), .Z(n36941) );
  XNOR U38136 ( .A(n38436), .B(n36068), .Z(n32619) );
  XNOR U38137 ( .A(n38437), .B(n38438), .Z(n36068) );
  NOR U38138 ( .A(n36484), .B(n36483), .Z(n38436) );
  XOR U38139 ( .A(n38439), .B(n38440), .Z(n36483) );
  XOR U38140 ( .A(n38441), .B(n35634), .Z(n36484) );
  XOR U38141 ( .A(n38442), .B(n36050), .Z(n33019) );
  XOR U38142 ( .A(n38443), .B(n38444), .Z(n36050) );
  ANDN U38143 ( .B(n36491), .A(n36492), .Z(n38442) );
  XOR U38144 ( .A(n38445), .B(n38446), .Z(n36492) );
  XOR U38145 ( .A(n38447), .B(n37176), .Z(n36491) );
  XNOR U38146 ( .A(n38448), .B(n38449), .Z(n37176) );
  XOR U38147 ( .A(n38450), .B(n38451), .Z(n35561) );
  XNOR U38148 ( .A(n30265), .B(n32594), .Z(n38451) );
  XNOR U38149 ( .A(n38452), .B(n36875), .Z(n32594) );
  NOR U38150 ( .A(n36876), .B(n36469), .Z(n38452) );
  XNOR U38151 ( .A(n37912), .B(n38453), .Z(n36469) );
  XOR U38152 ( .A(n38454), .B(n35297), .Z(n36876) );
  XNOR U38153 ( .A(n38455), .B(n36879), .Z(n30265) );
  ANDN U38154 ( .B(n36464), .A(n36463), .Z(n38455) );
  XNOR U38155 ( .A(n38456), .B(n38457), .Z(n36463) );
  XOR U38156 ( .A(n38458), .B(n36353), .Z(n36464) );
  XOR U38157 ( .A(n34788), .B(n38459), .Z(n38450) );
  XNOR U38158 ( .A(n32765), .B(n31259), .Z(n38459) );
  XNOR U38159 ( .A(n38460), .B(n36868), .Z(n31259) );
  ANDN U38160 ( .B(n36477), .A(n36476), .Z(n38460) );
  XNOR U38161 ( .A(n38461), .B(n35932), .Z(n36476) );
  XNOR U38162 ( .A(n35933), .B(n38462), .Z(n36477) );
  XOR U38163 ( .A(n38463), .B(n36883), .Z(n32765) );
  ANDN U38164 ( .B(n36882), .A(n38014), .Z(n38463) );
  XNOR U38165 ( .A(n38464), .B(n36871), .Z(n34788) );
  ANDN U38166 ( .B(n36474), .A(n36472), .Z(n38464) );
  XOR U38167 ( .A(n38465), .B(n38037), .Z(n36472) );
  XNOR U38168 ( .A(n38466), .B(n38467), .Z(n36474) );
  XOR U38169 ( .A(n38468), .B(n36882), .Z(n36461) );
  XOR U38170 ( .A(n38469), .B(n37061), .Z(n36882) );
  XOR U38171 ( .A(n38470), .B(n37326), .Z(n38014) );
  XNOR U38172 ( .A(n32142), .B(n34476), .Z(n27856) );
  XOR U38173 ( .A(n38471), .B(n37241), .Z(n34476) );
  ANDN U38174 ( .B(n35173), .A(n35175), .Z(n38471) );
  XNOR U38175 ( .A(n38472), .B(n38473), .Z(n35396) );
  XNOR U38176 ( .A(n33326), .B(n33193), .Z(n38473) );
  XOR U38177 ( .A(n38474), .B(n34757), .Z(n33193) );
  ANDN U38178 ( .B(n34758), .A(n38214), .Z(n38474) );
  XOR U38179 ( .A(n38475), .B(n36092), .Z(n33326) );
  NOR U38180 ( .A(n38476), .B(n36091), .Z(n38475) );
  XOR U38181 ( .A(n33716), .B(n38477), .Z(n38472) );
  XOR U38182 ( .A(n32515), .B(n30214), .Z(n38477) );
  XNOR U38183 ( .A(n38478), .B(n34763), .Z(n30214) );
  ANDN U38184 ( .B(n34764), .A(n38206), .Z(n38478) );
  XNOR U38185 ( .A(n38479), .B(n34754), .Z(n32515) );
  NOR U38186 ( .A(n34753), .B(n38211), .Z(n38479) );
  XNOR U38187 ( .A(n38480), .B(n34767), .Z(n33716) );
  ANDN U38188 ( .B(n34768), .A(n38233), .Z(n38480) );
  XOR U38189 ( .A(n38481), .B(n38482), .Z(n35149) );
  XOR U38190 ( .A(n28431), .B(n34747), .Z(n38482) );
  XOR U38191 ( .A(n38483), .B(n37251), .Z(n34747) );
  XNOR U38192 ( .A(n38484), .B(n35579), .Z(n34478) );
  XOR U38193 ( .A(n38485), .B(n38486), .Z(n34479) );
  XNOR U38194 ( .A(n38487), .B(n37243), .Z(n28431) );
  ANDN U38195 ( .B(n34473), .A(n34471), .Z(n38487) );
  IV U38196 ( .A(n37244), .Z(n34471) );
  XOR U38197 ( .A(n38488), .B(n38489), .Z(n37244) );
  XOR U38198 ( .A(n38490), .B(n38491), .Z(n34473) );
  XNOR U38199 ( .A(n29932), .B(n38492), .Z(n38481) );
  XOR U38200 ( .A(n32084), .B(n32974), .Z(n38492) );
  XNOR U38201 ( .A(n38493), .B(n37240), .Z(n32974) );
  ANDN U38202 ( .B(n37241), .A(n35173), .Z(n38493) );
  XNOR U38203 ( .A(n37018), .B(n38494), .Z(n35173) );
  XNOR U38204 ( .A(n38495), .B(n37623), .Z(n37241) );
  XNOR U38205 ( .A(n38496), .B(n38497), .Z(n32084) );
  NOR U38206 ( .A(n34467), .B(n34468), .Z(n38496) );
  XNOR U38207 ( .A(n38498), .B(n38499), .Z(n34468) );
  XOR U38208 ( .A(n38500), .B(n37249), .Z(n29932) );
  NOR U38209 ( .A(n37248), .B(n35182), .Z(n38500) );
  XOR U38210 ( .A(n35787), .B(n38501), .Z(n35182) );
  XOR U38211 ( .A(n35519), .B(n38502), .Z(n37248) );
  XNOR U38212 ( .A(n38503), .B(n27865), .Z(n24246) );
  XOR U38213 ( .A(n36571), .B(n30009), .Z(n27865) );
  IV U38214 ( .A(n29943), .Z(n30009) );
  XNOR U38215 ( .A(n38504), .B(n38505), .Z(n36243) );
  XOR U38216 ( .A(n34955), .B(n31546), .Z(n38505) );
  XOR U38217 ( .A(n38506), .B(n35258), .Z(n31546) );
  XNOR U38218 ( .A(n38507), .B(n38508), .Z(n35258) );
  ANDN U38219 ( .B(n35259), .A(n36574), .Z(n38506) );
  XOR U38220 ( .A(n38509), .B(n37331), .Z(n35259) );
  XOR U38221 ( .A(n38511), .B(n36359), .Z(n35255) );
  NOR U38222 ( .A(n38512), .B(n35254), .Z(n38510) );
  XOR U38223 ( .A(n33183), .B(n38513), .Z(n38504) );
  XNOR U38224 ( .A(n31106), .B(n33050), .Z(n38513) );
  XNOR U38225 ( .A(n38514), .B(n35267), .Z(n33050) );
  XOR U38226 ( .A(n38515), .B(n37968), .Z(n35267) );
  NOR U38227 ( .A(n36564), .B(n36565), .Z(n38514) );
  XOR U38228 ( .A(n38516), .B(n37076), .Z(n36564) );
  XOR U38229 ( .A(n38518), .B(n38519), .Z(n35263) );
  ANDN U38230 ( .B(n35264), .A(n36576), .Z(n38517) );
  XNOR U38231 ( .A(n38520), .B(n38521), .Z(n35264) );
  XNOR U38232 ( .A(n38522), .B(n35271), .Z(n33183) );
  XOR U38233 ( .A(n38523), .B(n38524), .Z(n35271) );
  ANDN U38234 ( .B(n35272), .A(n36568), .Z(n38522) );
  XOR U38235 ( .A(n38525), .B(n38526), .Z(n35272) );
  XOR U38236 ( .A(n38528), .B(n35254), .Z(n36571) );
  XOR U38237 ( .A(n38529), .B(n38530), .Z(n35254) );
  NOR U38238 ( .A(n27866), .B(n27770), .Z(n38503) );
  XOR U38239 ( .A(n37552), .B(n32191), .Z(n27770) );
  XOR U38240 ( .A(n38531), .B(n38532), .Z(n37810) );
  XNOR U38241 ( .A(n33327), .B(n28996), .Z(n38532) );
  XNOR U38242 ( .A(n38533), .B(n35196), .Z(n28996) );
  XOR U38243 ( .A(n38534), .B(n38535), .Z(n35196) );
  ANDN U38244 ( .B(n35197), .A(n37565), .Z(n38533) );
  XNOR U38245 ( .A(n38536), .B(n38537), .Z(n35197) );
  XNOR U38246 ( .A(n38538), .B(n35200), .Z(n33327) );
  XNOR U38247 ( .A(n38539), .B(n35522), .Z(n35200) );
  AND U38248 ( .A(n38540), .B(n35201), .Z(n38538) );
  XNOR U38249 ( .A(n30951), .B(n38541), .Z(n38531) );
  XOR U38250 ( .A(n30824), .B(n32540), .Z(n38541) );
  XOR U38251 ( .A(n38542), .B(n37743), .Z(n32540) );
  IV U38252 ( .A(n35210), .Z(n37743) );
  XOR U38253 ( .A(n38543), .B(n38544), .Z(n35210) );
  ANDN U38254 ( .B(n35211), .A(n37560), .Z(n38542) );
  XOR U38255 ( .A(n37449), .B(n38545), .Z(n35211) );
  XOR U38256 ( .A(n38546), .B(n35206), .Z(n30824) );
  XOR U38257 ( .A(n38131), .B(n38547), .Z(n35206) );
  ANDN U38258 ( .B(n35207), .A(n37562), .Z(n38546) );
  XOR U38259 ( .A(n38548), .B(n38248), .Z(n35207) );
  XNOR U38260 ( .A(n38549), .B(n37749), .Z(n30951) );
  XOR U38261 ( .A(n34628), .B(n38550), .Z(n37749) );
  ANDN U38262 ( .B(n37554), .A(n37556), .Z(n38549) );
  XNOR U38263 ( .A(n38551), .B(n38332), .Z(n37554) );
  XNOR U38264 ( .A(n38552), .B(n38553), .Z(n34526) );
  XNOR U38265 ( .A(n35560), .B(n33536), .Z(n38553) );
  XNOR U38266 ( .A(n38554), .B(n35567), .Z(n33536) );
  XNOR U38267 ( .A(n35510), .B(n38555), .Z(n35567) );
  ANDN U38268 ( .B(n35068), .A(n35066), .Z(n38554) );
  XNOR U38269 ( .A(n38556), .B(n38557), .Z(n35066) );
  XNOR U38270 ( .A(n38558), .B(n36151), .Z(n35560) );
  XOR U38271 ( .A(n38559), .B(n36423), .Z(n36151) );
  NOR U38272 ( .A(n35070), .B(n35071), .Z(n38558) );
  XOR U38273 ( .A(n38560), .B(n37848), .Z(n35070) );
  XNOR U38274 ( .A(n31667), .B(n38561), .Z(n38552) );
  XOR U38275 ( .A(n32749), .B(n32722), .Z(n38561) );
  XNOR U38276 ( .A(n38562), .B(n36886), .Z(n32722) );
  XOR U38277 ( .A(n38563), .B(n38564), .Z(n36886) );
  NOR U38278 ( .A(n35053), .B(n35054), .Z(n38562) );
  XNOR U38279 ( .A(n38565), .B(n35932), .Z(n35053) );
  XOR U38280 ( .A(n38566), .B(n38567), .Z(n32749) );
  ANDN U38281 ( .B(n35057), .A(n35058), .Z(n38566) );
  XNOR U38282 ( .A(n35586), .B(n38568), .Z(n35057) );
  XNOR U38283 ( .A(n38569), .B(n35572), .Z(n31667) );
  NOR U38284 ( .A(n35064), .B(n35062), .Z(n38569) );
  XOR U38285 ( .A(n36894), .B(n38570), .Z(n35062) );
  XOR U38286 ( .A(n38571), .B(n35201), .Z(n37552) );
  XNOR U38287 ( .A(n38572), .B(n38573), .Z(n35201) );
  ANDN U38288 ( .B(n37751), .A(n38540), .Z(n38571) );
  XOR U38289 ( .A(n36080), .B(n31467), .Z(n27866) );
  XOR U38290 ( .A(n33714), .B(n33365), .Z(n31467) );
  XNOR U38291 ( .A(n38574), .B(n38575), .Z(n33365) );
  XNOR U38292 ( .A(n29031), .B(n30545), .Z(n38575) );
  XNOR U38293 ( .A(n38576), .B(n36733), .Z(n30545) );
  XNOR U38294 ( .A(n38577), .B(n38096), .Z(n37135) );
  XOR U38295 ( .A(n38578), .B(n36737), .Z(n29031) );
  XNOR U38296 ( .A(n38579), .B(n36507), .Z(n37128) );
  XNOR U38297 ( .A(n33330), .B(n38580), .Z(n38574) );
  XOR U38298 ( .A(n32231), .B(n29405), .Z(n38580) );
  XOR U38299 ( .A(n38581), .B(n37155), .Z(n29405) );
  XOR U38300 ( .A(n38582), .B(n35078), .Z(n37131) );
  XOR U38301 ( .A(n38583), .B(n36728), .Z(n32231) );
  XNOR U38302 ( .A(n38584), .B(n37183), .Z(n37483) );
  XNOR U38303 ( .A(n38585), .B(n36723), .Z(n33330) );
  ANDN U38304 ( .B(n37478), .A(n37138), .Z(n38585) );
  XNOR U38305 ( .A(n38586), .B(n38587), .Z(n37138) );
  XOR U38306 ( .A(n38588), .B(n38589), .Z(n33714) );
  XNOR U38307 ( .A(n36818), .B(n33848), .Z(n38589) );
  XNOR U38308 ( .A(n38590), .B(n37280), .Z(n33848) );
  NOR U38309 ( .A(n36072), .B(n36073), .Z(n38590) );
  XOR U38310 ( .A(n37677), .B(n38591), .Z(n36073) );
  XNOR U38311 ( .A(n38592), .B(n38593), .Z(n36818) );
  XNOR U38312 ( .A(n4687), .B(n38594), .Z(n38593) );
  OR U38313 ( .A(n36077), .B(n36076), .Z(n38594) );
  XOR U38314 ( .A(n37172), .B(n38595), .Z(n36077) );
  XOR U38315 ( .A(n31055), .B(n38596), .Z(n38588) );
  XOR U38316 ( .A(n38597), .B(n32680), .Z(n38596) );
  XNOR U38317 ( .A(n38598), .B(n37285), .Z(n32680) );
  ANDN U38318 ( .B(n38337), .A(n38599), .Z(n38598) );
  XNOR U38319 ( .A(n38600), .B(n37289), .Z(n31055) );
  ANDN U38320 ( .B(n36082), .A(n36083), .Z(n38600) );
  XOR U38321 ( .A(n38601), .B(n38134), .Z(n36083) );
  IV U38322 ( .A(n36935), .Z(n38134) );
  XNOR U38323 ( .A(n38602), .B(n38599), .Z(n36080) );
  ANDN U38324 ( .B(n37284), .A(n38337), .Z(n38602) );
  XOR U38325 ( .A(n38498), .B(n38603), .Z(n38337) );
  XOR U38326 ( .A(n38604), .B(n38605), .Z(n37284) );
  XNOR U38327 ( .A(n38606), .B(n35889), .Z(n26235) );
  XOR U38328 ( .A(n33395), .B(n30505), .Z(n35889) );
  XNOR U38329 ( .A(n35709), .B(n33042), .Z(n30505) );
  XOR U38330 ( .A(n38607), .B(n38608), .Z(n33042) );
  XOR U38331 ( .A(n37094), .B(n34499), .Z(n38608) );
  XOR U38332 ( .A(n38609), .B(n36169), .Z(n34499) );
  XNOR U38333 ( .A(n38610), .B(n37272), .Z(n36169) );
  ANDN U38334 ( .B(n37100), .A(n34277), .Z(n38609) );
  XNOR U38335 ( .A(n38611), .B(n36167), .Z(n37094) );
  XNOR U38336 ( .A(n38612), .B(n33922), .Z(n36167) );
  ANDN U38337 ( .B(n37111), .A(n34282), .Z(n38611) );
  XOR U38338 ( .A(n32338), .B(n38613), .Z(n38607) );
  XOR U38339 ( .A(n33958), .B(n28820), .Z(n38613) );
  XNOR U38340 ( .A(n38614), .B(n36164), .Z(n28820) );
  XNOR U38341 ( .A(n38615), .B(n38616), .Z(n36164) );
  ANDN U38342 ( .B(n37107), .A(n38617), .Z(n38614) );
  XNOR U38343 ( .A(n38618), .B(n36171), .Z(n33958) );
  XNOR U38344 ( .A(n38619), .B(n38620), .Z(n36171) );
  NOR U38345 ( .A(n37115), .B(n34286), .Z(n38618) );
  XNOR U38346 ( .A(n38621), .B(n36160), .Z(n32338) );
  XOR U38347 ( .A(n38622), .B(n36955), .Z(n36160) );
  XOR U38348 ( .A(n38623), .B(n38624), .Z(n36955) );
  ANDN U38349 ( .B(n37104), .A(n34290), .Z(n38621) );
  XNOR U38350 ( .A(n38625), .B(n38626), .Z(n35709) );
  XOR U38351 ( .A(n34111), .B(n30169), .Z(n38626) );
  XOR U38352 ( .A(n38627), .B(n33783), .Z(n30169) );
  XNOR U38353 ( .A(n37720), .B(n38628), .Z(n33783) );
  AND U38354 ( .A(n38629), .B(n36232), .Z(n38627) );
  XNOR U38355 ( .A(n38630), .B(n33789), .Z(n34111) );
  XNOR U38356 ( .A(n38631), .B(n35782), .Z(n33789) );
  IV U38357 ( .A(n37069), .Z(n35782) );
  XNOR U38358 ( .A(n38632), .B(n36434), .Z(n33401) );
  XNOR U38359 ( .A(n31992), .B(n38633), .Z(n38625) );
  XOR U38360 ( .A(n31558), .B(n29746), .Z(n38633) );
  XOR U38361 ( .A(n38634), .B(n33793), .Z(n29746) );
  XOR U38362 ( .A(n38635), .B(n38432), .Z(n33793) );
  ANDN U38363 ( .B(n35356), .A(n35357), .Z(n38634) );
  XOR U38364 ( .A(n38636), .B(n38637), .Z(n35356) );
  XOR U38365 ( .A(n38638), .B(n33786), .Z(n31558) );
  XOR U38366 ( .A(n38639), .B(n38640), .Z(n33786) );
  XOR U38367 ( .A(n38641), .B(n38642), .Z(n33391) );
  XOR U38368 ( .A(n38643), .B(n33797), .Z(n31992) );
  XOR U38369 ( .A(n38644), .B(n37152), .Z(n33797) );
  ANDN U38370 ( .B(n33397), .A(n33398), .Z(n38643) );
  XOR U38371 ( .A(n37786), .B(n38645), .Z(n33397) );
  XNOR U38372 ( .A(n38646), .B(n36232), .Z(n33395) );
  XNOR U38373 ( .A(n37204), .B(n38647), .Z(n36232) );
  ANDN U38374 ( .B(n38648), .A(n38629), .Z(n38646) );
  ANDN U38375 ( .B(n27761), .A(n31424), .Z(n38606) );
  IV U38376 ( .A(n36178), .Z(n31424) );
  XOR U38377 ( .A(n35720), .B(n31834), .Z(n36178) );
  XNOR U38378 ( .A(n38649), .B(n37583), .Z(n35720) );
  NOR U38379 ( .A(n38650), .B(n37818), .Z(n38649) );
  XNOR U38380 ( .A(n32705), .B(n36026), .Z(n27761) );
  XNOR U38381 ( .A(n38651), .B(n34514), .Z(n36026) );
  ANDN U38382 ( .B(n36020), .A(n36021), .Z(n38651) );
  XOR U38383 ( .A(n32379), .B(n33063), .Z(n32705) );
  XOR U38384 ( .A(n38652), .B(n38653), .Z(n33063) );
  XNOR U38385 ( .A(n33600), .B(n36642), .Z(n38653) );
  XNOR U38386 ( .A(n38654), .B(n36646), .Z(n36642) );
  ANDN U38387 ( .B(n36274), .A(n34237), .Z(n38654) );
  XNOR U38388 ( .A(n38655), .B(n38656), .Z(n34237) );
  XNOR U38389 ( .A(n38657), .B(n38271), .Z(n36274) );
  XNOR U38390 ( .A(n38658), .B(n36653), .Z(n33600) );
  NOR U38391 ( .A(n36279), .B(n34232), .Z(n38658) );
  XNOR U38392 ( .A(n38659), .B(n36423), .Z(n34232) );
  XNOR U38393 ( .A(n38660), .B(n38174), .Z(n36279) );
  XOR U38394 ( .A(n34133), .B(n38661), .Z(n38652) );
  XOR U38395 ( .A(n32890), .B(n32992), .Z(n38661) );
  XOR U38396 ( .A(n38662), .B(n36651), .Z(n32992) );
  ANDN U38397 ( .B(n34241), .A(n36277), .Z(n38662) );
  XOR U38398 ( .A(n37071), .B(n38663), .Z(n36277) );
  XNOR U38399 ( .A(n38664), .B(n38537), .Z(n34241) );
  IV U38400 ( .A(n38352), .Z(n38537) );
  XNOR U38401 ( .A(n38665), .B(n36648), .Z(n32890) );
  ANDN U38402 ( .B(n36281), .A(n36282), .Z(n38665) );
  XNOR U38403 ( .A(n38666), .B(n38667), .Z(n36282) );
  XOR U38404 ( .A(n38668), .B(n37837), .Z(n36281) );
  XNOR U38405 ( .A(n38669), .B(n36656), .Z(n34133) );
  ANDN U38406 ( .B(n36272), .A(n34245), .Z(n38669) );
  XOR U38407 ( .A(n38671), .B(n38024), .Z(n36272) );
  XOR U38408 ( .A(n38672), .B(n38673), .Z(n32379) );
  XOR U38409 ( .A(n34502), .B(n31147), .Z(n38673) );
  XOR U38410 ( .A(n38674), .B(n34510), .Z(n31147) );
  NOR U38411 ( .A(n34509), .B(n35681), .Z(n38674) );
  XOR U38412 ( .A(n38675), .B(n37837), .Z(n35681) );
  IV U38413 ( .A(n36031), .Z(n34509) );
  XOR U38414 ( .A(n37592), .B(n38676), .Z(n36031) );
  IV U38415 ( .A(n37677), .Z(n37592) );
  XNOR U38416 ( .A(n38677), .B(n38678), .Z(n34502) );
  ANDN U38417 ( .B(n37378), .A(n35687), .Z(n38677) );
  XNOR U38418 ( .A(n38679), .B(n37646), .Z(n35687) );
  XOR U38419 ( .A(n32955), .B(n38680), .Z(n38672) );
  XNOR U38420 ( .A(n32936), .B(n33902), .Z(n38680) );
  XOR U38421 ( .A(n38681), .B(n38682), .Z(n33902) );
  NOR U38422 ( .A(n34514), .B(n36020), .Z(n38681) );
  XOR U38423 ( .A(n38685), .B(n38686), .Z(n34514) );
  XNOR U38424 ( .A(n38687), .B(n34518), .Z(n32936) );
  ANDN U38425 ( .B(n34519), .A(n35677), .Z(n38687) );
  XOR U38426 ( .A(n38688), .B(n36423), .Z(n35677) );
  XOR U38427 ( .A(n38691), .B(n38640), .Z(n34519) );
  XNOR U38428 ( .A(n38692), .B(n34522), .Z(n32955) );
  NOR U38429 ( .A(n36029), .B(n35684), .Z(n38692) );
  XNOR U38430 ( .A(n38616), .B(n38693), .Z(n35684) );
  XOR U38431 ( .A(n38694), .B(n38656), .Z(n36029) );
  XOR U38432 ( .A(n38695), .B(n38696), .Z(n29041) );
  XOR U38433 ( .A(n27850), .B(n25775), .Z(n38696) );
  XNOR U38434 ( .A(n38697), .B(n31774), .Z(n25775) );
  IV U38435 ( .A(n29484), .Z(n31774) );
  XNOR U38436 ( .A(n38698), .B(n30275), .Z(n29484) );
  XNOR U38437 ( .A(n36501), .B(n38699), .Z(n30275) );
  XOR U38438 ( .A(n38700), .B(n38701), .Z(n36501) );
  XOR U38439 ( .A(n37969), .B(n32848), .Z(n38701) );
  XNOR U38440 ( .A(n38702), .B(n38703), .Z(n32848) );
  NOR U38441 ( .A(n38007), .B(n38704), .Z(n38702) );
  XNOR U38442 ( .A(n38705), .B(n37991), .Z(n37969) );
  XNOR U38443 ( .A(n38706), .B(n37014), .Z(n37991) );
  IV U38444 ( .A(n35297), .Z(n37014) );
  ANDN U38445 ( .B(n37990), .A(n38709), .Z(n38705) );
  XOR U38446 ( .A(n31375), .B(n38710), .Z(n38700) );
  XOR U38447 ( .A(n33239), .B(n31552), .Z(n38710) );
  XNOR U38448 ( .A(n38711), .B(n38388), .Z(n31552) );
  XOR U38449 ( .A(n38712), .B(n36406), .Z(n38388) );
  NOR U38450 ( .A(n38713), .B(n37999), .Z(n38711) );
  XOR U38451 ( .A(n38714), .B(n37995), .Z(n33239) );
  XOR U38452 ( .A(n35926), .B(n38715), .Z(n37995) );
  ANDN U38453 ( .B(n38716), .A(n38717), .Z(n38714) );
  XNOR U38454 ( .A(n38718), .B(n38004), .Z(n31375) );
  XOR U38455 ( .A(n38719), .B(n38720), .Z(n38004) );
  ANDN U38456 ( .B(n38721), .A(n38722), .Z(n38718) );
  XOR U38457 ( .A(n38723), .B(n29470), .Z(n27850) );
  XNOR U38458 ( .A(n36138), .B(n31674), .Z(n29470) );
  IV U38459 ( .A(n29713), .Z(n31674) );
  XOR U38460 ( .A(n36222), .B(n37342), .Z(n29713) );
  XOR U38461 ( .A(n38724), .B(n38725), .Z(n37342) );
  XOR U38462 ( .A(n28813), .B(n31806), .Z(n38725) );
  XOR U38463 ( .A(n38726), .B(n36844), .Z(n31806) );
  ANDN U38464 ( .B(n36845), .A(n38727), .Z(n38726) );
  XNOR U38465 ( .A(n38728), .B(n36852), .Z(n28813) );
  IV U38466 ( .A(n38729), .Z(n36852) );
  ANDN U38467 ( .B(n36141), .A(n36142), .Z(n38728) );
  XNOR U38468 ( .A(n38730), .B(n37264), .Z(n36141) );
  XNOR U38469 ( .A(n33411), .B(n38731), .Z(n38724) );
  XOR U38470 ( .A(n30590), .B(n36820), .Z(n38731) );
  XOR U38471 ( .A(n38732), .B(n36849), .Z(n36820) );
  NOR U38472 ( .A(n36145), .B(n36146), .Z(n38732) );
  XOR U38473 ( .A(n38733), .B(n38734), .Z(n36145) );
  XNOR U38474 ( .A(n38735), .B(n36841), .Z(n30590) );
  AND U38475 ( .A(n36131), .B(n36132), .Z(n38735) );
  XOR U38476 ( .A(n38736), .B(n35155), .Z(n36131) );
  XOR U38477 ( .A(n38737), .B(n36855), .Z(n33411) );
  NOR U38478 ( .A(n36856), .B(n36136), .Z(n38737) );
  XOR U38479 ( .A(n37718), .B(n38738), .Z(n36856) );
  IV U38480 ( .A(n37625), .Z(n37718) );
  XOR U38481 ( .A(n38739), .B(n38740), .Z(n36222) );
  XOR U38482 ( .A(n30506), .B(n32197), .Z(n38740) );
  XOR U38483 ( .A(n38741), .B(n36833), .Z(n32197) );
  ANDN U38484 ( .B(n35901), .A(n35903), .Z(n38741) );
  XOR U38485 ( .A(n38742), .B(n36507), .Z(n35901) );
  XNOR U38486 ( .A(n38743), .B(n36825), .Z(n30506) );
  ANDN U38487 ( .B(n36235), .A(n36236), .Z(n38743) );
  XNOR U38488 ( .A(n38744), .B(n37491), .Z(n36235) );
  IV U38489 ( .A(n36946), .Z(n37491) );
  XOR U38490 ( .A(n33537), .B(n38745), .Z(n38739) );
  XNOR U38491 ( .A(n31363), .B(n32220), .Z(n38745) );
  XNOR U38492 ( .A(n38746), .B(n36828), .Z(n32220) );
  NOR U38493 ( .A(n35909), .B(n35907), .Z(n38746) );
  XNOR U38494 ( .A(n37635), .B(n38747), .Z(n35907) );
  XNOR U38495 ( .A(n38748), .B(n38749), .Z(n31363) );
  ANDN U38496 ( .B(n35897), .A(n35898), .Z(n38748) );
  XNOR U38497 ( .A(n38750), .B(n36836), .Z(n33537) );
  ANDN U38498 ( .B(n35911), .A(n35912), .Z(n38750) );
  XOR U38499 ( .A(n37786), .B(n38751), .Z(n35911) );
  XOR U38500 ( .A(n38753), .B(n35940), .Z(n36845) );
  NOR U38501 ( .A(n38754), .B(n38755), .Z(n38752) );
  IV U38502 ( .A(n38727), .Z(n38754) );
  ANDN U38503 ( .B(n31429), .A(n31446), .Z(n38723) );
  IV U38504 ( .A(n31430), .Z(n31446) );
  XOR U38505 ( .A(n35880), .B(n37465), .Z(n31430) );
  XOR U38506 ( .A(n38756), .B(n38757), .Z(n37465) );
  XOR U38507 ( .A(n38758), .B(n38759), .Z(n35880) );
  ANDN U38508 ( .B(n37973), .A(n38760), .Z(n38758) );
  XOR U38509 ( .A(n34672), .B(n30303), .Z(n31429) );
  IV U38510 ( .A(n30260), .Z(n30303) );
  XNOR U38511 ( .A(n38761), .B(n38762), .Z(n38527) );
  XNOR U38512 ( .A(n30668), .B(n33445), .Z(n38762) );
  XOR U38513 ( .A(n38763), .B(n34970), .Z(n33445) );
  XOR U38514 ( .A(n38764), .B(n36359), .Z(n34970) );
  XOR U38515 ( .A(n38765), .B(n38766), .Z(n34674) );
  XOR U38516 ( .A(n38767), .B(n38027), .Z(n34675) );
  XNOR U38517 ( .A(n38768), .B(n34973), .Z(n30668) );
  XOR U38518 ( .A(n37690), .B(n38769), .Z(n34973) );
  ANDN U38519 ( .B(n37337), .A(n38770), .Z(n38768) );
  XOR U38520 ( .A(n31938), .B(n38771), .Z(n38761) );
  XOR U38521 ( .A(n33238), .B(n30067), .Z(n38771) );
  XNOR U38522 ( .A(n38772), .B(n34965), .Z(n30067) );
  XNOR U38523 ( .A(n38773), .B(n36362), .Z(n34965) );
  ANDN U38524 ( .B(n34682), .A(n34680), .Z(n38772) );
  XOR U38525 ( .A(n38774), .B(n38775), .Z(n34680) );
  XNOR U38526 ( .A(n38776), .B(n38777), .Z(n34682) );
  XOR U38527 ( .A(n38779), .B(n36779), .Z(n34962) );
  ANDN U38528 ( .B(n35705), .A(n34961), .Z(n38778) );
  XOR U38529 ( .A(n38780), .B(n38781), .Z(n34961) );
  XNOR U38530 ( .A(n38782), .B(n37264), .Z(n35705) );
  XNOR U38531 ( .A(n38783), .B(n36126), .Z(n31938) );
  XNOR U38532 ( .A(n38784), .B(n38486), .Z(n36126) );
  AND U38533 ( .A(n34685), .B(n34684), .Z(n38783) );
  XOR U38534 ( .A(n38785), .B(n37851), .Z(n34684) );
  XOR U38535 ( .A(n38786), .B(n35792), .Z(n34685) );
  XNOR U38536 ( .A(n38787), .B(n38788), .Z(n34432) );
  XOR U38537 ( .A(n38789), .B(n32286), .Z(n38788) );
  XNOR U38538 ( .A(n38790), .B(n36133), .Z(n32286) );
  AND U38539 ( .A(n36841), .B(n36840), .Z(n38790) );
  XOR U38540 ( .A(n38791), .B(n38792), .Z(n36841) );
  XOR U38541 ( .A(n33196), .B(n38793), .Z(n38787) );
  XNOR U38542 ( .A(n30940), .B(n30751), .Z(n38793) );
  XNOR U38543 ( .A(n38794), .B(n36147), .Z(n30751) );
  NOR U38544 ( .A(n36849), .B(n36848), .Z(n38794) );
  XOR U38545 ( .A(n38795), .B(n37841), .Z(n36849) );
  XNOR U38546 ( .A(n38796), .B(n38755), .Z(n30940) );
  NOR U38547 ( .A(n38797), .B(n36844), .Z(n38796) );
  XNOR U38548 ( .A(n38798), .B(n33922), .Z(n36844) );
  XNOR U38549 ( .A(n38799), .B(n36143), .Z(n33196) );
  IV U38550 ( .A(n38800), .Z(n36143) );
  NOR U38551 ( .A(n38729), .B(n36851), .Z(n38799) );
  XOR U38552 ( .A(n38801), .B(n38802), .Z(n38729) );
  XNOR U38553 ( .A(n38803), .B(n34974), .Z(n34672) );
  IV U38554 ( .A(n38770), .Z(n34974) );
  XNOR U38555 ( .A(n38804), .B(n38805), .Z(n38770) );
  NOR U38556 ( .A(n37338), .B(n37337), .Z(n38803) );
  XNOR U38557 ( .A(n38806), .B(n38807), .Z(n37337) );
  XOR U38558 ( .A(n38808), .B(n36406), .Z(n37338) );
  IV U38559 ( .A(n36209), .Z(n36406) );
  XOR U38560 ( .A(n25970), .B(n38811), .Z(n38695) );
  XNOR U38561 ( .A(n27237), .B(n25765), .Z(n38811) );
  XNOR U38562 ( .A(n38812), .B(n29466), .Z(n25765) );
  XNOR U38563 ( .A(n37530), .B(n30662), .Z(n29466) );
  XNOR U38564 ( .A(n33881), .B(n34042), .Z(n30662) );
  XOR U38565 ( .A(n38813), .B(n38814), .Z(n34042) );
  XNOR U38566 ( .A(n33197), .B(n33005), .Z(n38814) );
  XNOR U38567 ( .A(n38815), .B(n35339), .Z(n33005) );
  XNOR U38568 ( .A(n38816), .B(n38277), .Z(n35339) );
  NOR U38569 ( .A(n35130), .B(n36305), .Z(n38815) );
  XOR U38570 ( .A(n38817), .B(n38818), .Z(n36305) );
  XNOR U38571 ( .A(n38819), .B(n38820), .Z(n35130) );
  XNOR U38572 ( .A(n38821), .B(n35350), .Z(n33197) );
  XNOR U38573 ( .A(n36442), .B(n38822), .Z(n35350) );
  ANDN U38574 ( .B(n36317), .A(n35144), .Z(n38821) );
  XOR U38575 ( .A(n32539), .B(n38823), .Z(n38813) );
  XOR U38576 ( .A(n32739), .B(n30294), .Z(n38823) );
  XOR U38577 ( .A(n38824), .B(n35345), .Z(n30294) );
  XOR U38578 ( .A(n38825), .B(n38826), .Z(n35345) );
  ANDN U38579 ( .B(n36313), .A(n35140), .Z(n38824) );
  XOR U38580 ( .A(n38827), .B(n38093), .Z(n35140) );
  XNOR U38581 ( .A(n38828), .B(n36779), .Z(n36313) );
  XNOR U38582 ( .A(n38829), .B(n35348), .Z(n32739) );
  XOR U38583 ( .A(n38830), .B(n38401), .Z(n35348) );
  ANDN U38584 ( .B(n35245), .A(n37531), .Z(n38829) );
  IV U38585 ( .A(n36321), .Z(n37531) );
  XOR U38586 ( .A(n38831), .B(n35526), .Z(n36321) );
  XNOR U38587 ( .A(n38832), .B(n37515), .Z(n35245) );
  XNOR U38588 ( .A(n38833), .B(n35342), .Z(n32539) );
  XNOR U38589 ( .A(n35378), .B(n38834), .Z(n35342) );
  NOR U38590 ( .A(n35134), .B(n36309), .Z(n38833) );
  XOR U38591 ( .A(n38835), .B(n38836), .Z(n36309) );
  XOR U38592 ( .A(n38837), .B(n38792), .Z(n35134) );
  IV U38593 ( .A(n38573), .Z(n38792) );
  XNOR U38594 ( .A(n38838), .B(n38839), .Z(n33881) );
  XNOR U38595 ( .A(n31592), .B(n32391), .Z(n38839) );
  XNOR U38596 ( .A(n38840), .B(n38841), .Z(n32391) );
  ANDN U38597 ( .B(n35232), .A(n33750), .Z(n38840) );
  XOR U38598 ( .A(n38842), .B(n38843), .Z(n33750) );
  XNOR U38599 ( .A(n38844), .B(n35654), .Z(n31592) );
  ANDN U38600 ( .B(n35234), .A(n33759), .Z(n38844) );
  IV U38601 ( .A(n35235), .Z(n33759) );
  XNOR U38602 ( .A(n38845), .B(n37027), .Z(n35235) );
  XNOR U38603 ( .A(n36979), .B(n38846), .Z(n35234) );
  XOR U38604 ( .A(n31453), .B(n38847), .Z(n38838) );
  XNOR U38605 ( .A(n32846), .B(n35635), .Z(n38847) );
  XNOR U38606 ( .A(n38848), .B(n38849), .Z(n35635) );
  ANDN U38607 ( .B(n35243), .A(n33755), .Z(n38848) );
  XNOR U38608 ( .A(n38850), .B(n35516), .Z(n33755) );
  XOR U38609 ( .A(n38851), .B(n38852), .Z(n35243) );
  XNOR U38610 ( .A(n38853), .B(n37586), .Z(n32846) );
  ANDN U38611 ( .B(n33746), .A(n35238), .Z(n38853) );
  XOR U38612 ( .A(n38854), .B(n38432), .Z(n35238) );
  XOR U38613 ( .A(n38855), .B(n35613), .Z(n33746) );
  XOR U38614 ( .A(n38856), .B(n35918), .Z(n31453) );
  ANDN U38615 ( .B(n35240), .A(n33763), .Z(n38856) );
  IV U38616 ( .A(n35241), .Z(n33763) );
  XOR U38617 ( .A(n38857), .B(n37011), .Z(n35241) );
  XNOR U38618 ( .A(n38858), .B(n38859), .Z(n35240) );
  XOR U38619 ( .A(n38860), .B(n36317), .Z(n37530) );
  XOR U38620 ( .A(n38861), .B(n38777), .Z(n36317) );
  XOR U38621 ( .A(n38862), .B(n38863), .Z(n35144) );
  XOR U38622 ( .A(n38864), .B(n38865), .Z(n35146) );
  ANDN U38623 ( .B(n30390), .A(n31438), .Z(n38812) );
  XNOR U38624 ( .A(n32302), .B(n37364), .Z(n31438) );
  XOR U38625 ( .A(n38866), .B(n35225), .Z(n37364) );
  ANDN U38626 ( .B(n33278), .A(n33279), .Z(n38866) );
  XOR U38627 ( .A(n38867), .B(n35078), .Z(n33279) );
  XNOR U38628 ( .A(n38868), .B(n38323), .Z(n32302) );
  XOR U38629 ( .A(n38869), .B(n38870), .Z(n38323) );
  XNOR U38630 ( .A(n30542), .B(n31012), .Z(n38870) );
  XNOR U38631 ( .A(n38871), .B(n33811), .Z(n31012) );
  XNOR U38632 ( .A(n38872), .B(n37630), .Z(n33811) );
  ANDN U38633 ( .B(n33810), .A(n33284), .Z(n38871) );
  XOR U38634 ( .A(n37110), .B(n38873), .Z(n33284) );
  XOR U38635 ( .A(n38874), .B(n37710), .Z(n33810) );
  XNOR U38636 ( .A(n38875), .B(n35226), .Z(n30542) );
  XOR U38637 ( .A(n38876), .B(n38158), .Z(n35226) );
  IV U38638 ( .A(n38318), .Z(n38158) );
  ANDN U38639 ( .B(n35225), .A(n33278), .Z(n38875) );
  XOR U38640 ( .A(n38877), .B(n35155), .Z(n33278) );
  IV U38641 ( .A(n38878), .Z(n35155) );
  XOR U38642 ( .A(n38851), .B(n38879), .Z(n35225) );
  XOR U38643 ( .A(n29162), .B(n38880), .Z(n38869) );
  XOR U38644 ( .A(n33801), .B(n32851), .Z(n38880) );
  XNOR U38645 ( .A(n38881), .B(n37459), .Z(n32851) );
  IV U38646 ( .A(n37438), .Z(n37459) );
  XOR U38647 ( .A(n38882), .B(n38438), .Z(n37438) );
  ANDN U38648 ( .B(n37366), .A(n33274), .Z(n38881) );
  XOR U38649 ( .A(n38883), .B(n38884), .Z(n33274) );
  XOR U38650 ( .A(n38885), .B(n38886), .Z(n37366) );
  XOR U38651 ( .A(n38887), .B(n33814), .Z(n33801) );
  XOR U38652 ( .A(n38888), .B(n36351), .Z(n33814) );
  ANDN U38653 ( .B(n33815), .A(n37373), .Z(n38887) );
  XOR U38654 ( .A(n38889), .B(n38890), .Z(n37373) );
  XOR U38655 ( .A(n38891), .B(n38892), .Z(n33815) );
  XOR U38656 ( .A(n38893), .B(n36035), .Z(n29162) );
  XOR U38657 ( .A(n38894), .B(n38895), .Z(n36035) );
  NOR U38658 ( .A(n36036), .B(n33288), .Z(n38893) );
  XOR U38659 ( .A(n38896), .B(n38897), .Z(n33288) );
  XOR U38660 ( .A(n38898), .B(n38781), .Z(n36036) );
  IV U38661 ( .A(n37152), .Z(n38781) );
  XOR U38662 ( .A(n38899), .B(n38900), .Z(n37152) );
  XOR U38663 ( .A(n30822), .B(n37245), .Z(n30390) );
  XNOR U38664 ( .A(n38901), .B(n35180), .Z(n37245) );
  AND U38665 ( .A(n34467), .B(n38497), .Z(n38901) );
  XOR U38666 ( .A(n37328), .B(n38902), .Z(n34467) );
  XOR U38667 ( .A(n37492), .B(n36116), .Z(n30822) );
  XNOR U38668 ( .A(n38903), .B(n38904), .Z(n36116) );
  XNOR U38669 ( .A(n32869), .B(n32145), .Z(n38904) );
  XOR U38670 ( .A(n38905), .B(n38215), .Z(n32145) );
  XOR U38671 ( .A(n38906), .B(n38907), .Z(n34756) );
  XOR U38672 ( .A(n38908), .B(n36367), .Z(n34757) );
  XOR U38673 ( .A(n38909), .B(n38212), .Z(n32869) );
  ANDN U38674 ( .B(n34752), .A(n34754), .Z(n38909) );
  XOR U38675 ( .A(n38910), .B(n37623), .Z(n34754) );
  XNOR U38676 ( .A(n38911), .B(n38912), .Z(n34752) );
  XNOR U38677 ( .A(n31267), .B(n38913), .Z(n38903) );
  XOR U38678 ( .A(n38201), .B(n29936), .Z(n38913) );
  XNOR U38679 ( .A(n38914), .B(n38915), .Z(n29936) );
  ANDN U38680 ( .B(n36092), .A(n38916), .Z(n38914) );
  XOR U38681 ( .A(n37005), .B(n38917), .Z(n36092) );
  XOR U38682 ( .A(n38918), .B(n38234), .Z(n38201) );
  NOR U38683 ( .A(n34766), .B(n34767), .Z(n38918) );
  XNOR U38684 ( .A(n38684), .B(n38919), .Z(n34767) );
  XNOR U38685 ( .A(n38920), .B(n33922), .Z(n34766) );
  XNOR U38686 ( .A(n38921), .B(n38207), .Z(n31267) );
  XNOR U38687 ( .A(n36513), .B(n38922), .Z(n34763) );
  XNOR U38688 ( .A(n37018), .B(n38923), .Z(n34762) );
  XNOR U38689 ( .A(n38924), .B(n38925), .Z(n37492) );
  XNOR U38690 ( .A(n32950), .B(n35169), .Z(n38925) );
  XNOR U38691 ( .A(n38926), .B(n35183), .Z(n35169) );
  XOR U38692 ( .A(n38927), .B(n37954), .Z(n35183) );
  XOR U38693 ( .A(n38928), .B(n38929), .Z(n37249) );
  XOR U38694 ( .A(n38556), .B(n38930), .Z(n35184) );
  XNOR U38695 ( .A(n38931), .B(n34480), .Z(n32950) );
  XNOR U38696 ( .A(n38932), .B(n35159), .Z(n34480) );
  XNOR U38697 ( .A(n38933), .B(n38934), .Z(n37251) );
  XOR U38698 ( .A(n38935), .B(n35792), .Z(n35186) );
  XOR U38699 ( .A(n34424), .B(n38936), .Z(n38924) );
  XOR U38700 ( .A(n31321), .B(n34999), .Z(n38936) );
  XNOR U38701 ( .A(n38937), .B(n34469), .Z(n34999) );
  XOR U38702 ( .A(n38938), .B(n37437), .Z(n34469) );
  NOR U38703 ( .A(n38497), .B(n35180), .Z(n38937) );
  XOR U38704 ( .A(n38939), .B(n37802), .Z(n35180) );
  XOR U38705 ( .A(n38940), .B(n37804), .Z(n38497) );
  XNOR U38706 ( .A(n38941), .B(n35175), .Z(n31321) );
  XOR U38707 ( .A(n38942), .B(n37497), .Z(n35175) );
  NOR U38708 ( .A(n35174), .B(n37240), .Z(n38941) );
  XOR U38709 ( .A(n38943), .B(n35308), .Z(n37240) );
  XOR U38710 ( .A(n38944), .B(n38945), .Z(n35174) );
  XOR U38711 ( .A(n38947), .B(n37776), .Z(n34472) );
  ANDN U38712 ( .B(n35177), .A(n37243), .Z(n38946) );
  XNOR U38713 ( .A(n38948), .B(n38949), .Z(n37243) );
  XOR U38714 ( .A(n38950), .B(n38951), .Z(n35177) );
  XNOR U38715 ( .A(n38952), .B(n29475), .Z(n27237) );
  XOR U38716 ( .A(n31960), .B(n35084), .Z(n29475) );
  XNOR U38717 ( .A(n38953), .B(n35599), .Z(n35084) );
  NOR U38718 ( .A(n34142), .B(n35108), .Z(n38953) );
  IV U38719 ( .A(n31359), .Z(n31960) );
  XNOR U38720 ( .A(n38955), .B(n34066), .Z(n31359) );
  XNOR U38721 ( .A(n38956), .B(n38957), .Z(n34066) );
  XOR U38722 ( .A(n32794), .B(n30763), .Z(n38957) );
  XNOR U38723 ( .A(n38958), .B(n34144), .Z(n30763) );
  XNOR U38724 ( .A(n38959), .B(n38960), .Z(n34144) );
  AND U38725 ( .A(n35108), .B(n35599), .Z(n38958) );
  XOR U38726 ( .A(n38961), .B(n38962), .Z(n35599) );
  XNOR U38727 ( .A(n38963), .B(n38637), .Z(n35108) );
  XNOR U38728 ( .A(n38964), .B(n34152), .Z(n32794) );
  XNOR U38729 ( .A(n38906), .B(n38965), .Z(n34152) );
  NOR U38730 ( .A(n33458), .B(n35086), .Z(n38964) );
  XOR U38731 ( .A(n38966), .B(n37187), .Z(n35086) );
  IV U38732 ( .A(n35087), .Z(n33458) );
  XOR U38733 ( .A(n38967), .B(n38619), .Z(n35087) );
  XOR U38734 ( .A(n31529), .B(n38968), .Z(n38956) );
  XNOR U38735 ( .A(n32586), .B(n33511), .Z(n38968) );
  XNOR U38736 ( .A(n38969), .B(n34149), .Z(n33511) );
  XNOR U38737 ( .A(n38719), .B(n38970), .Z(n34149) );
  ANDN U38738 ( .B(n35076), .A(n33320), .Z(n38969) );
  XOR U38739 ( .A(n38971), .B(n38972), .Z(n33320) );
  XNOR U38740 ( .A(n38973), .B(n36439), .Z(n35076) );
  XNOR U38741 ( .A(n38974), .B(n34146), .Z(n32586) );
  XOR U38742 ( .A(n38817), .B(n38975), .Z(n34146) );
  ANDN U38743 ( .B(n33313), .A(n35592), .Z(n38974) );
  XOR U38744 ( .A(n38976), .B(n38977), .Z(n35592) );
  XNOR U38745 ( .A(n38978), .B(n38530), .Z(n33313) );
  XNOR U38746 ( .A(n38979), .B(n34154), .Z(n31529) );
  XOR U38747 ( .A(n38980), .B(n35320), .Z(n34154) );
  XNOR U38748 ( .A(n38981), .B(n38982), .Z(n35320) );
  ANDN U38749 ( .B(n33546), .A(n35588), .Z(n38979) );
  XOR U38750 ( .A(n38983), .B(n36779), .Z(n35588) );
  XOR U38751 ( .A(n38984), .B(n38985), .Z(n33546) );
  XNOR U38752 ( .A(n30644), .B(n38986), .Z(n30396) );
  XNOR U38753 ( .A(n35656), .B(n38987), .Z(n30644) );
  XOR U38754 ( .A(n38988), .B(n38989), .Z(n35656) );
  XNOR U38755 ( .A(n33959), .B(n33471), .Z(n38989) );
  XNOR U38756 ( .A(n38990), .B(n36574), .Z(n33471) );
  XOR U38757 ( .A(n38991), .B(n38090), .Z(n36574) );
  IV U38758 ( .A(n37008), .Z(n38090) );
  ANDN U38759 ( .B(n35257), .A(n36573), .Z(n38990) );
  XOR U38760 ( .A(n38992), .B(n35627), .Z(n36573) );
  XNOR U38761 ( .A(n38993), .B(n37114), .Z(n35257) );
  XNOR U38762 ( .A(n38994), .B(n36576), .Z(n33959) );
  XOR U38763 ( .A(n38995), .B(n36557), .Z(n36576) );
  IV U38764 ( .A(n38082), .Z(n36557) );
  XOR U38765 ( .A(n38996), .B(n38997), .Z(n36577) );
  XOR U38766 ( .A(n38998), .B(n38401), .Z(n35262) );
  XOR U38767 ( .A(n33358), .B(n38999), .Z(n38988) );
  XOR U38768 ( .A(n32553), .B(n30650), .Z(n38999) );
  XNOR U38769 ( .A(n39000), .B(n36568), .Z(n30650) );
  XNOR U38770 ( .A(n39001), .B(n39002), .Z(n36568) );
  ANDN U38771 ( .B(n35270), .A(n37760), .Z(n39000) );
  XOR U38772 ( .A(n39003), .B(n37776), .Z(n37760) );
  XOR U38773 ( .A(n39004), .B(n37000), .Z(n35270) );
  XNOR U38774 ( .A(n39005), .B(n38512), .Z(n32553) );
  XOR U38775 ( .A(n39006), .B(n37510), .Z(n38512) );
  IV U38776 ( .A(n38843), .Z(n37510) );
  XOR U38777 ( .A(n39007), .B(n37859), .Z(n37762) );
  IV U38778 ( .A(n36996), .Z(n37859) );
  XOR U38779 ( .A(n39008), .B(n37267), .Z(n35253) );
  XNOR U38780 ( .A(n39009), .B(n36565), .Z(n33358) );
  NOR U38781 ( .A(n35266), .B(n36566), .Z(n39009) );
  XNOR U38782 ( .A(n39011), .B(n39012), .Z(n36566) );
  XOR U38783 ( .A(n39013), .B(n39014), .Z(n35266) );
  XOR U38784 ( .A(n36605), .B(n32449), .Z(n31442) );
  IV U38785 ( .A(n28982), .Z(n32449) );
  XNOR U38786 ( .A(n39015), .B(n39016), .Z(n38226) );
  XNOR U38787 ( .A(n30782), .B(n31832), .Z(n39016) );
  XNOR U38788 ( .A(n39017), .B(n35405), .Z(n31832) );
  IV U38789 ( .A(n39018), .Z(n35405) );
  ANDN U38790 ( .B(n35406), .A(n36599), .Z(n39017) );
  XOR U38791 ( .A(n39019), .B(n39020), .Z(n36599) );
  XNOR U38792 ( .A(n39021), .B(n39022), .Z(n35406) );
  XOR U38793 ( .A(n39023), .B(n35418), .Z(n30782) );
  AND U38794 ( .A(n36611), .B(n35419), .Z(n39023) );
  XOR U38795 ( .A(n39024), .B(n39025), .Z(n35419) );
  XNOR U38796 ( .A(n39026), .B(n38997), .Z(n36611) );
  XNOR U38797 ( .A(n34175), .B(n39027), .Z(n39015) );
  XOR U38798 ( .A(n30812), .B(n30993), .Z(n39027) );
  XOR U38799 ( .A(n39028), .B(n37387), .Z(n30993) );
  ANDN U38800 ( .B(n37388), .A(n38198), .Z(n39028) );
  XOR U38801 ( .A(n39029), .B(n35414), .Z(n30812) );
  ANDN U38802 ( .B(n35415), .A(n38196), .Z(n39029) );
  IV U38803 ( .A(n36608), .Z(n38196) );
  XNOR U38804 ( .A(n39030), .B(n36434), .Z(n36608) );
  XOR U38805 ( .A(n39031), .B(n39032), .Z(n35415) );
  XOR U38806 ( .A(n39033), .B(n35410), .Z(n34175) );
  ANDN U38807 ( .B(n35411), .A(n38192), .Z(n39033) );
  IV U38808 ( .A(n36603), .Z(n38192) );
  XOR U38809 ( .A(n39034), .B(n38865), .Z(n36603) );
  XOR U38810 ( .A(n39035), .B(n36946), .Z(n35411) );
  XNOR U38811 ( .A(n39036), .B(n39037), .Z(n33736) );
  XNOR U38812 ( .A(n32991), .B(n33370), .Z(n39037) );
  XNOR U38813 ( .A(n39038), .B(n37225), .Z(n33370) );
  ANDN U38814 ( .B(n36632), .A(n36633), .Z(n39038) );
  XNOR U38815 ( .A(n39039), .B(n38896), .Z(n36632) );
  XOR U38816 ( .A(n39040), .B(n37228), .Z(n32991) );
  ANDN U38817 ( .B(n36628), .A(n36629), .Z(n39040) );
  XOR U38818 ( .A(n39041), .B(n39031), .Z(n36628) );
  XNOR U38819 ( .A(n33264), .B(n39042), .Z(n39036) );
  XOR U38820 ( .A(n35845), .B(n37199), .Z(n39042) );
  XOR U38821 ( .A(n39043), .B(n39044), .Z(n37199) );
  ANDN U38822 ( .B(n36619), .A(n39045), .Z(n39043) );
  XNOR U38823 ( .A(n39046), .B(n37233), .Z(n35845) );
  ANDN U38824 ( .B(n36615), .A(n36616), .Z(n39046) );
  XNOR U38825 ( .A(n39047), .B(n37172), .Z(n36615) );
  XOR U38826 ( .A(n39048), .B(n37236), .Z(n33264) );
  ANDN U38827 ( .B(n36624), .A(n39049), .Z(n39048) );
  XOR U38828 ( .A(n39050), .B(n39051), .Z(n36624) );
  XNOR U38829 ( .A(n39052), .B(n37388), .Z(n36605) );
  XOR U38830 ( .A(n39053), .B(n36390), .Z(n37388) );
  ANDN U38831 ( .B(n38198), .A(n38199), .Z(n39052) );
  XNOR U38832 ( .A(n39054), .B(n39055), .Z(n38198) );
  XNOR U38833 ( .A(n39056), .B(n29479), .Z(n25970) );
  XOR U38834 ( .A(n31588), .B(n38109), .Z(n29479) );
  XOR U38835 ( .A(n39057), .B(n37597), .Z(n38109) );
  ANDN U38836 ( .B(n32637), .A(n33257), .Z(n39057) );
  XOR U38837 ( .A(n39058), .B(n36794), .Z(n32637) );
  XOR U38838 ( .A(n34770), .B(n34799), .Z(n31588) );
  XNOR U38839 ( .A(n39059), .B(n39060), .Z(n34799) );
  XNOR U38840 ( .A(n34438), .B(n31245), .Z(n39060) );
  XNOR U38841 ( .A(n39061), .B(n37598), .Z(n31245) );
  XOR U38842 ( .A(n39062), .B(n35366), .Z(n37598) );
  ANDN U38843 ( .B(n33257), .A(n37597), .Z(n39061) );
  XNOR U38844 ( .A(n38985), .B(n39063), .Z(n37597) );
  XOR U38845 ( .A(n36550), .B(n39064), .Z(n33257) );
  XNOR U38846 ( .A(n39065), .B(n32433), .Z(n34438) );
  XOR U38847 ( .A(n39066), .B(n37144), .Z(n32433) );
  XOR U38848 ( .A(n39067), .B(n39068), .Z(n37594) );
  XOR U38849 ( .A(n39069), .B(n38820), .Z(n33248) );
  XOR U38850 ( .A(n37588), .B(n39070), .Z(n39059) );
  XNOR U38851 ( .A(n31126), .B(n31231), .Z(n39070) );
  XNOR U38852 ( .A(n39071), .B(n37604), .Z(n31231) );
  XOR U38853 ( .A(n39072), .B(n37800), .Z(n37604) );
  IV U38854 ( .A(n38526), .Z(n37800) );
  ANDN U38855 ( .B(n33255), .A(n37603), .Z(n39071) );
  XOR U38856 ( .A(n39073), .B(n38491), .Z(n37603) );
  XNOR U38857 ( .A(n39074), .B(n37776), .Z(n33255) );
  XOR U38858 ( .A(n39075), .B(n39076), .Z(n37776) );
  XNOR U38859 ( .A(n39077), .B(n32857), .Z(n31126) );
  XOR U38860 ( .A(n39078), .B(n36717), .Z(n32857) );
  ANDN U38861 ( .B(n37607), .A(n33253), .Z(n39077) );
  XNOR U38862 ( .A(n39079), .B(n37646), .Z(n33253) );
  XNOR U38863 ( .A(n39080), .B(n37027), .Z(n37607) );
  XNOR U38864 ( .A(n39081), .B(n33120), .Z(n37588) );
  XOR U38865 ( .A(n35519), .B(n39082), .Z(n33120) );
  ANDN U38866 ( .B(n33250), .A(n37611), .Z(n39081) );
  XOR U38867 ( .A(n37431), .B(n39083), .Z(n37611) );
  XOR U38868 ( .A(n39084), .B(n37848), .Z(n33250) );
  XOR U38869 ( .A(n39085), .B(n39086), .Z(n34770) );
  XOR U38870 ( .A(n34527), .B(n32010), .Z(n39086) );
  XNOR U38871 ( .A(n39087), .B(n35973), .Z(n32010) );
  IV U38872 ( .A(n37619), .Z(n35973) );
  XOR U38873 ( .A(n39088), .B(n39089), .Z(n37619) );
  NOR U38874 ( .A(n36991), .B(n36990), .Z(n39087) );
  XNOR U38875 ( .A(n39090), .B(n37714), .Z(n36990) );
  XOR U38876 ( .A(n38113), .B(n39091), .Z(n36991) );
  XNOR U38877 ( .A(n39092), .B(n35967), .Z(n34527) );
  XNOR U38878 ( .A(n39093), .B(n37789), .Z(n35967) );
  NOR U38879 ( .A(n33110), .B(n36974), .Z(n39092) );
  XNOR U38880 ( .A(n39094), .B(n37000), .Z(n36974) );
  XNOR U38881 ( .A(n39095), .B(n37525), .Z(n33110) );
  XOR U38882 ( .A(n33182), .B(n39096), .Z(n39085) );
  XOR U38883 ( .A(n33205), .B(n31679), .Z(n39096) );
  XNOR U38884 ( .A(n39097), .B(n35964), .Z(n31679) );
  XOR U38885 ( .A(n39098), .B(n39099), .Z(n35964) );
  NOR U38886 ( .A(n36983), .B(n33104), .Z(n39097) );
  XNOR U38887 ( .A(n39100), .B(n37707), .Z(n33104) );
  IV U38888 ( .A(n37627), .Z(n36983) );
  XOR U38889 ( .A(n39101), .B(n39102), .Z(n37627) );
  XNOR U38890 ( .A(n39103), .B(n35961), .Z(n33205) );
  XOR U38891 ( .A(n39104), .B(n36996), .Z(n35961) );
  XOR U38892 ( .A(n39105), .B(n39106), .Z(n36996) );
  ANDN U38893 ( .B(n35214), .A(n36986), .Z(n39103) );
  XNOR U38894 ( .A(n39107), .B(n35778), .Z(n36986) );
  XOR U38895 ( .A(n39108), .B(n38878), .Z(n35214) );
  XNOR U38896 ( .A(n39111), .B(n35969), .Z(n33182) );
  XOR U38897 ( .A(n39112), .B(n39113), .Z(n35969) );
  NOR U38898 ( .A(n36978), .B(n33114), .Z(n39111) );
  XOR U38899 ( .A(n34628), .B(n39114), .Z(n33114) );
  IV U38900 ( .A(n37616), .Z(n36978) );
  XOR U38901 ( .A(n39115), .B(n38248), .Z(n37616) );
  ANDN U38902 ( .B(n30392), .A(n31432), .Z(n39056) );
  XOR U38903 ( .A(n34561), .B(n31169), .Z(n31432) );
  IV U38904 ( .A(n29519), .Z(n31169) );
  XNOR U38905 ( .A(n32712), .B(n32986), .Z(n29519) );
  XNOR U38906 ( .A(n39116), .B(n39117), .Z(n32986) );
  XNOR U38907 ( .A(n31993), .B(n31569), .Z(n39117) );
  XOR U38908 ( .A(n39118), .B(n34340), .Z(n31569) );
  XNOR U38909 ( .A(n39119), .B(n35940), .Z(n34340) );
  AND U38910 ( .A(n34568), .B(n34341), .Z(n39118) );
  XNOR U38911 ( .A(n39120), .B(n38352), .Z(n34341) );
  XOR U38912 ( .A(n39121), .B(n39122), .Z(n34568) );
  XOR U38913 ( .A(n39123), .B(n34331), .Z(n31993) );
  XOR U38914 ( .A(n39124), .B(n39125), .Z(n34331) );
  ANDN U38915 ( .B(n34332), .A(n36773), .Z(n39123) );
  XOR U38916 ( .A(n28991), .B(n39126), .Z(n39116) );
  XNOR U38917 ( .A(n34116), .B(n31070), .Z(n39126) );
  XNOR U38918 ( .A(n39127), .B(n34344), .Z(n31070) );
  XOR U38919 ( .A(n39128), .B(n35778), .Z(n34344) );
  ANDN U38920 ( .B(n34345), .A(n34564), .Z(n39127) );
  XOR U38921 ( .A(n39129), .B(n38374), .Z(n34564) );
  XOR U38922 ( .A(n35583), .B(n39130), .Z(n34345) );
  XOR U38923 ( .A(n39131), .B(n34348), .Z(n34116) );
  XOR U38924 ( .A(n34618), .B(n39132), .Z(n34348) );
  AND U38925 ( .A(n34571), .B(n34349), .Z(n39131) );
  XOR U38926 ( .A(n39133), .B(n37331), .Z(n34349) );
  XOR U38927 ( .A(n39134), .B(n35938), .Z(n34571) );
  XNOR U38928 ( .A(n39135), .B(n34335), .Z(n28991) );
  XNOR U38929 ( .A(n39136), .B(n33917), .Z(n34335) );
  ANDN U38930 ( .B(n34336), .A(n36766), .Z(n39135) );
  IV U38931 ( .A(n34574), .Z(n36766) );
  XOR U38932 ( .A(n39137), .B(n37789), .Z(n34574) );
  XNOR U38933 ( .A(n39138), .B(n38096), .Z(n34336) );
  XOR U38934 ( .A(n39139), .B(n39140), .Z(n32712) );
  XOR U38935 ( .A(n31961), .B(n30001), .Z(n39140) );
  XNOR U38936 ( .A(n39141), .B(n35223), .Z(n30001) );
  AND U38937 ( .A(n34546), .B(n34544), .Z(n39141) );
  XNOR U38938 ( .A(n39142), .B(n38544), .Z(n34544) );
  XOR U38939 ( .A(n39143), .B(n34123), .Z(n31961) );
  XNOR U38940 ( .A(n39144), .B(n38149), .Z(n34123) );
  ANDN U38941 ( .B(n34124), .A(n39145), .Z(n39143) );
  XOR U38942 ( .A(n39146), .B(n35625), .Z(n34124) );
  XOR U38943 ( .A(n32460), .B(n39147), .Z(n39139) );
  XNOR U38944 ( .A(n30819), .B(n31387), .Z(n39147) );
  XOR U38945 ( .A(n39148), .B(n35982), .Z(n31387) );
  XOR U38946 ( .A(n38801), .B(n39149), .Z(n35982) );
  XNOR U38947 ( .A(n39121), .B(n39150), .Z(n34556) );
  XOR U38948 ( .A(n39151), .B(n34130), .Z(n30819) );
  XOR U38949 ( .A(n39152), .B(n39153), .Z(n34130) );
  XNOR U38950 ( .A(n39154), .B(n36946), .Z(n34131) );
  XNOR U38951 ( .A(n39157), .B(n34902), .Z(n32460) );
  XOR U38952 ( .A(n39158), .B(n39159), .Z(n34902) );
  AND U38953 ( .A(n34553), .B(n34552), .Z(n39157) );
  XOR U38954 ( .A(n39160), .B(n39161), .Z(n34552) );
  XNOR U38955 ( .A(n39162), .B(n34332), .Z(n34561) );
  XOR U38956 ( .A(n39163), .B(n36417), .Z(n34332) );
  ANDN U38957 ( .B(n36773), .A(n36774), .Z(n39162) );
  XOR U38958 ( .A(n37786), .B(n39164), .Z(n36774) );
  IV U38959 ( .A(n39165), .Z(n37786) );
  XNOR U38960 ( .A(n39166), .B(n36976), .Z(n36773) );
  XOR U38961 ( .A(n35492), .B(n30671), .Z(n30392) );
  IV U38962 ( .A(n32018), .Z(n30671) );
  XNOR U38963 ( .A(n39167), .B(n39168), .Z(n33270) );
  XNOR U38964 ( .A(n34362), .B(n35750), .Z(n39168) );
  XOR U38965 ( .A(n39169), .B(n35763), .Z(n35750) );
  XOR U38966 ( .A(n39170), .B(n38642), .Z(n35763) );
  ANDN U38967 ( .B(n35485), .A(n34315), .Z(n39169) );
  XNOR U38968 ( .A(n39171), .B(n39172), .Z(n34315) );
  XNOR U38969 ( .A(n39173), .B(n35579), .Z(n35485) );
  XOR U38970 ( .A(n39174), .B(n35756), .Z(n34362) );
  XNOR U38971 ( .A(n39175), .B(n39176), .Z(n35756) );
  NOR U38972 ( .A(n34302), .B(n35487), .Z(n39174) );
  XOR U38973 ( .A(n39177), .B(n37535), .Z(n35487) );
  XNOR U38974 ( .A(n39178), .B(n36359), .Z(n34302) );
  XOR U38975 ( .A(n33943), .B(n39181), .Z(n39167) );
  XOR U38976 ( .A(n32730), .B(n32035), .Z(n39181) );
  XNOR U38977 ( .A(n39182), .B(n35761), .Z(n32035) );
  XOR U38978 ( .A(n35933), .B(n39183), .Z(n35761) );
  IV U38979 ( .A(n39184), .Z(n35933) );
  ANDN U38980 ( .B(n35482), .A(n34298), .Z(n39182) );
  XOR U38981 ( .A(n39185), .B(n39186), .Z(n34298) );
  XOR U38982 ( .A(n39187), .B(n38777), .Z(n35482) );
  XNOR U38983 ( .A(n39188), .B(n35759), .Z(n32730) );
  XNOR U38984 ( .A(n38126), .B(n39189), .Z(n35759) );
  ANDN U38985 ( .B(n35480), .A(n34307), .Z(n39188) );
  XNOR U38986 ( .A(n39190), .B(n35613), .Z(n34307) );
  IV U38987 ( .A(n38637), .Z(n35613) );
  XOR U38988 ( .A(n39191), .B(n39156), .Z(n38637) );
  XOR U38989 ( .A(n39192), .B(n39193), .Z(n39156) );
  XOR U38990 ( .A(n37938), .B(n38138), .Z(n39193) );
  XOR U38991 ( .A(n39194), .B(n39195), .Z(n38138) );
  XNOR U38992 ( .A(n39198), .B(n39199), .Z(n37938) );
  ANDN U38993 ( .B(n39200), .A(n39201), .Z(n39198) );
  XOR U38994 ( .A(n39202), .B(n39203), .Z(n39192) );
  XOR U38995 ( .A(n39204), .B(n37024), .Z(n39203) );
  XNOR U38996 ( .A(n39205), .B(n39206), .Z(n37024) );
  ANDN U38997 ( .B(n39207), .A(n39208), .Z(n39205) );
  XOR U38998 ( .A(n39209), .B(n37851), .Z(n35480) );
  XOR U38999 ( .A(n39210), .B(n38322), .Z(n33943) );
  XOR U39000 ( .A(n38242), .B(n39211), .Z(n38322) );
  ANDN U39001 ( .B(n35489), .A(n34311), .Z(n39210) );
  XOR U39002 ( .A(n39212), .B(n39213), .Z(n34311) );
  XOR U39003 ( .A(n39011), .B(n39214), .Z(n35489) );
  XNOR U39004 ( .A(n39215), .B(n39216), .Z(n35957) );
  XNOR U39005 ( .A(n33605), .B(n28804), .Z(n39216) );
  XOR U39006 ( .A(n39217), .B(n33686), .Z(n28804) );
  XOR U39007 ( .A(n39218), .B(n39219), .Z(n33686) );
  NOR U39008 ( .A(n34782), .B(n33687), .Z(n39217) );
  XOR U39009 ( .A(n39220), .B(n37272), .Z(n33687) );
  XOR U39010 ( .A(n39221), .B(n35617), .Z(n34782) );
  IV U39011 ( .A(n38093), .Z(n35617) );
  XOR U39012 ( .A(n39222), .B(n39223), .Z(n38093) );
  XNOR U39013 ( .A(n39224), .B(n34183), .Z(n33605) );
  XNOR U39014 ( .A(n38176), .B(n39225), .Z(n34183) );
  ANDN U39015 ( .B(n34182), .A(n34779), .Z(n39224) );
  XOR U39016 ( .A(n39226), .B(n39227), .Z(n34779) );
  XOR U39017 ( .A(n39228), .B(n39176), .Z(n34182) );
  XNOR U39018 ( .A(n32227), .B(n39229), .Z(n39215) );
  XOR U39019 ( .A(n33674), .B(n32155), .Z(n39229) );
  XOR U39020 ( .A(n39230), .B(n33690), .Z(n32155) );
  XNOR U39021 ( .A(n39231), .B(n37040), .Z(n33690) );
  ANDN U39022 ( .B(n34785), .A(n39232), .Z(n39230) );
  XOR U39023 ( .A(n39233), .B(n33695), .Z(n33674) );
  XOR U39024 ( .A(n39234), .B(n37851), .Z(n33695) );
  XOR U39025 ( .A(n39235), .B(n39236), .Z(n37851) );
  ANDN U39026 ( .B(n33694), .A(n35475), .Z(n39233) );
  XOR U39027 ( .A(n39237), .B(n39238), .Z(n35475) );
  XOR U39028 ( .A(n39240), .B(n33681), .Z(n32227) );
  XOR U39029 ( .A(n38033), .B(n39241), .Z(n33681) );
  ANDN U39030 ( .B(n33682), .A(n34775), .Z(n39240) );
  XOR U39031 ( .A(n39243), .B(n35625), .Z(n33682) );
  XNOR U39032 ( .A(n39244), .B(n33691), .Z(n35492) );
  IV U39033 ( .A(n39232), .Z(n33691) );
  XOR U39034 ( .A(n39245), .B(n38777), .Z(n39232) );
  ANDN U39035 ( .B(n34786), .A(n34785), .Z(n39244) );
  XOR U39036 ( .A(n39246), .B(n39247), .Z(n34785) );
  XOR U39037 ( .A(n38604), .B(n39248), .Z(n34786) );
  IV U39038 ( .A(n38801), .Z(n38604) );
  XNOR U39039 ( .A(n39249), .B(n31773), .Z(n31436) );
  XOR U39040 ( .A(n38597), .B(n31054), .Z(n31773) );
  XOR U39041 ( .A(n33993), .B(n33331), .Z(n31054) );
  XNOR U39042 ( .A(n39250), .B(n39251), .Z(n33331) );
  XNOR U39043 ( .A(n36694), .B(n29926), .Z(n39251) );
  XNOR U39044 ( .A(n39252), .B(n36724), .Z(n29926) );
  XOR U39045 ( .A(n39253), .B(n37434), .Z(n36724) );
  IV U39046 ( .A(n36219), .Z(n37434) );
  NOR U39047 ( .A(n37478), .B(n36723), .Z(n39252) );
  XNOR U39048 ( .A(n39254), .B(n39255), .Z(n36723) );
  XNOR U39049 ( .A(n39256), .B(n38080), .Z(n37478) );
  XOR U39050 ( .A(n39257), .B(n37132), .Z(n36694) );
  XOR U39051 ( .A(n39258), .B(n39259), .Z(n37132) );
  ANDN U39052 ( .B(n37470), .A(n37155), .Z(n39257) );
  XOR U39053 ( .A(n37890), .B(n39260), .Z(n37155) );
  XOR U39054 ( .A(n39261), .B(n39262), .Z(n37470) );
  XOR U39055 ( .A(n32092), .B(n39263), .Z(n39250) );
  XOR U39056 ( .A(n36152), .B(n30737), .Z(n39263) );
  XNOR U39057 ( .A(n39264), .B(n36729), .Z(n30737) );
  XNOR U39058 ( .A(n38858), .B(n39265), .Z(n36729) );
  NOR U39059 ( .A(n37482), .B(n36728), .Z(n39264) );
  XOR U39060 ( .A(n39266), .B(n39267), .Z(n36728) );
  XOR U39061 ( .A(n39268), .B(n39269), .Z(n37482) );
  XNOR U39062 ( .A(n39270), .B(n36732), .Z(n36152) );
  XNOR U39063 ( .A(n38181), .B(n39271), .Z(n36732) );
  ANDN U39064 ( .B(n36733), .A(n37485), .Z(n39270) );
  XOR U39065 ( .A(n39011), .B(n39272), .Z(n37485) );
  XOR U39066 ( .A(n38684), .B(n39273), .Z(n36733) );
  XNOR U39067 ( .A(n39274), .B(n36736), .Z(n32092) );
  XOR U39068 ( .A(n39275), .B(n36907), .Z(n36736) );
  NOR U39069 ( .A(n37474), .B(n36737), .Z(n39274) );
  XOR U39070 ( .A(n39276), .B(n38457), .Z(n36737) );
  IV U39071 ( .A(n39219), .Z(n38457) );
  XOR U39072 ( .A(n39277), .B(n39278), .Z(n37474) );
  XOR U39073 ( .A(n39279), .B(n39280), .Z(n33993) );
  XOR U39074 ( .A(n32246), .B(n32825), .Z(n39280) );
  XOR U39075 ( .A(n39281), .B(n37288), .Z(n32825) );
  XNOR U39076 ( .A(n38181), .B(n39282), .Z(n37288) );
  ANDN U39077 ( .B(n37289), .A(n36082), .Z(n39281) );
  XOR U39078 ( .A(n39283), .B(n39284), .Z(n36082) );
  XOR U39079 ( .A(n38891), .B(n39285), .Z(n37289) );
  IV U39080 ( .A(n38906), .Z(n38891) );
  XNOR U39081 ( .A(n39286), .B(n37286), .Z(n32246) );
  XOR U39082 ( .A(n39287), .B(n37055), .Z(n37286) );
  AND U39083 ( .A(n38599), .B(n37285), .Z(n39286) );
  XNOR U39084 ( .A(n39288), .B(n37887), .Z(n37285) );
  XNOR U39085 ( .A(n39289), .B(n35516), .Z(n38599) );
  IV U39086 ( .A(n38024), .Z(n35516) );
  XOR U39087 ( .A(n39290), .B(n39291), .Z(n38024) );
  XOR U39088 ( .A(n29257), .B(n39292), .Z(n39279) );
  XOR U39089 ( .A(n33375), .B(n32204), .Z(n39292) );
  XOR U39090 ( .A(n39293), .B(n37281), .Z(n32204) );
  XOR U39091 ( .A(n39294), .B(n37081), .Z(n37281) );
  IV U39092 ( .A(n39295), .Z(n37081) );
  XOR U39093 ( .A(n38948), .B(n39296), .Z(n36072) );
  XNOR U39094 ( .A(n37431), .B(n39297), .Z(n37280) );
  IV U39095 ( .A(n39031), .Z(n37431) );
  XNOR U39096 ( .A(n39298), .B(n39299), .Z(n39031) );
  XOR U39097 ( .A(n39300), .B(n37292), .Z(n33375) );
  XNOR U39098 ( .A(n39301), .B(n35627), .Z(n37292) );
  ANDN U39099 ( .B(n36076), .A(n38592), .Z(n39300) );
  IV U39100 ( .A(n37293), .Z(n38592) );
  XNOR U39101 ( .A(n39302), .B(n38169), .Z(n37293) );
  XOR U39102 ( .A(n39303), .B(n39304), .Z(n36076) );
  XOR U39103 ( .A(n39305), .B(n37277), .Z(n29257) );
  XOR U39104 ( .A(n39306), .B(n39307), .Z(n37277) );
  ANDN U39105 ( .B(n37278), .A(n36086), .Z(n39305) );
  XNOR U39106 ( .A(n39308), .B(n37278), .Z(n38597) );
  XNOR U39107 ( .A(n38030), .B(n39309), .Z(n37278) );
  IV U39108 ( .A(n36413), .Z(n38030) );
  ANDN U39109 ( .B(n36086), .A(n36087), .Z(n39308) );
  XNOR U39110 ( .A(n39310), .B(n39099), .Z(n36087) );
  XOR U39111 ( .A(n39311), .B(n39312), .Z(n36086) );
  ANDN U39112 ( .B(n30399), .A(n30398), .Z(n39249) );
  XNOR U39113 ( .A(n28807), .B(n36830), .Z(n30398) );
  XOR U39114 ( .A(n39313), .B(n39314), .Z(n36830) );
  ANDN U39115 ( .B(n38749), .A(n35897), .Z(n39313) );
  XNOR U39116 ( .A(n39315), .B(n39316), .Z(n35897) );
  XNOR U39117 ( .A(n34431), .B(n32864), .Z(n28807) );
  XOR U39118 ( .A(n39317), .B(n39318), .Z(n32864) );
  XOR U39119 ( .A(n31110), .B(n32695), .Z(n39318) );
  XNOR U39120 ( .A(n39319), .B(n33392), .Z(n32695) );
  XOR U39121 ( .A(n39320), .B(n36353), .Z(n33392) );
  ANDN U39122 ( .B(n33393), .A(n33785), .Z(n39319) );
  XOR U39123 ( .A(n39321), .B(n38343), .Z(n33785) );
  XOR U39124 ( .A(n39322), .B(n36701), .Z(n33393) );
  XOR U39125 ( .A(n39323), .B(n35357), .Z(n31110) );
  ANDN U39126 ( .B(n33794), .A(n33792), .Z(n39323) );
  XOR U39127 ( .A(n39325), .B(n39326), .Z(n33792) );
  XNOR U39128 ( .A(n39327), .B(n39328), .Z(n33794) );
  XNOR U39129 ( .A(n33385), .B(n39329), .Z(n39317) );
  XNOR U39130 ( .A(n33129), .B(n30783), .Z(n39329) );
  XNOR U39131 ( .A(n39330), .B(n33398), .Z(n30783) );
  XOR U39132 ( .A(n39331), .B(n37427), .Z(n33398) );
  ANDN U39133 ( .B(n33399), .A(n36226), .Z(n39330) );
  XOR U39134 ( .A(n37679), .B(n39332), .Z(n36226) );
  XNOR U39135 ( .A(n39333), .B(n38997), .Z(n33399) );
  XNOR U39136 ( .A(n39334), .B(n38629), .Z(n33129) );
  XOR U39137 ( .A(n39335), .B(n35093), .Z(n38629) );
  ANDN U39138 ( .B(n33782), .A(n38648), .Z(n39334) );
  IV U39139 ( .A(n33781), .Z(n38648) );
  XOR U39140 ( .A(n39336), .B(n39337), .Z(n33781) );
  IV U39141 ( .A(n36231), .Z(n33782) );
  XOR U39142 ( .A(n39338), .B(n36351), .Z(n36231) );
  XNOR U39143 ( .A(n39339), .B(n33403), .Z(n33385) );
  XNOR U39144 ( .A(n39340), .B(n38176), .Z(n33403) );
  XOR U39145 ( .A(n39341), .B(n39342), .Z(n33402) );
  XNOR U39146 ( .A(n39343), .B(n39344), .Z(n33790) );
  XOR U39147 ( .A(n39345), .B(n39346), .Z(n34431) );
  XOR U39148 ( .A(n31974), .B(n32740), .Z(n39346) );
  XNOR U39149 ( .A(n39347), .B(n35913), .Z(n32740) );
  NOR U39150 ( .A(n36835), .B(n36836), .Z(n39347) );
  XOR U39151 ( .A(n39348), .B(n39113), .Z(n36836) );
  XOR U39152 ( .A(n39349), .B(n35908), .Z(n31974) );
  NOR U39153 ( .A(n36827), .B(n36828), .Z(n39349) );
  XOR U39154 ( .A(n39160), .B(n39350), .Z(n36828) );
  IV U39155 ( .A(n38320), .Z(n39160) );
  IV U39156 ( .A(n39351), .Z(n36827) );
  XNOR U39157 ( .A(n31708), .B(n39352), .Z(n39345) );
  XOR U39158 ( .A(n31582), .B(n30104), .Z(n39352) );
  XNOR U39159 ( .A(n39353), .B(n35899), .Z(n30104) );
  ANDN U39160 ( .B(n39314), .A(n38749), .Z(n39353) );
  XNOR U39161 ( .A(n39354), .B(n35619), .Z(n38749) );
  XNOR U39162 ( .A(n39357), .B(n35902), .Z(n31582) );
  ANDN U39163 ( .B(n36832), .A(n36833), .Z(n39357) );
  XOR U39164 ( .A(n39358), .B(n36393), .Z(n36833) );
  XOR U39165 ( .A(n39359), .B(n36237), .Z(n31708) );
  IV U39166 ( .A(n39360), .Z(n36237) );
  ANDN U39167 ( .B(n36824), .A(n36825), .Z(n39359) );
  XOR U39168 ( .A(n39361), .B(n37497), .Z(n36825) );
  IV U39169 ( .A(n37076), .Z(n37497) );
  XOR U39170 ( .A(n39362), .B(n39363), .Z(n37076) );
  IV U39171 ( .A(n29482), .Z(n30399) );
  XNOR U39172 ( .A(n30253), .B(n37942), .Z(n29482) );
  XNOR U39173 ( .A(n39364), .B(n33662), .Z(n37942) );
  ANDN U39174 ( .B(n34895), .A(n34896), .Z(n39364) );
  XNOR U39175 ( .A(n35304), .B(n39365), .Z(n34896) );
  XOR U39176 ( .A(n35191), .B(n39366), .Z(n30253) );
  XOR U39177 ( .A(n39367), .B(n39368), .Z(n35191) );
  XNOR U39178 ( .A(n30529), .B(n33456), .Z(n39368) );
  XOR U39179 ( .A(n39369), .B(n35724), .Z(n33456) );
  IV U39180 ( .A(n39370), .Z(n35724) );
  NOR U39181 ( .A(n37578), .B(n35723), .Z(n39369) );
  XNOR U39182 ( .A(n39371), .B(n39372), .Z(n35723) );
  XNOR U39183 ( .A(n37868), .B(n39373), .Z(n37578) );
  XNOR U39184 ( .A(n39374), .B(n35728), .Z(n30529) );
  ANDN U39185 ( .B(n37570), .A(n35727), .Z(n39374) );
  XOR U39186 ( .A(n39375), .B(n36212), .Z(n35727) );
  XOR U39187 ( .A(n39376), .B(n37349), .Z(n37570) );
  XNOR U39188 ( .A(n35000), .B(n39377), .Z(n39367) );
  XNOR U39189 ( .A(n35710), .B(n34360), .Z(n39377) );
  XNOR U39190 ( .A(n39378), .B(n38650), .Z(n34360) );
  IV U39191 ( .A(n39379), .Z(n38650) );
  ANDN U39192 ( .B(n37818), .A(n37581), .Z(n39378) );
  XNOR U39193 ( .A(n35620), .B(n39380), .Z(n37581) );
  IV U39194 ( .A(n39315), .Z(n35620) );
  XNOR U39195 ( .A(n39381), .B(n39382), .Z(n37818) );
  XNOR U39196 ( .A(n39383), .B(n39384), .Z(n35710) );
  ANDN U39197 ( .B(n37821), .A(n37822), .Z(n39383) );
  XOR U39198 ( .A(n39385), .B(n35304), .Z(n37822) );
  XNOR U39199 ( .A(n39386), .B(n35718), .Z(n35000) );
  IV U39200 ( .A(n39387), .Z(n35718) );
  NOR U39201 ( .A(n35717), .B(n37573), .Z(n39386) );
  XOR U39202 ( .A(n39388), .B(n39389), .Z(n37573) );
  XNOR U39203 ( .A(n39390), .B(n39278), .Z(n35717) );
  XOR U39204 ( .A(n31293), .B(n27228), .Z(n23680) );
  XOR U39205 ( .A(n32346), .B(n29954), .Z(n27228) );
  XNOR U39206 ( .A(n39391), .B(n39392), .Z(n29954) );
  XNOR U39207 ( .A(n25578), .B(n28176), .Z(n39392) );
  XOR U39208 ( .A(n39393), .B(n28209), .Z(n28176) );
  XOR U39209 ( .A(n37653), .B(n32875), .Z(n28209) );
  IV U39210 ( .A(n30798), .Z(n32875) );
  XOR U39211 ( .A(n35920), .B(n34136), .Z(n30798) );
  XNOR U39212 ( .A(n39394), .B(n39395), .Z(n34136) );
  XNOR U39213 ( .A(n33773), .B(n34249), .Z(n39395) );
  XOR U39214 ( .A(n39396), .B(n34266), .Z(n34249) );
  ANDN U39215 ( .B(n33987), .A(n34265), .Z(n39396) );
  IV U39216 ( .A(n35698), .Z(n34265) );
  XOR U39217 ( .A(n39398), .B(n39399), .Z(n35698) );
  XNOR U39218 ( .A(n38176), .B(n39400), .Z(n33987) );
  XNOR U39219 ( .A(n39401), .B(n34262), .Z(n33773) );
  XOR U39220 ( .A(n39402), .B(n34623), .Z(n34262) );
  AND U39221 ( .A(n34263), .B(n33615), .Z(n39401) );
  XOR U39222 ( .A(n39403), .B(n39404), .Z(n33615) );
  XOR U39223 ( .A(n39405), .B(n39406), .Z(n34263) );
  XOR U39224 ( .A(n32632), .B(n39407), .Z(n39394) );
  XNOR U39225 ( .A(n31952), .B(n31460), .Z(n39407) );
  XNOR U39226 ( .A(n39408), .B(n34260), .Z(n31460) );
  XNOR U39227 ( .A(n39409), .B(n36907), .Z(n34260) );
  ANDN U39228 ( .B(n33625), .A(n34259), .Z(n39408) );
  XOR U39229 ( .A(n39410), .B(n36555), .Z(n34259) );
  XOR U39230 ( .A(n39411), .B(n37602), .Z(n33625) );
  XNOR U39231 ( .A(n39412), .B(n36348), .Z(n31952) );
  XOR U39232 ( .A(n39413), .B(n39414), .Z(n36348) );
  AND U39233 ( .A(n35700), .B(n34162), .Z(n39412) );
  XNOR U39234 ( .A(n38804), .B(n39415), .Z(n34162) );
  XNOR U39235 ( .A(n39416), .B(n37909), .Z(n35700) );
  IV U39236 ( .A(n37521), .Z(n37909) );
  XNOR U39237 ( .A(n39417), .B(n39418), .Z(n37521) );
  XNOR U39238 ( .A(n39419), .B(n34255), .Z(n32632) );
  XOR U39239 ( .A(n36987), .B(n39420), .Z(n34255) );
  AND U39240 ( .A(n34256), .B(n33621), .Z(n39419) );
  XOR U39241 ( .A(n38619), .B(n39421), .Z(n33621) );
  XNOR U39242 ( .A(n36303), .B(n39422), .Z(n34256) );
  XOR U39243 ( .A(n39423), .B(n39424), .Z(n35920) );
  XNOR U39244 ( .A(n32546), .B(n30664), .Z(n39424) );
  XNOR U39245 ( .A(n39425), .B(n34918), .Z(n30664) );
  XOR U39246 ( .A(n39426), .B(n38642), .Z(n34918) );
  AND U39247 ( .A(n37663), .B(n34919), .Z(n39425) );
  XOR U39248 ( .A(n39427), .B(n36393), .Z(n34919) );
  XNOR U39249 ( .A(n39428), .B(n34927), .Z(n32546) );
  XOR U39250 ( .A(n39001), .B(n39429), .Z(n34927) );
  AND U39251 ( .A(n34926), .B(n37659), .Z(n39428) );
  XOR U39252 ( .A(n39430), .B(n39431), .Z(n34926) );
  XNOR U39253 ( .A(n32932), .B(n39432), .Z(n39423) );
  XNOR U39254 ( .A(n30013), .B(n33219), .Z(n39432) );
  XOR U39255 ( .A(n39433), .B(n34923), .Z(n33219) );
  XOR U39256 ( .A(n39434), .B(n38807), .Z(n34923) );
  IV U39257 ( .A(n37797), .Z(n38807) );
  ANDN U39258 ( .B(n34922), .A(n39435), .Z(n39433) );
  XOR U39259 ( .A(n39436), .B(n34909), .Z(n30013) );
  XOR U39260 ( .A(n39437), .B(n37948), .Z(n34909) );
  IV U39261 ( .A(n38486), .Z(n37948) );
  ANDN U39262 ( .B(n34910), .A(n39438), .Z(n39436) );
  XNOR U39263 ( .A(n38619), .B(n39439), .Z(n34910) );
  XNOR U39264 ( .A(n39440), .B(n34914), .Z(n32932) );
  XNOR U39265 ( .A(n39441), .B(n38298), .Z(n34914) );
  ANDN U39266 ( .B(n37661), .A(n34913), .Z(n39440) );
  XOR U39267 ( .A(n39442), .B(n37008), .Z(n34913) );
  XNOR U39268 ( .A(n39443), .B(n34922), .Z(n37653) );
  XOR U39269 ( .A(n37875), .B(n39444), .Z(n34922) );
  NOR U39270 ( .A(n39445), .B(n36685), .Z(n39443) );
  ANDN U39271 ( .B(n28210), .A(n27598), .Z(n39393) );
  XNOR U39272 ( .A(n30961), .B(n35096), .Z(n27598) );
  XNOR U39273 ( .A(n39446), .B(n35953), .Z(n35096) );
  ANDN U39274 ( .B(n33441), .A(n39447), .Z(n39446) );
  XOR U39275 ( .A(n39448), .B(n39449), .Z(n33441) );
  XNOR U39276 ( .A(n38955), .B(n37829), .Z(n30961) );
  XNOR U39277 ( .A(n39450), .B(n39451), .Z(n37829) );
  XOR U39278 ( .A(n32218), .B(n32892), .Z(n39451) );
  XOR U39279 ( .A(n39452), .B(n35554), .Z(n32892) );
  XOR U39280 ( .A(n39453), .B(n39454), .Z(n35554) );
  XNOR U39281 ( .A(n39455), .B(n37051), .Z(n35555) );
  XOR U39282 ( .A(n39456), .B(n38912), .Z(n38289) );
  XNOR U39283 ( .A(n39457), .B(n35558), .Z(n32218) );
  XOR U39284 ( .A(n39458), .B(n38037), .Z(n35558) );
  XOR U39285 ( .A(n39459), .B(n35632), .Z(n35559) );
  XOR U39286 ( .A(n39460), .B(n37834), .Z(n35816) );
  XNOR U39287 ( .A(n32505), .B(n39461), .Z(n39450) );
  XNOR U39288 ( .A(n31854), .B(n32852), .Z(n39461) );
  XOR U39289 ( .A(n39462), .B(n35545), .Z(n32852) );
  XOR U39290 ( .A(n39463), .B(n35952), .Z(n35545) );
  ANDN U39291 ( .B(n35812), .A(n38281), .Z(n39462) );
  IV U39292 ( .A(n35546), .Z(n38281) );
  XOR U39293 ( .A(n39464), .B(n39025), .Z(n35546) );
  XNOR U39294 ( .A(n39465), .B(n35301), .Z(n35812) );
  XNOR U39295 ( .A(n39466), .B(n35550), .Z(n31854) );
  XOR U39296 ( .A(n39467), .B(n39468), .Z(n35550) );
  ANDN U39297 ( .B(n35551), .A(n35808), .Z(n39466) );
  XOR U39298 ( .A(n39469), .B(n39470), .Z(n35808) );
  XOR U39299 ( .A(n39471), .B(n38360), .Z(n35551) );
  XOR U39300 ( .A(n39472), .B(n36400), .Z(n32505) );
  XNOR U39301 ( .A(n39473), .B(n36537), .Z(n36400) );
  NOR U39302 ( .A(n38293), .B(n35819), .Z(n39472) );
  XNOR U39303 ( .A(n39474), .B(n39475), .Z(n35819) );
  XOR U39304 ( .A(n38518), .B(n39476), .Z(n38293) );
  XOR U39305 ( .A(n39477), .B(n39478), .Z(n38955) );
  XNOR U39306 ( .A(n31334), .B(n29716), .Z(n39478) );
  XOR U39307 ( .A(n39479), .B(n35533), .Z(n29716) );
  XOR U39308 ( .A(n39480), .B(n36369), .Z(n35533) );
  ANDN U39309 ( .B(n35103), .A(n33425), .Z(n39479) );
  XNOR U39310 ( .A(n39481), .B(n39482), .Z(n33425) );
  XOR U39311 ( .A(n39483), .B(n39484), .Z(n35103) );
  XNOR U39312 ( .A(n39485), .B(n35537), .Z(n31334) );
  XNOR U39313 ( .A(n39486), .B(n36541), .Z(n35537) );
  NOR U39314 ( .A(n33435), .B(n35098), .Z(n39485) );
  XNOR U39315 ( .A(n39487), .B(n35308), .Z(n35098) );
  XOR U39316 ( .A(n38961), .B(n39488), .Z(n33435) );
  XNOR U39317 ( .A(n35527), .B(n39489), .Z(n39477) );
  XOR U39318 ( .A(n32177), .B(n31735), .Z(n39489) );
  XNOR U39319 ( .A(n39490), .B(n35539), .Z(n31735) );
  XOR U39320 ( .A(n39491), .B(n37630), .Z(n35539) );
  ANDN U39321 ( .B(n35106), .A(n33429), .Z(n39490) );
  XOR U39322 ( .A(n39492), .B(n36522), .Z(n33429) );
  XNOR U39323 ( .A(n38619), .B(n39493), .Z(n35106) );
  XNOR U39324 ( .A(n39290), .B(n39494), .Z(n38619) );
  XOR U39325 ( .A(n39495), .B(n39496), .Z(n39290) );
  XOR U39326 ( .A(n38786), .B(n39497), .Z(n39496) );
  XNOR U39327 ( .A(n39498), .B(n39499), .Z(n38786) );
  ANDN U39328 ( .B(n39500), .A(n39501), .Z(n39498) );
  XOR U39329 ( .A(n38935), .B(n39502), .Z(n39495) );
  XOR U39330 ( .A(n37941), .B(n35791), .Z(n39502) );
  XOR U39331 ( .A(n39503), .B(n39504), .Z(n35791) );
  ANDN U39332 ( .B(n39505), .A(n39506), .Z(n39503) );
  XNOR U39333 ( .A(n39507), .B(n39508), .Z(n37941) );
  ANDN U39334 ( .B(n39509), .A(n39510), .Z(n39507) );
  XNOR U39335 ( .A(n39511), .B(n39512), .Z(n38935) );
  ANDN U39336 ( .B(n39513), .A(n39514), .Z(n39511) );
  XOR U39337 ( .A(n39515), .B(n35531), .Z(n32177) );
  XOR U39338 ( .A(n39516), .B(n39454), .Z(n35531) );
  ANDN U39339 ( .B(n35101), .A(n34172), .Z(n39515) );
  XOR U39340 ( .A(n39517), .B(n37420), .Z(n34172) );
  XOR U39341 ( .A(n36704), .B(n39518), .Z(n35101) );
  IV U39342 ( .A(n38535), .Z(n36704) );
  XNOR U39343 ( .A(n39519), .B(n35947), .Z(n35527) );
  XNOR U39344 ( .A(n37110), .B(n39520), .Z(n35947) );
  ANDN U39345 ( .B(n35953), .A(n33439), .Z(n39519) );
  IV U39346 ( .A(n39447), .Z(n33439) );
  XNOR U39347 ( .A(n39521), .B(n39278), .Z(n39447) );
  XOR U39348 ( .A(n39522), .B(n39523), .Z(n35953) );
  XOR U39349 ( .A(n34275), .B(n30559), .Z(n28210) );
  XNOR U39350 ( .A(n37065), .B(n33386), .Z(n30559) );
  XNOR U39351 ( .A(n39524), .B(n39525), .Z(n33386) );
  XNOR U39352 ( .A(n32606), .B(n33041), .Z(n39525) );
  XNOR U39353 ( .A(n39526), .B(n37111), .Z(n33041) );
  XOR U39354 ( .A(n39527), .B(n39528), .Z(n37111) );
  XOR U39355 ( .A(n39529), .B(n39530), .Z(n34282) );
  XNOR U39356 ( .A(n39531), .B(n38343), .Z(n34284) );
  XNOR U39357 ( .A(n39532), .B(n37104), .Z(n32606) );
  XNOR U39358 ( .A(n34633), .B(n39534), .Z(n34291) );
  XOR U39359 ( .A(n39535), .B(n39536), .Z(n34290) );
  XOR U39360 ( .A(n31296), .B(n39537), .Z(n39524) );
  XOR U39361 ( .A(n31046), .B(n32030), .Z(n39537) );
  XNOR U39362 ( .A(n39538), .B(n37100), .Z(n32030) );
  XOR U39363 ( .A(n35799), .B(n39539), .Z(n37100) );
  ANDN U39364 ( .B(n34277), .A(n34279), .Z(n39538) );
  XOR U39365 ( .A(n39540), .B(n38422), .Z(n34279) );
  XOR U39366 ( .A(n39541), .B(n39542), .Z(n34277) );
  XOR U39367 ( .A(n39543), .B(n37115), .Z(n31046) );
  XOR U39368 ( .A(n39544), .B(n39545), .Z(n37115) );
  ANDN U39369 ( .B(n34286), .A(n34287), .Z(n39543) );
  XOR U39370 ( .A(n39546), .B(n39547), .Z(n34287) );
  XOR U39371 ( .A(n39548), .B(n37270), .Z(n34286) );
  XNOR U39372 ( .A(n39549), .B(n37107), .Z(n31296) );
  XOR U39373 ( .A(n38804), .B(n39550), .Z(n37107) );
  AND U39374 ( .A(n36162), .B(n38617), .Z(n39549) );
  XOR U39375 ( .A(n39551), .B(n39552), .Z(n37065) );
  XOR U39376 ( .A(n30778), .B(n32451), .Z(n39552) );
  XNOR U39377 ( .A(n39553), .B(n33085), .Z(n32451) );
  XNOR U39378 ( .A(n39554), .B(n38977), .Z(n33085) );
  XNOR U39379 ( .A(n35604), .B(n39555), .Z(n33086) );
  XOR U39380 ( .A(n39556), .B(n39557), .Z(n30778) );
  AND U39381 ( .A(n34744), .B(n34746), .Z(n39556) );
  XOR U39382 ( .A(n39158), .B(n39558), .Z(n34744) );
  XNOR U39383 ( .A(n30266), .B(n39559), .Z(n39551) );
  XNOR U39384 ( .A(n33071), .B(n30532), .Z(n39559) );
  XOR U39385 ( .A(n39561), .B(n35598), .Z(n33480) );
  XNOR U39386 ( .A(n39562), .B(n39563), .Z(n38448) );
  XNOR U39387 ( .A(n39172), .B(n39564), .Z(n39563) );
  XOR U39388 ( .A(n39565), .B(n39566), .Z(n39172) );
  ANDN U39389 ( .B(n39567), .A(n39568), .Z(n39565) );
  XOR U39390 ( .A(n39569), .B(n39570), .Z(n39562) );
  XOR U39391 ( .A(n39050), .B(n39571), .Z(n39570) );
  XOR U39392 ( .A(n39572), .B(n39573), .Z(n39050) );
  NOR U39393 ( .A(n39574), .B(n39575), .Z(n39572) );
  AND U39394 ( .A(n36862), .B(n33481), .Z(n39560) );
  XNOR U39395 ( .A(n39577), .B(n38027), .Z(n33481) );
  XNOR U39396 ( .A(n39578), .B(n34997), .Z(n33071) );
  XOR U39397 ( .A(n37172), .B(n39579), .Z(n34997) );
  XNOR U39398 ( .A(n39580), .B(n37270), .Z(n34733) );
  XOR U39399 ( .A(n39582), .B(n38080), .Z(n33082) );
  IV U39400 ( .A(n39542), .Z(n38080) );
  NOR U39401 ( .A(n33081), .B(n34738), .Z(n39581) );
  IV U39402 ( .A(n34737), .Z(n33081) );
  XOR U39403 ( .A(n39583), .B(n38295), .Z(n34737) );
  IV U39404 ( .A(n39484), .Z(n38295) );
  XOR U39405 ( .A(n39584), .B(n38617), .Z(n34275) );
  XNOR U39406 ( .A(n35772), .B(n39585), .Z(n38617) );
  ANDN U39407 ( .B(n36163), .A(n36162), .Z(n39584) );
  XNOR U39408 ( .A(n39586), .B(n37646), .Z(n36162) );
  XNOR U39409 ( .A(n39587), .B(n39341), .Z(n36163) );
  IV U39410 ( .A(n39121), .Z(n39341) );
  XOR U39411 ( .A(n39588), .B(n36238), .Z(n25578) );
  XOR U39412 ( .A(n30491), .B(n35429), .Z(n36238) );
  XOR U39413 ( .A(n39589), .B(n34196), .Z(n35429) );
  ANDN U39414 ( .B(n39590), .A(n35640), .Z(n39589) );
  XNOR U39415 ( .A(n37383), .B(n33598), .Z(n30491) );
  XNOR U39416 ( .A(n39591), .B(n39592), .Z(n33598) );
  XNOR U39417 ( .A(n29921), .B(n34187), .Z(n39592) );
  XNOR U39418 ( .A(n39593), .B(n34210), .Z(n34187) );
  XOR U39419 ( .A(n39594), .B(n37036), .Z(n34210) );
  IV U39420 ( .A(n36347), .Z(n37036) );
  ANDN U39421 ( .B(n34209), .A(n35431), .Z(n39593) );
  XOR U39422 ( .A(n39595), .B(n39596), .Z(n34209) );
  XOR U39423 ( .A(n39597), .B(n34197), .Z(n29921) );
  XOR U39424 ( .A(n39598), .B(n37318), .Z(n34197) );
  NOR U39425 ( .A(n34196), .B(n39590), .Z(n39597) );
  XOR U39426 ( .A(n39599), .B(n38667), .Z(n34196) );
  XNOR U39427 ( .A(n32352), .B(n39600), .Z(n39591) );
  XOR U39428 ( .A(n31358), .B(n33263), .Z(n39600) );
  XNOR U39429 ( .A(n39601), .B(n34205), .Z(n33263) );
  XOR U39430 ( .A(n39602), .B(n35308), .Z(n34205) );
  ANDN U39431 ( .B(n34206), .A(n35426), .Z(n39601) );
  XNOR U39432 ( .A(n39603), .B(n39604), .Z(n34206) );
  XNOR U39433 ( .A(n39605), .B(n34192), .Z(n31358) );
  XOR U39434 ( .A(n39606), .B(n38305), .Z(n34192) );
  ANDN U39435 ( .B(n34193), .A(n35434), .Z(n39605) );
  XOR U39436 ( .A(n39607), .B(n39608), .Z(n34193) );
  XNOR U39437 ( .A(n39609), .B(n34201), .Z(n32352) );
  XOR U39438 ( .A(n35926), .B(n39610), .Z(n34201) );
  ANDN U39439 ( .B(n34202), .A(n35423), .Z(n39609) );
  XOR U39440 ( .A(n37428), .B(n39611), .Z(n34202) );
  XOR U39441 ( .A(n39612), .B(n39613), .Z(n37383) );
  XNOR U39442 ( .A(n38187), .B(n32305), .Z(n39613) );
  XNOR U39443 ( .A(n39614), .B(n38199), .Z(n32305) );
  XNOR U39444 ( .A(n39615), .B(n39616), .Z(n38199) );
  XOR U39445 ( .A(n39617), .B(n37002), .Z(n37387) );
  XNOR U39446 ( .A(n39618), .B(n38777), .Z(n37386) );
  XOR U39447 ( .A(n39619), .B(n39620), .Z(n38777) );
  XNOR U39448 ( .A(n39621), .B(n36610), .Z(n38187) );
  XNOR U39449 ( .A(n39622), .B(n33927), .Z(n36610) );
  ANDN U39450 ( .B(n35417), .A(n35418), .Z(n39621) );
  XOR U39451 ( .A(n38896), .B(n39623), .Z(n35418) );
  XOR U39452 ( .A(n39624), .B(n38526), .Z(n35417) );
  XOR U39453 ( .A(n32098), .B(n39625), .Z(n39612) );
  XNOR U39454 ( .A(n30851), .B(n32771), .Z(n39625) );
  XNOR U39455 ( .A(n39626), .B(n36602), .Z(n32771) );
  XOR U39456 ( .A(n39627), .B(n39213), .Z(n36602) );
  ANDN U39457 ( .B(n35409), .A(n35410), .Z(n39626) );
  XOR U39458 ( .A(n39628), .B(n37183), .Z(n35410) );
  XOR U39459 ( .A(n38339), .B(n39629), .Z(n35409) );
  XNOR U39460 ( .A(n39630), .B(n36600), .Z(n30851) );
  XOR U39461 ( .A(n39631), .B(n38305), .Z(n36600) );
  IV U39462 ( .A(n38118), .Z(n38305) );
  XNOR U39463 ( .A(n39632), .B(n39633), .Z(n38118) );
  NOR U39464 ( .A(n39018), .B(n35404), .Z(n39630) );
  XOR U39465 ( .A(n39634), .B(n37848), .Z(n35404) );
  XOR U39466 ( .A(n39635), .B(n39636), .Z(n37848) );
  XOR U39467 ( .A(n39637), .B(n36367), .Z(n39018) );
  XOR U39468 ( .A(n39638), .B(n36607), .Z(n32098) );
  XNOR U39469 ( .A(n38285), .B(n39639), .Z(n36607) );
  NOR U39470 ( .A(n35414), .B(n35413), .Z(n39638) );
  XNOR U39471 ( .A(n39640), .B(n39542), .Z(n35413) );
  XNOR U39472 ( .A(n39641), .B(n39642), .Z(n39542) );
  XOR U39473 ( .A(n39643), .B(n39484), .Z(n35414) );
  ANDN U39474 ( .B(n31284), .A(n27606), .Z(n39588) );
  XOR U39475 ( .A(n31566), .B(n35976), .Z(n27606) );
  XOR U39476 ( .A(n39644), .B(n34545), .Z(n35976) );
  NOR U39477 ( .A(n35223), .B(n35222), .Z(n39644) );
  XOR U39478 ( .A(n39645), .B(n37040), .Z(n35223) );
  IV U39479 ( .A(n32300), .Z(n31566) );
  XNOR U39480 ( .A(n33048), .B(n39646), .Z(n32300) );
  XOR U39481 ( .A(n39647), .B(n39648), .Z(n33048) );
  XNOR U39482 ( .A(n33602), .B(n29931), .Z(n39648) );
  XNOR U39483 ( .A(n39649), .B(n34553), .Z(n29931) );
  XOR U39484 ( .A(n39650), .B(n35938), .Z(n34553) );
  AND U39485 ( .A(n34901), .B(n34554), .Z(n39649) );
  XOR U39486 ( .A(n39653), .B(n39608), .Z(n34554) );
  XOR U39487 ( .A(n39654), .B(n38169), .Z(n34901) );
  XNOR U39488 ( .A(n39655), .B(n34557), .Z(n33602) );
  XOR U39489 ( .A(n39656), .B(n39657), .Z(n34557) );
  ANDN U39490 ( .B(n34558), .A(n35994), .Z(n39655) );
  IV U39491 ( .A(n35981), .Z(n35994) );
  XNOR U39492 ( .A(n39658), .B(n37525), .Z(n35981) );
  XOR U39493 ( .A(n39659), .B(n37928), .Z(n34558) );
  XNOR U39494 ( .A(n31217), .B(n39660), .Z(n39647) );
  XOR U39495 ( .A(n31994), .B(n31981), .Z(n39660) );
  XNOR U39496 ( .A(n39661), .B(n34549), .Z(n31981) );
  XNOR U39497 ( .A(n39662), .B(n39389), .Z(n34549) );
  AND U39498 ( .A(n34550), .B(n34129), .Z(n39661) );
  XOR U39499 ( .A(n37323), .B(n39663), .Z(n34129) );
  XNOR U39500 ( .A(n39664), .B(n39665), .Z(n34550) );
  XNOR U39501 ( .A(n39666), .B(n34546), .Z(n31994) );
  XNOR U39502 ( .A(n39667), .B(n36970), .Z(n34546) );
  ANDN U39503 ( .B(n35222), .A(n34545), .Z(n39666) );
  XOR U39504 ( .A(n39668), .B(n39468), .Z(n34545) );
  XOR U39505 ( .A(n39669), .B(n37610), .Z(n35222) );
  IV U39506 ( .A(n36437), .Z(n37610) );
  XOR U39507 ( .A(n39670), .B(n39145), .Z(n31217) );
  IV U39508 ( .A(n34541), .Z(n39145) );
  XOR U39509 ( .A(n39671), .B(n38096), .Z(n34541) );
  AND U39510 ( .A(n34542), .B(n34122), .Z(n39670) );
  XNOR U39511 ( .A(n39672), .B(n38972), .Z(n34122) );
  XOR U39512 ( .A(n34628), .B(n39673), .Z(n34542) );
  XOR U39513 ( .A(n39674), .B(n39675), .Z(n34628) );
  XOR U39514 ( .A(n39676), .B(n30371), .Z(n31284) );
  XOR U39515 ( .A(n26348), .B(n39677), .Z(n39391) );
  XNOR U39516 ( .A(n26100), .B(n27666), .Z(n39677) );
  XNOR U39517 ( .A(n39678), .B(n28212), .Z(n27666) );
  XOR U39518 ( .A(n37392), .B(n31299), .Z(n28212) );
  IV U39519 ( .A(n31542), .Z(n31299) );
  XNOR U39520 ( .A(n39679), .B(n39680), .Z(n33717) );
  XOR U39521 ( .A(n30526), .B(n33207), .Z(n39680) );
  XNOR U39522 ( .A(n39681), .B(n36110), .Z(n33207) );
  XNOR U39523 ( .A(n39682), .B(n35376), .Z(n36110) );
  ANDN U39524 ( .B(n36111), .A(n39683), .Z(n39681) );
  XOR U39525 ( .A(n39315), .B(n39684), .Z(n36111) );
  XOR U39526 ( .A(n39685), .B(n36106), .Z(n30526) );
  XNOR U39527 ( .A(n39686), .B(n37040), .Z(n36106) );
  ANDN U39528 ( .B(n36107), .A(n39687), .Z(n39685) );
  XOR U39529 ( .A(n39688), .B(n37523), .Z(n36107) );
  XOR U39530 ( .A(n33188), .B(n39689), .Z(n39679) );
  XOR U39531 ( .A(n28746), .B(n35731), .Z(n39689) );
  XNOR U39532 ( .A(n39690), .B(n36097), .Z(n35731) );
  XOR U39533 ( .A(n39691), .B(n39692), .Z(n36097) );
  ANDN U39534 ( .B(n36098), .A(n39693), .Z(n39690) );
  XNOR U39535 ( .A(n39694), .B(n38027), .Z(n36098) );
  XNOR U39536 ( .A(n39695), .B(n36114), .Z(n28746) );
  XNOR U39537 ( .A(n37698), .B(n39696), .Z(n36114) );
  ANDN U39538 ( .B(n36115), .A(n39697), .Z(n39695) );
  XNOR U39539 ( .A(n39121), .B(n39698), .Z(n36115) );
  XNOR U39540 ( .A(n39699), .B(n39700), .Z(n39121) );
  XNOR U39541 ( .A(n39701), .B(n36102), .Z(n33188) );
  XNOR U39542 ( .A(n39702), .B(n33922), .Z(n36102) );
  ANDN U39543 ( .B(n36101), .A(n39705), .Z(n39701) );
  XNOR U39544 ( .A(n39706), .B(n39707), .Z(n34020) );
  XOR U39545 ( .A(n31472), .B(n29054), .Z(n39707) );
  XOR U39546 ( .A(n39708), .B(n39709), .Z(n29054) );
  ANDN U39547 ( .B(n37411), .A(n36804), .Z(n39708) );
  XOR U39548 ( .A(n38556), .B(n39710), .Z(n36804) );
  IV U39549 ( .A(n37204), .Z(n38556) );
  XOR U39550 ( .A(n39711), .B(n39652), .Z(n37204) );
  XNOR U39551 ( .A(n39712), .B(n39713), .Z(n39652) );
  XNOR U39552 ( .A(n38765), .B(n38867), .Z(n39713) );
  XNOR U39553 ( .A(n39714), .B(n39715), .Z(n38867) );
  ANDN U39554 ( .B(n39716), .A(n39717), .Z(n39714) );
  XNOR U39555 ( .A(n39718), .B(n39719), .Z(n38765) );
  ANDN U39556 ( .B(n39720), .A(n39721), .Z(n39718) );
  XOR U39557 ( .A(n39722), .B(n39723), .Z(n39712) );
  XOR U39558 ( .A(n38582), .B(n35077), .Z(n39723) );
  XNOR U39559 ( .A(n39724), .B(n39725), .Z(n35077) );
  XNOR U39560 ( .A(n39728), .B(n39729), .Z(n38582) );
  NOR U39561 ( .A(n39730), .B(n39731), .Z(n39728) );
  XNOR U39562 ( .A(n39732), .B(n39733), .Z(n31472) );
  NOR U39563 ( .A(n36816), .B(n35738), .Z(n39732) );
  XOR U39564 ( .A(n39734), .B(n39735), .Z(n35738) );
  XNOR U39565 ( .A(n39736), .B(n39213), .Z(n36816) );
  XOR U39566 ( .A(n30566), .B(n39737), .Z(n39706) );
  XNOR U39567 ( .A(n32526), .B(n31073), .Z(n39737) );
  XNOR U39568 ( .A(n39738), .B(n36528), .Z(n31073) );
  ANDN U39569 ( .B(n36529), .A(n36812), .Z(n39738) );
  XOR U39570 ( .A(n38851), .B(n39739), .Z(n36812) );
  XNOR U39571 ( .A(n39741), .B(n36640), .Z(n32526) );
  ANDN U39572 ( .B(n36641), .A(n36809), .Z(n39741) );
  IV U39573 ( .A(n37409), .Z(n36809) );
  XNOR U39574 ( .A(n39742), .B(n37027), .Z(n37409) );
  XNOR U39575 ( .A(n39743), .B(n39744), .Z(n37027) );
  XOR U39576 ( .A(n37069), .B(n39745), .Z(n36641) );
  XNOR U39577 ( .A(n39746), .B(n39747), .Z(n37069) );
  XNOR U39578 ( .A(n39748), .B(n35745), .Z(n30566) );
  ANDN U39579 ( .B(n35746), .A(n36801), .Z(n39748) );
  XNOR U39580 ( .A(n35583), .B(n39749), .Z(n36801) );
  XNOR U39581 ( .A(n39750), .B(n37535), .Z(n35746) );
  XOR U39582 ( .A(n39751), .B(n36101), .Z(n37392) );
  XOR U39583 ( .A(n39752), .B(n38863), .Z(n36101) );
  ANDN U39584 ( .B(n38223), .A(n39753), .Z(n39751) );
  ANDN U39585 ( .B(n28213), .A(n27589), .Z(n39678) );
  XOR U39586 ( .A(n37229), .B(n30583), .Z(n27589) );
  XOR U39587 ( .A(n37384), .B(n37753), .Z(n30583) );
  XNOR U39588 ( .A(n39754), .B(n39755), .Z(n37753) );
  XNOR U39589 ( .A(n30645), .B(n34425), .Z(n39755) );
  XOR U39590 ( .A(n39756), .B(n36590), .Z(n34425) );
  ANDN U39591 ( .B(n37218), .A(n36264), .Z(n39756) );
  XOR U39592 ( .A(n39757), .B(n38801), .Z(n36264) );
  XOR U39593 ( .A(n39760), .B(n36586), .Z(n30645) );
  XOR U39594 ( .A(n39761), .B(n39762), .Z(n36256) );
  XOR U39595 ( .A(n32954), .B(n39763), .Z(n39754) );
  XOR U39596 ( .A(n38986), .B(n33824), .Z(n39763) );
  XNOR U39597 ( .A(n39764), .B(n36588), .Z(n33824) );
  ANDN U39598 ( .B(n37207), .A(n36251), .Z(n39764) );
  IV U39599 ( .A(n37208), .Z(n36251) );
  XOR U39600 ( .A(n39765), .B(n37428), .Z(n37208) );
  IV U39601 ( .A(n37635), .Z(n37428) );
  XNOR U39602 ( .A(n39766), .B(n39767), .Z(n37635) );
  XOR U39603 ( .A(n39768), .B(n36581), .Z(n38986) );
  ANDN U39604 ( .B(n37765), .A(n36260), .Z(n39768) );
  XOR U39605 ( .A(n39769), .B(n39770), .Z(n36260) );
  XOR U39606 ( .A(n39771), .B(n36583), .Z(n32954) );
  ANDN U39607 ( .B(n36247), .A(n37203), .Z(n39771) );
  XOR U39608 ( .A(n39772), .B(n37715), .Z(n36247) );
  XOR U39609 ( .A(n39773), .B(n39774), .Z(n37384) );
  XNOR U39610 ( .A(n30761), .B(n39775), .Z(n39774) );
  XNOR U39611 ( .A(n39776), .B(n36621), .Z(n30761) );
  ANDN U39612 ( .B(n39777), .A(n39044), .Z(n39776) );
  XOR U39613 ( .A(n32488), .B(n39778), .Z(n39773) );
  XOR U39614 ( .A(n32192), .B(n32906), .Z(n39778) );
  XOR U39615 ( .A(n39779), .B(n36617), .Z(n32906) );
  XNOR U39616 ( .A(n39780), .B(n36899), .Z(n37233) );
  XOR U39617 ( .A(n39781), .B(n36630), .Z(n32192) );
  ANDN U39618 ( .B(n37227), .A(n37228), .Z(n39781) );
  XOR U39619 ( .A(n39782), .B(n39783), .Z(n37228) );
  XNOR U39620 ( .A(n39784), .B(n36634), .Z(n32488) );
  XOR U39621 ( .A(n38858), .B(n39785), .Z(n37225) );
  XNOR U39622 ( .A(n39786), .B(n39777), .Z(n37229) );
  ANDN U39623 ( .B(n39044), .A(n36619), .Z(n39786) );
  XOR U39624 ( .A(n39787), .B(n39788), .Z(n36619) );
  XOR U39625 ( .A(n39789), .B(n38804), .Z(n39044) );
  XOR U39626 ( .A(n37121), .B(n30746), .Z(n28213) );
  XNOR U39627 ( .A(n36155), .B(n33852), .Z(n30746) );
  XNOR U39628 ( .A(n39790), .B(n39791), .Z(n33852) );
  XNOR U39629 ( .A(n32396), .B(n33052), .Z(n39791) );
  XNOR U39630 ( .A(n39792), .B(n36559), .Z(n33052) );
  XOR U39631 ( .A(n39794), .B(n39795), .Z(n36779) );
  XOR U39632 ( .A(n36519), .B(n39796), .Z(n34876) );
  XOR U39633 ( .A(n38176), .B(n39797), .Z(n36385) );
  XOR U39634 ( .A(n39798), .B(n39799), .Z(n38176) );
  XNOR U39635 ( .A(n39800), .B(n34719), .Z(n32396) );
  XOR U39636 ( .A(n39770), .B(n39801), .Z(n34719) );
  IV U39637 ( .A(n36550), .Z(n39770) );
  XNOR U39638 ( .A(n39802), .B(n39803), .Z(n36550) );
  ANDN U39639 ( .B(n34873), .A(n34718), .Z(n39800) );
  XOR U39640 ( .A(n37890), .B(n39804), .Z(n34718) );
  XOR U39641 ( .A(n38950), .B(n39805), .Z(n34873) );
  XOR U39642 ( .A(n31347), .B(n39806), .Z(n39790) );
  XOR U39643 ( .A(n33409), .B(n34000), .Z(n39806) );
  XNOR U39644 ( .A(n39807), .B(n34724), .Z(n34000) );
  XNOR U39645 ( .A(n39808), .B(n38169), .Z(n34724) );
  XOR U39646 ( .A(n39809), .B(n38298), .Z(n34861) );
  XOR U39647 ( .A(n39810), .B(n37144), .Z(n34725) );
  XNOR U39648 ( .A(n39811), .B(n34715), .Z(n33409) );
  XNOR U39649 ( .A(n39812), .B(n36555), .Z(n34715) );
  ANDN U39650 ( .B(n34870), .A(n34714), .Z(n39811) );
  XNOR U39651 ( .A(n39813), .B(n39278), .Z(n34714) );
  XOR U39652 ( .A(n39814), .B(n39307), .Z(n34870) );
  XNOR U39653 ( .A(n39815), .B(n37090), .Z(n31347) );
  XNOR U39654 ( .A(n37172), .B(n39816), .Z(n37090) );
  XNOR U39655 ( .A(n39817), .B(n39818), .Z(n37172) );
  NOR U39656 ( .A(n34865), .B(n34728), .Z(n39815) );
  XNOR U39657 ( .A(n39819), .B(n35929), .Z(n34728) );
  XOR U39658 ( .A(n39820), .B(n39821), .Z(n34865) );
  XNOR U39659 ( .A(n39822), .B(n39823), .Z(n36155) );
  XOR U39660 ( .A(n34399), .B(n34709), .Z(n39823) );
  XNOR U39661 ( .A(n39824), .B(n34735), .Z(n34709) );
  XOR U39662 ( .A(n39825), .B(n38948), .Z(n34735) );
  NOR U39663 ( .A(n34734), .B(n34996), .Z(n39824) );
  XOR U39664 ( .A(n39826), .B(n39827), .Z(n34996) );
  XOR U39665 ( .A(n39828), .B(n37030), .Z(n34734) );
  XNOR U39666 ( .A(n39829), .B(n34738), .Z(n34399) );
  XOR U39667 ( .A(n37672), .B(n39830), .Z(n34738) );
  XOR U39668 ( .A(n39831), .B(n38863), .Z(n34739) );
  XOR U39669 ( .A(n39832), .B(n38352), .Z(n33080) );
  XOR U39670 ( .A(n39833), .B(n39834), .Z(n38352) );
  XOR U39671 ( .A(n31690), .B(n39835), .Z(n39822) );
  XNOR U39672 ( .A(n29170), .B(n33008), .Z(n39835) );
  XNOR U39673 ( .A(n39836), .B(n34746), .Z(n33008) );
  XOR U39674 ( .A(n39837), .B(n39838), .Z(n34746) );
  XOR U39675 ( .A(n39839), .B(n36862), .Z(n29170) );
  XOR U39676 ( .A(n39840), .B(n37512), .Z(n36862) );
  IV U39677 ( .A(n36369), .Z(n37512) );
  XOR U39678 ( .A(n39841), .B(n39842), .Z(n36369) );
  ANDN U39679 ( .B(n33479), .A(n36861), .Z(n39839) );
  XOR U39680 ( .A(n39843), .B(n38037), .Z(n36861) );
  XNOR U39681 ( .A(n38950), .B(n39844), .Z(n33479) );
  XNOR U39682 ( .A(n39845), .B(n37093), .Z(n31690) );
  XOR U39683 ( .A(n39846), .B(n39847), .Z(n37093) );
  ANDN U39684 ( .B(n33084), .A(n37092), .Z(n39845) );
  XOR U39685 ( .A(n39848), .B(n39849), .Z(n37092) );
  XOR U39686 ( .A(n39850), .B(n38422), .Z(n33084) );
  IV U39687 ( .A(n39616), .Z(n38422) );
  XOR U39688 ( .A(n39851), .B(n34745), .Z(n37121) );
  XOR U39689 ( .A(n39852), .B(n37517), .Z(n34745) );
  ANDN U39690 ( .B(n36373), .A(n39557), .Z(n39851) );
  IV U39691 ( .A(n36374), .Z(n39557) );
  XOR U39692 ( .A(n39853), .B(n39113), .Z(n36374) );
  XOR U39693 ( .A(n34638), .B(n39854), .Z(n36373) );
  XNOR U39694 ( .A(n39855), .B(n28207), .Z(n26100) );
  XNOR U39695 ( .A(n39856), .B(n39857), .Z(n37771) );
  XNOR U39696 ( .A(n30212), .B(n30587), .Z(n39857) );
  XNOR U39697 ( .A(n39858), .B(n38047), .Z(n30587) );
  XOR U39698 ( .A(n39859), .B(n37802), .Z(n33845) );
  XOR U39699 ( .A(n39860), .B(n38054), .Z(n30212) );
  AND U39700 ( .A(n33228), .B(n33230), .Z(n39860) );
  XOR U39701 ( .A(n39861), .B(n38564), .Z(n33230) );
  XNOR U39702 ( .A(n31269), .B(n39862), .Z(n39856) );
  XOR U39703 ( .A(n33640), .B(n32720), .Z(n39862) );
  XOR U39704 ( .A(n39863), .B(n38057), .Z(n32720) );
  AND U39705 ( .A(n36042), .B(n36044), .Z(n39863) );
  XOR U39706 ( .A(n39864), .B(n37791), .Z(n36044) );
  XOR U39707 ( .A(n39865), .B(n38044), .Z(n33640) );
  ANDN U39708 ( .B(n33937), .A(n33938), .Z(n39865) );
  XNOR U39709 ( .A(n37148), .B(n39866), .Z(n33938) );
  XOR U39710 ( .A(n39867), .B(n38051), .Z(n31269) );
  ANDN U39711 ( .B(n37806), .A(n37807), .Z(n39867) );
  XOR U39712 ( .A(n39868), .B(n38895), .Z(n37807) );
  XNOR U39713 ( .A(n39869), .B(n39870), .Z(n35871) );
  XOR U39714 ( .A(n33029), .B(n32633), .Z(n39870) );
  XOR U39715 ( .A(n39871), .B(n38074), .Z(n32633) );
  ANDN U39716 ( .B(n36743), .A(n39872), .Z(n39871) );
  XOR U39717 ( .A(n39873), .B(n38062), .Z(n33029) );
  ANDN U39718 ( .B(n36748), .A(n36747), .Z(n39873) );
  XNOR U39719 ( .A(n39874), .B(n39875), .Z(n39869) );
  XNOR U39720 ( .A(n31118), .B(n31967), .Z(n39875) );
  XOR U39721 ( .A(n39876), .B(n38414), .Z(n31967) );
  AND U39722 ( .A(n36754), .B(n36753), .Z(n39876) );
  XNOR U39723 ( .A(n39877), .B(n38070), .Z(n31118) );
  ANDN U39724 ( .B(n39878), .A(n39879), .Z(n39877) );
  XOR U39725 ( .A(n39880), .B(n39879), .Z(n36751) );
  NOR U39726 ( .A(n39878), .B(n38069), .Z(n39880) );
  ANDN U39727 ( .B(n27602), .A(n28206), .Z(n39855) );
  XNOR U39728 ( .A(n35742), .B(n32456), .Z(n28206) );
  XOR U39729 ( .A(n33669), .B(n34222), .Z(n32456) );
  XNOR U39730 ( .A(n39881), .B(n39882), .Z(n34222) );
  XOR U39731 ( .A(n32086), .B(n32040), .Z(n39882) );
  XOR U39732 ( .A(n39883), .B(n36509), .Z(n32040) );
  XNOR U39733 ( .A(n39884), .B(n38950), .Z(n36509) );
  ANDN U39734 ( .B(n36523), .A(n34025), .Z(n39883) );
  IV U39735 ( .A(n38376), .Z(n34025) );
  XNOR U39736 ( .A(n39885), .B(n37114), .Z(n38376) );
  XNOR U39737 ( .A(n39886), .B(n36417), .Z(n36523) );
  IV U39738 ( .A(n37602), .Z(n36417) );
  XNOR U39739 ( .A(n39887), .B(n39888), .Z(n37602) );
  XNOR U39740 ( .A(n39889), .B(n35855), .Z(n32086) );
  XOR U39741 ( .A(n39890), .B(n36987), .Z(n35855) );
  IV U39742 ( .A(n39891), .Z(n36987) );
  ANDN U39743 ( .B(n35856), .A(n34030), .Z(n39889) );
  IV U39744 ( .A(n38369), .Z(n34030) );
  XOR U39745 ( .A(n38896), .B(n39892), .Z(n38369) );
  XOR U39746 ( .A(n39893), .B(n38690), .Z(n38896) );
  XOR U39747 ( .A(n39894), .B(n39895), .Z(n38690) );
  XOR U39748 ( .A(n39003), .B(n37775), .Z(n39895) );
  XNOR U39749 ( .A(n39896), .B(n39897), .Z(n37775) );
  ANDN U39750 ( .B(n39898), .A(n39899), .Z(n39896) );
  XOR U39751 ( .A(n39900), .B(n39901), .Z(n39003) );
  ANDN U39752 ( .B(n39902), .A(n39903), .Z(n39900) );
  XOR U39753 ( .A(n38947), .B(n39904), .Z(n39894) );
  XNOR U39754 ( .A(n39074), .B(n38408), .Z(n39904) );
  XOR U39755 ( .A(n39905), .B(n39906), .Z(n38408) );
  ANDN U39756 ( .B(n39907), .A(n39908), .Z(n39905) );
  XNOR U39757 ( .A(n39909), .B(n39910), .Z(n39074) );
  NOR U39758 ( .A(n39911), .B(n39912), .Z(n39909) );
  XOR U39759 ( .A(n39913), .B(n39914), .Z(n38947) );
  ANDN U39760 ( .B(n39915), .A(n39916), .Z(n39913) );
  XNOR U39761 ( .A(n37912), .B(n39917), .Z(n35856) );
  XNOR U39762 ( .A(n31593), .B(n39918), .Z(n39881) );
  XOR U39763 ( .A(n31926), .B(n31564), .Z(n39918) );
  XOR U39764 ( .A(n39919), .B(n36505), .Z(n31564) );
  IV U39765 ( .A(n35864), .Z(n36505) );
  XOR U39766 ( .A(n39920), .B(n39381), .Z(n35864) );
  IV U39767 ( .A(n34626), .Z(n39381) );
  ANDN U39768 ( .B(n35865), .A(n34038), .Z(n39919) );
  IV U39769 ( .A(n38372), .Z(n34038) );
  XOR U39770 ( .A(n39921), .B(n39482), .Z(n38372) );
  XOR U39771 ( .A(n38851), .B(n39922), .Z(n35865) );
  XNOR U39772 ( .A(n39924), .B(n38817), .Z(n35861) );
  ANDN U39773 ( .B(n35862), .A(n34034), .Z(n39923) );
  XNOR U39774 ( .A(n39925), .B(n36970), .Z(n34034) );
  XOR U39775 ( .A(n39926), .B(n34633), .Z(n35862) );
  XOR U39776 ( .A(n39927), .B(n35852), .Z(n31593) );
  XOR U39777 ( .A(n39928), .B(n37794), .Z(n35852) );
  ANDN U39778 ( .B(n35853), .A(n38366), .Z(n39927) );
  XOR U39779 ( .A(n39929), .B(n38446), .Z(n38366) );
  XNOR U39780 ( .A(n39930), .B(n39931), .Z(n35853) );
  XOR U39781 ( .A(n39932), .B(n39933), .Z(n33669) );
  XNOR U39782 ( .A(n33639), .B(n33552), .Z(n39933) );
  XOR U39783 ( .A(n39934), .B(n36813), .Z(n33552) );
  XOR U39784 ( .A(n39935), .B(n37672), .Z(n36813) );
  IV U39785 ( .A(n39936), .Z(n37672) );
  NOR U39786 ( .A(n36814), .B(n36528), .Z(n39934) );
  XOR U39787 ( .A(n39937), .B(n39938), .Z(n36528) );
  XNOR U39788 ( .A(n39939), .B(n37071), .Z(n36814) );
  XNOR U39789 ( .A(n39940), .B(n36805), .Z(n33639) );
  XOR U39790 ( .A(n39941), .B(n36215), .Z(n36805) );
  ANDN U39791 ( .B(n36806), .A(n39709), .Z(n39940) );
  XNOR U39792 ( .A(n30912), .B(n39942), .Z(n39932) );
  XOR U39793 ( .A(n35846), .B(n33826), .Z(n39942) );
  XNOR U39794 ( .A(n39943), .B(n36802), .Z(n33826) );
  XOR U39795 ( .A(n39944), .B(n39945), .Z(n36802) );
  NOR U39796 ( .A(n35745), .B(n35744), .Z(n39943) );
  XNOR U39797 ( .A(n39946), .B(n39947), .Z(n35744) );
  XOR U39798 ( .A(n35304), .B(n39948), .Z(n35745) );
  XOR U39799 ( .A(n39949), .B(n39619), .Z(n35304) );
  XNOR U39800 ( .A(n39950), .B(n39951), .Z(n39619) );
  XOR U39801 ( .A(n37080), .B(n38357), .Z(n39951) );
  XOR U39802 ( .A(n39952), .B(n39953), .Z(n38357) );
  ANDN U39803 ( .B(n39954), .A(n39955), .Z(n39952) );
  XNOR U39804 ( .A(n39956), .B(n39957), .Z(n37080) );
  ANDN U39805 ( .B(n39958), .A(n39959), .Z(n39956) );
  XOR U39806 ( .A(n39960), .B(n39961), .Z(n39950) );
  XNOR U39807 ( .A(n39294), .B(n39962), .Z(n39961) );
  XOR U39808 ( .A(n39963), .B(n39964), .Z(n39294) );
  NOR U39809 ( .A(n39965), .B(n39966), .Z(n39963) );
  XNOR U39810 ( .A(n39967), .B(n36810), .Z(n35846) );
  XOR U39811 ( .A(n39968), .B(n35378), .Z(n36810) );
  XNOR U39812 ( .A(n39969), .B(n39970), .Z(n35378) );
  AND U39813 ( .A(n36640), .B(n36639), .Z(n39967) );
  XOR U39814 ( .A(n39158), .B(n39971), .Z(n36639) );
  XOR U39815 ( .A(n39972), .B(n34631), .Z(n36640) );
  XNOR U39816 ( .A(n39973), .B(n36817), .Z(n30912) );
  XOR U39817 ( .A(n39974), .B(n38320), .Z(n36817) );
  ANDN U39818 ( .B(n35737), .A(n39733), .Z(n39973) );
  IV U39819 ( .A(n35739), .Z(n39733) );
  XOR U39820 ( .A(n39975), .B(n39976), .Z(n35739) );
  XNOR U39821 ( .A(n35787), .B(n39977), .Z(n35737) );
  XNOR U39822 ( .A(n39978), .B(n36806), .Z(n35742) );
  XNOR U39823 ( .A(n35586), .B(n39979), .Z(n36806) );
  ANDN U39824 ( .B(n39709), .A(n37411), .Z(n39978) );
  XNOR U39825 ( .A(n39980), .B(n37051), .Z(n37411) );
  XNOR U39826 ( .A(n39981), .B(n39982), .Z(n39709) );
  XNOR U39827 ( .A(n32203), .B(n37353), .Z(n27602) );
  ANDN U39828 ( .B(n34945), .A(n34946), .Z(n39983) );
  XOR U39829 ( .A(n39984), .B(n37270), .Z(n34946) );
  IV U39830 ( .A(n39982), .Z(n37270) );
  IV U39831 ( .A(n29060), .Z(n32203) );
  XNOR U39832 ( .A(n39987), .B(n28203), .Z(n26348) );
  XOR U39833 ( .A(n34991), .B(n31050), .Z(n28203) );
  IV U39834 ( .A(n29286), .Z(n31050) );
  XNOR U39835 ( .A(n39988), .B(n39989), .Z(n35335) );
  XOR U39836 ( .A(n32102), .B(n35111), .Z(n39989) );
  XNOR U39837 ( .A(n39990), .B(n35117), .Z(n35111) );
  ANDN U39838 ( .B(n34056), .A(n35116), .Z(n39990) );
  XNOR U39839 ( .A(n39413), .B(n39991), .Z(n35116) );
  XNOR U39840 ( .A(n37005), .B(n39992), .Z(n34056) );
  XNOR U39841 ( .A(n39993), .B(n35123), .Z(n32102) );
  ANDN U39842 ( .B(n36287), .A(n35122), .Z(n39993) );
  XNOR U39843 ( .A(n39994), .B(n39255), .Z(n35122) );
  IV U39844 ( .A(n37707), .Z(n39255) );
  XOR U39845 ( .A(n39995), .B(n37326), .Z(n36287) );
  IV U39846 ( .A(n39996), .Z(n37326) );
  XOR U39847 ( .A(n33985), .B(n39997), .Z(n39988) );
  XOR U39848 ( .A(n33638), .B(n33267), .Z(n39997) );
  XNOR U39849 ( .A(n39998), .B(n35126), .Z(n33267) );
  ANDN U39850 ( .B(n34050), .A(n35125), .Z(n39998) );
  XOR U39851 ( .A(n39999), .B(n40000), .Z(n35125) );
  XOR U39852 ( .A(n40001), .B(n38444), .Z(n34050) );
  XNOR U39853 ( .A(n40002), .B(n36457), .Z(n33638) );
  ANDN U39854 ( .B(n36296), .A(n34060), .Z(n40002) );
  XOR U39855 ( .A(n40003), .B(n39547), .Z(n34060) );
  IV U39856 ( .A(n35634), .Z(n39547) );
  XNOR U39857 ( .A(n40004), .B(n40005), .Z(n36296) );
  XNOR U39858 ( .A(n40006), .B(n37547), .Z(n33985) );
  ANDN U39859 ( .B(n34046), .A(n37548), .Z(n40006) );
  XOR U39860 ( .A(n37323), .B(n40007), .Z(n37548) );
  XNOR U39861 ( .A(n40008), .B(n37183), .Z(n34046) );
  XOR U39862 ( .A(n38809), .B(n40009), .Z(n37183) );
  XNOR U39863 ( .A(n40010), .B(n40011), .Z(n38809) );
  XOR U39864 ( .A(n40012), .B(n40013), .Z(n40011) );
  XNOR U39865 ( .A(n35773), .B(n40014), .Z(n40010) );
  XNOR U39866 ( .A(n40015), .B(n39585), .Z(n40014) );
  XOR U39867 ( .A(n40016), .B(n40017), .Z(n39585) );
  AND U39868 ( .A(n40018), .B(n40019), .Z(n40016) );
  XOR U39869 ( .A(n40020), .B(n40021), .Z(n35773) );
  AND U39870 ( .A(n40022), .B(n40023), .Z(n40020) );
  XNOR U39871 ( .A(n40024), .B(n40025), .Z(n35506) );
  XOR U39872 ( .A(n29725), .B(n32506), .Z(n40025) );
  XOR U39873 ( .A(n40026), .B(n40027), .Z(n32506) );
  NOR U39874 ( .A(n34987), .B(n34986), .Z(n40026) );
  XNOR U39875 ( .A(n40028), .B(n33896), .Z(n29725) );
  NOR U39876 ( .A(n40029), .B(n33897), .Z(n40028) );
  XOR U39877 ( .A(n30134), .B(n40030), .Z(n40024) );
  XOR U39878 ( .A(n32753), .B(n29412), .Z(n40030) );
  XNOR U39879 ( .A(n40031), .B(n35438), .Z(n29412) );
  NOR U39880 ( .A(n34982), .B(n34983), .Z(n40031) );
  XOR U39881 ( .A(n40032), .B(n39186), .Z(n34982) );
  XNOR U39882 ( .A(n40033), .B(n33891), .Z(n32753) );
  NOR U39883 ( .A(n37894), .B(n33890), .Z(n40033) );
  XNOR U39884 ( .A(n35315), .B(n40034), .Z(n33890) );
  XOR U39885 ( .A(n40035), .B(n33901), .Z(n30134) );
  NOR U39886 ( .A(n34993), .B(n33900), .Z(n40035) );
  XNOR U39887 ( .A(n40036), .B(n37044), .Z(n33900) );
  XNOR U39888 ( .A(n40037), .B(n33897), .Z(n34991) );
  XNOR U39889 ( .A(n40038), .B(n39664), .Z(n33897) );
  ANDN U39890 ( .B(n40029), .A(n40039), .Z(n40037) );
  ANDN U39891 ( .B(n28202), .A(n27593), .Z(n39987) );
  IV U39892 ( .A(n31279), .Z(n27593) );
  XOR U39893 ( .A(n33295), .B(n37732), .Z(n31279) );
  XNOR U39894 ( .A(n40040), .B(n35059), .Z(n37732) );
  ANDN U39895 ( .B(n35575), .A(n40041), .Z(n40040) );
  IV U39896 ( .A(n38567), .Z(n35575) );
  XOR U39897 ( .A(n40042), .B(n39996), .Z(n38567) );
  XOR U39898 ( .A(n30793), .B(n40043), .Z(n28202) );
  IV U39899 ( .A(n31659), .Z(n30793) );
  XNOR U39900 ( .A(n34358), .B(n32088), .Z(n31659) );
  XNOR U39901 ( .A(n40044), .B(n40045), .Z(n32088) );
  XOR U39902 ( .A(n30274), .B(n31867), .Z(n40045) );
  XNOR U39903 ( .A(n40046), .B(n37994), .Z(n31867) );
  IV U39904 ( .A(n38717), .Z(n37994) );
  XOR U39905 ( .A(n40047), .B(n38977), .Z(n38717) );
  NOR U39906 ( .A(n38716), .B(n38385), .Z(n40046) );
  XOR U39907 ( .A(n40048), .B(n37990), .Z(n30274) );
  XOR U39908 ( .A(n40049), .B(n39596), .Z(n37990) );
  XOR U39909 ( .A(n38698), .B(n40050), .Z(n40044) );
  XNOR U39910 ( .A(n34353), .B(n32579), .Z(n40050) );
  XNOR U39911 ( .A(n40052), .B(n37525), .Z(n38007) );
  ANDN U39912 ( .B(n38704), .A(n40053), .Z(n40051) );
  XOR U39913 ( .A(n40054), .B(n37999), .Z(n34353) );
  XOR U39914 ( .A(n39001), .B(n40055), .Z(n37999) );
  ANDN U39915 ( .B(n38387), .A(n40056), .Z(n40054) );
  XNOR U39916 ( .A(n40057), .B(n38003), .Z(n38698) );
  IV U39917 ( .A(n38722), .Z(n38003) );
  XOR U39918 ( .A(n40058), .B(n38446), .Z(n38722) );
  NOR U39919 ( .A(n38721), .B(n38382), .Z(n40057) );
  XOR U39920 ( .A(n40059), .B(n40060), .Z(n34358) );
  XOR U39921 ( .A(n39676), .B(n32341), .Z(n40060) );
  XNOR U39922 ( .A(n40061), .B(n37985), .Z(n32341) );
  ANDN U39923 ( .B(n35886), .A(n40062), .Z(n40061) );
  XNOR U39924 ( .A(n40063), .B(n37980), .Z(n39676) );
  ANDN U39925 ( .B(n40064), .A(n35876), .Z(n40063) );
  XNOR U39926 ( .A(n30370), .B(n40065), .Z(n40059) );
  XOR U39927 ( .A(n40066), .B(n33516), .Z(n40065) );
  XNOR U39928 ( .A(n40067), .B(n37975), .Z(n33516) );
  NOR U39929 ( .A(n40068), .B(n38759), .Z(n40067) );
  XOR U39930 ( .A(n40069), .B(n37977), .Z(n30370) );
  ANDN U39931 ( .B(n40070), .A(n37462), .Z(n40069) );
  IV U39932 ( .A(n40071), .Z(n37462) );
  XOR U39933 ( .A(n40072), .B(n40073), .Z(n32346) );
  XNOR U39934 ( .A(n25545), .B(n24845), .Z(n40073) );
  XNOR U39935 ( .A(n40074), .B(n28050), .Z(n24845) );
  IV U39936 ( .A(n27378), .Z(n28050) );
  XOR U39937 ( .A(n28811), .B(n38264), .Z(n27378) );
  XNOR U39938 ( .A(n40075), .B(n36008), .Z(n38264) );
  XNOR U39939 ( .A(n39960), .B(n39295), .Z(n35840) );
  XNOR U39940 ( .A(n40076), .B(n40077), .Z(n39960) );
  ANDN U39941 ( .B(n40078), .A(n40079), .Z(n40076) );
  XNOR U39942 ( .A(n32923), .B(n37828), .Z(n28811) );
  XNOR U39943 ( .A(n40080), .B(n40081), .Z(n37828) );
  XNOR U39944 ( .A(n27658), .B(n35999), .Z(n40081) );
  XOR U39945 ( .A(n40082), .B(n36011), .Z(n35999) );
  IV U39946 ( .A(n36415), .Z(n36011) );
  XOR U39947 ( .A(n38131), .B(n40083), .Z(n36415) );
  ANDN U39948 ( .B(n36012), .A(n38266), .Z(n40082) );
  XOR U39949 ( .A(n36356), .B(n40084), .Z(n38266) );
  XOR U39950 ( .A(n40085), .B(n40086), .Z(n36356) );
  XNOR U39951 ( .A(n40087), .B(n37884), .Z(n36012) );
  XNOR U39952 ( .A(n40088), .B(n36017), .Z(n27658) );
  XNOR U39953 ( .A(n39603), .B(n40089), .Z(n36017) );
  ANDN U39954 ( .B(n36018), .A(n35834), .Z(n40088) );
  XNOR U39955 ( .A(n40090), .B(n38163), .Z(n35834) );
  XOR U39956 ( .A(n40091), .B(n38298), .Z(n36018) );
  XNOR U39957 ( .A(n33135), .B(n40092), .Z(n40080) );
  XNOR U39958 ( .A(n35747), .B(n30675), .Z(n40092) );
  XNOR U39959 ( .A(n40093), .B(n36007), .Z(n30675) );
  XNOR U39960 ( .A(n40094), .B(n36434), .Z(n36007) );
  ANDN U39961 ( .B(n36008), .A(n35838), .Z(n40093) );
  XNOR U39962 ( .A(n40097), .B(n35159), .Z(n35838) );
  XNOR U39963 ( .A(n40098), .B(n40009), .Z(n35159) );
  XNOR U39964 ( .A(n40099), .B(n40100), .Z(n40009) );
  XNOR U39965 ( .A(n39684), .B(n39380), .Z(n40100) );
  XNOR U39966 ( .A(n40101), .B(n40102), .Z(n39380) );
  NOR U39967 ( .A(n40103), .B(n40104), .Z(n40101) );
  XNOR U39968 ( .A(n40105), .B(n40106), .Z(n39684) );
  AND U39969 ( .A(n40107), .B(n40108), .Z(n40105) );
  XOR U39970 ( .A(n35621), .B(n40109), .Z(n40099) );
  XNOR U39971 ( .A(n40110), .B(n39316), .Z(n40109) );
  XOR U39972 ( .A(n40111), .B(n40112), .Z(n39316) );
  ANDN U39973 ( .B(n40113), .A(n40114), .Z(n40111) );
  XNOR U39974 ( .A(n40115), .B(n40116), .Z(n35621) );
  NOR U39975 ( .A(n40117), .B(n40118), .Z(n40115) );
  XOR U39976 ( .A(n39051), .B(n39569), .Z(n36008) );
  XOR U39977 ( .A(n40119), .B(n40120), .Z(n39569) );
  XNOR U39978 ( .A(n40123), .B(n36015), .Z(n35747) );
  XNOR U39979 ( .A(n40124), .B(n39312), .Z(n36015) );
  XOR U39980 ( .A(n40125), .B(n36353), .Z(n35842) );
  IV U39981 ( .A(n39102), .Z(n36353) );
  XOR U39982 ( .A(n40126), .B(n40127), .Z(n39102) );
  XOR U39983 ( .A(n40128), .B(n39125), .Z(n36014) );
  XOR U39984 ( .A(n40129), .B(n36004), .Z(n33135) );
  XOR U39985 ( .A(n40130), .B(n34637), .Z(n36004) );
  IV U39986 ( .A(n37791), .Z(n34637) );
  XNOR U39987 ( .A(n40131), .B(n40132), .Z(n37791) );
  ANDN U39988 ( .B(n36005), .A(n35825), .Z(n40129) );
  XOR U39989 ( .A(n40133), .B(n40134), .Z(n35825) );
  XNOR U39990 ( .A(n35510), .B(n40135), .Z(n36005) );
  XOR U39991 ( .A(n40136), .B(n40137), .Z(n32923) );
  XNOR U39992 ( .A(n37898), .B(n32976), .Z(n40137) );
  XNOR U39993 ( .A(n40138), .B(n37924), .Z(n32976) );
  IV U39994 ( .A(n37319), .Z(n37924) );
  XNOR U39995 ( .A(n38124), .B(n40139), .Z(n37319) );
  ANDN U39996 ( .B(n33563), .A(n33564), .Z(n40138) );
  XOR U39997 ( .A(n40140), .B(n39389), .Z(n33564) );
  XOR U39998 ( .A(n40141), .B(n35323), .Z(n33563) );
  XOR U39999 ( .A(n40142), .B(n36194), .Z(n37898) );
  XOR U40000 ( .A(n40143), .B(n39938), .Z(n36194) );
  ANDN U40001 ( .B(n33567), .A(n33568), .Z(n40142) );
  XOR U40002 ( .A(n38146), .B(n40144), .Z(n33568) );
  IV U40003 ( .A(n39782), .Z(n38146) );
  XNOR U40004 ( .A(n40145), .B(n39603), .Z(n33567) );
  XOR U40005 ( .A(n32624), .B(n40146), .Z(n40136) );
  XNOR U40006 ( .A(n33408), .B(n30816), .Z(n40146) );
  XNOR U40007 ( .A(n40147), .B(n36188), .Z(n30816) );
  XOR U40008 ( .A(n40148), .B(n37272), .Z(n36188) );
  XOR U40009 ( .A(n40149), .B(n39075), .Z(n37272) );
  XNOR U40010 ( .A(n40150), .B(n40151), .Z(n39075) );
  XOR U40011 ( .A(n40152), .B(n40090), .Z(n40151) );
  XOR U40012 ( .A(n40153), .B(n40154), .Z(n40090) );
  ANDN U40013 ( .B(n40155), .A(n40156), .Z(n40153) );
  XOR U40014 ( .A(n40157), .B(n40158), .Z(n40150) );
  XOR U40015 ( .A(n38162), .B(n40159), .Z(n40158) );
  XNOR U40016 ( .A(n40160), .B(n40161), .Z(n38162) );
  NOR U40017 ( .A(n40162), .B(n40163), .Z(n40160) );
  ANDN U40018 ( .B(n33572), .A(n33573), .Z(n40147) );
  XOR U40019 ( .A(n40164), .B(n37055), .Z(n33573) );
  IV U40020 ( .A(n37032), .Z(n37055) );
  XNOR U40021 ( .A(n40165), .B(n39363), .Z(n37032) );
  XNOR U40022 ( .A(n40166), .B(n40167), .Z(n39363) );
  XOR U40023 ( .A(n36438), .B(n38314), .Z(n40167) );
  XNOR U40024 ( .A(n40168), .B(n40169), .Z(n38314) );
  NOR U40025 ( .A(n40170), .B(n40171), .Z(n40168) );
  XNOR U40026 ( .A(n40172), .B(n40173), .Z(n36438) );
  NOR U40027 ( .A(n40174), .B(n40175), .Z(n40172) );
  XNOR U40028 ( .A(n39226), .B(n40176), .Z(n40166) );
  XNOR U40029 ( .A(n38973), .B(n40177), .Z(n40176) );
  XNOR U40030 ( .A(n40178), .B(n40179), .Z(n38973) );
  ANDN U40031 ( .B(n40180), .A(n40181), .Z(n40178) );
  XOR U40032 ( .A(n40182), .B(n40183), .Z(n39226) );
  NOR U40033 ( .A(n40184), .B(n40185), .Z(n40182) );
  XNOR U40034 ( .A(n40187), .B(n36673), .Z(n33408) );
  XNOR U40035 ( .A(n40188), .B(n40189), .Z(n36673) );
  ANDN U40036 ( .B(n33578), .A(n33576), .Z(n40187) );
  XOR U40037 ( .A(n40190), .B(n38686), .Z(n33576) );
  IV U40038 ( .A(n37310), .Z(n33578) );
  XOR U40039 ( .A(n40191), .B(n37525), .Z(n37310) );
  XOR U40040 ( .A(n40192), .B(n40193), .Z(n37525) );
  XNOR U40041 ( .A(n40194), .B(n36196), .Z(n32624) );
  IV U40042 ( .A(n37921), .Z(n36196) );
  XOR U40043 ( .A(n40195), .B(n38929), .Z(n37921) );
  IV U40044 ( .A(n37884), .Z(n38929) );
  XOR U40045 ( .A(n40196), .B(n38255), .Z(n33581) );
  XOR U40046 ( .A(n40197), .B(n38587), .Z(n33580) );
  NOR U40047 ( .A(n28049), .B(n28986), .Z(n40074) );
  XOR U40048 ( .A(n40066), .B(n30371), .Z(n28986) );
  XNOR U40049 ( .A(n40198), .B(n40199), .Z(n38396) );
  XNOR U40050 ( .A(n29740), .B(n31234), .Z(n40199) );
  XNOR U40051 ( .A(n40200), .B(n39878), .Z(n31234) );
  XOR U40052 ( .A(n40201), .B(n40013), .Z(n39878) );
  XNOR U40053 ( .A(n40202), .B(n40203), .Z(n40013) );
  ANDN U40054 ( .B(n40204), .A(n40205), .Z(n40202) );
  ANDN U40055 ( .B(n38069), .A(n40206), .Z(n40200) );
  XOR U40056 ( .A(n40207), .B(n37964), .Z(n38069) );
  XNOR U40057 ( .A(n40208), .B(n36759), .Z(n29740) );
  XOR U40058 ( .A(n38906), .B(n40209), .Z(n36758) );
  XOR U40059 ( .A(n40210), .B(n40211), .Z(n38906) );
  XNOR U40060 ( .A(n29933), .B(n40212), .Z(n40198) );
  XOR U40061 ( .A(n30525), .B(n33208), .Z(n40212) );
  XOR U40062 ( .A(n40213), .B(n39872), .Z(n33208) );
  IV U40063 ( .A(n36744), .Z(n39872) );
  XOR U40064 ( .A(n40214), .B(n37030), .Z(n36744) );
  IV U40065 ( .A(n37714), .Z(n37030) );
  XOR U40066 ( .A(n40217), .B(n38360), .Z(n36745) );
  XNOR U40067 ( .A(n40218), .B(n36754), .Z(n30525) );
  XOR U40068 ( .A(n40219), .B(n33931), .Z(n36754) );
  ANDN U40069 ( .B(n36755), .A(n38413), .Z(n40218) );
  XNOR U40070 ( .A(n39019), .B(n40220), .Z(n36755) );
  XNOR U40071 ( .A(n40221), .B(n36748), .Z(n29933) );
  XNOR U40072 ( .A(n40222), .B(n38587), .Z(n36748) );
  IV U40073 ( .A(n37887), .Z(n38587) );
  XOR U40074 ( .A(n40095), .B(n40223), .Z(n37887) );
  XNOR U40075 ( .A(n40224), .B(n40225), .Z(n40095) );
  XNOR U40076 ( .A(n39611), .B(n37636), .Z(n40225) );
  XNOR U40077 ( .A(n40226), .B(n40227), .Z(n37636) );
  ANDN U40078 ( .B(n40228), .A(n40229), .Z(n40226) );
  XOR U40079 ( .A(n40230), .B(n40231), .Z(n39611) );
  ANDN U40080 ( .B(n40232), .A(n40233), .Z(n40230) );
  XOR U40081 ( .A(n37429), .B(n40234), .Z(n40224) );
  XOR U40082 ( .A(n39765), .B(n38747), .Z(n40234) );
  XNOR U40083 ( .A(n40235), .B(n40236), .Z(n38747) );
  AND U40084 ( .A(n40237), .B(n40238), .Z(n40235) );
  XOR U40085 ( .A(n40239), .B(n40240), .Z(n39765) );
  XNOR U40086 ( .A(n40243), .B(n40244), .Z(n37429) );
  ANDN U40087 ( .B(n40245), .A(n40246), .Z(n40243) );
  ANDN U40088 ( .B(n36749), .A(n38061), .Z(n40221) );
  XOR U40089 ( .A(n35787), .B(n40247), .Z(n36749) );
  XOR U40090 ( .A(n40248), .B(n39759), .Z(n35787) );
  XNOR U40091 ( .A(n40249), .B(n40250), .Z(n39759) );
  XOR U40092 ( .A(n40251), .B(n40252), .Z(n40250) );
  XOR U40093 ( .A(n37777), .B(n40253), .Z(n40249) );
  XOR U40094 ( .A(n36307), .B(n38086), .Z(n40253) );
  XNOR U40095 ( .A(n40254), .B(n40255), .Z(n38086) );
  ANDN U40096 ( .B(n40256), .A(n40257), .Z(n40254) );
  XNOR U40097 ( .A(n40258), .B(n40259), .Z(n36307) );
  ANDN U40098 ( .B(n40260), .A(n40261), .Z(n40258) );
  XNOR U40099 ( .A(n40262), .B(n40263), .Z(n37777) );
  AND U40100 ( .A(n40264), .B(n40265), .Z(n40262) );
  XOR U40101 ( .A(n40266), .B(n40267), .Z(n38699) );
  XOR U40102 ( .A(n36738), .B(n36496), .Z(n40267) );
  XNOR U40103 ( .A(n40268), .B(n35878), .Z(n36496) );
  XNOR U40104 ( .A(n40269), .B(n39307), .Z(n35878) );
  ANDN U40105 ( .B(n37980), .A(n40064), .Z(n40268) );
  XOR U40106 ( .A(n38719), .B(n40270), .Z(n37980) );
  XOR U40107 ( .A(n40271), .B(n35884), .Z(n36738) );
  IV U40108 ( .A(n37982), .Z(n35884) );
  XOR U40109 ( .A(n40272), .B(n39404), .Z(n37982) );
  ANDN U40110 ( .B(n37983), .A(n40273), .Z(n40271) );
  XNOR U40111 ( .A(n30199), .B(n40274), .Z(n40266) );
  XNOR U40112 ( .A(n32351), .B(n30770), .Z(n40274) );
  XNOR U40113 ( .A(n40275), .B(n35887), .Z(n30770) );
  XNOR U40114 ( .A(n40276), .B(n36783), .Z(n35887) );
  XNOR U40115 ( .A(n40277), .B(n38623), .Z(n36783) );
  XOR U40116 ( .A(n40278), .B(n40279), .Z(n38623) );
  XNOR U40117 ( .A(n38670), .B(n38998), .Z(n40279) );
  XNOR U40118 ( .A(n40280), .B(n40281), .Z(n38998) );
  NOR U40119 ( .A(n40282), .B(n40283), .Z(n40280) );
  XOR U40120 ( .A(n40284), .B(n40285), .Z(n38670) );
  NOR U40121 ( .A(n40286), .B(n40287), .Z(n40284) );
  XNOR U40122 ( .A(n38400), .B(n40288), .Z(n40278) );
  XNOR U40123 ( .A(n40289), .B(n38830), .Z(n40288) );
  XNOR U40124 ( .A(n40290), .B(n40291), .Z(n38830) );
  ANDN U40125 ( .B(n40292), .A(n40293), .Z(n40290) );
  XNOR U40126 ( .A(n40294), .B(n40295), .Z(n38400) );
  ANDN U40127 ( .B(n40296), .A(n40297), .Z(n40294) );
  XOR U40128 ( .A(n40298), .B(n37500), .Z(n37985) );
  XOR U40129 ( .A(n40299), .B(n37464), .Z(n32351) );
  XOR U40130 ( .A(n39001), .B(n40300), .Z(n37464) );
  IV U40131 ( .A(n37219), .Z(n39001) );
  XOR U40132 ( .A(n40302), .B(n40303), .Z(n40127) );
  XOR U40133 ( .A(n40304), .B(n36534), .Z(n40303) );
  XOR U40134 ( .A(n40305), .B(n40162), .Z(n36534) );
  ANDN U40135 ( .B(n40306), .A(n40307), .Z(n40305) );
  XOR U40136 ( .A(n36506), .B(n40308), .Z(n40302) );
  XNOR U40137 ( .A(n38579), .B(n38742), .Z(n40308) );
  XNOR U40138 ( .A(n40309), .B(n40310), .Z(n38742) );
  AND U40139 ( .A(n40311), .B(n40312), .Z(n40309) );
  XOR U40140 ( .A(n40313), .B(n40314), .Z(n38579) );
  ANDN U40141 ( .B(n40315), .A(n40316), .Z(n40313) );
  XNOR U40142 ( .A(n40317), .B(n40318), .Z(n36506) );
  ANDN U40143 ( .B(n40319), .A(n40320), .Z(n40317) );
  XOR U40144 ( .A(n40321), .B(n39431), .Z(n37977) );
  IV U40145 ( .A(n39838), .Z(n39431) );
  XOR U40146 ( .A(n40322), .B(n38760), .Z(n30199) );
  IV U40147 ( .A(n37974), .Z(n38760) );
  XNOR U40148 ( .A(n40323), .B(n39186), .Z(n37974) );
  ANDN U40149 ( .B(n37975), .A(n40324), .Z(n40322) );
  XOR U40150 ( .A(n40325), .B(n36390), .Z(n37975) );
  IV U40151 ( .A(n34617), .Z(n36390) );
  XNOR U40152 ( .A(n40326), .B(n37983), .Z(n40066) );
  XOR U40153 ( .A(n40327), .B(n35369), .Z(n37983) );
  IV U40154 ( .A(n38977), .Z(n35369) );
  XOR U40155 ( .A(n40328), .B(n40329), .Z(n38977) );
  ANDN U40156 ( .B(n40273), .A(n40330), .Z(n40326) );
  XOR U40157 ( .A(n37958), .B(n29722), .Z(n28049) );
  IV U40158 ( .A(n29941), .Z(n29722) );
  XOR U40159 ( .A(n39366), .B(n37299), .Z(n29941) );
  XNOR U40160 ( .A(n40331), .B(n40332), .Z(n37299) );
  XNOR U40161 ( .A(n29969), .B(n33366), .Z(n40332) );
  XOR U40162 ( .A(n40333), .B(n34435), .Z(n33366) );
  XOR U40163 ( .A(n40334), .B(n37267), .Z(n34435) );
  IV U40164 ( .A(n40189), .Z(n37267) );
  XNOR U40165 ( .A(n40335), .B(n40336), .Z(n40189) );
  ANDN U40166 ( .B(n34436), .A(n37903), .Z(n40333) );
  XNOR U40167 ( .A(n37715), .B(n40337), .Z(n37903) );
  IV U40168 ( .A(n38033), .Z(n37715) );
  XNOR U40169 ( .A(n40338), .B(n40339), .Z(n38033) );
  XOR U40170 ( .A(n40340), .B(n38332), .Z(n34436) );
  XOR U40171 ( .A(n40341), .B(n35288), .Z(n29969) );
  XNOR U40172 ( .A(n40342), .B(n38843), .Z(n35288) );
  XOR U40173 ( .A(n40343), .B(n37931), .Z(n35291) );
  IV U40174 ( .A(n35376), .Z(n37931) );
  XOR U40175 ( .A(n40344), .B(n36710), .Z(n37915) );
  IV U40176 ( .A(n34368), .Z(n36710) );
  XNOR U40177 ( .A(n30249), .B(n40345), .Z(n40331) );
  XOR U40178 ( .A(n32264), .B(n31170), .Z(n40345) );
  XNOR U40179 ( .A(n40346), .B(n33596), .Z(n31170) );
  XOR U40180 ( .A(n40347), .B(n35634), .Z(n33596) );
  XNOR U40181 ( .A(n40348), .B(n40349), .Z(n35634) );
  XOR U40182 ( .A(n38518), .B(n40350), .Z(n33595) );
  IV U40183 ( .A(n37794), .Z(n38518) );
  XNOR U40184 ( .A(n40351), .B(n40352), .Z(n37794) );
  XNOR U40185 ( .A(n40353), .B(n37318), .Z(n37961) );
  IV U40186 ( .A(n39055), .Z(n37318) );
  XNOR U40187 ( .A(n40354), .B(n33726), .Z(n32264) );
  XOR U40188 ( .A(n40355), .B(n37163), .Z(n33726) );
  ANDN U40189 ( .B(n33727), .A(n37907), .Z(n40354) );
  IV U40190 ( .A(n40356), .Z(n37907) );
  XOR U40191 ( .A(n40357), .B(n33588), .Z(n30249) );
  XOR U40192 ( .A(n40358), .B(n36215), .Z(n33588) );
  IV U40193 ( .A(n37683), .Z(n36215) );
  ANDN U40194 ( .B(n37911), .A(n37952), .Z(n40357) );
  XOR U40195 ( .A(n40359), .B(n40360), .Z(n35792) );
  XOR U40196 ( .A(n40361), .B(n40362), .Z(n39497) );
  ANDN U40197 ( .B(n40363), .A(n40364), .Z(n40361) );
  XNOR U40198 ( .A(n40365), .B(n37928), .Z(n37911) );
  XOR U40199 ( .A(n40366), .B(n40367), .Z(n39366) );
  XNOR U40200 ( .A(n31395), .B(n32560), .Z(n40367) );
  XOR U40201 ( .A(n40368), .B(n36207), .Z(n32560) );
  XOR U40202 ( .A(n39021), .B(n40369), .Z(n36207) );
  IV U40203 ( .A(n36899), .Z(n39021) );
  XNOR U40204 ( .A(n40370), .B(n40371), .Z(n36899) );
  ANDN U40205 ( .B(n33657), .A(n34892), .Z(n40368) );
  XOR U40206 ( .A(n40372), .B(n39153), .Z(n34892) );
  IV U40207 ( .A(n35632), .Z(n39153) );
  XOR U40208 ( .A(n40375), .B(n37331), .Z(n33657) );
  XOR U40209 ( .A(n40376), .B(n33667), .Z(n31395) );
  XNOR U40210 ( .A(n40377), .B(n37687), .Z(n33667) );
  IV U40211 ( .A(n36794), .Z(n37687) );
  XNOR U40212 ( .A(n40379), .B(n40380), .Z(n39834) );
  XNOR U40213 ( .A(n38359), .B(n40381), .Z(n40380) );
  XNOR U40214 ( .A(n40382), .B(n40383), .Z(n38359) );
  NOR U40215 ( .A(n40384), .B(n40385), .Z(n40382) );
  XOR U40216 ( .A(n39471), .B(n40386), .Z(n40379) );
  XOR U40217 ( .A(n40387), .B(n40217), .Z(n40386) );
  XNOR U40218 ( .A(n40388), .B(n40389), .Z(n40217) );
  XOR U40219 ( .A(n40392), .B(n40393), .Z(n39471) );
  ANDN U40220 ( .B(n40394), .A(n40395), .Z(n40392) );
  ANDN U40221 ( .B(n33666), .A(n34888), .Z(n40376) );
  XNOR U40222 ( .A(n40396), .B(n38530), .Z(n34888) );
  XOR U40223 ( .A(n40152), .B(n38163), .Z(n33666) );
  XOR U40224 ( .A(n40397), .B(n40398), .Z(n40152) );
  NOR U40225 ( .A(n40318), .B(n40399), .Z(n40397) );
  XOR U40226 ( .A(n33628), .B(n40400), .Z(n40366) );
  XOR U40227 ( .A(n33646), .B(n32118), .Z(n40400) );
  XNOR U40228 ( .A(n40401), .B(n33663), .Z(n32118) );
  XOR U40229 ( .A(n40402), .B(n37163), .Z(n33663) );
  XOR U40230 ( .A(n39802), .B(n40403), .Z(n37163) );
  XOR U40231 ( .A(n40404), .B(n40405), .Z(n39802) );
  XNOR U40232 ( .A(n35612), .B(n38636), .Z(n40405) );
  XNOR U40233 ( .A(n40406), .B(n40407), .Z(n38636) );
  ANDN U40234 ( .B(n40408), .A(n40409), .Z(n40406) );
  XNOR U40235 ( .A(n40410), .B(n40411), .Z(n35612) );
  ANDN U40236 ( .B(n40412), .A(n40413), .Z(n40410) );
  XNOR U40237 ( .A(n39190), .B(n40414), .Z(n40404) );
  XOR U40238 ( .A(n38963), .B(n38855), .Z(n40414) );
  XOR U40239 ( .A(n40415), .B(n40416), .Z(n38855) );
  NOR U40240 ( .A(n40417), .B(n40418), .Z(n40415) );
  ANDN U40241 ( .B(n40421), .A(n40422), .Z(n40419) );
  XNOR U40242 ( .A(n40423), .B(n40424), .Z(n39190) );
  ANDN U40243 ( .B(n40425), .A(n40426), .Z(n40423) );
  ANDN U40244 ( .B(n33662), .A(n34895), .Z(n40401) );
  XOR U40245 ( .A(n40427), .B(n38444), .Z(n34895) );
  IV U40246 ( .A(n39596), .Z(n38444) );
  XNOR U40247 ( .A(n38242), .B(n40430), .Z(n33662) );
  XNOR U40248 ( .A(n40431), .B(n33653), .Z(n33646) );
  XOR U40249 ( .A(n40432), .B(n35627), .Z(n33653) );
  XNOR U40250 ( .A(n40433), .B(n40434), .Z(n35627) );
  NOR U40251 ( .A(n33652), .B(n34898), .Z(n40431) );
  XOR U40252 ( .A(n40435), .B(n40436), .Z(n34898) );
  XOR U40253 ( .A(n40437), .B(n39328), .Z(n33652) );
  XOR U40254 ( .A(n40438), .B(n36204), .Z(n33628) );
  XNOR U40255 ( .A(n35944), .B(n40439), .Z(n36204) );
  ANDN U40256 ( .B(n36220), .A(n34884), .Z(n40438) );
  XNOR U40257 ( .A(n35519), .B(n40440), .Z(n34884) );
  XNOR U40258 ( .A(n40441), .B(n40442), .Z(n35519) );
  XOR U40259 ( .A(n40443), .B(n36437), .Z(n36220) );
  XOR U40260 ( .A(n40444), .B(n39703), .Z(n36437) );
  XNOR U40261 ( .A(n40445), .B(n40446), .Z(n39703) );
  XOR U40262 ( .A(n40447), .B(n40448), .Z(n40446) );
  XNOR U40263 ( .A(n38437), .B(n40449), .Z(n40445) );
  XNOR U40264 ( .A(n39469), .B(n38882), .Z(n40449) );
  XNOR U40265 ( .A(n40450), .B(n40451), .Z(n38882) );
  NOR U40266 ( .A(n40452), .B(n40453), .Z(n40450) );
  XNOR U40267 ( .A(n40454), .B(n40455), .Z(n39469) );
  XOR U40268 ( .A(n40458), .B(n40459), .Z(n38437) );
  NOR U40269 ( .A(n40460), .B(n40461), .Z(n40458) );
  XNOR U40270 ( .A(n40462), .B(n33727), .Z(n37958) );
  XNOR U40271 ( .A(n38948), .B(n40463), .Z(n33727) );
  IV U40272 ( .A(n38306), .Z(n38948) );
  ANDN U40273 ( .B(n35279), .A(n40356), .Z(n40462) );
  XNOR U40274 ( .A(n40466), .B(n37187), .Z(n40356) );
  XOR U40275 ( .A(n40467), .B(n38096), .Z(n35279) );
  XNOR U40276 ( .A(n40470), .B(n27611), .Z(n25545) );
  XOR U40277 ( .A(n38789), .B(n30752), .Z(n27611) );
  XNOR U40278 ( .A(n32741), .B(n33446), .Z(n30752) );
  XOR U40279 ( .A(n40471), .B(n40472), .Z(n33446) );
  XNOR U40280 ( .A(n35892), .B(n31841), .Z(n40472) );
  XOR U40281 ( .A(n40473), .B(n36132), .Z(n31841) );
  XOR U40282 ( .A(n38535), .B(n40474), .Z(n36132) );
  ANDN U40283 ( .B(n36133), .A(n36840), .Z(n40473) );
  XOR U40284 ( .A(n40475), .B(n38419), .Z(n36840) );
  XOR U40285 ( .A(n40476), .B(n39307), .Z(n36133) );
  IV U40286 ( .A(n39947), .Z(n39307) );
  XOR U40287 ( .A(n40477), .B(n40478), .Z(n39947) );
  XNOR U40288 ( .A(n40479), .B(n36136), .Z(n35892) );
  XOR U40289 ( .A(n40480), .B(n37517), .Z(n36136) );
  AND U40290 ( .A(n36137), .B(n36854), .Z(n40479) );
  XOR U40291 ( .A(n32003), .B(n40481), .Z(n40471) );
  XOR U40292 ( .A(n33775), .B(n32307), .Z(n40481) );
  XNOR U40293 ( .A(n40482), .B(n36146), .Z(n32307) );
  XOR U40294 ( .A(n40483), .B(n37710), .Z(n36146) );
  XNOR U40295 ( .A(n40484), .B(n40485), .Z(n39155) );
  XOR U40296 ( .A(n35379), .B(n38834), .Z(n40485) );
  XNOR U40297 ( .A(n40486), .B(n40487), .Z(n38834) );
  XOR U40298 ( .A(n40490), .B(n40491), .Z(n35379) );
  ANDN U40299 ( .B(n40492), .A(n40493), .Z(n40490) );
  XOR U40300 ( .A(n35607), .B(n40494), .Z(n40484) );
  XOR U40301 ( .A(n39968), .B(n36371), .Z(n40494) );
  XNOR U40302 ( .A(n40495), .B(n40496), .Z(n36371) );
  ANDN U40303 ( .B(n40497), .A(n40498), .Z(n40495) );
  XNOR U40304 ( .A(n40499), .B(n40500), .Z(n39968) );
  ANDN U40305 ( .B(n40501), .A(n40502), .Z(n40499) );
  XNOR U40306 ( .A(n40503), .B(n40504), .Z(n35607) );
  AND U40307 ( .A(n36147), .B(n36848), .Z(n40482) );
  XOR U40308 ( .A(n40508), .B(n38934), .Z(n36848) );
  XOR U40309 ( .A(n40509), .B(n36212), .Z(n36147) );
  XNOR U40310 ( .A(n40510), .B(n38727), .Z(n33775) );
  XOR U40311 ( .A(n40511), .B(n37646), .Z(n38727) );
  XOR U40312 ( .A(n40512), .B(n40513), .Z(n37646) );
  ANDN U40313 ( .B(n38755), .A(n36843), .Z(n40510) );
  IV U40314 ( .A(n38797), .Z(n36843) );
  XOR U40315 ( .A(n40514), .B(n40515), .Z(n38797) );
  XNOR U40316 ( .A(n40516), .B(n37802), .Z(n38755) );
  XNOR U40317 ( .A(n40517), .B(n36142), .Z(n32003) );
  XOR U40318 ( .A(n40518), .B(n37040), .Z(n36142) );
  XNOR U40319 ( .A(n40519), .B(n40520), .Z(n37040) );
  ANDN U40320 ( .B(n36851), .A(n38800), .Z(n40517) );
  XOR U40321 ( .A(n38325), .B(n40521), .Z(n38800) );
  XOR U40322 ( .A(n40522), .B(n38171), .Z(n36851) );
  XOR U40323 ( .A(n40523), .B(n40524), .Z(n32741) );
  XNOR U40324 ( .A(n33838), .B(n32360), .Z(n40524) );
  XOR U40325 ( .A(n40525), .B(n35909), .Z(n32360) );
  XNOR U40326 ( .A(n40526), .B(n33927), .Z(n35909) );
  NOR U40327 ( .A(n39351), .B(n35908), .Z(n40525) );
  XOR U40328 ( .A(n40527), .B(n39011), .Z(n35908) );
  XNOR U40329 ( .A(n40528), .B(n37802), .Z(n39351) );
  XNOR U40330 ( .A(n40531), .B(n35903), .Z(n33838) );
  XOR U40331 ( .A(n40532), .B(n39304), .Z(n35903) );
  IV U40332 ( .A(n38432), .Z(n39304) );
  XOR U40333 ( .A(n40533), .B(n40534), .Z(n38432) );
  NOR U40334 ( .A(n36832), .B(n35902), .Z(n40531) );
  XOR U40335 ( .A(n40535), .B(n39344), .Z(n35902) );
  XOR U40336 ( .A(n40536), .B(n39238), .Z(n36832) );
  XOR U40337 ( .A(n29316), .B(n40537), .Z(n40523) );
  XOR U40338 ( .A(n35707), .B(n34270), .Z(n40537) );
  XNOR U40339 ( .A(n40538), .B(n36236), .Z(n34270) );
  XNOR U40340 ( .A(n40539), .B(n40540), .Z(n36236) );
  NOR U40341 ( .A(n39360), .B(n36824), .Z(n40538) );
  XNOR U40342 ( .A(n40541), .B(n35630), .Z(n36824) );
  XNOR U40343 ( .A(n40543), .B(n40544), .Z(n38624) );
  XNOR U40344 ( .A(n36551), .B(n36984), .Z(n40544) );
  XNOR U40345 ( .A(n40545), .B(n40546), .Z(n36984) );
  ANDN U40346 ( .B(n40547), .A(n40548), .Z(n40545) );
  XNOR U40347 ( .A(n40549), .B(n40550), .Z(n36551) );
  AND U40348 ( .A(n40551), .B(n40552), .Z(n40549) );
  XOR U40349 ( .A(n39064), .B(n40553), .Z(n40543) );
  XOR U40350 ( .A(n39769), .B(n39801), .Z(n40553) );
  XNOR U40351 ( .A(n40554), .B(n40555), .Z(n39801) );
  ANDN U40352 ( .B(n40556), .A(n40557), .Z(n40554) );
  XNOR U40353 ( .A(n40558), .B(n40559), .Z(n39769) );
  ANDN U40354 ( .B(n40560), .A(n40561), .Z(n40558) );
  XNOR U40355 ( .A(n40562), .B(n40563), .Z(n39064) );
  ANDN U40356 ( .B(n40564), .A(n40565), .Z(n40562) );
  XOR U40357 ( .A(n40566), .B(n38419), .Z(n39360) );
  XNOR U40358 ( .A(n40567), .B(n35898), .Z(n35707) );
  XOR U40359 ( .A(n40568), .B(n40569), .Z(n35898) );
  NOR U40360 ( .A(n39314), .B(n35899), .Z(n40567) );
  XNOR U40361 ( .A(n40570), .B(n35510), .Z(n35899) );
  XOR U40362 ( .A(n40571), .B(n40572), .Z(n35510) );
  XOR U40363 ( .A(n40573), .B(n37258), .Z(n39314) );
  XNOR U40364 ( .A(n40574), .B(n35912), .Z(n29316) );
  XOR U40365 ( .A(n40575), .B(n38573), .Z(n35912) );
  ANDN U40366 ( .B(n36835), .A(n35913), .Z(n40574) );
  XOR U40367 ( .A(n39936), .B(n40576), .Z(n35913) );
  XOR U40368 ( .A(n40577), .B(n37834), .Z(n36835) );
  IV U40369 ( .A(n39608), .Z(n37834) );
  XNOR U40370 ( .A(n40578), .B(n40579), .Z(n39608) );
  XNOR U40371 ( .A(n40580), .B(n36137), .Z(n38789) );
  XOR U40372 ( .A(n40581), .B(n36347), .Z(n36137) );
  XNOR U40373 ( .A(n40582), .B(n40583), .Z(n40542) );
  XOR U40374 ( .A(n40355), .B(n37162), .Z(n40583) );
  XOR U40375 ( .A(n40584), .B(n40418), .Z(n37162) );
  AND U40376 ( .A(n40585), .B(n40417), .Z(n40584) );
  XOR U40377 ( .A(n40586), .B(n40421), .Z(n40355) );
  AND U40378 ( .A(n40587), .B(n40422), .Z(n40586) );
  XOR U40379 ( .A(n40402), .B(n40588), .Z(n40582) );
  XNOR U40380 ( .A(n36444), .B(n37778), .Z(n40588) );
  XOR U40381 ( .A(n40589), .B(n40412), .Z(n37778) );
  AND U40382 ( .A(n40590), .B(n40413), .Z(n40589) );
  XNOR U40383 ( .A(n40591), .B(n40425), .Z(n36444) );
  ANDN U40384 ( .B(n40426), .A(n40592), .Z(n40591) );
  XNOR U40385 ( .A(n40593), .B(n40408), .Z(n40402) );
  XNOR U40386 ( .A(n40595), .B(n40596), .Z(n39236) );
  XOR U40387 ( .A(n39696), .B(n37876), .Z(n40596) );
  XNOR U40388 ( .A(n40597), .B(n40598), .Z(n37876) );
  XNOR U40389 ( .A(n40601), .B(n40602), .Z(n39696) );
  ANDN U40390 ( .B(n40603), .A(n40604), .Z(n40601) );
  XNOR U40391 ( .A(n37699), .B(n40605), .Z(n40595) );
  XOR U40392 ( .A(n40606), .B(n39444), .Z(n40605) );
  XNOR U40393 ( .A(n40607), .B(n39196), .Z(n39444) );
  AND U40394 ( .A(n40608), .B(n40609), .Z(n40607) );
  XNOR U40395 ( .A(n40610), .B(n39207), .Z(n37699) );
  AND U40396 ( .A(n40611), .B(n40612), .Z(n40610) );
  NOR U40397 ( .A(n36855), .B(n36854), .Z(n40580) );
  XNOR U40398 ( .A(n40613), .B(n39389), .Z(n36854) );
  XNOR U40399 ( .A(n40614), .B(n39996), .Z(n36855) );
  XOR U40400 ( .A(n40615), .B(n40616), .Z(n39996) );
  NOR U40401 ( .A(n28053), .B(n28990), .Z(n40470) );
  XNOR U40402 ( .A(n28038), .B(n40617), .Z(n40072) );
  XOR U40403 ( .A(n24524), .B(n26503), .Z(n40617) );
  XNOR U40404 ( .A(n40618), .B(n27371), .Z(n26503) );
  XOR U40405 ( .A(n35714), .B(n31783), .Z(n27371) );
  IV U40406 ( .A(n31834), .Z(n31783) );
  XNOR U40407 ( .A(n40619), .B(n40620), .Z(n36216) );
  XOR U40408 ( .A(n32285), .B(n31643), .Z(n40620) );
  XNOR U40409 ( .A(n40621), .B(n37574), .Z(n31643) );
  XOR U40410 ( .A(n40435), .B(n40622), .Z(n37574) );
  ANDN U40411 ( .B(n35716), .A(n39387), .Z(n40621) );
  XOR U40412 ( .A(n40623), .B(n36420), .Z(n39387) );
  XOR U40413 ( .A(n37323), .B(n40624), .Z(n35716) );
  IV U40414 ( .A(n40514), .Z(n37323) );
  XNOR U40415 ( .A(n40625), .B(n40626), .Z(n40514) );
  XOR U40416 ( .A(n40627), .B(n37823), .Z(n32285) );
  XOR U40417 ( .A(n40628), .B(n35778), .Z(n37823) );
  XNOR U40418 ( .A(n40629), .B(n40630), .Z(n35778) );
  NOR U40419 ( .A(n40631), .B(n39384), .Z(n40627) );
  XNOR U40420 ( .A(n32059), .B(n40632), .Z(n40619) );
  XOR U40421 ( .A(n32356), .B(n37549), .Z(n40632) );
  XOR U40422 ( .A(n40633), .B(n37582), .Z(n37549) );
  XOR U40423 ( .A(n39202), .B(n37025), .Z(n37582) );
  IV U40424 ( .A(n37939), .Z(n37025) );
  XNOR U40425 ( .A(n40634), .B(n40635), .Z(n39202) );
  ANDN U40426 ( .B(n37583), .A(n39379), .Z(n40633) );
  XOR U40427 ( .A(n40637), .B(n39284), .Z(n39379) );
  XOR U40428 ( .A(n40638), .B(n38895), .Z(n37583) );
  IV U40429 ( .A(n39692), .Z(n38895) );
  XNOR U40430 ( .A(n40639), .B(n37571), .Z(n32356) );
  XOR U40431 ( .A(n39722), .B(n35078), .Z(n37571) );
  IV U40432 ( .A(n38766), .Z(n35078) );
  XNOR U40433 ( .A(n40642), .B(n40643), .Z(n39722) );
  NOR U40434 ( .A(n40644), .B(n40645), .Z(n40642) );
  ANDN U40435 ( .B(n35726), .A(n35728), .Z(n40639) );
  XOR U40436 ( .A(n35522), .B(n40646), .Z(n35728) );
  XOR U40437 ( .A(n40647), .B(n39530), .Z(n35726) );
  XNOR U40438 ( .A(n40648), .B(n37579), .Z(n32059) );
  IV U40439 ( .A(n37814), .Z(n37579) );
  XOR U40440 ( .A(n40649), .B(n38184), .Z(n37814) );
  NOR U40441 ( .A(n39370), .B(n35722), .Z(n40648) );
  XNOR U40442 ( .A(n40650), .B(n38113), .Z(n35722) );
  XNOR U40443 ( .A(n37018), .B(n40651), .Z(n39370) );
  XOR U40444 ( .A(n40652), .B(n40653), .Z(n35501) );
  XNOR U40445 ( .A(n33798), .B(n31697), .Z(n40653) );
  XOR U40446 ( .A(n40654), .B(n37562), .Z(n31697) );
  XNOR U40447 ( .A(n37005), .B(n40655), .Z(n37562) );
  ANDN U40448 ( .B(n37563), .A(n35205), .Z(n40654) );
  XNOR U40449 ( .A(n40656), .B(n35366), .Z(n35205) );
  IV U40450 ( .A(n39976), .Z(n35366) );
  XNOR U40451 ( .A(n40657), .B(n40658), .Z(n37563) );
  XOR U40452 ( .A(n40659), .B(n37556), .Z(n33798) );
  XOR U40453 ( .A(n40660), .B(n38283), .Z(n37556) );
  IV U40454 ( .A(n37841), .Z(n38283) );
  XNOR U40455 ( .A(n40661), .B(n40662), .Z(n37841) );
  ANDN U40456 ( .B(n37555), .A(n37748), .Z(n40659) );
  XOR U40457 ( .A(n34626), .B(n40663), .Z(n37748) );
  XNOR U40458 ( .A(n40664), .B(n37258), .Z(n37555) );
  XOR U40459 ( .A(n32700), .B(n40665), .Z(n40652) );
  XOR U40460 ( .A(n29283), .B(n35048), .Z(n40665) );
  XNOR U40461 ( .A(n40666), .B(n38540), .Z(n35048) );
  XOR U40462 ( .A(n40667), .B(n39523), .Z(n38540) );
  IV U40463 ( .A(n38255), .Z(n39523) );
  NOR U40464 ( .A(n35199), .B(n37751), .Z(n40666) );
  XOR U40465 ( .A(n40668), .B(n38120), .Z(n37751) );
  IV U40466 ( .A(n36537), .Z(n38120) );
  XNOR U40467 ( .A(n40669), .B(n37964), .Z(n35199) );
  IV U40468 ( .A(n40540), .Z(n37964) );
  XOR U40469 ( .A(n40670), .B(n37560), .Z(n29283) );
  XOR U40470 ( .A(n40671), .B(n40672), .Z(n37560) );
  NOR U40471 ( .A(n37559), .B(n35209), .Z(n40670) );
  XOR U40472 ( .A(n39336), .B(n40673), .Z(n35209) );
  IV U40473 ( .A(n35586), .Z(n39336) );
  XOR U40474 ( .A(n40351), .B(n40674), .Z(n35586) );
  XOR U40475 ( .A(n40675), .B(n40676), .Z(n40351) );
  XNOR U40476 ( .A(n40343), .B(n39682), .Z(n40676) );
  XNOR U40477 ( .A(n40677), .B(n40678), .Z(n39682) );
  NOR U40478 ( .A(n40679), .B(n40680), .Z(n40677) );
  XNOR U40479 ( .A(n40681), .B(n40682), .Z(n40343) );
  ANDN U40480 ( .B(n40683), .A(n40684), .Z(n40681) );
  XNOR U40481 ( .A(n35375), .B(n40685), .Z(n40675) );
  XOR U40482 ( .A(n37930), .B(n40686), .Z(n40685) );
  XNOR U40483 ( .A(n40687), .B(n40018), .Z(n37930) );
  ANDN U40484 ( .B(n40688), .A(n40689), .Z(n40687) );
  XNOR U40485 ( .A(n40690), .B(n40204), .Z(n35375) );
  NOR U40486 ( .A(n40691), .B(n40692), .Z(n40690) );
  XOR U40487 ( .A(n40693), .B(n38719), .Z(n37559) );
  XNOR U40488 ( .A(n40694), .B(n37565), .Z(n32700) );
  XNOR U40489 ( .A(n37344), .B(n40695), .Z(n37565) );
  ANDN U40490 ( .B(n37566), .A(n35195), .Z(n40694) );
  XNOR U40491 ( .A(n40696), .B(n38440), .Z(n35195) );
  XOR U40492 ( .A(n40110), .B(n39315), .Z(n37566) );
  XNOR U40493 ( .A(n40697), .B(n40698), .Z(n39315) );
  XNOR U40494 ( .A(n40699), .B(n40700), .Z(n40110) );
  XNOR U40495 ( .A(n40703), .B(n37825), .Z(n35714) );
  IV U40496 ( .A(n40631), .Z(n37825) );
  XNOR U40497 ( .A(n40704), .B(n38124), .Z(n40631) );
  XNOR U40498 ( .A(n40706), .B(n40707), .Z(n40301) );
  XOR U40499 ( .A(n39231), .B(n40518), .Z(n40707) );
  XOR U40500 ( .A(n40708), .B(n40709), .Z(n40518) );
  ANDN U40501 ( .B(n40710), .A(n40711), .Z(n40708) );
  XNOR U40502 ( .A(n40712), .B(n40713), .Z(n39231) );
  NOR U40503 ( .A(n40714), .B(n40715), .Z(n40712) );
  XOR U40504 ( .A(n37039), .B(n40716), .Z(n40706) );
  XNOR U40505 ( .A(n39686), .B(n39645), .Z(n40716) );
  XOR U40506 ( .A(n40717), .B(n40718), .Z(n39645) );
  NOR U40507 ( .A(n40719), .B(n40720), .Z(n40717) );
  XNOR U40508 ( .A(n40721), .B(n40722), .Z(n39686) );
  NOR U40509 ( .A(n40723), .B(n40724), .Z(n40721) );
  XNOR U40510 ( .A(n40725), .B(n40726), .Z(n37039) );
  NOR U40511 ( .A(n40727), .B(n40728), .Z(n40725) );
  ANDN U40512 ( .B(n39384), .A(n37821), .Z(n40703) );
  XNOR U40513 ( .A(n40729), .B(n38734), .Z(n37821) );
  IV U40514 ( .A(n36367), .Z(n38734) );
  XOR U40515 ( .A(n40730), .B(n40132), .Z(n36367) );
  XNOR U40516 ( .A(n40731), .B(n40732), .Z(n40132) );
  XNOR U40517 ( .A(n40337), .B(n39241), .Z(n40732) );
  XOR U40518 ( .A(n40733), .B(n40734), .Z(n39241) );
  ANDN U40519 ( .B(n40735), .A(n40736), .Z(n40733) );
  XOR U40520 ( .A(n40737), .B(n40738), .Z(n40337) );
  AND U40521 ( .A(n40739), .B(n40740), .Z(n40737) );
  XNOR U40522 ( .A(n37716), .B(n40741), .Z(n40731) );
  XOR U40523 ( .A(n39772), .B(n38034), .Z(n40741) );
  XOR U40524 ( .A(n40742), .B(n40743), .Z(n38034) );
  ANDN U40525 ( .B(n40744), .A(n40745), .Z(n40742) );
  XOR U40526 ( .A(n40746), .B(n40747), .Z(n39772) );
  XOR U40527 ( .A(n40750), .B(n40751), .Z(n37716) );
  ANDN U40528 ( .B(n40752), .A(n40753), .Z(n40750) );
  XNOR U40529 ( .A(n40754), .B(n36541), .Z(n39384) );
  XNOR U40530 ( .A(n39674), .B(n40444), .Z(n36541) );
  XOR U40531 ( .A(n40755), .B(n40756), .Z(n40444) );
  XNOR U40532 ( .A(n39100), .B(n39994), .Z(n40756) );
  XNOR U40533 ( .A(n40757), .B(n40758), .Z(n39994) );
  ANDN U40534 ( .B(n40759), .A(n40760), .Z(n40757) );
  XNOR U40535 ( .A(n40761), .B(n40762), .Z(n39100) );
  ANDN U40536 ( .B(n40763), .A(n40764), .Z(n40761) );
  XNOR U40537 ( .A(n39254), .B(n40765), .Z(n40755) );
  XOR U40538 ( .A(n37706), .B(n40766), .Z(n40765) );
  XNOR U40539 ( .A(n40767), .B(n40768), .Z(n37706) );
  XNOR U40540 ( .A(n40771), .B(n40772), .Z(n39254) );
  ANDN U40541 ( .B(n40773), .A(n40774), .Z(n40771) );
  XOR U40542 ( .A(n40775), .B(n40776), .Z(n39674) );
  XNOR U40543 ( .A(n39361), .B(n38516), .Z(n40776) );
  XOR U40544 ( .A(n40777), .B(n40185), .Z(n38516) );
  ANDN U40545 ( .B(n40184), .A(n40778), .Z(n40777) );
  XOR U40546 ( .A(n40779), .B(n40175), .Z(n39361) );
  ANDN U40547 ( .B(n40174), .A(n40780), .Z(n40779) );
  XOR U40548 ( .A(n38942), .B(n40781), .Z(n40775) );
  XNOR U40549 ( .A(n37075), .B(n37496), .Z(n40781) );
  XOR U40550 ( .A(n40782), .B(n40171), .Z(n37496) );
  ANDN U40551 ( .B(n40170), .A(n40783), .Z(n40782) );
  XOR U40552 ( .A(n40784), .B(n40180), .Z(n37075) );
  ANDN U40553 ( .B(n40181), .A(n40785), .Z(n40784) );
  XOR U40554 ( .A(n40786), .B(n40787), .Z(n38942) );
  ANDN U40555 ( .B(n40788), .A(n40789), .Z(n40786) );
  NOR U40556 ( .A(n28046), .B(n28994), .Z(n40618) );
  XOR U40557 ( .A(n36932), .B(n29409), .Z(n28994) );
  XOR U40558 ( .A(n32256), .B(n34950), .Z(n29409) );
  XNOR U40559 ( .A(n40790), .B(n40791), .Z(n34950) );
  XNOR U40560 ( .A(n33442), .B(n34373), .Z(n40791) );
  XNOR U40561 ( .A(n40792), .B(n35219), .Z(n34373) );
  XOR U40562 ( .A(n40793), .B(n39372), .Z(n35219) );
  IV U40563 ( .A(n38544), .Z(n39372) );
  NOR U40564 ( .A(n35220), .B(n34410), .Z(n40792) );
  XOR U40565 ( .A(n38488), .B(n40794), .Z(n34410) );
  IV U40566 ( .A(n35944), .Z(n38488) );
  XOR U40567 ( .A(n40795), .B(n36450), .Z(n35220) );
  IV U40568 ( .A(n37002), .Z(n36450) );
  XNOR U40569 ( .A(n40796), .B(n35512), .Z(n33442) );
  XOR U40570 ( .A(n40797), .B(n37630), .Z(n35512) );
  NOR U40571 ( .A(n34418), .B(n35504), .Z(n40796) );
  XOR U40572 ( .A(n30904), .B(n40798), .Z(n40790) );
  XOR U40573 ( .A(n31685), .B(n31862), .Z(n40798) );
  XNOR U40574 ( .A(n40799), .B(n34386), .Z(n31862) );
  XNOR U40575 ( .A(n40800), .B(n38082), .Z(n34386) );
  XOR U40576 ( .A(n40801), .B(n40513), .Z(n38082) );
  XNOR U40577 ( .A(n40802), .B(n40803), .Z(n40513) );
  XNOR U40578 ( .A(n40804), .B(n39321), .Z(n40803) );
  XNOR U40579 ( .A(n40805), .B(n40806), .Z(n39321) );
  XOR U40580 ( .A(n39531), .B(n40809), .Z(n40802) );
  XOR U40581 ( .A(n38342), .B(n39258), .Z(n40809) );
  XOR U40582 ( .A(n40810), .B(n40811), .Z(n39258) );
  ANDN U40583 ( .B(n40812), .A(n40813), .Z(n40810) );
  XOR U40584 ( .A(n40814), .B(n40815), .Z(n38342) );
  ANDN U40585 ( .B(n40816), .A(n40817), .Z(n40814) );
  XNOR U40586 ( .A(n40818), .B(n40819), .Z(n39531) );
  ANDN U40587 ( .B(n40820), .A(n40821), .Z(n40818) );
  ANDN U40588 ( .B(n34387), .A(n34415), .Z(n40799) );
  XOR U40589 ( .A(n39787), .B(n40822), .Z(n34415) );
  XOR U40590 ( .A(n40823), .B(n39262), .Z(n34387) );
  IV U40591 ( .A(n36202), .Z(n39262) );
  XNOR U40592 ( .A(n40824), .B(n34390), .Z(n31685) );
  XOR U40593 ( .A(n40825), .B(n39406), .Z(n34390) );
  NOR U40594 ( .A(n36944), .B(n34407), .Z(n40824) );
  XOR U40595 ( .A(n40826), .B(n40827), .Z(n34407) );
  XOR U40596 ( .A(n40828), .B(n35373), .Z(n36944) );
  IV U40597 ( .A(n37804), .Z(n35373) );
  XOR U40598 ( .A(n40829), .B(n40830), .Z(n37804) );
  XNOR U40599 ( .A(n40831), .B(n34380), .Z(n30904) );
  XNOR U40600 ( .A(n40832), .B(n37500), .Z(n34380) );
  ANDN U40601 ( .B(n34422), .A(n34381), .Z(n40831) );
  XOR U40602 ( .A(n40833), .B(n39847), .Z(n34381) );
  IV U40603 ( .A(n37437), .Z(n39847) );
  XOR U40604 ( .A(n39191), .B(n40834), .Z(n37437) );
  XOR U40605 ( .A(n40835), .B(n40836), .Z(n39191) );
  XNOR U40606 ( .A(n39007), .B(n37872), .Z(n40836) );
  XNOR U40607 ( .A(n40837), .B(n40838), .Z(n37872) );
  NOR U40608 ( .A(n40420), .B(n40421), .Z(n40837) );
  XNOR U40609 ( .A(n40839), .B(n40840), .Z(n40421) );
  XNOR U40610 ( .A(n40841), .B(n40842), .Z(n39007) );
  NOR U40611 ( .A(n40424), .B(n40425), .Z(n40841) );
  XNOR U40612 ( .A(n40843), .B(n40844), .Z(n40425) );
  XOR U40613 ( .A(n36995), .B(n40845), .Z(n40835) );
  XOR U40614 ( .A(n39104), .B(n37858), .Z(n40845) );
  XNOR U40615 ( .A(n40846), .B(n40847), .Z(n37858) );
  NOR U40616 ( .A(n40412), .B(n40411), .Z(n40846) );
  XOR U40617 ( .A(n40848), .B(n40849), .Z(n40412) );
  XNOR U40618 ( .A(n40850), .B(n40851), .Z(n39104) );
  XNOR U40619 ( .A(n40852), .B(n40853), .Z(n40418) );
  XNOR U40620 ( .A(n40854), .B(n40855), .Z(n36995) );
  NOR U40621 ( .A(n40407), .B(n40408), .Z(n40854) );
  XOR U40622 ( .A(n40856), .B(n40857), .Z(n40408) );
  IV U40623 ( .A(n40858), .Z(n40407) );
  XOR U40624 ( .A(n40859), .B(n35606), .Z(n34422) );
  XNOR U40625 ( .A(n39888), .B(n39110), .Z(n35606) );
  XOR U40626 ( .A(n40860), .B(n40861), .Z(n39110) );
  XNOR U40627 ( .A(n40862), .B(n39610), .Z(n40861) );
  XNOR U40628 ( .A(n40863), .B(n40864), .Z(n39610) );
  ANDN U40629 ( .B(n40865), .A(n40866), .Z(n40863) );
  XOR U40630 ( .A(n38715), .B(n40867), .Z(n40860) );
  XOR U40631 ( .A(n35927), .B(n40868), .Z(n40867) );
  XNOR U40632 ( .A(n40869), .B(n40870), .Z(n35927) );
  ANDN U40633 ( .B(n40871), .A(n40872), .Z(n40869) );
  XOR U40634 ( .A(n40873), .B(n40874), .Z(n38715) );
  AND U40635 ( .A(n40875), .B(n40876), .Z(n40873) );
  XNOR U40636 ( .A(n40877), .B(n40878), .Z(n39888) );
  XNOR U40637 ( .A(n39456), .B(n38183), .Z(n40878) );
  XNOR U40638 ( .A(n40879), .B(n40880), .Z(n38183) );
  ANDN U40639 ( .B(n40881), .A(n40882), .Z(n40879) );
  XOR U40640 ( .A(n40883), .B(n40884), .Z(n39456) );
  ANDN U40641 ( .B(n40885), .A(n40886), .Z(n40883) );
  XNOR U40642 ( .A(n40887), .B(n40888), .Z(n40877) );
  XOR U40643 ( .A(n40649), .B(n38911), .Z(n40888) );
  XNOR U40644 ( .A(n40889), .B(n40890), .Z(n38911) );
  ANDN U40645 ( .B(n40891), .A(n40892), .Z(n40889) );
  XNOR U40646 ( .A(n40893), .B(n40894), .Z(n40649) );
  ANDN U40647 ( .B(n40895), .A(n40896), .Z(n40893) );
  XNOR U40648 ( .A(n40897), .B(n40898), .Z(n32256) );
  XNOR U40649 ( .A(n33833), .B(n33555), .Z(n40898) );
  XNOR U40650 ( .A(n40899), .B(n40029), .Z(n33555) );
  XNOR U40651 ( .A(n40900), .B(n39657), .Z(n40029) );
  IV U40652 ( .A(n35311), .Z(n39657) );
  ANDN U40653 ( .B(n40039), .A(n33895), .Z(n40899) );
  XNOR U40654 ( .A(n40901), .B(n37894), .Z(n33833) );
  XOR U40655 ( .A(n34618), .B(n40902), .Z(n37894) );
  XOR U40656 ( .A(n33323), .B(n40903), .Z(n40897) );
  XOR U40657 ( .A(n32582), .B(n34977), .Z(n40903) );
  XNOR U40658 ( .A(n40904), .B(n34983), .Z(n34977) );
  XOR U40659 ( .A(n40887), .B(n38184), .Z(n34983) );
  IV U40660 ( .A(n38912), .Z(n38184) );
  XOR U40661 ( .A(n40907), .B(n40908), .Z(n40887) );
  ANDN U40662 ( .B(n40909), .A(n40910), .Z(n40907) );
  XNOR U40663 ( .A(n40911), .B(n34987), .Z(n32582) );
  XOR U40664 ( .A(n40201), .B(n40012), .Z(n34987) );
  XOR U40665 ( .A(n40912), .B(n40913), .Z(n40012) );
  IV U40666 ( .A(n35772), .Z(n40201) );
  NOR U40667 ( .A(n40915), .B(n40916), .Z(n40911) );
  XNOR U40668 ( .A(n40917), .B(n34993), .Z(n33323) );
  XNOR U40669 ( .A(n37216), .B(n40918), .Z(n34993) );
  IV U40670 ( .A(n36979), .Z(n37216) );
  XNOR U40671 ( .A(n40919), .B(n40920), .Z(n36979) );
  ANDN U40672 ( .B(n34994), .A(n33899), .Z(n40917) );
  IV U40673 ( .A(n40921), .Z(n33899) );
  XNOR U40674 ( .A(n40922), .B(n35504), .Z(n36932) );
  XNOR U40675 ( .A(n34618), .B(n40923), .Z(n35504) );
  XNOR U40676 ( .A(n40193), .B(n40924), .Z(n34618) );
  XNOR U40677 ( .A(n40925), .B(n40926), .Z(n40193) );
  XOR U40678 ( .A(n40083), .B(n38132), .Z(n40926) );
  XNOR U40679 ( .A(n40927), .B(n40928), .Z(n38132) );
  ANDN U40680 ( .B(n40929), .A(n40870), .Z(n40927) );
  IV U40681 ( .A(n40930), .Z(n40870) );
  XOR U40682 ( .A(n40931), .B(n40932), .Z(n40083) );
  ANDN U40683 ( .B(n40874), .A(n40933), .Z(n40931) );
  XOR U40684 ( .A(n40934), .B(n40935), .Z(n40925) );
  XNOR U40685 ( .A(n40936), .B(n38547), .Z(n40935) );
  XNOR U40686 ( .A(n40937), .B(n40938), .Z(n38547) );
  ANDN U40687 ( .B(n40939), .A(n40940), .Z(n40937) );
  XOR U40688 ( .A(n40941), .B(n37044), .Z(n34418) );
  XOR U40689 ( .A(n40942), .B(n36963), .Z(n34420) );
  IV U40690 ( .A(n38332), .Z(n36963) );
  XOR U40691 ( .A(n40944), .B(n40945), .Z(n40215) );
  XNOR U40692 ( .A(n39373), .B(n38091), .Z(n40945) );
  XNOR U40693 ( .A(n40946), .B(n40947), .Z(n38091) );
  ANDN U40694 ( .B(n40948), .A(n40949), .Z(n40946) );
  XNOR U40695 ( .A(n40950), .B(n40951), .Z(n39373) );
  ANDN U40696 ( .B(n40952), .A(n40953), .Z(n40950) );
  XOR U40697 ( .A(n37869), .B(n40954), .Z(n40944) );
  XOR U40698 ( .A(n40955), .B(n40956), .Z(n40954) );
  XNOR U40699 ( .A(n40957), .B(n40958), .Z(n37869) );
  ANDN U40700 ( .B(n40959), .A(n40960), .Z(n40957) );
  XOR U40701 ( .A(n32193), .B(n39775), .Z(n28046) );
  XOR U40702 ( .A(n40961), .B(n36625), .Z(n39775) );
  ANDN U40703 ( .B(n37235), .A(n37236), .Z(n40961) );
  XOR U40704 ( .A(n40962), .B(n37314), .Z(n37236) );
  IV U40705 ( .A(n30760), .Z(n32193) );
  XOR U40706 ( .A(n38188), .B(n38987), .Z(n30760) );
  XNOR U40707 ( .A(n40963), .B(n40964), .Z(n38987) );
  XOR U40708 ( .A(n31589), .B(n32937), .Z(n40964) );
  XOR U40709 ( .A(n40965), .B(n36258), .Z(n32937) );
  XOR U40710 ( .A(n40966), .B(n39528), .Z(n36258) );
  NOR U40711 ( .A(n37214), .B(n36586), .Z(n40965) );
  XNOR U40712 ( .A(n40967), .B(n38100), .Z(n36586) );
  IV U40713 ( .A(n38564), .Z(n38100) );
  XNOR U40714 ( .A(n40968), .B(n39930), .Z(n37214) );
  XOR U40715 ( .A(n40969), .B(n36248), .Z(n31589) );
  XOR U40716 ( .A(n38520), .B(n40970), .Z(n36248) );
  IV U40717 ( .A(n35522), .Z(n38520) );
  XOR U40718 ( .A(n40971), .B(n40972), .Z(n35522) );
  ANDN U40719 ( .B(n37203), .A(n36583), .Z(n40969) );
  XOR U40720 ( .A(n40973), .B(n37968), .Z(n36583) );
  XOR U40721 ( .A(n40974), .B(n40428), .Z(n37968) );
  XNOR U40722 ( .A(n40975), .B(n40976), .Z(n40428) );
  XNOR U40723 ( .A(n39604), .B(n40977), .Z(n40976) );
  XOR U40724 ( .A(n40978), .B(n40979), .Z(n39604) );
  ANDN U40725 ( .B(n40980), .A(n40981), .Z(n40978) );
  XOR U40726 ( .A(n40982), .B(n40983), .Z(n40975) );
  XOR U40727 ( .A(n40145), .B(n40089), .Z(n40983) );
  XNOR U40728 ( .A(n40984), .B(n40985), .Z(n40089) );
  AND U40729 ( .A(n40986), .B(n40987), .Z(n40984) );
  XNOR U40730 ( .A(n40988), .B(n40989), .Z(n40145) );
  ANDN U40731 ( .B(n40990), .A(n40991), .Z(n40988) );
  XOR U40732 ( .A(n36560), .B(n40993), .Z(n40963) );
  XOR U40733 ( .A(n29165), .B(n30497), .Z(n40993) );
  XNOR U40734 ( .A(n40994), .B(n36252), .Z(n30497) );
  XOR U40735 ( .A(n40995), .B(n39938), .Z(n36252) );
  XNOR U40736 ( .A(n38899), .B(n40997), .Z(n37890) );
  XOR U40737 ( .A(n40998), .B(n40999), .Z(n38899) );
  XNOR U40738 ( .A(n38854), .B(n40532), .Z(n40999) );
  XOR U40739 ( .A(n41000), .B(n41001), .Z(n40532) );
  ANDN U40740 ( .B(n41002), .A(n41003), .Z(n41000) );
  XOR U40741 ( .A(n41004), .B(n41005), .Z(n38854) );
  ANDN U40742 ( .B(n41006), .A(n41007), .Z(n41004) );
  XOR U40743 ( .A(n39303), .B(n41008), .Z(n40998) );
  XNOR U40744 ( .A(n38431), .B(n38635), .Z(n41008) );
  XNOR U40745 ( .A(n41009), .B(n41010), .Z(n38635) );
  ANDN U40746 ( .B(n41011), .A(n41012), .Z(n41009) );
  XOR U40747 ( .A(n41013), .B(n41014), .Z(n38431) );
  ANDN U40748 ( .B(n41015), .A(n41016), .Z(n41013) );
  XNOR U40749 ( .A(n41017), .B(n41018), .Z(n39303) );
  AND U40750 ( .A(n41019), .B(n41020), .Z(n41017) );
  XOR U40751 ( .A(n40435), .B(n41021), .Z(n36588) );
  XNOR U40752 ( .A(n41022), .B(n36262), .Z(n29165) );
  XNOR U40753 ( .A(n41023), .B(n37008), .Z(n36262) );
  XNOR U40754 ( .A(n41025), .B(n41026), .Z(n40905) );
  XOR U40755 ( .A(n40052), .B(n39095), .Z(n41026) );
  XOR U40756 ( .A(n41027), .B(n41028), .Z(n39095) );
  ANDN U40757 ( .B(n40908), .A(n40909), .Z(n41027) );
  XOR U40758 ( .A(n41029), .B(n41030), .Z(n40052) );
  NOR U40759 ( .A(n40891), .B(n40890), .Z(n41029) );
  XOR U40760 ( .A(n40191), .B(n41031), .Z(n41025) );
  XOR U40761 ( .A(n37524), .B(n39658), .Z(n41031) );
  XNOR U40762 ( .A(n41032), .B(n41033), .Z(n39658) );
  ANDN U40763 ( .B(n40884), .A(n40885), .Z(n41032) );
  XOR U40764 ( .A(n41034), .B(n41035), .Z(n37524) );
  ANDN U40765 ( .B(n40896), .A(n40894), .Z(n41034) );
  XNOR U40766 ( .A(n41036), .B(n41037), .Z(n40191) );
  ANDN U40767 ( .B(n40882), .A(n40880), .Z(n41036) );
  NOR U40768 ( .A(n37765), .B(n36581), .Z(n41022) );
  XOR U40769 ( .A(n35604), .B(n41038), .Z(n36581) );
  XNOR U40770 ( .A(n41039), .B(n38889), .Z(n37765) );
  IV U40771 ( .A(n36303), .Z(n38889) );
  XNOR U40772 ( .A(n40328), .B(n41040), .Z(n36303) );
  XOR U40773 ( .A(n41041), .B(n41042), .Z(n40328) );
  XOR U40774 ( .A(n41043), .B(n38119), .Z(n41042) );
  XOR U40775 ( .A(n41044), .B(n41045), .Z(n38119) );
  ANDN U40776 ( .B(n41046), .A(n41047), .Z(n41044) );
  XNOR U40777 ( .A(n39473), .B(n41048), .Z(n41041) );
  XOR U40778 ( .A(n40668), .B(n36536), .Z(n41048) );
  XNOR U40779 ( .A(n41049), .B(n41050), .Z(n36536) );
  NOR U40780 ( .A(n41051), .B(n41052), .Z(n41049) );
  XNOR U40781 ( .A(n41053), .B(n41054), .Z(n40668) );
  NOR U40782 ( .A(n41055), .B(n41056), .Z(n41053) );
  XOR U40783 ( .A(n41057), .B(n41058), .Z(n39473) );
  ANDN U40784 ( .B(n41059), .A(n41060), .Z(n41057) );
  XNOR U40785 ( .A(n41061), .B(n36266), .Z(n36560) );
  XNOR U40786 ( .A(n39782), .B(n41062), .Z(n36266) );
  NOR U40787 ( .A(n36590), .B(n37218), .Z(n41061) );
  XOR U40788 ( .A(n40015), .B(n35772), .Z(n37218) );
  XNOR U40789 ( .A(n41063), .B(n40697), .Z(n35772) );
  XOR U40790 ( .A(n41064), .B(n41065), .Z(n40697) );
  XOR U40791 ( .A(n37540), .B(n41066), .Z(n41065) );
  XNOR U40792 ( .A(n41067), .B(n40692), .Z(n37540) );
  AND U40793 ( .A(n40205), .B(n40203), .Z(n41067) );
  XOR U40794 ( .A(n39078), .B(n41068), .Z(n41064) );
  XOR U40795 ( .A(n40826), .B(n36716), .Z(n41068) );
  XNOR U40796 ( .A(n41069), .B(n40689), .Z(n36716) );
  ANDN U40797 ( .B(n40017), .A(n40019), .Z(n41069) );
  XNOR U40798 ( .A(n41070), .B(n40684), .Z(n40826) );
  AND U40799 ( .A(n40914), .B(n40913), .Z(n41070) );
  XNOR U40800 ( .A(n41071), .B(n40680), .Z(n39078) );
  ANDN U40801 ( .B(n41072), .A(n41073), .Z(n41071) );
  XNOR U40802 ( .A(n41074), .B(n41072), .Z(n40015) );
  ANDN U40803 ( .B(n41073), .A(n40678), .Z(n41074) );
  IV U40804 ( .A(n41075), .Z(n40678) );
  XOR U40805 ( .A(n41076), .B(n37517), .Z(n36590) );
  XOR U40806 ( .A(n41079), .B(n41080), .Z(n38188) );
  XNOR U40807 ( .A(n31225), .B(n32524), .Z(n41080) );
  XOR U40808 ( .A(n41081), .B(n36616), .Z(n32524) );
  XOR U40809 ( .A(n41082), .B(n38885), .Z(n36616) );
  IV U40810 ( .A(n38325), .Z(n38885) );
  ANDN U40811 ( .B(n36617), .A(n37232), .Z(n41081) );
  XOR U40812 ( .A(n40133), .B(n41083), .Z(n37232) );
  IV U40813 ( .A(n38959), .Z(n40133) );
  XOR U40814 ( .A(n41084), .B(n39186), .Z(n36617) );
  XOR U40815 ( .A(n41085), .B(n39049), .Z(n31225) );
  IV U40816 ( .A(n36626), .Z(n39049) );
  XOR U40817 ( .A(n41086), .B(n37144), .Z(n36626) );
  IV U40818 ( .A(n39827), .Z(n37144) );
  XNOR U40819 ( .A(n41087), .B(n41088), .Z(n39827) );
  NOR U40820 ( .A(n36625), .B(n37235), .Z(n41085) );
  XOR U40821 ( .A(n41089), .B(n37479), .Z(n37235) );
  XNOR U40822 ( .A(n41090), .B(n38298), .Z(n36625) );
  XNOR U40823 ( .A(n41092), .B(n41093), .Z(n39970) );
  XOR U40824 ( .A(n39354), .B(n37701), .Z(n41093) );
  XOR U40825 ( .A(n41094), .B(n41095), .Z(n37701) );
  ANDN U40826 ( .B(n41096), .A(n41097), .Z(n41094) );
  XNOR U40827 ( .A(n41098), .B(n41099), .Z(n39354) );
  AND U40828 ( .A(n41100), .B(n41101), .Z(n41098) );
  XNOR U40829 ( .A(n37643), .B(n41102), .Z(n41092) );
  XNOR U40830 ( .A(n37422), .B(n35618), .Z(n41102) );
  XOR U40831 ( .A(n41103), .B(n41104), .Z(n35618) );
  AND U40832 ( .A(n41105), .B(n41106), .Z(n41103) );
  XNOR U40833 ( .A(n41107), .B(n41108), .Z(n37422) );
  ANDN U40834 ( .B(n41109), .A(n41110), .Z(n41107) );
  XOR U40835 ( .A(n41111), .B(n41112), .Z(n37643) );
  AND U40836 ( .A(n41113), .B(n41114), .Z(n41111) );
  XNOR U40837 ( .A(n35351), .B(n41115), .Z(n41079) );
  XOR U40838 ( .A(n30074), .B(n31681), .Z(n41115) );
  XNOR U40839 ( .A(n41116), .B(n36629), .Z(n31681) );
  XOR U40840 ( .A(n35323), .B(n41117), .Z(n36629) );
  IV U40841 ( .A(n39088), .Z(n35323) );
  ANDN U40842 ( .B(n36630), .A(n37227), .Z(n41116) );
  XOR U40843 ( .A(n41118), .B(n40435), .Z(n37227) );
  IV U40844 ( .A(n38142), .Z(n40435) );
  XNOR U40845 ( .A(n40248), .B(n41119), .Z(n38142) );
  XOR U40846 ( .A(n41120), .B(n41121), .Z(n40248) );
  XOR U40847 ( .A(n41122), .B(n39343), .Z(n41121) );
  XNOR U40848 ( .A(n41123), .B(n41124), .Z(n39343) );
  ANDN U40849 ( .B(n41125), .A(n41126), .Z(n41123) );
  XNOR U40850 ( .A(n41127), .B(n41128), .Z(n41120) );
  XNOR U40851 ( .A(n38252), .B(n40535), .Z(n41128) );
  XNOR U40852 ( .A(n41129), .B(n41130), .Z(n40535) );
  AND U40853 ( .A(n41131), .B(n41132), .Z(n41129) );
  XOR U40854 ( .A(n41133), .B(n41134), .Z(n38252) );
  ANDN U40855 ( .B(n41135), .A(n41136), .Z(n41133) );
  XNOR U40856 ( .A(n41137), .B(n37258), .Z(n36630) );
  XNOR U40857 ( .A(n41138), .B(n36633), .Z(n30074) );
  XOR U40858 ( .A(n41139), .B(n39269), .Z(n36633) );
  IV U40859 ( .A(n39404), .Z(n39269) );
  ANDN U40860 ( .B(n36634), .A(n37224), .Z(n41138) );
  XOR U40861 ( .A(n41140), .B(n38944), .Z(n37224) );
  XOR U40862 ( .A(n41066), .B(n36717), .Z(n36634) );
  IV U40863 ( .A(n40827), .Z(n36717) );
  XNOR U40864 ( .A(n41143), .B(n41144), .Z(n41066) );
  ANDN U40865 ( .B(n40021), .A(n40022), .Z(n41143) );
  XOR U40866 ( .A(n41145), .B(n39045), .Z(n35351) );
  IV U40867 ( .A(n36620), .Z(n39045) );
  XOR U40868 ( .A(n41146), .B(n36976), .Z(n36620) );
  ANDN U40869 ( .B(n36621), .A(n39777), .Z(n41145) );
  XOR U40870 ( .A(n39019), .B(n41149), .Z(n39777) );
  IV U40871 ( .A(n36408), .Z(n39019) );
  XNOR U40872 ( .A(n41150), .B(n41151), .Z(n36408) );
  XNOR U40873 ( .A(n39930), .B(n41152), .Z(n36621) );
  XOR U40874 ( .A(n41153), .B(n27382), .Z(n24524) );
  XOR U40875 ( .A(n34506), .B(n31560), .Z(n27382) );
  IV U40876 ( .A(n30768), .Z(n31560) );
  XNOR U40877 ( .A(n36173), .B(n38235), .Z(n30768) );
  XNOR U40878 ( .A(n41154), .B(n41155), .Z(n38235) );
  XNOR U40879 ( .A(n31329), .B(n31465), .Z(n41155) );
  XNOR U40880 ( .A(n41156), .B(n35685), .Z(n31465) );
  XOR U40881 ( .A(n41157), .B(n36320), .Z(n35685) );
  IV U40882 ( .A(n38151), .Z(n36320) );
  ANDN U40883 ( .B(n34521), .A(n34522), .Z(n41156) );
  XNOR U40884 ( .A(n41158), .B(n37187), .Z(n34522) );
  XNOR U40885 ( .A(n39299), .B(n41159), .Z(n37187) );
  XOR U40886 ( .A(n41160), .B(n41161), .Z(n39299) );
  XOR U40887 ( .A(n37050), .B(n38098), .Z(n41161) );
  XNOR U40888 ( .A(n41162), .B(n41163), .Z(n38098) );
  ANDN U40889 ( .B(n41164), .A(n41165), .Z(n41162) );
  XNOR U40890 ( .A(n41166), .B(n41167), .Z(n37050) );
  ANDN U40891 ( .B(n41168), .A(n41169), .Z(n41166) );
  XNOR U40892 ( .A(n41170), .B(n41171), .Z(n41160) );
  XOR U40893 ( .A(n39980), .B(n39455), .Z(n41171) );
  XNOR U40894 ( .A(n41172), .B(n41173), .Z(n39455) );
  ANDN U40895 ( .B(n41174), .A(n41175), .Z(n41172) );
  XNOR U40896 ( .A(n41176), .B(n41177), .Z(n39980) );
  AND U40897 ( .A(n41178), .B(n41179), .Z(n41176) );
  XOR U40898 ( .A(n38883), .B(n41180), .Z(n34521) );
  XOR U40899 ( .A(n41181), .B(n36021), .Z(n31329) );
  XOR U40900 ( .A(n41182), .B(n37725), .Z(n36021) );
  IV U40901 ( .A(n39468), .Z(n37725) );
  ANDN U40902 ( .B(n34513), .A(n38682), .Z(n41181) );
  IV U40903 ( .A(n34515), .Z(n38682) );
  XOR U40904 ( .A(n40447), .B(n38438), .Z(n34515) );
  XNOR U40905 ( .A(n41183), .B(n41184), .Z(n40447) );
  XOR U40906 ( .A(n41187), .B(n38248), .Z(n34513) );
  XOR U40907 ( .A(n40572), .B(n39747), .Z(n38248) );
  XNOR U40908 ( .A(n41188), .B(n41189), .Z(n39747) );
  XOR U40909 ( .A(n36906), .B(n39409), .Z(n41189) );
  XNOR U40910 ( .A(n41190), .B(n41191), .Z(n39409) );
  ANDN U40911 ( .B(n41192), .A(n41193), .Z(n41190) );
  XOR U40912 ( .A(n41194), .B(n41195), .Z(n36906) );
  ANDN U40913 ( .B(n41196), .A(n41197), .Z(n41194) );
  XOR U40914 ( .A(n37308), .B(n41198), .Z(n41188) );
  XOR U40915 ( .A(n41199), .B(n39275), .Z(n41198) );
  XNOR U40916 ( .A(n41200), .B(n41201), .Z(n39275) );
  NOR U40917 ( .A(n41202), .B(n41203), .Z(n41200) );
  XNOR U40918 ( .A(n41204), .B(n41205), .Z(n37308) );
  NOR U40919 ( .A(n41206), .B(n41207), .Z(n41204) );
  XNOR U40920 ( .A(n41208), .B(n41209), .Z(n40572) );
  XOR U40921 ( .A(n39189), .B(n41210), .Z(n41209) );
  XNOR U40922 ( .A(n41211), .B(n41212), .Z(n39189) );
  NOR U40923 ( .A(n41213), .B(n41214), .Z(n41211) );
  XNOR U40924 ( .A(n39063), .B(n41215), .Z(n41208) );
  XOR U40925 ( .A(n38984), .B(n38127), .Z(n41215) );
  XNOR U40926 ( .A(n41216), .B(n41217), .Z(n38127) );
  ANDN U40927 ( .B(n41218), .A(n41219), .Z(n41216) );
  XNOR U40928 ( .A(n41220), .B(n41221), .Z(n38984) );
  NOR U40929 ( .A(n41222), .B(n41223), .Z(n41220) );
  XNOR U40930 ( .A(n41224), .B(n41225), .Z(n39063) );
  NOR U40931 ( .A(n41226), .B(n41227), .Z(n41224) );
  XNOR U40932 ( .A(n31241), .B(n41228), .Z(n41154) );
  XOR U40933 ( .A(n32276), .B(n34226), .Z(n41228) );
  XNOR U40934 ( .A(n41229), .B(n35682), .Z(n34226) );
  XOR U40935 ( .A(n41230), .B(n39838), .Z(n35682) );
  AND U40936 ( .A(n34510), .B(n34508), .Z(n41229) );
  XOR U40937 ( .A(n41231), .B(n38255), .Z(n34508) );
  XOR U40938 ( .A(n41232), .B(n40478), .Z(n38255) );
  XNOR U40939 ( .A(n41233), .B(n41234), .Z(n40478) );
  XOR U40940 ( .A(n39320), .B(n36352), .Z(n41234) );
  XOR U40941 ( .A(n41235), .B(n39912), .Z(n36352) );
  ANDN U40942 ( .B(n41236), .A(n41237), .Z(n41235) );
  XNOR U40943 ( .A(n41238), .B(n39903), .Z(n39320) );
  ANDN U40944 ( .B(n41239), .A(n41240), .Z(n41238) );
  XOR U40945 ( .A(n40125), .B(n41241), .Z(n41233) );
  XOR U40946 ( .A(n39101), .B(n38458), .Z(n41241) );
  NOR U40947 ( .A(n41243), .B(n41244), .Z(n41242) );
  XNOR U40948 ( .A(n41245), .B(n39899), .Z(n39101) );
  ANDN U40949 ( .B(n41246), .A(n41247), .Z(n41245) );
  XNOR U40950 ( .A(n41248), .B(n39908), .Z(n40125) );
  IV U40951 ( .A(n41249), .Z(n39908) );
  ANDN U40952 ( .B(n41250), .A(n41251), .Z(n41248) );
  XOR U40953 ( .A(n41252), .B(n35604), .Z(n34510) );
  XNOR U40954 ( .A(n40165), .B(n40378), .Z(n35604) );
  XNOR U40955 ( .A(n41253), .B(n41254), .Z(n40378) );
  XNOR U40956 ( .A(n39415), .B(n38805), .Z(n41254) );
  XNOR U40957 ( .A(n41255), .B(n41256), .Z(n38805) );
  ANDN U40958 ( .B(n41257), .A(n41258), .Z(n41255) );
  XOR U40959 ( .A(n41259), .B(n41260), .Z(n39415) );
  ANDN U40960 ( .B(n41261), .A(n41262), .Z(n41259) );
  XOR U40961 ( .A(n41263), .B(n41264), .Z(n41253) );
  XOR U40962 ( .A(n39789), .B(n39550), .Z(n41264) );
  XNOR U40963 ( .A(n41265), .B(n41266), .Z(n39550) );
  ANDN U40964 ( .B(n41267), .A(n41268), .Z(n41265) );
  XNOR U40965 ( .A(n41269), .B(n41270), .Z(n39789) );
  AND U40966 ( .A(n41271), .B(n41272), .Z(n41269) );
  XOR U40967 ( .A(n41273), .B(n41274), .Z(n40165) );
  XNOR U40968 ( .A(n38078), .B(n36942), .Z(n41274) );
  XNOR U40969 ( .A(n41275), .B(n41276), .Z(n36942) );
  XOR U40970 ( .A(n41279), .B(n41280), .Z(n38078) );
  NOR U40971 ( .A(n41281), .B(n41282), .Z(n41279) );
  XNOR U40972 ( .A(n38433), .B(n41283), .Z(n41273) );
  XOR U40973 ( .A(n37856), .B(n38257), .Z(n41283) );
  XOR U40974 ( .A(n41284), .B(n41285), .Z(n38257) );
  ANDN U40975 ( .B(n41286), .A(n41287), .Z(n41284) );
  XOR U40976 ( .A(n41288), .B(n41289), .Z(n37856) );
  XNOR U40977 ( .A(n41292), .B(n41293), .Z(n38433) );
  ANDN U40978 ( .B(n41294), .A(n41295), .Z(n41292) );
  XOR U40979 ( .A(n41296), .B(n35678), .Z(n32276) );
  XOR U40980 ( .A(n41297), .B(n38863), .Z(n35678) );
  IV U40981 ( .A(n38524), .Z(n38863) );
  XOR U40982 ( .A(n39494), .B(n41091), .Z(n38524) );
  XNOR U40983 ( .A(n41298), .B(n41299), .Z(n41091) );
  XNOR U40984 ( .A(n38570), .B(n36895), .Z(n41299) );
  XNOR U40985 ( .A(n41300), .B(n41301), .Z(n36895) );
  AND U40986 ( .A(n41302), .B(n41303), .Z(n41300) );
  XNOR U40987 ( .A(n41304), .B(n41305), .Z(n38570) );
  ANDN U40988 ( .B(n41306), .A(n41307), .Z(n41304) );
  XNOR U40989 ( .A(n38467), .B(n41308), .Z(n41298) );
  XOR U40990 ( .A(n41309), .B(n41310), .Z(n41308) );
  XNOR U40991 ( .A(n41311), .B(n41312), .Z(n38467) );
  ANDN U40992 ( .B(n41313), .A(n41314), .Z(n41311) );
  XNOR U40993 ( .A(n41315), .B(n41316), .Z(n39494) );
  XNOR U40994 ( .A(n34616), .B(n36389), .Z(n41316) );
  NOR U40995 ( .A(n41319), .B(n41320), .Z(n41317) );
  XNOR U40996 ( .A(n41321), .B(n41322), .Z(n34616) );
  ANDN U40997 ( .B(n41323), .A(n41324), .Z(n41321) );
  XNOR U40998 ( .A(n39053), .B(n41325), .Z(n41315) );
  XOR U40999 ( .A(n41326), .B(n40325), .Z(n41325) );
  XOR U41000 ( .A(n41327), .B(n41328), .Z(n40325) );
  ANDN U41001 ( .B(n41329), .A(n41330), .Z(n41327) );
  XNOR U41002 ( .A(n41331), .B(n41332), .Z(n39053) );
  ANDN U41003 ( .B(n41333), .A(n41334), .Z(n41331) );
  NOR U41004 ( .A(n34518), .B(n34517), .Z(n41296) );
  XNOR U41005 ( .A(n41335), .B(n39530), .Z(n34517) );
  IV U41006 ( .A(n37061), .Z(n39530) );
  XOR U41007 ( .A(n41336), .B(n39620), .Z(n37061) );
  XNOR U41008 ( .A(n41337), .B(n41338), .Z(n39620) );
  XNOR U41009 ( .A(n39607), .B(n39460), .Z(n41338) );
  XNOR U41010 ( .A(n41339), .B(n41340), .Z(n39460) );
  ANDN U41011 ( .B(n41341), .A(n41342), .Z(n41339) );
  XNOR U41012 ( .A(n41343), .B(n41344), .Z(n39607) );
  ANDN U41013 ( .B(n41345), .A(n41346), .Z(n41343) );
  XOR U41014 ( .A(n37833), .B(n41347), .Z(n41337) );
  XOR U41015 ( .A(n40577), .B(n39653), .Z(n41347) );
  XNOR U41016 ( .A(n41348), .B(n41349), .Z(n39653) );
  ANDN U41017 ( .B(n41350), .A(n41351), .Z(n41348) );
  XNOR U41018 ( .A(n41352), .B(n41353), .Z(n40577) );
  ANDN U41019 ( .B(n41354), .A(n41355), .Z(n41352) );
  XNOR U41020 ( .A(n41356), .B(n41357), .Z(n37833) );
  ANDN U41021 ( .B(n41358), .A(n41359), .Z(n41356) );
  XNOR U41022 ( .A(n39603), .B(n40982), .Z(n34518) );
  XNOR U41023 ( .A(n41360), .B(n41361), .Z(n40982) );
  ANDN U41024 ( .B(n41362), .A(n41363), .Z(n41360) );
  XNOR U41025 ( .A(n41364), .B(n35689), .Z(n31241) );
  XOR U41026 ( .A(n41365), .B(n37089), .Z(n35689) );
  IV U41027 ( .A(n36547), .Z(n37089) );
  ANDN U41028 ( .B(n38678), .A(n41366), .Z(n41364) );
  XOR U41029 ( .A(n41367), .B(n41368), .Z(n36173) );
  XOR U41030 ( .A(n29945), .B(n31384), .Z(n41368) );
  XNOR U41031 ( .A(n41369), .B(n36283), .Z(n31384) );
  XNOR U41032 ( .A(n40657), .B(n41370), .Z(n36283) );
  ANDN U41033 ( .B(n36285), .A(n36648), .Z(n41369) );
  XNOR U41034 ( .A(n41371), .B(n39113), .Z(n36648) );
  IV U41035 ( .A(n41372), .Z(n39113) );
  XNOR U41036 ( .A(n39945), .B(n41373), .Z(n36285) );
  IV U41037 ( .A(n37449), .Z(n39945) );
  XOR U41038 ( .A(n41151), .B(n41374), .Z(n37449) );
  XNOR U41039 ( .A(n41375), .B(n41376), .Z(n41151) );
  XNOR U41040 ( .A(n39338), .B(n41377), .Z(n41376) );
  XNOR U41041 ( .A(n41378), .B(n41379), .Z(n39338) );
  ANDN U41042 ( .B(n41380), .A(n41381), .Z(n41378) );
  XOR U41043 ( .A(n37098), .B(n41382), .Z(n41375) );
  XOR U41044 ( .A(n36350), .B(n38888), .Z(n41382) );
  XNOR U41045 ( .A(n41383), .B(n41384), .Z(n38888) );
  NOR U41046 ( .A(n41385), .B(n41386), .Z(n41383) );
  XNOR U41047 ( .A(n41387), .B(n41388), .Z(n36350) );
  ANDN U41048 ( .B(n41389), .A(n41390), .Z(n41387) );
  XNOR U41049 ( .A(n41391), .B(n41392), .Z(n37098) );
  ANDN U41050 ( .B(n41393), .A(n41394), .Z(n41391) );
  XOR U41051 ( .A(n41395), .B(n34246), .Z(n29945) );
  XOR U41052 ( .A(n35944), .B(n41396), .Z(n34246) );
  NOR U41053 ( .A(n36655), .B(n36656), .Z(n41395) );
  XNOR U41054 ( .A(n41399), .B(n39838), .Z(n36656) );
  XOR U41055 ( .A(n41400), .B(n38707), .Z(n39838) );
  XNOR U41056 ( .A(n41401), .B(n41402), .Z(n38707) );
  XOR U41057 ( .A(n39098), .B(n39310), .Z(n41402) );
  XOR U41058 ( .A(n41403), .B(n41404), .Z(n39310) );
  NOR U41059 ( .A(n41405), .B(n41406), .Z(n41403) );
  XNOR U41060 ( .A(n41407), .B(n41408), .Z(n39098) );
  NOR U41061 ( .A(n41409), .B(n41410), .Z(n41407) );
  XNOR U41062 ( .A(n41411), .B(n41412), .Z(n41401) );
  XOR U41063 ( .A(n38825), .B(n41413), .Z(n41412) );
  XNOR U41064 ( .A(n41414), .B(n41415), .Z(n38825) );
  IV U41065 ( .A(n34247), .Z(n36655) );
  XOR U41066 ( .A(n41418), .B(n38318), .Z(n34247) );
  XNOR U41067 ( .A(n33179), .B(n41419), .Z(n41367) );
  XNOR U41068 ( .A(n30681), .B(n31173), .Z(n41419) );
  XNOR U41069 ( .A(n41420), .B(n34234), .Z(n31173) );
  XOR U41070 ( .A(n41421), .B(n38530), .Z(n34234) );
  IV U41071 ( .A(n39821), .Z(n38530) );
  XOR U41072 ( .A(n40629), .B(n40469), .Z(n39821) );
  XNOR U41073 ( .A(n41422), .B(n41423), .Z(n40469) );
  XOR U41074 ( .A(n38676), .B(n37593), .Z(n41423) );
  XNOR U41075 ( .A(n41424), .B(n40778), .Z(n37593) );
  ANDN U41076 ( .B(n41425), .A(n40183), .Z(n41424) );
  XOR U41077 ( .A(n41426), .B(n40785), .Z(n38676) );
  AND U41078 ( .A(n40179), .B(n41427), .Z(n41426) );
  XOR U41079 ( .A(n37678), .B(n41428), .Z(n41422) );
  XNOR U41080 ( .A(n41429), .B(n38591), .Z(n41428) );
  XNOR U41081 ( .A(n41430), .B(n40780), .Z(n38591) );
  ANDN U41082 ( .B(n41431), .A(n40173), .Z(n41430) );
  IV U41083 ( .A(n41432), .Z(n40173) );
  XNOR U41084 ( .A(n41433), .B(n40783), .Z(n37678) );
  XOR U41085 ( .A(n41435), .B(n41436), .Z(n40629) );
  XOR U41086 ( .A(n40480), .B(n41076), .Z(n41436) );
  XOR U41087 ( .A(n41437), .B(n41438), .Z(n41076) );
  NOR U41088 ( .A(n41280), .B(n41439), .Z(n41437) );
  XNOR U41089 ( .A(n41440), .B(n41441), .Z(n40480) );
  XOR U41090 ( .A(n37516), .B(n41443), .Z(n41435) );
  XOR U41091 ( .A(n39852), .B(n39397), .Z(n41443) );
  XNOR U41092 ( .A(n41444), .B(n41445), .Z(n39397) );
  ANDN U41093 ( .B(n41446), .A(n41289), .Z(n41444) );
  XNOR U41094 ( .A(n41447), .B(n41448), .Z(n39852) );
  NOR U41095 ( .A(n41285), .B(n41449), .Z(n41447) );
  XNOR U41096 ( .A(n41450), .B(n41451), .Z(n37516) );
  AND U41097 ( .A(n41452), .B(n41276), .Z(n41450) );
  ANDN U41098 ( .B(n34233), .A(n36653), .Z(n41420) );
  XOR U41099 ( .A(n41453), .B(n35796), .Z(n36653) );
  IV U41100 ( .A(n33931), .Z(n35796) );
  XOR U41101 ( .A(n41454), .B(n41024), .Z(n33931) );
  XNOR U41102 ( .A(n41455), .B(n41456), .Z(n41024) );
  XNOR U41103 ( .A(n34632), .B(n38822), .Z(n41456) );
  XOR U41104 ( .A(n41457), .B(n41458), .Z(n38822) );
  NOR U41105 ( .A(n41459), .B(n41460), .Z(n41457) );
  XOR U41106 ( .A(n41461), .B(n41462), .Z(n34632) );
  XOR U41107 ( .A(n36443), .B(n41465), .Z(n41455) );
  XOR U41108 ( .A(n39972), .B(n41466), .Z(n41465) );
  XNOR U41109 ( .A(n41467), .B(n41468), .Z(n39972) );
  NOR U41110 ( .A(n41469), .B(n41470), .Z(n41467) );
  XOR U41111 ( .A(n41471), .B(n41472), .Z(n36443) );
  NOR U41112 ( .A(n41473), .B(n41474), .Z(n41471) );
  XNOR U41113 ( .A(n40766), .B(n37707), .Z(n34233) );
  XNOR U41114 ( .A(n41475), .B(n41476), .Z(n39362) );
  XOR U41115 ( .A(n38128), .B(n40660), .Z(n41476) );
  XNOR U41116 ( .A(n41477), .B(n41478), .Z(n40660) );
  NOR U41117 ( .A(n41479), .B(n41480), .Z(n41477) );
  ANDN U41118 ( .B(n40774), .A(n40772), .Z(n41481) );
  XOR U41119 ( .A(n37840), .B(n41483), .Z(n41475) );
  XOR U41120 ( .A(n38282), .B(n38795), .Z(n41483) );
  XNOR U41121 ( .A(n41484), .B(n41485), .Z(n38795) );
  NOR U41122 ( .A(n40763), .B(n40762), .Z(n41484) );
  XNOR U41123 ( .A(n41486), .B(n41487), .Z(n38282) );
  NOR U41124 ( .A(n40768), .B(n40769), .Z(n41486) );
  NOR U41125 ( .A(n40758), .B(n40759), .Z(n41488) );
  ANDN U41126 ( .B(n41480), .A(n41492), .Z(n41491) );
  XNOR U41127 ( .A(n41493), .B(n34239), .Z(n30681) );
  XOR U41128 ( .A(n41494), .B(n39312), .Z(n34239) );
  ANDN U41129 ( .B(n34238), .A(n36646), .Z(n41493) );
  XOR U41130 ( .A(n40251), .B(n36308), .Z(n36646) );
  XNOR U41131 ( .A(n41495), .B(n41496), .Z(n40251) );
  XOR U41132 ( .A(n41499), .B(n38411), .Z(n34238) );
  IV U41133 ( .A(n37928), .Z(n38411) );
  XNOR U41134 ( .A(n41500), .B(n41501), .Z(n41088) );
  XNOR U41135 ( .A(n37703), .B(n40541), .Z(n41501) );
  XNOR U41136 ( .A(n41502), .B(n40547), .Z(n40541) );
  ANDN U41137 ( .B(n40548), .A(n41503), .Z(n41502) );
  XNOR U41138 ( .A(n41504), .B(n40552), .Z(n37703) );
  ANDN U41139 ( .B(n41505), .A(n40551), .Z(n41504) );
  XOR U41140 ( .A(n36997), .B(n41506), .Z(n41500) );
  XOR U41141 ( .A(n35629), .B(n36312), .Z(n41506) );
  XNOR U41142 ( .A(n41507), .B(n40564), .Z(n36312) );
  ANDN U41143 ( .B(n40565), .A(n41508), .Z(n41507) );
  XNOR U41144 ( .A(n41509), .B(n40556), .Z(n35629) );
  ANDN U41145 ( .B(n40557), .A(n41510), .Z(n41509) );
  XNOR U41146 ( .A(n41511), .B(n40560), .Z(n36997) );
  AND U41147 ( .A(n41512), .B(n40561), .Z(n41511) );
  XOR U41148 ( .A(n41514), .B(n34242), .Z(n33179) );
  XNOR U41149 ( .A(n41515), .B(n39055), .Z(n34242) );
  XNOR U41150 ( .A(n41516), .B(n41517), .Z(n39055) );
  ANDN U41151 ( .B(n36651), .A(n34243), .Z(n41514) );
  XOR U41152 ( .A(n41518), .B(n39616), .Z(n34243) );
  XOR U41153 ( .A(n39758), .B(n41519), .Z(n39616) );
  XOR U41154 ( .A(n41520), .B(n41521), .Z(n39758) );
  XOR U41155 ( .A(n39995), .B(n37325), .Z(n41521) );
  XOR U41156 ( .A(n41522), .B(n41523), .Z(n37325) );
  ANDN U41157 ( .B(n41524), .A(n41525), .Z(n41522) );
  XNOR U41158 ( .A(n41526), .B(n41527), .Z(n39995) );
  ANDN U41159 ( .B(n41528), .A(n41529), .Z(n41526) );
  XNOR U41160 ( .A(n40614), .B(n41530), .Z(n41520) );
  XOR U41161 ( .A(n40042), .B(n38470), .Z(n41530) );
  XOR U41162 ( .A(n41531), .B(n41532), .Z(n38470) );
  NOR U41163 ( .A(n41533), .B(n41534), .Z(n41531) );
  XNOR U41164 ( .A(n41535), .B(n41536), .Z(n40042) );
  ANDN U41165 ( .B(n41537), .A(n41538), .Z(n41535) );
  XNOR U41166 ( .A(n41539), .B(n41540), .Z(n40614) );
  ANDN U41167 ( .B(n41541), .A(n41542), .Z(n41539) );
  XNOR U41168 ( .A(n41543), .B(n41544), .Z(n40157) );
  NOR U41169 ( .A(n40314), .B(n41545), .Z(n41543) );
  XNOR U41170 ( .A(n41546), .B(n35688), .Z(n34506) );
  IV U41171 ( .A(n41366), .Z(n35688) );
  XOR U41172 ( .A(n35926), .B(n40868), .Z(n41366) );
  XNOR U41173 ( .A(n41547), .B(n40940), .Z(n40868) );
  ANDN U41174 ( .B(n41548), .A(n41549), .Z(n41547) );
  NOR U41175 ( .A(n37378), .B(n38678), .Z(n41546) );
  XOR U41176 ( .A(n41550), .B(n38544), .Z(n38678) );
  XOR U41177 ( .A(n39235), .B(n41551), .Z(n38544) );
  XOR U41178 ( .A(n41552), .B(n41553), .Z(n39235) );
  XOR U41179 ( .A(n38294), .B(n39583), .Z(n41553) );
  XOR U41180 ( .A(n41554), .B(n40502), .Z(n39583) );
  ANDN U41181 ( .B(n41555), .A(n41556), .Z(n41554) );
  NOR U41182 ( .A(n41558), .B(n41559), .Z(n41557) );
  XOR U41183 ( .A(n41560), .B(n41561), .Z(n41552) );
  XOR U41184 ( .A(n39483), .B(n39643), .Z(n41561) );
  XNOR U41185 ( .A(n41562), .B(n40498), .Z(n39643) );
  NOR U41186 ( .A(n41563), .B(n41564), .Z(n41562) );
  XNOR U41187 ( .A(n41565), .B(n40505), .Z(n39483) );
  NOR U41188 ( .A(n41566), .B(n41567), .Z(n41565) );
  XOR U41189 ( .A(n41568), .B(n39692), .Z(n37378) );
  NOR U41190 ( .A(n31272), .B(n28055), .Z(n41153) );
  XOR U41191 ( .A(n30865), .B(n33893), .Z(n28055) );
  XOR U41192 ( .A(n41571), .B(n40916), .Z(n33893) );
  AND U41193 ( .A(n34986), .B(n40027), .Z(n41571) );
  XOR U41194 ( .A(n41572), .B(n40005), .Z(n34986) );
  XOR U41195 ( .A(n33174), .B(n37544), .Z(n30865) );
  XOR U41196 ( .A(n41573), .B(n41574), .Z(n37544) );
  XOR U41197 ( .A(n29303), .B(n34041), .Z(n41574) );
  XNOR U41198 ( .A(n41575), .B(n34047), .Z(n34041) );
  XOR U41199 ( .A(n41576), .B(n38684), .Z(n34047) );
  NOR U41200 ( .A(n37546), .B(n37547), .Z(n41575) );
  XNOR U41201 ( .A(n39664), .B(n41577), .Z(n37547) );
  IV U41202 ( .A(n38961), .Z(n39664) );
  XOR U41203 ( .A(n40606), .B(n37698), .Z(n37546) );
  IV U41204 ( .A(n37875), .Z(n37698) );
  XNOR U41205 ( .A(n41580), .B(n40403), .Z(n37875) );
  XNOR U41206 ( .A(n41581), .B(n41582), .Z(n40403) );
  XOR U41207 ( .A(n38744), .B(n39154), .Z(n41582) );
  XOR U41208 ( .A(n41583), .B(n39208), .Z(n39154) );
  NOR U41209 ( .A(n39207), .B(n40612), .Z(n41583) );
  XOR U41210 ( .A(n41584), .B(n41585), .Z(n39207) );
  XOR U41211 ( .A(n41586), .B(n39197), .Z(n38744) );
  NOR U41212 ( .A(n39196), .B(n40609), .Z(n41586) );
  XOR U41213 ( .A(n41587), .B(n41588), .Z(n39196) );
  XOR U41214 ( .A(n37490), .B(n41589), .Z(n41581) );
  XOR U41215 ( .A(n36945), .B(n39035), .Z(n41589) );
  XNOR U41216 ( .A(n41590), .B(n39201), .Z(n39035) );
  NOR U41217 ( .A(n39200), .B(n41591), .Z(n41590) );
  XOR U41218 ( .A(n41592), .B(n40636), .Z(n36945) );
  NOR U41219 ( .A(n40602), .B(n40603), .Z(n41592) );
  XOR U41220 ( .A(n41593), .B(n41594), .Z(n40602) );
  XOR U41221 ( .A(n41595), .B(n41596), .Z(n37490) );
  ANDN U41222 ( .B(n40598), .A(n40599), .Z(n41595) );
  XNOR U41223 ( .A(n41597), .B(n39200), .Z(n40606) );
  XNOR U41224 ( .A(n41598), .B(n41599), .Z(n39200) );
  AND U41225 ( .A(n41591), .B(n41600), .Z(n41597) );
  XOR U41226 ( .A(n41601), .B(n34058), .Z(n29303) );
  IV U41227 ( .A(n36299), .Z(n34058) );
  XOR U41228 ( .A(n38466), .B(n41309), .Z(n36299) );
  XOR U41229 ( .A(n41602), .B(n41603), .Z(n41309) );
  AND U41230 ( .A(n41604), .B(n41605), .Z(n41602) );
  IV U41231 ( .A(n36894), .Z(n38466) );
  NOR U41232 ( .A(n34057), .B(n35117), .Z(n41601) );
  XOR U41233 ( .A(n40936), .B(n41606), .Z(n35117) );
  XNOR U41234 ( .A(n41607), .B(n41608), .Z(n40936) );
  ANDN U41235 ( .B(n41609), .A(n41610), .Z(n41607) );
  XOR U41236 ( .A(n37209), .B(n41611), .Z(n34057) );
  XOR U41237 ( .A(n30196), .B(n41612), .Z(n41573) );
  XOR U41238 ( .A(n32942), .B(n31655), .Z(n41612) );
  XNOR U41239 ( .A(n41613), .B(n34061), .Z(n31655) );
  XOR U41240 ( .A(n39051), .B(n39571), .Z(n34061) );
  XOR U41241 ( .A(n41614), .B(n41615), .Z(n39571) );
  ANDN U41242 ( .B(n41616), .A(n41617), .Z(n41614) );
  IV U41243 ( .A(n39171), .Z(n39051) );
  ANDN U41244 ( .B(n34062), .A(n36457), .Z(n41613) );
  XOR U41245 ( .A(n36442), .B(n41466), .Z(n36457) );
  XOR U41246 ( .A(n41618), .B(n41619), .Z(n41466) );
  ANDN U41247 ( .B(n41620), .A(n41621), .Z(n41618) );
  IV U41248 ( .A(n34631), .Z(n36442) );
  XOR U41249 ( .A(n40192), .B(n41159), .Z(n34631) );
  XNOR U41250 ( .A(n41622), .B(n41623), .Z(n41159) );
  XOR U41251 ( .A(n41624), .B(n38160), .Z(n41623) );
  XOR U41252 ( .A(n41625), .B(n41626), .Z(n38160) );
  ANDN U41253 ( .B(n41459), .A(n41458), .Z(n41625) );
  IV U41254 ( .A(n41627), .Z(n41458) );
  XOR U41255 ( .A(n37697), .B(n41628), .Z(n41622) );
  XOR U41256 ( .A(n37692), .B(n37196), .Z(n41628) );
  XNOR U41257 ( .A(n41629), .B(n41630), .Z(n37196) );
  ANDN U41258 ( .B(n41619), .A(n41620), .Z(n41629) );
  XNOR U41259 ( .A(n41631), .B(n41632), .Z(n37692) );
  ANDN U41260 ( .B(n41469), .A(n41468), .Z(n41631) );
  XNOR U41261 ( .A(n41633), .B(n41634), .Z(n37697) );
  ANDN U41262 ( .B(n41473), .A(n41472), .Z(n41633) );
  XOR U41263 ( .A(n41635), .B(n41636), .Z(n40192) );
  XOR U41264 ( .A(n38511), .B(n36358), .Z(n41636) );
  XOR U41265 ( .A(n41637), .B(n41638), .Z(n36358) );
  ANDN U41266 ( .B(n41033), .A(n40884), .Z(n41637) );
  XNOR U41267 ( .A(n41639), .B(n41640), .Z(n40884) );
  XNOR U41268 ( .A(n41641), .B(n41642), .Z(n38511) );
  ANDN U41269 ( .B(n40890), .A(n41030), .Z(n41641) );
  XOR U41270 ( .A(n41643), .B(n41644), .Z(n40890) );
  XOR U41271 ( .A(n38764), .B(n41645), .Z(n41635) );
  XNOR U41272 ( .A(n39178), .B(n37596), .Z(n41645) );
  XOR U41273 ( .A(n41646), .B(n41647), .Z(n37596) );
  ANDN U41274 ( .B(n41028), .A(n40908), .Z(n41646) );
  XOR U41275 ( .A(n41648), .B(n41649), .Z(n40908) );
  XNOR U41276 ( .A(n41650), .B(n41651), .Z(n39178) );
  AND U41277 ( .A(n40880), .B(n41037), .Z(n41650) );
  XOR U41278 ( .A(n41652), .B(n41653), .Z(n40880) );
  XNOR U41279 ( .A(n41654), .B(n41655), .Z(n38764) );
  ANDN U41280 ( .B(n40894), .A(n41035), .Z(n41654) );
  XNOR U41281 ( .A(n41656), .B(n41657), .Z(n40894) );
  XOR U41282 ( .A(n41658), .B(n38836), .Z(n34062) );
  IV U41283 ( .A(n35952), .Z(n38836) );
  XNOR U41284 ( .A(n41659), .B(n41660), .Z(n35952) );
  XNOR U41285 ( .A(n41661), .B(n36288), .Z(n32942) );
  XOR U41286 ( .A(n41662), .B(n37625), .Z(n36288) );
  XNOR U41287 ( .A(n39798), .B(n41663), .Z(n37625) );
  XOR U41288 ( .A(n41664), .B(n41665), .Z(n39798) );
  XNOR U41289 ( .A(n41086), .B(n39826), .Z(n41665) );
  XOR U41290 ( .A(n41666), .B(n40293), .Z(n39826) );
  AND U41291 ( .A(n41667), .B(n41668), .Z(n41666) );
  XOR U41292 ( .A(n41669), .B(n41670), .Z(n41086) );
  AND U41293 ( .A(n41671), .B(n41672), .Z(n41669) );
  XOR U41294 ( .A(n39810), .B(n41673), .Z(n41664) );
  XOR U41295 ( .A(n39066), .B(n37143), .Z(n41673) );
  XNOR U41296 ( .A(n41674), .B(n40282), .Z(n37143) );
  ANDN U41297 ( .B(n41675), .A(n41676), .Z(n41674) );
  XNOR U41298 ( .A(n41677), .B(n40287), .Z(n39066) );
  AND U41299 ( .A(n41678), .B(n41679), .Z(n41677) );
  XNOR U41300 ( .A(n41680), .B(n40297), .Z(n39810) );
  AND U41301 ( .A(n41681), .B(n41682), .Z(n41680) );
  XNOR U41302 ( .A(n41683), .B(n38440), .Z(n35121) );
  IV U41303 ( .A(n38820), .Z(n38440) );
  XOR U41304 ( .A(n41684), .B(n41685), .Z(n38820) );
  XOR U41305 ( .A(n41686), .B(n34638), .Z(n35123) );
  XOR U41306 ( .A(n41687), .B(n34052), .Z(n30196) );
  XNOR U41307 ( .A(n41688), .B(n38491), .Z(n34052) );
  IV U41308 ( .A(n37515), .Z(n38491) );
  XOR U41309 ( .A(n41689), .B(n39651), .Z(n37515) );
  XNOR U41310 ( .A(n41690), .B(n41691), .Z(n39651) );
  XOR U41311 ( .A(n38445), .B(n40058), .Z(n41691) );
  XOR U41312 ( .A(n41692), .B(n41693), .Z(n40058) );
  ANDN U41313 ( .B(n41694), .A(n41695), .Z(n41692) );
  XNOR U41314 ( .A(n41696), .B(n41697), .Z(n38445) );
  AND U41315 ( .A(n41698), .B(n41699), .Z(n41696) );
  XOR U41316 ( .A(n39929), .B(n41700), .Z(n41690) );
  XOR U41317 ( .A(n37639), .B(n41701), .Z(n41700) );
  XOR U41318 ( .A(n41702), .B(n41703), .Z(n37639) );
  AND U41319 ( .A(n41704), .B(n41705), .Z(n41702) );
  XNOR U41320 ( .A(n41706), .B(n41707), .Z(n39929) );
  NOR U41321 ( .A(n41708), .B(n41709), .Z(n41706) );
  XOR U41322 ( .A(n41710), .B(n35311), .Z(n34051) );
  XNOR U41323 ( .A(n41711), .B(n37000), .Z(n35126) );
  XOR U41324 ( .A(n41712), .B(n41713), .Z(n33174) );
  XNOR U41325 ( .A(n32255), .B(n28886), .Z(n41713) );
  XNOR U41326 ( .A(n41714), .B(n37895), .Z(n28886) );
  XOR U41327 ( .A(n41715), .B(n37331), .Z(n37895) );
  NOR U41328 ( .A(n33889), .B(n33891), .Z(n41714) );
  XNOR U41329 ( .A(n41718), .B(n38260), .Z(n33891) );
  XOR U41330 ( .A(n38181), .B(n41719), .Z(n33889) );
  XNOR U41331 ( .A(n41720), .B(n34988), .Z(n32255) );
  IV U41332 ( .A(n40915), .Z(n34988) );
  XOR U41333 ( .A(n37677), .B(n41429), .Z(n40915) );
  XNOR U41334 ( .A(n41721), .B(n41722), .Z(n41429) );
  ANDN U41335 ( .B(n41723), .A(n41724), .Z(n41721) );
  XOR U41336 ( .A(n41725), .B(n41078), .Z(n37677) );
  XNOR U41337 ( .A(n41726), .B(n41727), .Z(n41078) );
  XNOR U41338 ( .A(n36891), .B(n40754), .Z(n41727) );
  XOR U41339 ( .A(n41728), .B(n40181), .Z(n40754) );
  XOR U41340 ( .A(n41729), .B(n41657), .Z(n40181) );
  ANDN U41341 ( .B(n40785), .A(n41427), .Z(n41728) );
  XNOR U41342 ( .A(n41730), .B(n41731), .Z(n40785) );
  XOR U41343 ( .A(n41732), .B(n40174), .Z(n36891) );
  XOR U41344 ( .A(n41733), .B(n41734), .Z(n40174) );
  ANDN U41345 ( .B(n40780), .A(n41431), .Z(n41732) );
  XNOR U41346 ( .A(n41735), .B(n41736), .Z(n40780) );
  XOR U41347 ( .A(n36540), .B(n41737), .Z(n41726) );
  XOR U41348 ( .A(n39486), .B(n37340), .Z(n41737) );
  XNOR U41349 ( .A(n41738), .B(n40184), .Z(n37340) );
  XNOR U41350 ( .A(n41739), .B(n41740), .Z(n40184) );
  ANDN U41351 ( .B(n40778), .A(n41425), .Z(n41738) );
  XNOR U41352 ( .A(n41741), .B(n41742), .Z(n40778) );
  XNOR U41353 ( .A(n41743), .B(n40170), .Z(n39486) );
  XOR U41354 ( .A(n41744), .B(n41745), .Z(n40170) );
  ANDN U41355 ( .B(n40783), .A(n41434), .Z(n41743) );
  XNOR U41356 ( .A(n41746), .B(n41747), .Z(n40783) );
  XNOR U41357 ( .A(n41748), .B(n40788), .Z(n36540) );
  ANDN U41358 ( .B(n41724), .A(n41722), .Z(n41748) );
  IV U41359 ( .A(n40789), .Z(n41722) );
  XOR U41360 ( .A(n41749), .B(n41750), .Z(n40789) );
  ANDN U41361 ( .B(n40916), .A(n40027), .Z(n41720) );
  XOR U41362 ( .A(n41751), .B(n37690), .Z(n40027) );
  IV U41363 ( .A(n39067), .Z(n37690) );
  XNOR U41364 ( .A(n41752), .B(n41753), .Z(n39067) );
  XOR U41365 ( .A(n41754), .B(n37344), .Z(n40916) );
  IV U41366 ( .A(n38507), .Z(n37344) );
  XOR U41367 ( .A(n31165), .B(n41755), .Z(n41712) );
  XOR U41368 ( .A(n29096), .B(n31135), .Z(n41755) );
  XNOR U41369 ( .A(n41756), .B(n40039), .Z(n31135) );
  XOR U41370 ( .A(n41757), .B(n36202), .Z(n40039) );
  XNOR U41371 ( .A(n41758), .B(n37015), .Z(n33896) );
  IV U41372 ( .A(n38285), .Z(n37015) );
  XNOR U41373 ( .A(n40441), .B(n39746), .Z(n38285) );
  XOR U41374 ( .A(n41759), .B(n41760), .Z(n39746) );
  XOR U41375 ( .A(n35597), .B(n37538), .Z(n41760) );
  XOR U41376 ( .A(n41761), .B(n41762), .Z(n37538) );
  ANDN U41377 ( .B(n41763), .A(n41764), .Z(n41761) );
  XNOR U41378 ( .A(n41765), .B(n41766), .Z(n35597) );
  ANDN U41379 ( .B(n41767), .A(n41768), .Z(n41765) );
  XOR U41380 ( .A(n37945), .B(n41769), .Z(n41759) );
  XOR U41381 ( .A(n38334), .B(n39561), .Z(n41769) );
  XNOR U41382 ( .A(n41770), .B(n41771), .Z(n39561) );
  NOR U41383 ( .A(n41772), .B(n41773), .Z(n41770) );
  XNOR U41384 ( .A(n41774), .B(n41775), .Z(n38334) );
  ANDN U41385 ( .B(n41776), .A(n41777), .Z(n41774) );
  XNOR U41386 ( .A(n41778), .B(n41779), .Z(n37945) );
  XOR U41387 ( .A(n41782), .B(n41783), .Z(n40441) );
  XNOR U41388 ( .A(n38447), .B(n37458), .Z(n41783) );
  XOR U41389 ( .A(n41784), .B(n40121), .Z(n37458) );
  NOR U41390 ( .A(n40122), .B(n41785), .Z(n41784) );
  XOR U41391 ( .A(n41786), .B(n39567), .Z(n38447) );
  XNOR U41392 ( .A(n38137), .B(n41788), .Z(n41782) );
  XOR U41393 ( .A(n37175), .B(n37455), .Z(n41788) );
  XOR U41394 ( .A(n41789), .B(n41790), .Z(n37455) );
  NOR U41395 ( .A(n41791), .B(n41792), .Z(n41789) );
  XNOR U41396 ( .A(n41793), .B(n41617), .Z(n37175) );
  NOR U41397 ( .A(n41794), .B(n41616), .Z(n41793) );
  XNOR U41398 ( .A(n41795), .B(n39575), .Z(n38137) );
  ANDN U41399 ( .B(n39574), .A(n41796), .Z(n41795) );
  XOR U41400 ( .A(n37720), .B(n41797), .Z(n33895) );
  XNOR U41401 ( .A(n41798), .B(n34994), .Z(n29096) );
  XOR U41402 ( .A(n38944), .B(n41799), .Z(n34994) );
  ANDN U41403 ( .B(n33901), .A(n40921), .Z(n41798) );
  XOR U41404 ( .A(n37912), .B(n41800), .Z(n40921) );
  IV U41405 ( .A(n41801), .Z(n37912) );
  XOR U41406 ( .A(n37503), .B(n41802), .Z(n33901) );
  IV U41407 ( .A(n39413), .Z(n37503) );
  XNOR U41408 ( .A(n39635), .B(n38981), .Z(n39413) );
  XOR U41409 ( .A(n41803), .B(n41804), .Z(n38981) );
  XNOR U41410 ( .A(n41805), .B(n38852), .Z(n41804) );
  XOR U41411 ( .A(n41806), .B(n41807), .Z(n38852) );
  NOR U41412 ( .A(n40747), .B(n41808), .Z(n41806) );
  XOR U41413 ( .A(n38879), .B(n41809), .Z(n41803) );
  XOR U41414 ( .A(n39922), .B(n39739), .Z(n41809) );
  XNOR U41415 ( .A(n41810), .B(n41811), .Z(n39739) );
  NOR U41416 ( .A(n40751), .B(n41812), .Z(n41810) );
  XNOR U41417 ( .A(n41813), .B(n41814), .Z(n39922) );
  NOR U41418 ( .A(n40743), .B(n41815), .Z(n41813) );
  XNOR U41419 ( .A(n41816), .B(n41817), .Z(n38879) );
  NOR U41420 ( .A(n41818), .B(n40738), .Z(n41816) );
  XOR U41421 ( .A(n41819), .B(n41820), .Z(n39635) );
  XNOR U41422 ( .A(n38485), .B(n38784), .Z(n41820) );
  XNOR U41423 ( .A(n41821), .B(n41822), .Z(n38784) );
  NOR U41424 ( .A(n41823), .B(n41824), .Z(n41821) );
  XNOR U41425 ( .A(n41825), .B(n41826), .Z(n38485) );
  ANDN U41426 ( .B(n41827), .A(n41828), .Z(n41825) );
  XOR U41427 ( .A(n39437), .B(n41829), .Z(n41819) );
  XOR U41428 ( .A(n37947), .B(n41830), .Z(n41829) );
  XNOR U41429 ( .A(n41831), .B(n41832), .Z(n37947) );
  NOR U41430 ( .A(n41833), .B(n41834), .Z(n41831) );
  XNOR U41431 ( .A(n41835), .B(n41836), .Z(n39437) );
  NOR U41432 ( .A(n41837), .B(n41838), .Z(n41835) );
  XNOR U41433 ( .A(n41839), .B(n34984), .Z(n31165) );
  XOR U41434 ( .A(n41840), .B(n39267), .Z(n34984) );
  IV U41435 ( .A(n39406), .Z(n39267) );
  NOR U41436 ( .A(n35437), .B(n35438), .Z(n41839) );
  XNOR U41437 ( .A(n40657), .B(n41841), .Z(n35438) );
  XOR U41438 ( .A(n41842), .B(n37018), .Z(n35437) );
  XNOR U41439 ( .A(n41843), .B(n41844), .Z(n39636) );
  XOR U41440 ( .A(n41845), .B(n41846), .Z(n41844) );
  XOR U41441 ( .A(n35300), .B(n41847), .Z(n41843) );
  XOR U41442 ( .A(n37892), .B(n39465), .Z(n41847) );
  XOR U41443 ( .A(n41848), .B(n41849), .Z(n39465) );
  ANDN U41444 ( .B(n41850), .A(n41851), .Z(n41848) );
  XOR U41445 ( .A(n41852), .B(n41853), .Z(n37892) );
  ANDN U41446 ( .B(n41854), .A(n41855), .Z(n41852) );
  XNOR U41447 ( .A(n41856), .B(n41857), .Z(n35300) );
  ANDN U41448 ( .B(n41858), .A(n41859), .Z(n41856) );
  XNOR U41449 ( .A(n29060), .B(n37352), .Z(n31272) );
  XNOR U41450 ( .A(n41861), .B(n37637), .Z(n37352) );
  ANDN U41451 ( .B(n34941), .A(n34943), .Z(n41861) );
  XOR U41452 ( .A(n41862), .B(n39312), .Z(n34943) );
  XNOR U41453 ( .A(n38868), .B(n33464), .Z(n29060) );
  XNOR U41454 ( .A(n41863), .B(n41864), .Z(n33464) );
  XOR U41455 ( .A(n28832), .B(n29522), .Z(n41864) );
  XOR U41456 ( .A(n41865), .B(n37659), .Z(n29522) );
  XNOR U41457 ( .A(n38804), .B(n41263), .Z(n37659) );
  XNOR U41458 ( .A(n41866), .B(n41867), .Z(n41263) );
  XOR U41459 ( .A(n41870), .B(n38434), .Z(n38804) );
  XNOR U41460 ( .A(n41871), .B(n41872), .Z(n38434) );
  XNOR U41461 ( .A(n41421), .B(n40396), .Z(n41872) );
  XOR U41462 ( .A(n41873), .B(n41449), .Z(n40396) );
  XNOR U41463 ( .A(n41874), .B(n41875), .Z(n41285) );
  XNOR U41464 ( .A(n41876), .B(n41442), .Z(n41421) );
  ANDN U41465 ( .B(n41295), .A(n41293), .Z(n41876) );
  XOR U41466 ( .A(n41877), .B(n41878), .Z(n41293) );
  IV U41467 ( .A(n41879), .Z(n41295) );
  XOR U41468 ( .A(n38529), .B(n41880), .Z(n41871) );
  XNOR U41469 ( .A(n38978), .B(n39820), .Z(n41880) );
  XNOR U41470 ( .A(n41881), .B(n41452), .Z(n39820) );
  NOR U41471 ( .A(n41277), .B(n41276), .Z(n41881) );
  XNOR U41472 ( .A(n41882), .B(n41883), .Z(n41276) );
  XOR U41473 ( .A(n41884), .B(n41446), .Z(n38978) );
  ANDN U41474 ( .B(n41289), .A(n41291), .Z(n41884) );
  XOR U41475 ( .A(n41885), .B(n40853), .Z(n41289) );
  XOR U41476 ( .A(n41886), .B(n41439), .Z(n38529) );
  ANDN U41477 ( .B(n41280), .A(n41887), .Z(n41886) );
  XOR U41478 ( .A(n41888), .B(n41889), .Z(n41280) );
  ANDN U41479 ( .B(n36689), .A(n34925), .Z(n41865) );
  XOR U41480 ( .A(n41890), .B(n41372), .Z(n34925) );
  XNOR U41481 ( .A(n41752), .B(n41891), .Z(n41372) );
  XOR U41482 ( .A(n41892), .B(n41893), .Z(n41752) );
  XNOR U41483 ( .A(n39640), .B(n39541), .Z(n41893) );
  XNOR U41484 ( .A(n41894), .B(n41895), .Z(n39541) );
  AND U41485 ( .A(n41896), .B(n41897), .Z(n41894) );
  XNOR U41486 ( .A(n41898), .B(n41899), .Z(n39640) );
  AND U41487 ( .A(n41900), .B(n41901), .Z(n41898) );
  XNOR U41488 ( .A(n38079), .B(n41902), .Z(n41892) );
  XOR U41489 ( .A(n39256), .B(n39582), .Z(n41902) );
  XNOR U41490 ( .A(n41903), .B(n41904), .Z(n39582) );
  AND U41491 ( .A(n41905), .B(n41906), .Z(n41903) );
  XOR U41492 ( .A(n41907), .B(n41908), .Z(n39256) );
  XOR U41493 ( .A(n41911), .B(n41912), .Z(n38079) );
  ANDN U41494 ( .B(n41913), .A(n41914), .Z(n41911) );
  XOR U41495 ( .A(n41915), .B(n38374), .Z(n36689) );
  XNOR U41496 ( .A(n41916), .B(n37661), .Z(n28832) );
  XOR U41497 ( .A(n41917), .B(n39976), .Z(n37661) );
  XNOR U41498 ( .A(n39699), .B(n41918), .Z(n39976) );
  XOR U41499 ( .A(n41919), .B(n41920), .Z(n39699) );
  XOR U41500 ( .A(n41921), .B(n35594), .Z(n41920) );
  XNOR U41501 ( .A(n41922), .B(n41923), .Z(n35594) );
  NOR U41502 ( .A(n41924), .B(n41925), .Z(n41922) );
  XNOR U41503 ( .A(n36790), .B(n41926), .Z(n41919) );
  XOR U41504 ( .A(n38310), .B(n37870), .Z(n41926) );
  XNOR U41505 ( .A(n41927), .B(n41928), .Z(n37870) );
  AND U41506 ( .A(n41929), .B(n41930), .Z(n41927) );
  XNOR U41507 ( .A(n41931), .B(n41932), .Z(n38310) );
  ANDN U41508 ( .B(n41933), .A(n41934), .Z(n41931) );
  XOR U41509 ( .A(n41935), .B(n41936), .Z(n36790) );
  ANDN U41510 ( .B(n41937), .A(n41938), .Z(n41935) );
  ANDN U41511 ( .B(n36681), .A(n34912), .Z(n41916) );
  IV U41512 ( .A(n36682), .Z(n34912) );
  XNOR U41513 ( .A(n41939), .B(n35093), .Z(n36682) );
  XNOR U41514 ( .A(n39171), .B(n39564), .Z(n36681) );
  XOR U41515 ( .A(n41940), .B(n41941), .Z(n39564) );
  ANDN U41516 ( .B(n41790), .A(n41942), .Z(n41940) );
  XOR U41517 ( .A(n41943), .B(n41860), .Z(n39171) );
  XOR U41518 ( .A(n41944), .B(n41945), .Z(n41860) );
  XOR U41519 ( .A(n38601), .B(n41946), .Z(n41945) );
  XNOR U41520 ( .A(n41947), .B(n41948), .Z(n38601) );
  NOR U41521 ( .A(n41949), .B(n41950), .Z(n41947) );
  XOR U41522 ( .A(n36934), .B(n41951), .Z(n41944) );
  XOR U41523 ( .A(n38133), .B(n41952), .Z(n41951) );
  XNOR U41524 ( .A(n41953), .B(n41047), .Z(n38133) );
  ANDN U41525 ( .B(n41954), .A(n41955), .Z(n41953) );
  XNOR U41526 ( .A(n41956), .B(n41060), .Z(n36934) );
  ANDN U41527 ( .B(n41957), .A(n41958), .Z(n41956) );
  XNOR U41528 ( .A(n33356), .B(n41959), .Z(n41863) );
  XOR U41529 ( .A(n35690), .B(n32623), .Z(n41959) );
  XNOR U41530 ( .A(n41960), .B(n39438), .Z(n32623) );
  IV U41531 ( .A(n37656), .Z(n39438) );
  XOR U41532 ( .A(n41961), .B(n39312), .Z(n37656) );
  XNOR U41533 ( .A(n41962), .B(n41963), .Z(n40348) );
  XOR U41534 ( .A(n38393), .B(n37070), .Z(n41963) );
  XNOR U41535 ( .A(n41964), .B(n41196), .Z(n37070) );
  AND U41536 ( .A(n41197), .B(n41965), .Z(n41964) );
  XNOR U41537 ( .A(n41966), .B(n41203), .Z(n38393) );
  ANDN U41538 ( .B(n41202), .A(n41967), .Z(n41966) );
  XNOR U41539 ( .A(n39745), .B(n41968), .Z(n41962) );
  XOR U41540 ( .A(n38631), .B(n35783), .Z(n41968) );
  XNOR U41541 ( .A(n41969), .B(n41206), .Z(n35783) );
  ANDN U41542 ( .B(n41207), .A(n41970), .Z(n41969) );
  XNOR U41543 ( .A(n41971), .B(n41972), .Z(n38631) );
  ANDN U41544 ( .B(n41973), .A(n41974), .Z(n41971) );
  XOR U41545 ( .A(n41975), .B(n41976), .Z(n39745) );
  ANDN U41546 ( .B(n41977), .A(n41192), .Z(n41975) );
  XOR U41547 ( .A(n41978), .B(n41979), .Z(n39223) );
  XNOR U41548 ( .A(n39242), .B(n41187), .Z(n41979) );
  XNOR U41549 ( .A(n41980), .B(n41981), .Z(n41187) );
  ANDN U41550 ( .B(n41982), .A(n41983), .Z(n41980) );
  ANDN U41551 ( .B(n41214), .A(n41985), .Z(n41984) );
  XNOR U41552 ( .A(n38548), .B(n41986), .Z(n41978) );
  XNOR U41553 ( .A(n39115), .B(n38247), .Z(n41986) );
  XNOR U41554 ( .A(n41987), .B(n41218), .Z(n38247) );
  ANDN U41555 ( .B(n41219), .A(n41988), .Z(n41987) );
  XNOR U41556 ( .A(n41989), .B(n41222), .Z(n39115) );
  ANDN U41557 ( .B(n41223), .A(n41990), .Z(n41989) );
  XNOR U41558 ( .A(n41991), .B(n41226), .Z(n38548) );
  ANDN U41559 ( .B(n41227), .A(n41992), .Z(n41991) );
  ANDN U41560 ( .B(n34908), .A(n37655), .Z(n41960) );
  IV U41561 ( .A(n36679), .Z(n37655) );
  XOR U41562 ( .A(n38950), .B(n41993), .Z(n36679) );
  XOR U41563 ( .A(n41994), .B(n41995), .Z(n38950) );
  XOR U41564 ( .A(n41170), .B(n37051), .Z(n34908) );
  XNOR U41565 ( .A(n41998), .B(n41999), .Z(n41170) );
  AND U41566 ( .A(n42000), .B(n42001), .Z(n41998) );
  XOR U41567 ( .A(n42002), .B(n37663), .Z(n35690) );
  XOR U41568 ( .A(n35769), .B(n42003), .Z(n37663) );
  IV U41569 ( .A(n38271), .Z(n35769) );
  XOR U41570 ( .A(n42004), .B(n42005), .Z(n38271) );
  XOR U41571 ( .A(n41952), .B(n36935), .Z(n36687) );
  XNOR U41572 ( .A(n42006), .B(n41051), .Z(n41952) );
  ANDN U41573 ( .B(n42007), .A(n42008), .Z(n42006) );
  XOR U41574 ( .A(n42009), .B(n38339), .Z(n34917) );
  XNOR U41575 ( .A(n42010), .B(n39445), .Z(n33356) );
  IV U41576 ( .A(n39435), .Z(n39445) );
  XOR U41577 ( .A(n42011), .B(n39406), .Z(n39435) );
  XNOR U41578 ( .A(n40131), .B(n42012), .Z(n39406) );
  XOR U41579 ( .A(n42013), .B(n42014), .Z(n40131) );
  XNOR U41580 ( .A(n37534), .B(n39750), .Z(n42014) );
  XOR U41581 ( .A(n42015), .B(n41833), .Z(n39750) );
  ANDN U41582 ( .B(n42016), .A(n42017), .Z(n42015) );
  XOR U41583 ( .A(n42018), .B(n41837), .Z(n37534) );
  ANDN U41584 ( .B(n42019), .A(n42020), .Z(n42018) );
  XNOR U41585 ( .A(n39177), .B(n42021), .Z(n42013) );
  XOR U41586 ( .A(n42022), .B(n42023), .Z(n42021) );
  XOR U41587 ( .A(n42024), .B(n41823), .Z(n39177) );
  ANDN U41588 ( .B(n42025), .A(n42026), .Z(n42024) );
  ANDN U41589 ( .B(n36685), .A(n34921), .Z(n42010) );
  XOR U41590 ( .A(n42027), .B(n38997), .Z(n34921) );
  XOR U41591 ( .A(n41199), .B(n36907), .Z(n36685) );
  XNOR U41592 ( .A(n42028), .B(n39576), .Z(n36907) );
  XOR U41593 ( .A(n42029), .B(n42030), .Z(n39576) );
  XOR U41594 ( .A(n37878), .B(n42031), .Z(n42030) );
  XOR U41595 ( .A(n42032), .B(n42033), .Z(n37878) );
  ANDN U41596 ( .B(n41762), .A(n41763), .Z(n42032) );
  XOR U41597 ( .A(n34634), .B(n42034), .Z(n42029) );
  XNOR U41598 ( .A(n39926), .B(n39534), .Z(n42034) );
  XNOR U41599 ( .A(n42035), .B(n42036), .Z(n39534) );
  AND U41600 ( .A(n41771), .B(n41773), .Z(n42035) );
  XOR U41601 ( .A(n42037), .B(n42038), .Z(n39926) );
  ANDN U41602 ( .B(n41779), .A(n41781), .Z(n42037) );
  XNOR U41603 ( .A(n42039), .B(n42040), .Z(n34634) );
  ANDN U41604 ( .B(n41775), .A(n42041), .Z(n42039) );
  XNOR U41605 ( .A(n42042), .B(n42043), .Z(n41199) );
  NOR U41606 ( .A(n41973), .B(n41972), .Z(n42042) );
  XOR U41607 ( .A(n42044), .B(n42045), .Z(n38868) );
  XNOR U41608 ( .A(n34440), .B(n37631), .Z(n42045) );
  XNOR U41609 ( .A(n42046), .B(n37451), .Z(n37631) );
  XOR U41610 ( .A(n39930), .B(n42047), .Z(n37451) );
  ANDN U41611 ( .B(n37356), .A(n36691), .Z(n42046) );
  XOR U41612 ( .A(n42048), .B(n38997), .Z(n36691) );
  XOR U41613 ( .A(n42049), .B(n42050), .Z(n38997) );
  XOR U41614 ( .A(n38616), .B(n42051), .Z(n37356) );
  XOR U41615 ( .A(n42052), .B(n37650), .Z(n34440) );
  XOR U41616 ( .A(n42053), .B(n38843), .Z(n37650) );
  NOR U41617 ( .A(n37649), .B(n34945), .Z(n42052) );
  XNOR U41618 ( .A(n40448), .B(n39470), .Z(n34945) );
  IV U41619 ( .A(n38438), .Z(n39470) );
  XNOR U41620 ( .A(n42056), .B(n42057), .Z(n41490) );
  XNOR U41621 ( .A(n39091), .B(n42058), .Z(n42057) );
  XOR U41622 ( .A(n42059), .B(n42060), .Z(n39091) );
  ANDN U41623 ( .B(n40452), .A(n42061), .Z(n42059) );
  XOR U41624 ( .A(n42062), .B(n42063), .Z(n42056) );
  XOR U41625 ( .A(n40650), .B(n38114), .Z(n42063) );
  XOR U41626 ( .A(n42064), .B(n42065), .Z(n38114) );
  ANDN U41627 ( .B(n42066), .A(n42067), .Z(n42064) );
  XNOR U41628 ( .A(n42068), .B(n42069), .Z(n40650) );
  NOR U41629 ( .A(n41186), .B(n41184), .Z(n42068) );
  XNOR U41630 ( .A(n42071), .B(n42072), .Z(n40448) );
  NOR U41631 ( .A(n42066), .B(n42073), .Z(n42071) );
  XOR U41632 ( .A(n42074), .B(n35093), .Z(n37649) );
  XNOR U41633 ( .A(n42075), .B(n42076), .Z(n35093) );
  XOR U41634 ( .A(n32925), .B(n42077), .Z(n42044) );
  XNOR U41635 ( .A(n31879), .B(n33951), .Z(n42077) );
  XNOR U41636 ( .A(n42078), .B(n37456), .Z(n33951) );
  XOR U41637 ( .A(n42079), .B(n39238), .Z(n37456) );
  IV U41638 ( .A(n38934), .Z(n39238) );
  XOR U41639 ( .A(n42080), .B(n40924), .Z(n38934) );
  XNOR U41640 ( .A(n42081), .B(n42082), .Z(n40924) );
  XNOR U41641 ( .A(n39464), .B(n39024), .Z(n42082) );
  XNOR U41642 ( .A(n42083), .B(n42084), .Z(n39024) );
  ANDN U41643 ( .B(n42085), .A(n42086), .Z(n42083) );
  XNOR U41644 ( .A(n42087), .B(n42088), .Z(n39464) );
  ANDN U41645 ( .B(n42089), .A(n42090), .Z(n42087) );
  XNOR U41646 ( .A(n39599), .B(n42091), .Z(n42081) );
  XOR U41647 ( .A(n38666), .B(n42092), .Z(n42091) );
  XOR U41648 ( .A(n42093), .B(n42094), .Z(n38666) );
  XOR U41649 ( .A(n42097), .B(n42098), .Z(n39599) );
  ANDN U41650 ( .B(n42099), .A(n42100), .Z(n42097) );
  NOR U41651 ( .A(n37360), .B(n34932), .Z(n42078) );
  XNOR U41652 ( .A(n42101), .B(n39468), .Z(n34932) );
  XNOR U41653 ( .A(n42102), .B(n42103), .Z(n40830) );
  XNOR U41654 ( .A(n42104), .B(n38258), .Z(n42103) );
  XNOR U41655 ( .A(n42105), .B(n42106), .Z(n38258) );
  NOR U41656 ( .A(n42107), .B(n42108), .Z(n42105) );
  XOR U41657 ( .A(n36546), .B(n42109), .Z(n42102) );
  XOR U41658 ( .A(n37088), .B(n41365), .Z(n42109) );
  XOR U41659 ( .A(n42110), .B(n42111), .Z(n41365) );
  NOR U41660 ( .A(n42112), .B(n42113), .Z(n42110) );
  XNOR U41661 ( .A(n42114), .B(n42115), .Z(n37088) );
  NOR U41662 ( .A(n42120), .B(n42121), .Z(n42118) );
  XOR U41663 ( .A(n38535), .B(n42123), .Z(n37360) );
  XNOR U41664 ( .A(n39893), .B(n42124), .Z(n38535) );
  XOR U41665 ( .A(n42125), .B(n42126), .Z(n39893) );
  XNOR U41666 ( .A(n42127), .B(n39577), .Z(n42126) );
  XNOR U41667 ( .A(n42128), .B(n42129), .Z(n39577) );
  ANDN U41668 ( .B(n42130), .A(n42131), .Z(n42128) );
  XOR U41669 ( .A(n39694), .B(n42132), .Z(n42125) );
  XOR U41670 ( .A(n38026), .B(n38767), .Z(n42132) );
  XNOR U41671 ( .A(n42133), .B(n42134), .Z(n38767) );
  ANDN U41672 ( .B(n42135), .A(n42136), .Z(n42133) );
  XOR U41673 ( .A(n42137), .B(n42138), .Z(n38026) );
  ANDN U41674 ( .B(n42139), .A(n42140), .Z(n42137) );
  XNOR U41675 ( .A(n42141), .B(n42142), .Z(n39694) );
  NOR U41676 ( .A(n42143), .B(n42144), .Z(n42141) );
  XNOR U41677 ( .A(n42145), .B(n37445), .Z(n31879) );
  XNOR U41678 ( .A(n41560), .B(n39484), .Z(n37445) );
  XOR U41679 ( .A(n41580), .B(n42146), .Z(n39484) );
  XOR U41680 ( .A(n42147), .B(n42148), .Z(n41580) );
  XNOR U41681 ( .A(n38313), .B(n40483), .Z(n42148) );
  XNOR U41682 ( .A(n42149), .B(n40492), .Z(n40483) );
  AND U41683 ( .A(n40493), .B(n42150), .Z(n42149) );
  XNOR U41684 ( .A(n42151), .B(n40497), .Z(n38313) );
  AND U41685 ( .A(n41564), .B(n40498), .Z(n42151) );
  XNOR U41686 ( .A(n42152), .B(n42153), .Z(n40498) );
  XOR U41687 ( .A(n37709), .B(n42154), .Z(n42147) );
  XOR U41688 ( .A(n38874), .B(n37726), .Z(n42154) );
  XNOR U41689 ( .A(n42155), .B(n40489), .Z(n37726) );
  ANDN U41690 ( .B(n41558), .A(n40488), .Z(n42155) );
  XNOR U41691 ( .A(n42156), .B(n42157), .Z(n40488) );
  XNOR U41692 ( .A(n42158), .B(n40501), .Z(n38874) );
  ANDN U41693 ( .B(n40502), .A(n41555), .Z(n42158) );
  XOR U41694 ( .A(n42159), .B(n42160), .Z(n40502) );
  XNOR U41695 ( .A(n42161), .B(n40506), .Z(n37709) );
  AND U41696 ( .A(n41567), .B(n40505), .Z(n42161) );
  XOR U41697 ( .A(n42162), .B(n42163), .Z(n40505) );
  XNOR U41698 ( .A(n42164), .B(n40493), .Z(n41560) );
  XNOR U41699 ( .A(n42165), .B(n42166), .Z(n40493) );
  NOR U41700 ( .A(n42167), .B(n42150), .Z(n42164) );
  NOR U41701 ( .A(n34937), .B(n37358), .Z(n42145) );
  XNOR U41702 ( .A(n37479), .B(n42168), .Z(n37358) );
  XOR U41703 ( .A(n42169), .B(n41398), .Z(n37479) );
  XNOR U41704 ( .A(n42170), .B(n42171), .Z(n41398) );
  XOR U41705 ( .A(n39886), .B(n37601), .Z(n42171) );
  XNOR U41706 ( .A(n42172), .B(n41621), .Z(n37601) );
  NOR U41707 ( .A(n42173), .B(n41630), .Z(n42172) );
  XOR U41708 ( .A(n42174), .B(n41460), .Z(n39886) );
  ANDN U41709 ( .B(n42175), .A(n41626), .Z(n42174) );
  XOR U41710 ( .A(n39411), .B(n42176), .Z(n42170) );
  XNOR U41711 ( .A(n39163), .B(n36416), .Z(n42176) );
  XOR U41712 ( .A(n42177), .B(n41463), .Z(n36416) );
  ANDN U41713 ( .B(n42178), .A(n42179), .Z(n42177) );
  XNOR U41714 ( .A(n42180), .B(n41470), .Z(n39163) );
  ANDN U41715 ( .B(n42181), .A(n41632), .Z(n42180) );
  XNOR U41716 ( .A(n42182), .B(n41474), .Z(n39411) );
  ANDN U41717 ( .B(n42183), .A(n41634), .Z(n42182) );
  IV U41718 ( .A(n42184), .Z(n41634) );
  XNOR U41719 ( .A(n37868), .B(n40956), .Z(n34937) );
  XNOR U41720 ( .A(n42185), .B(n42186), .Z(n40956) );
  ANDN U41721 ( .B(n42187), .A(n42188), .Z(n42185) );
  XNOR U41722 ( .A(n42189), .B(n37453), .Z(n32925) );
  XNOR U41723 ( .A(n40289), .B(n38401), .Z(n37453) );
  XNOR U41724 ( .A(n39803), .B(n41753), .Z(n38401) );
  XNOR U41725 ( .A(n42190), .B(n42191), .Z(n41753) );
  XNOR U41726 ( .A(n40128), .B(n38685), .Z(n42191) );
  XNOR U41727 ( .A(n42192), .B(n41676), .Z(n38685) );
  ANDN U41728 ( .B(n40283), .A(n40281), .Z(n42192) );
  IV U41729 ( .A(n42193), .Z(n40281) );
  XOR U41730 ( .A(n42194), .B(n41667), .Z(n40128) );
  ANDN U41731 ( .B(n40291), .A(n40292), .Z(n42194) );
  XOR U41732 ( .A(n39124), .B(n42195), .Z(n42190) );
  XOR U41733 ( .A(n40190), .B(n42196), .Z(n42195) );
  XOR U41734 ( .A(n42197), .B(n41678), .Z(n40190) );
  XOR U41735 ( .A(n42198), .B(n41671), .Z(n39124) );
  NOR U41736 ( .A(n42199), .B(n42200), .Z(n42198) );
  XNOR U41737 ( .A(n42201), .B(n42202), .Z(n39803) );
  XNOR U41738 ( .A(n39846), .B(n40833), .Z(n42202) );
  XOR U41739 ( .A(n42203), .B(n42204), .Z(n40833) );
  ANDN U41740 ( .B(n40555), .A(n40556), .Z(n42203) );
  XOR U41741 ( .A(n42205), .B(n42206), .Z(n40556) );
  XOR U41742 ( .A(n42207), .B(n42208), .Z(n39846) );
  ANDN U41743 ( .B(n40559), .A(n40560), .Z(n42207) );
  XOR U41744 ( .A(n42209), .B(n42210), .Z(n40560) );
  XOR U41745 ( .A(n38938), .B(n42211), .Z(n42201) );
  XOR U41746 ( .A(n37436), .B(n37835), .Z(n42211) );
  XNOR U41747 ( .A(n42212), .B(n42213), .Z(n37835) );
  ANDN U41748 ( .B(n40550), .A(n40552), .Z(n42212) );
  XNOR U41749 ( .A(n42214), .B(n42215), .Z(n40552) );
  XNOR U41750 ( .A(n42216), .B(n42217), .Z(n37436) );
  ANDN U41751 ( .B(n40563), .A(n40564), .Z(n42216) );
  XOR U41752 ( .A(n42218), .B(n42219), .Z(n40564) );
  XNOR U41753 ( .A(n42220), .B(n42221), .Z(n38938) );
  ANDN U41754 ( .B(n40546), .A(n40547), .Z(n42220) );
  XOR U41755 ( .A(n42222), .B(n42223), .Z(n40547) );
  XNOR U41756 ( .A(n42224), .B(n42199), .Z(n40289) );
  ANDN U41757 ( .B(n42200), .A(n41670), .Z(n42224) );
  ANDN U41758 ( .B(n37637), .A(n34941), .Z(n42189) );
  XOR U41759 ( .A(n41946), .B(n36935), .Z(n34941) );
  XOR U41760 ( .A(n42225), .B(n42226), .Z(n36935) );
  XOR U41761 ( .A(n42227), .B(n41055), .Z(n41946) );
  ANDN U41762 ( .B(n42228), .A(n42229), .Z(n42227) );
  XOR U41763 ( .A(n35315), .B(n42230), .Z(n37637) );
  XNOR U41764 ( .A(n42231), .B(n27367), .Z(n28038) );
  XOR U41765 ( .A(n39874), .B(n31968), .Z(n27367) );
  XNOR U41766 ( .A(n42232), .B(n42233), .Z(n38757) );
  XNOR U41767 ( .A(n32222), .B(n30484), .Z(n42233) );
  XOR U41768 ( .A(n42234), .B(n38073), .Z(n30484) );
  XOR U41769 ( .A(n42235), .B(n39404), .Z(n38073) );
  XOR U41770 ( .A(n39711), .B(n42236), .Z(n39404) );
  XOR U41771 ( .A(n42237), .B(n42238), .Z(n39711) );
  XNOR U41772 ( .A(n39736), .B(n39627), .Z(n42238) );
  XOR U41773 ( .A(n42239), .B(n42240), .Z(n39627) );
  XOR U41774 ( .A(n42243), .B(n42244), .Z(n39736) );
  NOR U41775 ( .A(n42245), .B(n42246), .Z(n42243) );
  XOR U41776 ( .A(n39212), .B(n42247), .Z(n42237) );
  XNOR U41777 ( .A(n42248), .B(n42249), .Z(n42247) );
  XOR U41778 ( .A(n42250), .B(n42251), .Z(n39212) );
  ANDN U41779 ( .B(n42252), .A(n42253), .Z(n42250) );
  ANDN U41780 ( .B(n38074), .A(n36743), .Z(n42234) );
  XOR U41781 ( .A(n38498), .B(n42254), .Z(n36743) );
  IV U41782 ( .A(n38260), .Z(n38498) );
  XNOR U41783 ( .A(n40626), .B(n40972), .Z(n38260) );
  XNOR U41784 ( .A(n42255), .B(n42256), .Z(n40972) );
  XOR U41785 ( .A(n37334), .B(n36975), .Z(n42256) );
  XOR U41786 ( .A(n42257), .B(n42258), .Z(n36975) );
  XNOR U41787 ( .A(n42261), .B(n42262), .Z(n37334) );
  NOR U41788 ( .A(n42263), .B(n41130), .Z(n42261) );
  XOR U41789 ( .A(n41146), .B(n42264), .Z(n42255) );
  XOR U41790 ( .A(n39166), .B(n38427), .Z(n42264) );
  XNOR U41791 ( .A(n42265), .B(n42266), .Z(n38427) );
  NOR U41792 ( .A(n41134), .B(n42267), .Z(n42265) );
  IV U41793 ( .A(n42268), .Z(n41134) );
  XNOR U41794 ( .A(n42269), .B(n42270), .Z(n39166) );
  XNOR U41795 ( .A(n42272), .B(n42273), .Z(n41146) );
  NOR U41796 ( .A(n42274), .B(n42275), .Z(n42272) );
  XNOR U41797 ( .A(n42276), .B(n42277), .Z(n40626) );
  XNOR U41798 ( .A(n39688), .B(n37885), .Z(n42277) );
  XNOR U41799 ( .A(n42278), .B(n42279), .Z(n37885) );
  ANDN U41800 ( .B(n42280), .A(n42281), .Z(n42278) );
  XNOR U41801 ( .A(n42282), .B(n42283), .Z(n39688) );
  ANDN U41802 ( .B(n42284), .A(n42285), .Z(n42282) );
  XOR U41803 ( .A(n37522), .B(n42286), .Z(n42276) );
  XOR U41804 ( .A(n37853), .B(n42287), .Z(n42286) );
  XNOR U41805 ( .A(n42288), .B(n42289), .Z(n37853) );
  NOR U41806 ( .A(n42290), .B(n42291), .Z(n42288) );
  XNOR U41807 ( .A(n42292), .B(n42293), .Z(n37522) );
  NOR U41808 ( .A(n42294), .B(n42295), .Z(n42292) );
  XOR U41809 ( .A(n42196), .B(n39125), .Z(n38074) );
  IV U41810 ( .A(n38686), .Z(n39125) );
  XOR U41811 ( .A(n39641), .B(n40834), .Z(n38686) );
  XNOR U41812 ( .A(n42296), .B(n42297), .Z(n40834) );
  XNOR U41813 ( .A(n42298), .B(n37796), .Z(n42297) );
  XOR U41814 ( .A(n42299), .B(n41505), .Z(n37796) );
  NOR U41815 ( .A(n40550), .B(n42213), .Z(n42299) );
  XOR U41816 ( .A(n42300), .B(n42301), .Z(n40550) );
  XOR U41817 ( .A(n38185), .B(n42302), .Z(n42296) );
  XNOR U41818 ( .A(n38806), .B(n39434), .Z(n42302) );
  XOR U41819 ( .A(n42303), .B(n41512), .Z(n39434) );
  NOR U41820 ( .A(n42304), .B(n40559), .Z(n42303) );
  XOR U41821 ( .A(n42305), .B(n42306), .Z(n40559) );
  XOR U41822 ( .A(n42307), .B(n41508), .Z(n38806) );
  NOR U41823 ( .A(n40563), .B(n42217), .Z(n42307) );
  XNOR U41824 ( .A(n42308), .B(n42309), .Z(n40563) );
  XNOR U41825 ( .A(n42310), .B(n41503), .Z(n38185) );
  NOR U41826 ( .A(n42311), .B(n40546), .Z(n42310) );
  XNOR U41827 ( .A(n42312), .B(n42313), .Z(n40546) );
  XOR U41828 ( .A(n42314), .B(n42315), .Z(n39641) );
  XNOR U41829 ( .A(n37728), .B(n38738), .Z(n42315) );
  XNOR U41830 ( .A(n42316), .B(n41679), .Z(n38738) );
  NOR U41831 ( .A(n40285), .B(n41678), .Z(n42316) );
  XOR U41832 ( .A(n42317), .B(n42318), .Z(n41678) );
  XOR U41833 ( .A(n42319), .B(n42320), .Z(n40285) );
  XNOR U41834 ( .A(n42321), .B(n41681), .Z(n37728) );
  ANDN U41835 ( .B(n40295), .A(n41682), .Z(n42321) );
  XOR U41836 ( .A(n37626), .B(n42322), .Z(n42314) );
  XOR U41837 ( .A(n41662), .B(n37719), .Z(n42322) );
  XNOR U41838 ( .A(n42323), .B(n41668), .Z(n37719) );
  NOR U41839 ( .A(n40291), .B(n41667), .Z(n42323) );
  XNOR U41840 ( .A(n42324), .B(n42325), .Z(n41667) );
  XOR U41841 ( .A(n42326), .B(n42327), .Z(n40291) );
  XNOR U41842 ( .A(n42328), .B(n41675), .Z(n41662) );
  ANDN U41843 ( .B(n41676), .A(n42193), .Z(n42328) );
  XNOR U41844 ( .A(n42329), .B(n42330), .Z(n42193) );
  XOR U41845 ( .A(n42331), .B(n42332), .Z(n41676) );
  XNOR U41846 ( .A(n42333), .B(n41672), .Z(n37626) );
  ANDN U41847 ( .B(n42199), .A(n41671), .Z(n42333) );
  XOR U41848 ( .A(n42334), .B(n42335), .Z(n41671) );
  XOR U41849 ( .A(n42336), .B(n42337), .Z(n42199) );
  XOR U41850 ( .A(n42338), .B(n41682), .Z(n42196) );
  XNOR U41851 ( .A(n42339), .B(n42340), .Z(n41682) );
  NOR U41852 ( .A(n40295), .B(n40296), .Z(n42338) );
  XOR U41853 ( .A(n42341), .B(n42342), .Z(n40295) );
  XNOR U41854 ( .A(n42343), .B(n38064), .Z(n32222) );
  XOR U41855 ( .A(n40671), .B(n42344), .Z(n38064) );
  IV U41856 ( .A(n38858), .Z(n40671) );
  XOR U41857 ( .A(n40625), .B(n39986), .Z(n38858) );
  XOR U41858 ( .A(n42345), .B(n42346), .Z(n39986) );
  XNOR U41859 ( .A(n39144), .B(n39398), .Z(n42346) );
  XNOR U41860 ( .A(n42347), .B(n42348), .Z(n39398) );
  AND U41861 ( .A(n42349), .B(n42350), .Z(n42347) );
  AND U41862 ( .A(n42353), .B(n42354), .Z(n42351) );
  XOR U41863 ( .A(n42355), .B(n42356), .Z(n42345) );
  XNOR U41864 ( .A(n38148), .B(n42357), .Z(n42356) );
  XOR U41865 ( .A(n42358), .B(n42359), .Z(n38148) );
  AND U41866 ( .A(n42360), .B(n42361), .Z(n42358) );
  XOR U41867 ( .A(n42362), .B(n42363), .Z(n40625) );
  XNOR U41868 ( .A(n36900), .B(n39022), .Z(n42363) );
  XNOR U41869 ( .A(n42364), .B(n42365), .Z(n39022) );
  ANDN U41870 ( .B(n42366), .A(n42367), .Z(n42364) );
  XNOR U41871 ( .A(n42368), .B(n42369), .Z(n36900) );
  ANDN U41872 ( .B(n42370), .A(n42371), .Z(n42368) );
  XOR U41873 ( .A(n40369), .B(n42372), .Z(n42362) );
  XNOR U41874 ( .A(n39780), .B(n37904), .Z(n42372) );
  XOR U41875 ( .A(n42373), .B(n42374), .Z(n37904) );
  NOR U41876 ( .A(n42375), .B(n42376), .Z(n42373) );
  XNOR U41877 ( .A(n42377), .B(n42378), .Z(n39780) );
  AND U41878 ( .A(n42379), .B(n42380), .Z(n42377) );
  XNOR U41879 ( .A(n42381), .B(n42382), .Z(n40369) );
  ANDN U41880 ( .B(n42383), .A(n42384), .Z(n42381) );
  NOR U41881 ( .A(n42385), .B(n36757), .Z(n42343) );
  XOR U41882 ( .A(n32946), .B(n42386), .Z(n42232) );
  XOR U41883 ( .A(n32707), .B(n38039), .Z(n42386) );
  XNOR U41884 ( .A(n42387), .B(n38061), .Z(n38039) );
  XNOR U41885 ( .A(n38242), .B(n42388), .Z(n38061) );
  XNOR U41886 ( .A(n42389), .B(n35932), .Z(n36747) );
  XOR U41887 ( .A(n40304), .B(n36507), .Z(n38062) );
  IV U41888 ( .A(n36535), .Z(n36507) );
  XNOR U41889 ( .A(n40519), .B(n38689), .Z(n36535) );
  XNOR U41890 ( .A(n42390), .B(n42391), .Z(n38689) );
  XNOR U41891 ( .A(n38610), .B(n37271), .Z(n42391) );
  XNOR U41892 ( .A(n42392), .B(n42393), .Z(n37271) );
  ANDN U41893 ( .B(n40310), .A(n40312), .Z(n42392) );
  XNOR U41894 ( .A(n42394), .B(n40399), .Z(n38610) );
  ANDN U41895 ( .B(n40318), .A(n40319), .Z(n42394) );
  XOR U41896 ( .A(n42395), .B(n42396), .Z(n40318) );
  XNOR U41897 ( .A(n38430), .B(n42397), .Z(n42390) );
  XOR U41898 ( .A(n39220), .B(n40148), .Z(n42397) );
  XOR U41899 ( .A(n42398), .B(n40155), .Z(n40148) );
  XNOR U41900 ( .A(n42400), .B(n41545), .Z(n39220) );
  ANDN U41901 ( .B(n40314), .A(n40315), .Z(n42400) );
  XNOR U41902 ( .A(n42401), .B(n42402), .Z(n40314) );
  XNOR U41903 ( .A(n42403), .B(n40163), .Z(n38430) );
  ANDN U41904 ( .B(n40162), .A(n40306), .Z(n42403) );
  XNOR U41905 ( .A(n42404), .B(n42405), .Z(n40162) );
  XOR U41906 ( .A(n42406), .B(n42407), .Z(n40519) );
  XNOR U41907 ( .A(n42408), .B(n38773), .Z(n42407) );
  XNOR U41908 ( .A(n42409), .B(n42410), .Z(n38773) );
  AND U41909 ( .A(n40722), .B(n40724), .Z(n42409) );
  XOR U41910 ( .A(n39013), .B(n42411), .Z(n42406) );
  XOR U41911 ( .A(n36361), .B(n42412), .Z(n42411) );
  XOR U41912 ( .A(n42413), .B(n42414), .Z(n36361) );
  AND U41913 ( .A(n40711), .B(n40709), .Z(n42413) );
  XNOR U41914 ( .A(n42415), .B(n42416), .Z(n39013) );
  AND U41915 ( .A(n40713), .B(n40715), .Z(n42415) );
  XNOR U41916 ( .A(n42417), .B(n40156), .Z(n40304) );
  XOR U41917 ( .A(n42418), .B(n42419), .Z(n40156) );
  NOR U41918 ( .A(n42399), .B(n42420), .Z(n42417) );
  XNOR U41919 ( .A(n42421), .B(n40206), .Z(n32707) );
  IV U41920 ( .A(n38071), .Z(n40206) );
  XOR U41921 ( .A(n42422), .B(n37264), .Z(n38071) );
  XNOR U41922 ( .A(n42423), .B(n40464), .Z(n37264) );
  XNOR U41923 ( .A(n42424), .B(n42425), .Z(n40464) );
  XNOR U41924 ( .A(n42426), .B(n37783), .Z(n42425) );
  XNOR U41925 ( .A(n42427), .B(n42428), .Z(n37783) );
  ANDN U41926 ( .B(n42429), .A(n42430), .Z(n42427) );
  XOR U41927 ( .A(n39539), .B(n42431), .Z(n42424) );
  XOR U41928 ( .A(n35798), .B(n38105), .Z(n42431) );
  XNOR U41929 ( .A(n42432), .B(n42433), .Z(n38105) );
  NOR U41930 ( .A(n42434), .B(n42435), .Z(n42432) );
  XNOR U41931 ( .A(n42436), .B(n42437), .Z(n35798) );
  XNOR U41932 ( .A(n42440), .B(n42441), .Z(n39539) );
  ANDN U41933 ( .B(n42442), .A(n42443), .Z(n42440) );
  ANDN U41934 ( .B(n39879), .A(n38070), .Z(n42421) );
  XNOR U41935 ( .A(n39761), .B(n42444), .Z(n38070) );
  IV U41936 ( .A(n37148), .Z(n39761) );
  XNOR U41937 ( .A(n40126), .B(n42445), .Z(n37148) );
  XOR U41938 ( .A(n42446), .B(n42447), .Z(n40126) );
  XNOR U41939 ( .A(n37956), .B(n36422), .Z(n42447) );
  XOR U41940 ( .A(n42448), .B(n39907), .Z(n36422) );
  ANDN U41941 ( .B(n41251), .A(n41249), .Z(n42448) );
  XOR U41942 ( .A(n42449), .B(n42450), .Z(n41249) );
  XOR U41943 ( .A(n42451), .B(n39902), .Z(n37956) );
  AND U41944 ( .A(n41240), .B(n39903), .Z(n42451) );
  XOR U41945 ( .A(n42452), .B(n42453), .Z(n39903) );
  XOR U41946 ( .A(n38688), .B(n42454), .Z(n42446) );
  XNOR U41947 ( .A(n38559), .B(n38659), .Z(n42454) );
  XNOR U41948 ( .A(n42455), .B(n39916), .Z(n38659) );
  ANDN U41949 ( .B(n41244), .A(n39915), .Z(n42455) );
  XOR U41950 ( .A(n42456), .B(n42457), .Z(n39915) );
  XOR U41951 ( .A(n42458), .B(n42459), .Z(n38559) );
  ANDN U41952 ( .B(n39912), .A(n41236), .Z(n42458) );
  XOR U41953 ( .A(n42460), .B(n42461), .Z(n39912) );
  XNOR U41954 ( .A(n42462), .B(n39898), .Z(n38688) );
  ANDN U41955 ( .B(n39899), .A(n41246), .Z(n42462) );
  XOR U41956 ( .A(n42395), .B(n42463), .Z(n39899) );
  XOR U41957 ( .A(n42464), .B(n35929), .Z(n39879) );
  XNOR U41958 ( .A(n42465), .B(n38413), .Z(n32946) );
  XOR U41959 ( .A(n41845), .B(n35301), .Z(n38413) );
  XNOR U41960 ( .A(n42466), .B(n42467), .Z(n41845) );
  NOR U41961 ( .A(n42468), .B(n42469), .Z(n42466) );
  XNOR U41962 ( .A(n38959), .B(n42470), .Z(n36753) );
  XOR U41963 ( .A(n38883), .B(n42471), .Z(n38414) );
  IV U41964 ( .A(n37209), .Z(n38883) );
  XNOR U41965 ( .A(n41087), .B(n40801), .Z(n37209) );
  XNOR U41966 ( .A(n42472), .B(n42473), .Z(n40801) );
  XNOR U41967 ( .A(n38291), .B(n38239), .Z(n42473) );
  XNOR U41968 ( .A(n42474), .B(n41909), .Z(n38239) );
  ANDN U41969 ( .B(n42475), .A(n42476), .Z(n42474) );
  XNOR U41970 ( .A(n42477), .B(n41897), .Z(n38291) );
  XNOR U41971 ( .A(n38267), .B(n42480), .Z(n42472) );
  XNOR U41972 ( .A(n36782), .B(n40276), .Z(n42480) );
  XOR U41973 ( .A(n42481), .B(n41905), .Z(n40276) );
  ANDN U41974 ( .B(n42482), .A(n42483), .Z(n42481) );
  XNOR U41975 ( .A(n42484), .B(n41901), .Z(n36782) );
  AND U41976 ( .A(n42485), .B(n42486), .Z(n42484) );
  XNOR U41977 ( .A(n42487), .B(n41913), .Z(n38267) );
  NOR U41978 ( .A(n42488), .B(n42489), .Z(n42487) );
  XOR U41979 ( .A(n42490), .B(n42491), .Z(n41087) );
  XOR U41980 ( .A(n38622), .B(n36954), .Z(n42491) );
  XOR U41981 ( .A(n42492), .B(n40292), .Z(n36954) );
  XOR U41982 ( .A(n42493), .B(n42494), .Z(n40292) );
  ANDN U41983 ( .B(n40293), .A(n41668), .Z(n42492) );
  XNOR U41984 ( .A(n42495), .B(n42496), .Z(n41668) );
  XNOR U41985 ( .A(n42497), .B(n42498), .Z(n40293) );
  XNOR U41986 ( .A(n42499), .B(n42200), .Z(n38622) );
  XNOR U41987 ( .A(n42500), .B(n42501), .Z(n42200) );
  ANDN U41988 ( .B(n41670), .A(n41672), .Z(n42499) );
  XOR U41989 ( .A(n42502), .B(n42503), .Z(n41672) );
  XNOR U41990 ( .A(n42504), .B(n42505), .Z(n41670) );
  XNOR U41991 ( .A(n37498), .B(n42506), .Z(n42490) );
  XNOR U41992 ( .A(n38316), .B(n36544), .Z(n42506) );
  XNOR U41993 ( .A(n42507), .B(n40296), .Z(n36544) );
  XNOR U41994 ( .A(n42508), .B(n42509), .Z(n40296) );
  ANDN U41995 ( .B(n40297), .A(n41681), .Z(n42507) );
  XOR U41996 ( .A(n42510), .B(n42511), .Z(n41681) );
  XOR U41997 ( .A(n42512), .B(n42513), .Z(n40297) );
  XNOR U41998 ( .A(n42514), .B(n40283), .Z(n38316) );
  XNOR U41999 ( .A(n42515), .B(n42516), .Z(n40283) );
  ANDN U42000 ( .B(n40282), .A(n41675), .Z(n42514) );
  XOR U42001 ( .A(n42517), .B(n42518), .Z(n41675) );
  XNOR U42002 ( .A(n42520), .B(n40286), .Z(n37498) );
  XNOR U42003 ( .A(n42521), .B(n42522), .Z(n40286) );
  ANDN U42004 ( .B(n40287), .A(n41679), .Z(n42520) );
  XOR U42005 ( .A(n42523), .B(n42524), .Z(n41679) );
  XNOR U42006 ( .A(n42525), .B(n42526), .Z(n40287) );
  XNOR U42007 ( .A(n42527), .B(n42528), .Z(n33642) );
  XOR U42008 ( .A(n33040), .B(n30141), .Z(n42528) );
  XOR U42009 ( .A(n42529), .B(n38043), .Z(n30141) );
  XOR U42010 ( .A(n38684), .B(n42530), .Z(n38043) );
  XNOR U42011 ( .A(n42531), .B(n42532), .Z(n38684) );
  ANDN U42012 ( .B(n38044), .A(n33937), .Z(n42529) );
  XOR U42013 ( .A(n36413), .B(n42533), .Z(n33937) );
  XNOR U42014 ( .A(n42534), .B(n42535), .Z(n41077) );
  XNOR U42015 ( .A(n34629), .B(n39239), .Z(n42535) );
  XNOR U42016 ( .A(n42536), .B(n41290), .Z(n39239) );
  ANDN U42017 ( .B(n41445), .A(n41446), .Z(n42536) );
  XOR U42018 ( .A(n42537), .B(n42538), .Z(n41446) );
  XNOR U42019 ( .A(n42539), .B(n41287), .Z(n34629) );
  AND U42020 ( .A(n41449), .B(n41448), .Z(n42539) );
  XOR U42021 ( .A(n42540), .B(n42541), .Z(n41449) );
  XOR U42022 ( .A(n39114), .B(n42542), .Z(n42534) );
  XNOR U42023 ( .A(n38550), .B(n39673), .Z(n42542) );
  XOR U42024 ( .A(n42543), .B(n41294), .Z(n39673) );
  ANDN U42025 ( .B(n41441), .A(n41442), .Z(n42543) );
  XOR U42026 ( .A(n42544), .B(n42309), .Z(n41442) );
  XNOR U42027 ( .A(n42545), .B(n41278), .Z(n38550) );
  ANDN U42028 ( .B(n41451), .A(n41452), .Z(n42545) );
  XOR U42029 ( .A(n42546), .B(n42547), .Z(n41452) );
  XNOR U42030 ( .A(n42548), .B(n41282), .Z(n39114) );
  AND U42031 ( .A(n41439), .B(n41438), .Z(n42548) );
  XOR U42032 ( .A(n42549), .B(n42550), .Z(n41439) );
  XOR U42033 ( .A(n42552), .B(n35625), .Z(n38044) );
  IV U42034 ( .A(n37085), .Z(n35625) );
  XNOR U42035 ( .A(n42553), .B(n41400), .Z(n37085) );
  XNOR U42036 ( .A(n42554), .B(n42555), .Z(n41400) );
  XNOR U42037 ( .A(n39698), .B(n39122), .Z(n42555) );
  XNOR U42038 ( .A(n42556), .B(n41934), .Z(n39122) );
  ANDN U42039 ( .B(n42557), .A(n41933), .Z(n42556) );
  XOR U42040 ( .A(n42558), .B(n41937), .Z(n39698) );
  ANDN U42041 ( .B(n41938), .A(n42559), .Z(n42558) );
  XNOR U42042 ( .A(n39150), .B(n42560), .Z(n42554) );
  XOR U42043 ( .A(n39587), .B(n39342), .Z(n42560) );
  XOR U42044 ( .A(n42561), .B(n41929), .Z(n39342) );
  ANDN U42045 ( .B(n42562), .A(n41930), .Z(n42561) );
  XNOR U42046 ( .A(n42563), .B(n41925), .Z(n39587) );
  ANDN U42047 ( .B(n41924), .A(n42564), .Z(n42563) );
  XNOR U42048 ( .A(n42565), .B(n42566), .Z(n39150) );
  ANDN U42049 ( .B(n42567), .A(n42568), .Z(n42565) );
  XNOR U42050 ( .A(n42569), .B(n38050), .Z(n33040) );
  XOR U42051 ( .A(n40381), .B(n38360), .Z(n38050) );
  XNOR U42052 ( .A(n42570), .B(n42571), .Z(n40381) );
  NOR U42053 ( .A(n42572), .B(n42573), .Z(n42570) );
  ANDN U42054 ( .B(n38051), .A(n37806), .Z(n42569) );
  XOR U42055 ( .A(n37684), .B(n42574), .Z(n37806) );
  IV U42056 ( .A(n36513), .Z(n37684) );
  XNOR U42057 ( .A(n42575), .B(n40971), .Z(n36513) );
  XNOR U42058 ( .A(n42576), .B(n42577), .Z(n40971) );
  XOR U42059 ( .A(n38691), .B(n39535), .Z(n42577) );
  XOR U42060 ( .A(n42578), .B(n42579), .Z(n39535) );
  NOR U42061 ( .A(n41496), .B(n42580), .Z(n42578) );
  XNOR U42062 ( .A(n42581), .B(n42582), .Z(n38691) );
  NOR U42063 ( .A(n42583), .B(n40259), .Z(n42581) );
  XOR U42064 ( .A(n38639), .B(n42584), .Z(n42576) );
  XOR U42065 ( .A(n42585), .B(n42586), .Z(n42584) );
  XNOR U42066 ( .A(n42587), .B(n42588), .Z(n38639) );
  ANDN U42067 ( .B(n42589), .A(n42590), .Z(n42587) );
  XOR U42068 ( .A(n42591), .B(n34368), .Z(n38051) );
  XNOR U42069 ( .A(n42592), .B(n41336), .Z(n34368) );
  XOR U42070 ( .A(n42593), .B(n42594), .Z(n41336) );
  XNOR U42071 ( .A(n38461), .B(n42389), .Z(n42594) );
  XNOR U42072 ( .A(n42595), .B(n42596), .Z(n42389) );
  ANDN U42073 ( .B(n42597), .A(n40227), .Z(n42595) );
  XOR U42074 ( .A(n42598), .B(n42599), .Z(n38461) );
  AND U42075 ( .A(n40231), .B(n42600), .Z(n42598) );
  XOR U42076 ( .A(n42601), .B(n42602), .Z(n42593) );
  XNOR U42077 ( .A(n35931), .B(n38565), .Z(n42602) );
  XNOR U42078 ( .A(n42603), .B(n42604), .Z(n38565) );
  ANDN U42079 ( .B(n42605), .A(n40244), .Z(n42603) );
  IV U42080 ( .A(n42606), .Z(n40244) );
  XOR U42081 ( .A(n42607), .B(n42608), .Z(n35931) );
  ANDN U42082 ( .B(n42609), .A(n40240), .Z(n42607) );
  XOR U42083 ( .A(n32512), .B(n42610), .Z(n42527) );
  XOR U42084 ( .A(n36498), .B(n31706), .Z(n42610) );
  XNOR U42085 ( .A(n42611), .B(n38056), .Z(n31706) );
  XOR U42086 ( .A(n42612), .B(n39449), .Z(n38056) );
  IV U42087 ( .A(n39938), .Z(n39449) );
  XOR U42088 ( .A(n40698), .B(n39291), .Z(n39938) );
  XNOR U42089 ( .A(n42613), .B(n42614), .Z(n39291) );
  XNOR U42090 ( .A(n40526), .B(n39622), .Z(n42614) );
  XNOR U42091 ( .A(n42615), .B(n42616), .Z(n39622) );
  ANDN U42092 ( .B(n42617), .A(n42618), .Z(n42615) );
  XNOR U42093 ( .A(n42619), .B(n42620), .Z(n40526) );
  ANDN U42094 ( .B(n42621), .A(n42622), .Z(n42619) );
  XNOR U42095 ( .A(n33926), .B(n42623), .Z(n42613) );
  XOR U42096 ( .A(n37191), .B(n42624), .Z(n42623) );
  XNOR U42097 ( .A(n42625), .B(n42626), .Z(n37191) );
  NOR U42098 ( .A(n42627), .B(n42628), .Z(n42625) );
  XNOR U42099 ( .A(n42629), .B(n42630), .Z(n33926) );
  ANDN U42100 ( .B(n42631), .A(n42632), .Z(n42629) );
  XOR U42101 ( .A(n42633), .B(n42634), .Z(n40698) );
  XNOR U42102 ( .A(n40087), .B(n40195), .Z(n42634) );
  XOR U42103 ( .A(n42635), .B(n42636), .Z(n40195) );
  ANDN U42104 ( .B(n40102), .A(n42637), .Z(n42635) );
  XNOR U42105 ( .A(n42638), .B(n42639), .Z(n40087) );
  ANDN U42106 ( .B(n40700), .A(n40702), .Z(n42638) );
  XOR U42107 ( .A(n42640), .B(n42641), .Z(n42633) );
  XNOR U42108 ( .A(n37883), .B(n38928), .Z(n42641) );
  XNOR U42109 ( .A(n42642), .B(n42643), .Z(n38928) );
  ANDN U42110 ( .B(n40112), .A(n40113), .Z(n42642) );
  XNOR U42111 ( .A(n42644), .B(n42645), .Z(n37883) );
  ANDN U42112 ( .B(n40106), .A(n40108), .Z(n42644) );
  ANDN U42113 ( .B(n38057), .A(n36042), .Z(n42611) );
  XNOR U42114 ( .A(n39782), .B(n42646), .Z(n36042) );
  XNOR U42115 ( .A(n42647), .B(n42648), .Z(n39782) );
  XOR U42116 ( .A(n41624), .B(n37197), .Z(n38057) );
  IV U42117 ( .A(n38161), .Z(n37197) );
  XOR U42118 ( .A(n41996), .B(n39179), .Z(n38161) );
  XNOR U42119 ( .A(n42649), .B(n42650), .Z(n39179) );
  XNOR U42120 ( .A(n38975), .B(n42651), .Z(n42650) );
  XOR U42121 ( .A(n42652), .B(n40881), .Z(n38975) );
  ANDN U42122 ( .B(n41651), .A(n41037), .Z(n42652) );
  XOR U42123 ( .A(n42653), .B(n42654), .Z(n41037) );
  XNOR U42124 ( .A(n42655), .B(n42656), .Z(n42649) );
  XNOR U42125 ( .A(n39924), .B(n38818), .Z(n42656) );
  XNOR U42126 ( .A(n42657), .B(n40910), .Z(n38818) );
  XNOR U42127 ( .A(n42658), .B(n42659), .Z(n41028) );
  XOR U42128 ( .A(n42660), .B(n40886), .Z(n39924) );
  ANDN U42129 ( .B(n41638), .A(n41033), .Z(n42660) );
  XOR U42130 ( .A(n42661), .B(n42662), .Z(n41033) );
  XNOR U42131 ( .A(n42663), .B(n42664), .Z(n41996) );
  XOR U42132 ( .A(n40794), .B(n40439), .Z(n42664) );
  XNOR U42133 ( .A(n42665), .B(n42183), .Z(n40439) );
  ANDN U42134 ( .B(n41472), .A(n42184), .Z(n42665) );
  XOR U42135 ( .A(n42666), .B(n42667), .Z(n42184) );
  XOR U42136 ( .A(n42668), .B(n42669), .Z(n41472) );
  XNOR U42137 ( .A(n42670), .B(n42173), .Z(n40794) );
  ANDN U42138 ( .B(n41630), .A(n41619), .Z(n42670) );
  XOR U42139 ( .A(n42671), .B(n42672), .Z(n41619) );
  XNOR U42140 ( .A(n42673), .B(n42674), .Z(n41630) );
  XNOR U42141 ( .A(n38489), .B(n42675), .Z(n42663) );
  XNOR U42142 ( .A(n35945), .B(n41396), .Z(n42675) );
  XNOR U42143 ( .A(n42676), .B(n42178), .Z(n41396) );
  ANDN U42144 ( .B(n41462), .A(n42677), .Z(n42676) );
  XOR U42145 ( .A(n42678), .B(n42181), .Z(n35945) );
  XOR U42146 ( .A(n42679), .B(n41888), .Z(n41632) );
  XOR U42147 ( .A(n42680), .B(n42681), .Z(n41468) );
  XOR U42148 ( .A(n42682), .B(n42175), .Z(n38489) );
  ANDN U42149 ( .B(n41626), .A(n41627), .Z(n42682) );
  XOR U42150 ( .A(n42683), .B(n42684), .Z(n41627) );
  XOR U42151 ( .A(n42685), .B(n42686), .Z(n41626) );
  XNOR U42152 ( .A(n42687), .B(n42179), .Z(n41624) );
  IV U42153 ( .A(n42677), .Z(n42179) );
  XOR U42154 ( .A(n42688), .B(n42689), .Z(n42677) );
  NOR U42155 ( .A(n41464), .B(n41462), .Z(n42687) );
  XNOR U42156 ( .A(n42690), .B(n42691), .Z(n41462) );
  XNOR U42157 ( .A(n42692), .B(n38046), .Z(n36498) );
  XNOR U42158 ( .A(n41846), .B(n35301), .Z(n38046) );
  XNOR U42159 ( .A(n42694), .B(n42695), .Z(n42226) );
  XOR U42160 ( .A(n38917), .B(n39992), .Z(n42695) );
  XNOR U42161 ( .A(n42696), .B(n42697), .Z(n39992) );
  ANDN U42162 ( .B(n41857), .A(n41858), .Z(n42696) );
  XNOR U42163 ( .A(n42698), .B(n42699), .Z(n38917) );
  NOR U42164 ( .A(n41853), .B(n41854), .Z(n42698) );
  XNOR U42165 ( .A(n37006), .B(n42700), .Z(n42694) );
  XNOR U42166 ( .A(n42701), .B(n40655), .Z(n42700) );
  XOR U42167 ( .A(n42702), .B(n42703), .Z(n40655) );
  NOR U42168 ( .A(n41850), .B(n41849), .Z(n42702) );
  XNOR U42169 ( .A(n42704), .B(n42705), .Z(n37006) );
  AND U42170 ( .A(n42706), .B(n42707), .Z(n42704) );
  XOR U42171 ( .A(n42708), .B(n42706), .Z(n41846) );
  NOR U42172 ( .A(n42707), .B(n42709), .Z(n42708) );
  ANDN U42173 ( .B(n38047), .A(n33844), .Z(n42692) );
  XNOR U42174 ( .A(n42710), .B(n42711), .Z(n33844) );
  XOR U42175 ( .A(n34638), .B(n42712), .Z(n38047) );
  XNOR U42176 ( .A(n42713), .B(n42714), .Z(n39949) );
  XOR U42177 ( .A(n40669), .B(n42715), .Z(n42714) );
  ANDN U42178 ( .B(n42718), .A(n42719), .Z(n42716) );
  XNOR U42179 ( .A(n37963), .B(n42720), .Z(n42713) );
  XOR U42180 ( .A(n40539), .B(n40207), .Z(n42720) );
  AND U42181 ( .A(n42723), .B(n42724), .Z(n42721) );
  XOR U42182 ( .A(n42725), .B(n42726), .Z(n40539) );
  AND U42183 ( .A(n42727), .B(n42728), .Z(n42725) );
  AND U42184 ( .A(n42731), .B(n42732), .Z(n42729) );
  XNOR U42185 ( .A(n42733), .B(n42734), .Z(n40674) );
  XOR U42186 ( .A(n36980), .B(n38846), .Z(n42734) );
  XOR U42187 ( .A(n42735), .B(n42736), .Z(n38846) );
  ANDN U42188 ( .B(n42737), .A(n42738), .Z(n42735) );
  XNOR U42189 ( .A(n42739), .B(n42740), .Z(n36980) );
  NOR U42190 ( .A(n42741), .B(n42742), .Z(n42739) );
  XNOR U42191 ( .A(n40918), .B(n42743), .Z(n42733) );
  XOR U42192 ( .A(n37215), .B(n38107), .Z(n42743) );
  XOR U42193 ( .A(n42744), .B(n42745), .Z(n38107) );
  ANDN U42194 ( .B(n42746), .A(n42747), .Z(n42744) );
  XNOR U42195 ( .A(n42748), .B(n42749), .Z(n37215) );
  ANDN U42196 ( .B(n42750), .A(n42751), .Z(n42748) );
  XOR U42197 ( .A(n42752), .B(n42753), .Z(n40918) );
  ANDN U42198 ( .B(n42754), .A(n42755), .Z(n42752) );
  XNOR U42199 ( .A(n42756), .B(n38053), .Z(n32512) );
  XOR U42200 ( .A(n42757), .B(n36967), .Z(n38053) );
  XOR U42201 ( .A(n42758), .B(n40211), .Z(n36967) );
  XNOR U42202 ( .A(n42759), .B(n42760), .Z(n40211) );
  XOR U42203 ( .A(n38117), .B(n38347), .Z(n42760) );
  XOR U42204 ( .A(n42761), .B(n42113), .Z(n38347) );
  XNOR U42205 ( .A(n42764), .B(n42765), .Z(n38117) );
  ANDN U42206 ( .B(n42766), .A(n42767), .Z(n42764) );
  XOR U42207 ( .A(n39606), .B(n42768), .Z(n42759) );
  XOR U42208 ( .A(n38304), .B(n39631), .Z(n42768) );
  XNOR U42209 ( .A(n42769), .B(n42120), .Z(n39631) );
  ANDN U42210 ( .B(n42770), .A(n42771), .Z(n42769) );
  XNOR U42211 ( .A(n42772), .B(n42116), .Z(n38304) );
  ANDN U42212 ( .B(n42773), .A(n42774), .Z(n42772) );
  XNOR U42213 ( .A(n42775), .B(n42108), .Z(n39606) );
  ANDN U42214 ( .B(n42776), .A(n42777), .Z(n42775) );
  NOR U42215 ( .A(n33228), .B(n38054), .Z(n42756) );
  XNOR U42216 ( .A(n35943), .B(n42779), .Z(n33228) );
  XOR U42217 ( .A(n42780), .B(n38065), .Z(n39874) );
  IV U42218 ( .A(n42385), .Z(n38065) );
  XOR U42219 ( .A(n42412), .B(n36362), .Z(n42385) );
  XOR U42220 ( .A(n42781), .B(n42782), .Z(n42412) );
  AND U42221 ( .A(n36759), .B(n36757), .Z(n42780) );
  XOR U42222 ( .A(n42783), .B(n38174), .Z(n36757) );
  IV U42223 ( .A(n36364), .Z(n38174) );
  XOR U42224 ( .A(n42786), .B(n39482), .Z(n36759) );
  IV U42225 ( .A(n38972), .Z(n39482) );
  XNOR U42226 ( .A(n42787), .B(n42788), .Z(n41891) );
  XOR U42227 ( .A(n40032), .B(n40323), .Z(n42788) );
  XNOR U42228 ( .A(n42789), .B(n42790), .Z(n40323) );
  NOR U42229 ( .A(n42791), .B(n40819), .Z(n42789) );
  XOR U42230 ( .A(n42792), .B(n42793), .Z(n40032) );
  NOR U42231 ( .A(n40806), .B(n42794), .Z(n42792) );
  XNOR U42232 ( .A(n42795), .B(n42796), .Z(n42787) );
  XOR U42233 ( .A(n41084), .B(n39185), .Z(n42796) );
  XOR U42234 ( .A(n42797), .B(n42798), .Z(n39185) );
  AND U42235 ( .A(n42799), .B(n42800), .Z(n42797) );
  XOR U42236 ( .A(n42801), .B(n42802), .Z(n41084) );
  AND U42237 ( .A(n40815), .B(n42803), .Z(n42801) );
  NOR U42238 ( .A(n28981), .B(n28043), .Z(n42231) );
  XOR U42239 ( .A(n33295), .B(n37735), .Z(n28043) );
  XOR U42240 ( .A(n42805), .B(n35063), .Z(n37735) );
  ANDN U42241 ( .B(n35572), .A(n42806), .Z(n42805) );
  XOR U42242 ( .A(n42022), .B(n37535), .Z(n35572) );
  XOR U42243 ( .A(n42807), .B(n42808), .Z(n42022) );
  ANDN U42244 ( .B(n42809), .A(n42810), .Z(n42807) );
  XNOR U42245 ( .A(n35500), .B(n33998), .Z(n33295) );
  XNOR U42246 ( .A(n42811), .B(n42812), .Z(n33998) );
  XNOR U42247 ( .A(n34607), .B(n36858), .Z(n42812) );
  XOR U42248 ( .A(n42813), .B(n38015), .Z(n36858) );
  XOR U42249 ( .A(n42586), .B(n39536), .Z(n38015) );
  IV U42250 ( .A(n38640), .Z(n39536) );
  XOR U42251 ( .A(n42814), .B(n42815), .Z(n42586) );
  NOR U42252 ( .A(n42816), .B(n40255), .Z(n42814) );
  XOR U42253 ( .A(n40159), .B(n38163), .Z(n36881) );
  XOR U42254 ( .A(n42817), .B(n42818), .Z(n38163) );
  XOR U42255 ( .A(n42819), .B(n42820), .Z(n40159) );
  NOR U42256 ( .A(n40310), .B(n42393), .Z(n42819) );
  XOR U42257 ( .A(n42821), .B(n42822), .Z(n40310) );
  XOR U42258 ( .A(n39088), .B(n42823), .Z(n36883) );
  XNOR U42259 ( .A(n41689), .B(n42824), .Z(n39088) );
  XOR U42260 ( .A(n42825), .B(n42826), .Z(n41689) );
  XOR U42261 ( .A(n38908), .B(n38733), .Z(n42826) );
  XNOR U42262 ( .A(n42827), .B(n40740), .Z(n38733) );
  ANDN U42263 ( .B(n42828), .A(n40739), .Z(n42827) );
  XOR U42264 ( .A(n42829), .B(n40752), .Z(n38908) );
  ANDN U42265 ( .B(n40753), .A(n41811), .Z(n42829) );
  XNOR U42266 ( .A(n36366), .B(n42830), .Z(n42825) );
  XOR U42267 ( .A(n40729), .B(n39637), .Z(n42830) );
  XNOR U42268 ( .A(n42831), .B(n40735), .Z(n39637) );
  ANDN U42269 ( .B(n40736), .A(n42832), .Z(n42831) );
  XNOR U42270 ( .A(n42833), .B(n40744), .Z(n40729) );
  NOR U42271 ( .A(n42834), .B(n41814), .Z(n42833) );
  XOR U42272 ( .A(n42835), .B(n40749), .Z(n36366) );
  NOR U42273 ( .A(n42836), .B(n40748), .Z(n42835) );
  XNOR U42274 ( .A(n42837), .B(n36470), .Z(n34607) );
  XOR U42275 ( .A(n42838), .B(n38318), .Z(n36470) );
  XOR U42276 ( .A(n40349), .B(n40329), .Z(n38318) );
  XNOR U42277 ( .A(n42839), .B(n42840), .Z(n40329) );
  XNOR U42278 ( .A(n35520), .B(n38502), .Z(n42840) );
  XOR U42279 ( .A(n42841), .B(n40122), .Z(n38502) );
  XOR U42280 ( .A(n42842), .B(n42843), .Z(n40122) );
  ANDN U42281 ( .B(n41785), .A(n42844), .Z(n42841) );
  XNOR U42282 ( .A(n42845), .B(n39568), .Z(n35520) );
  XOR U42283 ( .A(n42846), .B(n42847), .Z(n39568) );
  ANDN U42284 ( .B(n41787), .A(n42848), .Z(n42845) );
  XNOR U42285 ( .A(n39082), .B(n42849), .Z(n42839) );
  XOR U42286 ( .A(n37518), .B(n40440), .Z(n42849) );
  XOR U42287 ( .A(n42850), .B(n41616), .Z(n40440) );
  XOR U42288 ( .A(n42851), .B(n42852), .Z(n41616) );
  ANDN U42289 ( .B(n41794), .A(n42853), .Z(n42850) );
  XNOR U42290 ( .A(n42854), .B(n41942), .Z(n37518) );
  IV U42291 ( .A(n41791), .Z(n41942) );
  XOR U42292 ( .A(n42855), .B(n42856), .Z(n41791) );
  ANDN U42293 ( .B(n41792), .A(n42857), .Z(n42854) );
  XOR U42294 ( .A(n42858), .B(n39574), .Z(n39082) );
  XOR U42295 ( .A(n42859), .B(n42860), .Z(n39574) );
  ANDN U42296 ( .B(n41796), .A(n42861), .Z(n42858) );
  XOR U42297 ( .A(n42862), .B(n42863), .Z(n40349) );
  XOR U42298 ( .A(n37444), .B(n39639), .Z(n42863) );
  XNOR U42299 ( .A(n42864), .B(n41767), .Z(n39639) );
  ANDN U42300 ( .B(n41768), .A(n42865), .Z(n42864) );
  XNOR U42301 ( .A(n42866), .B(n41773), .Z(n37444) );
  XNOR U42302 ( .A(n42867), .B(n42868), .Z(n41773) );
  XNOR U42303 ( .A(n37016), .B(n42870), .Z(n42862) );
  XOR U42304 ( .A(n41758), .B(n38286), .Z(n42870) );
  XNOR U42305 ( .A(n42871), .B(n41781), .Z(n38286) );
  XOR U42306 ( .A(n42872), .B(n42873), .Z(n41781) );
  AND U42307 ( .A(n41780), .B(n42874), .Z(n42871) );
  XNOR U42308 ( .A(n42875), .B(n42041), .Z(n41758) );
  IV U42309 ( .A(n41777), .Z(n42041) );
  XOR U42310 ( .A(n42876), .B(n42877), .Z(n41777) );
  ANDN U42311 ( .B(n42878), .A(n41776), .Z(n42875) );
  IV U42312 ( .A(n42879), .Z(n41776) );
  XOR U42313 ( .A(n42880), .B(n41763), .Z(n37016) );
  XOR U42314 ( .A(n42881), .B(n42882), .Z(n41763) );
  AND U42315 ( .A(n41764), .B(n42883), .Z(n42880) );
  NOR U42316 ( .A(n36875), .B(n36874), .Z(n42837) );
  XNOR U42317 ( .A(n38851), .B(n41805), .Z(n36874) );
  XNOR U42318 ( .A(n42884), .B(n42832), .Z(n41805) );
  NOR U42319 ( .A(n40734), .B(n42885), .Z(n42884) );
  XNOR U42320 ( .A(n40433), .B(n42886), .Z(n38851) );
  XOR U42321 ( .A(n42887), .B(n42888), .Z(n40433) );
  XNOR U42322 ( .A(n35937), .B(n37722), .Z(n42888) );
  XNOR U42323 ( .A(n42889), .B(n42890), .Z(n37722) );
  ANDN U42324 ( .B(n41709), .A(n42891), .Z(n42889) );
  XOR U42325 ( .A(n42892), .B(n42893), .Z(n35937) );
  ANDN U42326 ( .B(n42894), .A(n42895), .Z(n42892) );
  XOR U42327 ( .A(n39650), .B(n42896), .Z(n42887) );
  XOR U42328 ( .A(n37966), .B(n39134), .Z(n42896) );
  XNOR U42329 ( .A(n42897), .B(n42898), .Z(n39134) );
  NOR U42330 ( .A(n41694), .B(n42899), .Z(n42897) );
  XNOR U42331 ( .A(n42900), .B(n41698), .Z(n37966) );
  ANDN U42332 ( .B(n42901), .A(n41699), .Z(n42900) );
  XNOR U42333 ( .A(n42902), .B(n41705), .Z(n39650) );
  ANDN U42334 ( .B(n42903), .A(n41704), .Z(n42902) );
  XOR U42335 ( .A(n42904), .B(n38151), .Z(n36875) );
  XNOR U42336 ( .A(n42905), .B(n42075), .Z(n38151) );
  XOR U42337 ( .A(n42906), .B(n42907), .Z(n42075) );
  XNOR U42338 ( .A(n37266), .B(n40188), .Z(n42907) );
  XNOR U42339 ( .A(n42908), .B(n41320), .Z(n40188) );
  ANDN U42340 ( .B(n42909), .A(n42910), .Z(n42908) );
  XNOR U42341 ( .A(n42911), .B(n41324), .Z(n37266) );
  NOR U42342 ( .A(n42912), .B(n42913), .Z(n42911) );
  XOR U42343 ( .A(n40334), .B(n42914), .Z(n42906) );
  XOR U42344 ( .A(n39008), .B(n37860), .Z(n42914) );
  XOR U42345 ( .A(n42915), .B(n42916), .Z(n37860) );
  ANDN U42346 ( .B(n42917), .A(n42918), .Z(n42915) );
  XOR U42347 ( .A(n42919), .B(n42920), .Z(n39008) );
  ANDN U42348 ( .B(n42921), .A(n42922), .Z(n42919) );
  XOR U42349 ( .A(n42923), .B(n41333), .Z(n40334) );
  XOR U42350 ( .A(n31122), .B(n42926), .Z(n42811) );
  XNOR U42351 ( .A(n38009), .B(n33030), .Z(n42926) );
  XNOR U42352 ( .A(n42927), .B(n36478), .Z(n33030) );
  XNOR U42353 ( .A(n42928), .B(n37349), .Z(n36478) );
  IV U42354 ( .A(n40005), .Z(n37349) );
  XOR U42355 ( .A(n42929), .B(n40529), .Z(n40005) );
  XNOR U42356 ( .A(n42930), .B(n42931), .Z(n40529) );
  XNOR U42357 ( .A(n42932), .B(n42933), .Z(n42931) );
  XOR U42358 ( .A(n42051), .B(n42934), .Z(n42930) );
  XNOR U42359 ( .A(n38615), .B(n38693), .Z(n42934) );
  XNOR U42360 ( .A(n42935), .B(n42936), .Z(n38693) );
  ANDN U42361 ( .B(n42937), .A(n42938), .Z(n42935) );
  XNOR U42362 ( .A(n42939), .B(n42940), .Z(n38615) );
  XOR U42363 ( .A(n42943), .B(n42944), .Z(n42051) );
  XNOR U42364 ( .A(n42947), .B(n37114), .Z(n36868) );
  XOR U42365 ( .A(n37720), .B(n42948), .Z(n36867) );
  XOR U42366 ( .A(n42949), .B(n42950), .Z(n42070) );
  XNOR U42367 ( .A(n39830), .B(n40576), .Z(n42950) );
  XOR U42368 ( .A(n42951), .B(n42952), .Z(n40576) );
  ANDN U42369 ( .B(n41212), .A(n42953), .Z(n42951) );
  XNOR U42370 ( .A(n42954), .B(n41992), .Z(n39830) );
  XOR U42371 ( .A(n42956), .B(n42957), .Z(n42949) );
  XOR U42372 ( .A(n39935), .B(n37673), .Z(n42957) );
  XNOR U42373 ( .A(n42958), .B(n41988), .Z(n37673) );
  NOR U42374 ( .A(n42959), .B(n41217), .Z(n42958) );
  XNOR U42375 ( .A(n42960), .B(n41983), .Z(n39935) );
  ANDN U42376 ( .B(n42961), .A(n42962), .Z(n42960) );
  XNOR U42377 ( .A(n42964), .B(n36465), .Z(n38009) );
  XNOR U42378 ( .A(n42965), .B(n37472), .Z(n36465) );
  ANDN U42379 ( .B(n36878), .A(n36879), .Z(n42964) );
  XOR U42380 ( .A(n42966), .B(n36522), .Z(n36879) );
  XOR U42381 ( .A(n42967), .B(n37543), .Z(n36878) );
  IV U42382 ( .A(n38419), .Z(n37543) );
  XOR U42383 ( .A(n42968), .B(n42969), .Z(n42804) );
  XNOR U42384 ( .A(n39260), .B(n37891), .Z(n42969) );
  XNOR U42385 ( .A(n42970), .B(n41002), .Z(n37891) );
  ANDN U42386 ( .B(n41003), .A(n42971), .Z(n42970) );
  XOR U42387 ( .A(n42972), .B(n41007), .Z(n39260) );
  ANDN U42388 ( .B(n42973), .A(n41006), .Z(n42972) );
  XOR U42389 ( .A(n39804), .B(n42974), .Z(n42968) );
  XOR U42390 ( .A(n40996), .B(n38144), .Z(n42974) );
  XNOR U42391 ( .A(n42975), .B(n41015), .Z(n38144) );
  ANDN U42392 ( .B(n41016), .A(n42976), .Z(n42975) );
  XNOR U42393 ( .A(n42977), .B(n41019), .Z(n40996) );
  ANDN U42394 ( .B(n42978), .A(n41020), .Z(n42977) );
  XNOR U42395 ( .A(n42979), .B(n41011), .Z(n39804) );
  XNOR U42396 ( .A(n42981), .B(n42982), .Z(n39744) );
  XNOR U42397 ( .A(n38644), .B(n38898), .Z(n42982) );
  XNOR U42398 ( .A(n42983), .B(n42984), .Z(n38898) );
  NOR U42399 ( .A(n42985), .B(n42986), .Z(n42983) );
  XNOR U42400 ( .A(n42987), .B(n42988), .Z(n38644) );
  NOR U42401 ( .A(n42989), .B(n42990), .Z(n42987) );
  XOR U42402 ( .A(n38780), .B(n42991), .Z(n42981) );
  XOR U42403 ( .A(n38244), .B(n37151), .Z(n42991) );
  XNOR U42404 ( .A(n42992), .B(n42993), .Z(n37151) );
  XNOR U42405 ( .A(n42996), .B(n42997), .Z(n38244) );
  ANDN U42406 ( .B(n42998), .A(n42999), .Z(n42996) );
  XNOR U42407 ( .A(n43000), .B(n43001), .Z(n38780) );
  NOR U42408 ( .A(n43002), .B(n43003), .Z(n43000) );
  XOR U42409 ( .A(n43004), .B(n36473), .Z(n31122) );
  XOR U42410 ( .A(n42357), .B(n39399), .Z(n36473) );
  XNOR U42411 ( .A(n43005), .B(n43006), .Z(n42357) );
  AND U42412 ( .A(n43007), .B(n43008), .Z(n43005) );
  ANDN U42413 ( .B(n36870), .A(n36871), .Z(n43004) );
  XOR U42414 ( .A(n40387), .B(n38360), .Z(n36871) );
  XOR U42415 ( .A(n41870), .B(n40096), .Z(n38360) );
  XNOR U42416 ( .A(n43009), .B(n43010), .Z(n40096) );
  XNOR U42417 ( .A(n39302), .B(n38168), .Z(n43010) );
  XNOR U42418 ( .A(n43011), .B(n43012), .Z(n38168) );
  ANDN U42419 ( .B(n42572), .A(n43013), .Z(n43011) );
  XNOR U42420 ( .A(n43014), .B(n43015), .Z(n39302) );
  ANDN U42421 ( .B(n40384), .A(n43016), .Z(n43014) );
  XNOR U42422 ( .A(n43017), .B(n43018), .Z(n43009) );
  XOR U42423 ( .A(n39808), .B(n39654), .Z(n43018) );
  XOR U42424 ( .A(n43019), .B(n43020), .Z(n39654) );
  ANDN U42425 ( .B(n40389), .A(n40391), .Z(n43019) );
  XNOR U42426 ( .A(n43021), .B(n43022), .Z(n39808) );
  AND U42427 ( .A(n43023), .B(n43024), .Z(n43021) );
  XOR U42428 ( .A(n43025), .B(n43026), .Z(n41870) );
  XNOR U42429 ( .A(n39128), .B(n39107), .Z(n43026) );
  XNOR U42430 ( .A(n43027), .B(n43028), .Z(n39107) );
  ANDN U42431 ( .B(n41867), .A(n41869), .Z(n43027) );
  XNOR U42432 ( .A(n43029), .B(n43030), .Z(n39128) );
  ANDN U42433 ( .B(n41256), .A(n41257), .Z(n43029) );
  XNOR U42434 ( .A(n40628), .B(n43031), .Z(n43025) );
  XOR U42435 ( .A(n35777), .B(n37606), .Z(n43031) );
  XNOR U42436 ( .A(n43032), .B(n43033), .Z(n37606) );
  ANDN U42437 ( .B(n41270), .A(n41272), .Z(n43032) );
  XNOR U42438 ( .A(n43034), .B(n43035), .Z(n35777) );
  ANDN U42439 ( .B(n41266), .A(n41267), .Z(n43034) );
  XOR U42440 ( .A(n43036), .B(n43037), .Z(n40628) );
  NOR U42441 ( .A(n41260), .B(n41261), .Z(n43036) );
  XNOR U42442 ( .A(n43038), .B(n43023), .Z(n40387) );
  NOR U42443 ( .A(n43024), .B(n43039), .Z(n43038) );
  XOR U42444 ( .A(n43040), .B(n38526), .Z(n36870) );
  XOR U42445 ( .A(n43041), .B(n43042), .Z(n38526) );
  XOR U42446 ( .A(n43043), .B(n43044), .Z(n35500) );
  XNOR U42447 ( .A(n31553), .B(n31777), .Z(n43044) );
  XOR U42448 ( .A(n35071), .B(n43045), .Z(n31777) );
  XOR U42449 ( .A(n43046), .B(n4407), .Z(n43045) );
  NOR U42450 ( .A(n36150), .B(n35072), .Z(n43046) );
  XNOR U42451 ( .A(n38507), .B(n43047), .Z(n35072) );
  XNOR U42452 ( .A(n43048), .B(n42531), .Z(n38507) );
  XNOR U42453 ( .A(n43049), .B(n43050), .Z(n42531) );
  XNOR U42454 ( .A(n39248), .B(n38802), .Z(n43050) );
  XNOR U42455 ( .A(n43051), .B(n43052), .Z(n38802) );
  NOR U42456 ( .A(n43053), .B(n42588), .Z(n43051) );
  XNOR U42457 ( .A(n43054), .B(n40265), .Z(n39248) );
  ANDN U42458 ( .B(n43055), .A(n40264), .Z(n43054) );
  XOR U42459 ( .A(n38605), .B(n43056), .Z(n43049) );
  XOR U42460 ( .A(n39757), .B(n39149), .Z(n43056) );
  XNOR U42461 ( .A(n43057), .B(n41498), .Z(n39149) );
  NOR U42462 ( .A(n41497), .B(n42579), .Z(n43057) );
  XNOR U42463 ( .A(n43058), .B(n40256), .Z(n39757) );
  XNOR U42464 ( .A(n43059), .B(n40260), .Z(n38605) );
  ANDN U42465 ( .B(n40261), .A(n42582), .Z(n43059) );
  XOR U42466 ( .A(n41122), .B(n38253), .Z(n36150) );
  XNOR U42467 ( .A(n43060), .B(n42275), .Z(n41122) );
  ANDN U42468 ( .B(n43061), .A(n43062), .Z(n43060) );
  XOR U42469 ( .A(n43063), .B(n42711), .Z(n35071) );
  XOR U42470 ( .A(n43064), .B(n35058), .Z(n31553) );
  XOR U42471 ( .A(n41413), .B(n39099), .Z(n35058) );
  NOR U42472 ( .A(n43067), .B(n43068), .Z(n43065) );
  ANDN U42473 ( .B(n35059), .A(n35574), .Z(n43064) );
  IV U42474 ( .A(n40041), .Z(n35574) );
  XOR U42475 ( .A(n43017), .B(n38169), .Z(n40041) );
  XNOR U42476 ( .A(n39767), .B(n40630), .Z(n38169) );
  XNOR U42477 ( .A(n43069), .B(n43070), .Z(n40630) );
  XNOR U42478 ( .A(n37781), .B(n39309), .Z(n43070) );
  XOR U42479 ( .A(n43071), .B(n43072), .Z(n39309) );
  NOR U42480 ( .A(n41270), .B(n43033), .Z(n43071) );
  XOR U42481 ( .A(n43073), .B(n43074), .Z(n41270) );
  XNOR U42482 ( .A(n43075), .B(n43076), .Z(n37781) );
  ANDN U42483 ( .B(n41260), .A(n43077), .Z(n43075) );
  XOR U42484 ( .A(n43078), .B(n43079), .Z(n41260) );
  XOR U42485 ( .A(n42533), .B(n43080), .Z(n43069) );
  XOR U42486 ( .A(n36412), .B(n38031), .Z(n43080) );
  XNOR U42487 ( .A(n43081), .B(n43082), .Z(n38031) );
  NOR U42488 ( .A(n43028), .B(n41867), .Z(n43081) );
  XOR U42489 ( .A(n43083), .B(n43084), .Z(n41867) );
  XNOR U42490 ( .A(n43085), .B(n43086), .Z(n36412) );
  NOR U42491 ( .A(n43030), .B(n41256), .Z(n43085) );
  XOR U42492 ( .A(n43087), .B(n43088), .Z(n41256) );
  XNOR U42493 ( .A(n43089), .B(n43090), .Z(n42533) );
  NOR U42494 ( .A(n41266), .B(n43035), .Z(n43089) );
  XNOR U42495 ( .A(n43091), .B(n43092), .Z(n41266) );
  XNOR U42496 ( .A(n43093), .B(n43094), .Z(n39767) );
  XNOR U42497 ( .A(n37103), .B(n37315), .Z(n43094) );
  XNOR U42498 ( .A(n43095), .B(n43096), .Z(n37315) );
  NOR U42499 ( .A(n43097), .B(n40389), .Z(n43095) );
  XNOR U42500 ( .A(n43098), .B(n42453), .Z(n40389) );
  XNOR U42501 ( .A(n43099), .B(n43100), .Z(n37103) );
  NOR U42502 ( .A(n42571), .B(n43012), .Z(n43099) );
  IV U42503 ( .A(n43013), .Z(n42571) );
  XOR U42504 ( .A(n43101), .B(n43102), .Z(n43013) );
  XOR U42505 ( .A(n37696), .B(n43103), .Z(n43093) );
  XOR U42506 ( .A(n40962), .B(n43104), .Z(n43103) );
  XNOR U42507 ( .A(n43105), .B(n43106), .Z(n40962) );
  NOR U42508 ( .A(n40383), .B(n43015), .Z(n43105) );
  IV U42509 ( .A(n43016), .Z(n40383) );
  XOR U42510 ( .A(n43107), .B(n43108), .Z(n43016) );
  XNOR U42511 ( .A(n43109), .B(n43110), .Z(n37696) );
  NOR U42512 ( .A(n43023), .B(n43022), .Z(n43109) );
  XOR U42513 ( .A(n43111), .B(n42691), .Z(n43023) );
  XNOR U42514 ( .A(n43112), .B(n43113), .Z(n43017) );
  NOR U42515 ( .A(n40394), .B(n40393), .Z(n43112) );
  XOR U42516 ( .A(n43114), .B(n36393), .Z(n35059) );
  XNOR U42517 ( .A(n43115), .B(n43116), .Z(n42236) );
  XOR U42518 ( .A(n40196), .B(n39522), .Z(n43116) );
  XNOR U42519 ( .A(n43117), .B(n43118), .Z(n39522) );
  NOR U42520 ( .A(n43119), .B(n43120), .Z(n43117) );
  XNOR U42521 ( .A(n43121), .B(n43122), .Z(n40196) );
  NOR U42522 ( .A(n42142), .B(n43123), .Z(n43121) );
  IV U42523 ( .A(n43124), .Z(n42142) );
  XOR U42524 ( .A(n41231), .B(n43125), .Z(n43115) );
  XOR U42525 ( .A(n40667), .B(n38254), .Z(n43125) );
  XOR U42526 ( .A(n43126), .B(n43127), .Z(n38254) );
  XOR U42527 ( .A(n43129), .B(n43130), .Z(n40667) );
  NOR U42528 ( .A(n42134), .B(n43131), .Z(n43129) );
  IV U42529 ( .A(n43132), .Z(n42134) );
  XNOR U42530 ( .A(n43133), .B(n43134), .Z(n41231) );
  NOR U42531 ( .A(n42129), .B(n43135), .Z(n43133) );
  XOR U42532 ( .A(n32549), .B(n43137), .Z(n43043) );
  XOR U42533 ( .A(n30242), .B(n30732), .Z(n43137) );
  XNOR U42534 ( .A(n43138), .B(n35064), .Z(n30732) );
  XOR U42535 ( .A(n39891), .B(n43139), .Z(n35064) );
  XNOR U42536 ( .A(n43140), .B(n43141), .Z(n39891) );
  NOR U42537 ( .A(n35571), .B(n35063), .Z(n43138) );
  XOR U42538 ( .A(n43142), .B(n39735), .Z(n35063) );
  IV U42539 ( .A(n35526), .Z(n39735) );
  XOR U42540 ( .A(n41150), .B(n39109), .Z(n35526) );
  XNOR U42541 ( .A(n43143), .B(n43144), .Z(n39109) );
  XNOR U42542 ( .A(n42388), .B(n39211), .Z(n43144) );
  XNOR U42543 ( .A(n43145), .B(n42100), .Z(n39211) );
  ANDN U42544 ( .B(n43146), .A(n43147), .Z(n43145) );
  XOR U42545 ( .A(n43148), .B(n42085), .Z(n42388) );
  ANDN U42546 ( .B(n43149), .A(n43150), .Z(n43148) );
  XOR U42547 ( .A(n40430), .B(n43151), .Z(n43143) );
  XOR U42548 ( .A(n43152), .B(n38243), .Z(n43151) );
  XNOR U42549 ( .A(n43153), .B(n43154), .Z(n38243) );
  ANDN U42550 ( .B(n43155), .A(n43156), .Z(n43153) );
  XNOR U42551 ( .A(n43157), .B(n42090), .Z(n40430) );
  XOR U42552 ( .A(n43160), .B(n43161), .Z(n41150) );
  XOR U42553 ( .A(n36447), .B(n41658), .Z(n43161) );
  XOR U42554 ( .A(n43162), .B(n43163), .Z(n41658) );
  NOR U42555 ( .A(n43164), .B(n43165), .Z(n43162) );
  XNOR U42556 ( .A(n43166), .B(n43167), .Z(n36447) );
  NOR U42557 ( .A(n43168), .B(n43169), .Z(n43166) );
  XOR U42558 ( .A(n38835), .B(n43170), .Z(n43160) );
  XOR U42559 ( .A(n35951), .B(n39463), .Z(n43170) );
  XNOR U42560 ( .A(n43171), .B(n43172), .Z(n39463) );
  ANDN U42561 ( .B(n43173), .A(n43174), .Z(n43171) );
  XNOR U42562 ( .A(n43175), .B(n43176), .Z(n35951) );
  ANDN U42563 ( .B(n43177), .A(n43178), .Z(n43175) );
  XNOR U42564 ( .A(n43179), .B(n43180), .Z(n38835) );
  NOR U42565 ( .A(n43181), .B(n43182), .Z(n43179) );
  IV U42566 ( .A(n42806), .Z(n35571) );
  XOR U42567 ( .A(n43183), .B(n38656), .Z(n42806) );
  IV U42568 ( .A(n39176), .Z(n38656) );
  XOR U42569 ( .A(n43184), .B(n42963), .Z(n39176) );
  XNOR U42570 ( .A(n43185), .B(n43186), .Z(n42963) );
  XNOR U42571 ( .A(n38872), .B(n43187), .Z(n43186) );
  XNOR U42572 ( .A(n43188), .B(n41974), .Z(n38872) );
  IV U42573 ( .A(n43189), .Z(n41974) );
  NOR U42574 ( .A(n43190), .B(n42043), .Z(n43188) );
  XNOR U42575 ( .A(n37629), .B(n43191), .Z(n43185) );
  XNOR U42576 ( .A(n39491), .B(n40797), .Z(n43191) );
  XNOR U42577 ( .A(n43192), .B(n41970), .Z(n40797) );
  IV U42578 ( .A(n43193), .Z(n41970) );
  NOR U42579 ( .A(n41205), .B(n43194), .Z(n43192) );
  XNOR U42580 ( .A(n43195), .B(n41977), .Z(n39491) );
  NOR U42581 ( .A(n43196), .B(n41191), .Z(n43195) );
  XNOR U42582 ( .A(n43197), .B(n41965), .Z(n37629) );
  ANDN U42583 ( .B(n43198), .A(n41195), .Z(n43197) );
  XNOR U42584 ( .A(n43199), .B(n35054), .Z(n30242) );
  XOR U42585 ( .A(n43200), .B(n36522), .Z(n35054) );
  IV U42586 ( .A(n39545), .Z(n36522) );
  XOR U42587 ( .A(n39794), .B(n38810), .Z(n39545) );
  XOR U42588 ( .A(n43201), .B(n43202), .Z(n38810) );
  XOR U42589 ( .A(n36214), .B(n39941), .Z(n43202) );
  XOR U42590 ( .A(n43203), .B(n43204), .Z(n39941) );
  XOR U42591 ( .A(n43206), .B(n43207), .Z(n36214) );
  ANDN U42592 ( .B(n43208), .A(n42753), .Z(n43206) );
  XNOR U42593 ( .A(n37682), .B(n43209), .Z(n43201) );
  XOR U42594 ( .A(n40358), .B(n43210), .Z(n43209) );
  XNOR U42595 ( .A(n43211), .B(n43212), .Z(n40358) );
  AND U42596 ( .A(n43213), .B(n42745), .Z(n43211) );
  XOR U42597 ( .A(n43214), .B(n43215), .Z(n37682) );
  XOR U42598 ( .A(n43217), .B(n43218), .Z(n39794) );
  XOR U42599 ( .A(n43219), .B(n39004), .Z(n43218) );
  XOR U42600 ( .A(n43220), .B(n43221), .Z(n39004) );
  ANDN U42601 ( .B(n42722), .A(n43222), .Z(n43220) );
  XOR U42602 ( .A(n36999), .B(n43223), .Z(n43217) );
  XOR U42603 ( .A(n39094), .B(n41711), .Z(n43223) );
  XNOR U42604 ( .A(n43224), .B(n43225), .Z(n41711) );
  ANDN U42605 ( .B(n42717), .A(n43226), .Z(n43224) );
  XNOR U42606 ( .A(n43227), .B(n43228), .Z(n39094) );
  NOR U42607 ( .A(n42726), .B(n43229), .Z(n43227) );
  IV U42608 ( .A(n43230), .Z(n42726) );
  XNOR U42609 ( .A(n43231), .B(n43232), .Z(n36999) );
  ANDN U42610 ( .B(n35055), .A(n36885), .Z(n43199) );
  IV U42611 ( .A(n37738), .Z(n36885) );
  XOR U42612 ( .A(n43235), .B(n37166), .Z(n37738) );
  IV U42613 ( .A(n38374), .Z(n37166) );
  XOR U42614 ( .A(n42648), .B(n41517), .Z(n38374) );
  XNOR U42615 ( .A(n43236), .B(n43237), .Z(n41517) );
  XNOR U42616 ( .A(n39265), .B(n38859), .Z(n43237) );
  XNOR U42617 ( .A(n43238), .B(n43007), .Z(n38859) );
  ANDN U42618 ( .B(n43239), .A(n43008), .Z(n43238) );
  XNOR U42619 ( .A(n43240), .B(n43241), .Z(n39265) );
  NOR U42620 ( .A(n43242), .B(n43243), .Z(n43240) );
  XOR U42621 ( .A(n42344), .B(n43244), .Z(n43236) );
  XOR U42622 ( .A(n39785), .B(n40672), .Z(n43244) );
  XNOR U42623 ( .A(n43245), .B(n42360), .Z(n40672) );
  NOR U42624 ( .A(n43246), .B(n42361), .Z(n43245) );
  XNOR U42625 ( .A(n43247), .B(n42349), .Z(n39785) );
  NOR U42626 ( .A(n42350), .B(n43248), .Z(n43247) );
  XNOR U42627 ( .A(n43249), .B(n42353), .Z(n42344) );
  NOR U42628 ( .A(n43250), .B(n42354), .Z(n43249) );
  XNOR U42629 ( .A(n43251), .B(n43252), .Z(n42648) );
  XNOR U42630 ( .A(n39548), .B(n39981), .Z(n43252) );
  XOR U42631 ( .A(n43253), .B(n40986), .Z(n39981) );
  NOR U42632 ( .A(n43254), .B(n43255), .Z(n43253) );
  XNOR U42633 ( .A(n43256), .B(n43257), .Z(n39548) );
  NOR U42634 ( .A(n43258), .B(n43259), .Z(n43256) );
  XNOR U42635 ( .A(n39580), .B(n43260), .Z(n43251) );
  XOR U42636 ( .A(n37269), .B(n39984), .Z(n43260) );
  XNOR U42637 ( .A(n43261), .B(n40981), .Z(n39984) );
  ANDN U42638 ( .B(n43262), .A(n43263), .Z(n43261) );
  XNOR U42639 ( .A(n43264), .B(n41363), .Z(n37269) );
  XOR U42640 ( .A(n43267), .B(n40991), .Z(n39580) );
  IV U42641 ( .A(n43268), .Z(n40991) );
  NOR U42642 ( .A(n43269), .B(n43270), .Z(n43267) );
  XOR U42643 ( .A(n40657), .B(n43271), .Z(n35055) );
  XNOR U42644 ( .A(n43272), .B(n35068), .Z(n32549) );
  XNOR U42645 ( .A(n38719), .B(n43273), .Z(n35068) );
  XNOR U42646 ( .A(n39766), .B(n43274), .Z(n38719) );
  XOR U42647 ( .A(n43275), .B(n43276), .Z(n39766) );
  XOR U42648 ( .A(n42591), .B(n37486), .Z(n43276) );
  XOR U42649 ( .A(n43277), .B(n42600), .Z(n37486) );
  NOR U42650 ( .A(n43278), .B(n40231), .Z(n43277) );
  XOR U42651 ( .A(n43279), .B(n43280), .Z(n40231) );
  XNOR U42652 ( .A(n43281), .B(n42609), .Z(n42591) );
  ANDN U42653 ( .B(n40240), .A(n40242), .Z(n43281) );
  XOR U42654 ( .A(n43282), .B(n43283), .Z(n40240) );
  XOR U42655 ( .A(n40344), .B(n43284), .Z(n43275) );
  XNOR U42656 ( .A(n34367), .B(n36709), .Z(n43284) );
  XOR U42657 ( .A(n43285), .B(n42605), .Z(n36709) );
  ANDN U42658 ( .B(n40246), .A(n42606), .Z(n43285) );
  XOR U42659 ( .A(n43286), .B(n43287), .Z(n42606) );
  XNOR U42660 ( .A(n43288), .B(n43289), .Z(n34367) );
  NOR U42661 ( .A(n40236), .B(n40238), .Z(n43288) );
  XNOR U42662 ( .A(n43290), .B(n42597), .Z(n40344) );
  ANDN U42663 ( .B(n40227), .A(n43291), .Z(n43290) );
  XNOR U42664 ( .A(n43292), .B(n43108), .Z(n40227) );
  NOR U42665 ( .A(n35566), .B(n35067), .Z(n43272) );
  XOR U42666 ( .A(n40177), .B(n39227), .Z(n35067) );
  IV U42667 ( .A(n36439), .Z(n39227) );
  XOR U42668 ( .A(n38435), .B(n40662), .Z(n36439) );
  XNOR U42669 ( .A(n43293), .B(n43294), .Z(n40662) );
  XNOR U42670 ( .A(n38902), .B(n37329), .Z(n43294) );
  XNOR U42671 ( .A(n43295), .B(n43296), .Z(n37329) );
  ANDN U42672 ( .B(n40762), .A(n43297), .Z(n43295) );
  XOR U42673 ( .A(n43298), .B(n43299), .Z(n40762) );
  XNOR U42674 ( .A(n43300), .B(n43301), .Z(n38902) );
  AND U42675 ( .A(n41487), .B(n40768), .Z(n43300) );
  XOR U42676 ( .A(n43302), .B(n43303), .Z(n40768) );
  XOR U42677 ( .A(n37865), .B(n43304), .Z(n43293) );
  XOR U42678 ( .A(n39324), .B(n43305), .Z(n43304) );
  XNOR U42679 ( .A(n43306), .B(n43307), .Z(n39324) );
  ANDN U42680 ( .B(n40772), .A(n41482), .Z(n43306) );
  XNOR U42681 ( .A(n43308), .B(n41745), .Z(n40772) );
  XNOR U42682 ( .A(n43309), .B(n43310), .Z(n37865) );
  ANDN U42683 ( .B(n41479), .A(n41478), .Z(n43309) );
  XOR U42684 ( .A(n43311), .B(n43312), .Z(n41479) );
  XOR U42685 ( .A(n43313), .B(n43314), .Z(n38435) );
  XNOR U42686 ( .A(n38095), .B(n39671), .Z(n43314) );
  XOR U42687 ( .A(n43315), .B(n41724), .Z(n39671) );
  XOR U42688 ( .A(n43316), .B(n42206), .Z(n41724) );
  ANDN U42689 ( .B(n40787), .A(n41723), .Z(n43315) );
  XNOR U42690 ( .A(n43317), .B(n41425), .Z(n38095) );
  XOR U42691 ( .A(n43318), .B(n43319), .Z(n41425) );
  XOR U42692 ( .A(n43320), .B(n43321), .Z(n40183) );
  XOR U42693 ( .A(n43322), .B(n43323), .Z(n40185) );
  XOR U42694 ( .A(n40467), .B(n43324), .Z(n43313) );
  XOR U42695 ( .A(n38577), .B(n39138), .Z(n43324) );
  XNOR U42696 ( .A(n43325), .B(n41427), .Z(n39138) );
  XNOR U42697 ( .A(n43326), .B(n43327), .Z(n41427) );
  NOR U42698 ( .A(n40180), .B(n40179), .Z(n43325) );
  XNOR U42699 ( .A(n43328), .B(n43329), .Z(n40179) );
  XOR U42700 ( .A(n43330), .B(n43331), .Z(n40180) );
  XNOR U42701 ( .A(n43332), .B(n41434), .Z(n38577) );
  XOR U42702 ( .A(n42540), .B(n43333), .Z(n41434) );
  ANDN U42703 ( .B(n40171), .A(n40169), .Z(n43332) );
  XOR U42704 ( .A(n43334), .B(n43335), .Z(n40169) );
  XNOR U42705 ( .A(n43336), .B(n43337), .Z(n40171) );
  XNOR U42706 ( .A(n43338), .B(n41431), .Z(n40467) );
  XOR U42707 ( .A(n43339), .B(n42672), .Z(n41431) );
  ANDN U42708 ( .B(n40175), .A(n41432), .Z(n43338) );
  XOR U42709 ( .A(n43340), .B(n43341), .Z(n41432) );
  XNOR U42710 ( .A(n43342), .B(n43343), .Z(n40175) );
  XOR U42711 ( .A(n43344), .B(n41723), .Z(n40177) );
  NOR U42712 ( .A(n40788), .B(n40787), .Z(n43344) );
  XNOR U42713 ( .A(n43347), .B(n42501), .Z(n40787) );
  XOR U42714 ( .A(n43348), .B(n40853), .Z(n40788) );
  IV U42715 ( .A(n37734), .Z(n35566) );
  XOR U42716 ( .A(n43349), .B(n36202), .Z(n37734) );
  XNOR U42717 ( .A(n42423), .B(n42553), .Z(n36202) );
  XOR U42718 ( .A(n43350), .B(n43351), .Z(n42553) );
  XOR U42719 ( .A(n40656), .B(n39062), .Z(n43351) );
  XNOR U42720 ( .A(n43352), .B(n43353), .Z(n39062) );
  ANDN U42721 ( .B(n43354), .A(n43355), .Z(n43352) );
  XNOR U42722 ( .A(n43356), .B(n43357), .Z(n40656) );
  ANDN U42723 ( .B(n43358), .A(n43359), .Z(n43356) );
  XNOR U42724 ( .A(n41917), .B(n43360), .Z(n43350) );
  XOR U42725 ( .A(n39975), .B(n35365), .Z(n43360) );
  XNOR U42726 ( .A(n43361), .B(n42941), .Z(n35365) );
  ANDN U42727 ( .B(n43362), .A(n43363), .Z(n43361) );
  XNOR U42728 ( .A(n43364), .B(n42945), .Z(n39975) );
  ANDN U42729 ( .B(n43368), .A(n43369), .Z(n43367) );
  XOR U42730 ( .A(n43370), .B(n43371), .Z(n42423) );
  XNOR U42731 ( .A(n39331), .B(n38250), .Z(n43371) );
  XOR U42732 ( .A(n43372), .B(n43373), .Z(n38250) );
  NOR U42733 ( .A(n43374), .B(n42186), .Z(n43372) );
  XOR U42734 ( .A(n43375), .B(n43376), .Z(n39331) );
  ANDN U42735 ( .B(n43377), .A(n40958), .Z(n43375) );
  IV U42736 ( .A(n43378), .Z(n40958) );
  XOR U42737 ( .A(n38370), .B(n43379), .Z(n43370) );
  XOR U42738 ( .A(n37426), .B(n43380), .Z(n43379) );
  XNOR U42739 ( .A(n43381), .B(n43382), .Z(n37426) );
  ANDN U42740 ( .B(n43383), .A(n43384), .Z(n43381) );
  XNOR U42741 ( .A(n43385), .B(n43386), .Z(n38370) );
  XOR U42742 ( .A(n32362), .B(n38204), .Z(n28981) );
  XNOR U42743 ( .A(n43388), .B(n38476), .Z(n38204) );
  ANDN U42744 ( .B(n38916), .A(n43389), .Z(n43388) );
  IV U42745 ( .A(n36090), .Z(n38916) );
  XOR U42746 ( .A(n43390), .B(n37011), .Z(n36090) );
  XOR U42747 ( .A(n33771), .B(n36797), .Z(n32362) );
  XNOR U42748 ( .A(n43391), .B(n43392), .Z(n36797) );
  XNOR U42749 ( .A(n32610), .B(n32258), .Z(n43392) );
  XNOR U42750 ( .A(n43393), .B(n39683), .Z(n32258) );
  IV U42751 ( .A(n37399), .Z(n39683) );
  XOR U42752 ( .A(n41377), .B(n37099), .Z(n37399) );
  IV U42753 ( .A(n36351), .Z(n37099) );
  XOR U42754 ( .A(n41660), .B(n43394), .Z(n36351) );
  XOR U42755 ( .A(n43395), .B(n43396), .Z(n41660) );
  XNOR U42756 ( .A(n41062), .B(n42646), .Z(n43396) );
  XNOR U42757 ( .A(n43397), .B(n43398), .Z(n42646) );
  AND U42758 ( .A(n43399), .B(n43400), .Z(n43397) );
  XNOR U42759 ( .A(n43401), .B(n43402), .Z(n41062) );
  ANDN U42760 ( .B(n41379), .A(n41380), .Z(n43401) );
  XOR U42761 ( .A(n38147), .B(n43403), .Z(n43395) );
  XNOR U42762 ( .A(n39783), .B(n40144), .Z(n43403) );
  XNOR U42763 ( .A(n43404), .B(n43405), .Z(n40144) );
  ANDN U42764 ( .B(n41388), .A(n41389), .Z(n43404) );
  XOR U42765 ( .A(n43406), .B(n43407), .Z(n39783) );
  AND U42766 ( .A(n41384), .B(n41385), .Z(n43406) );
  XNOR U42767 ( .A(n43408), .B(n43409), .Z(n38147) );
  ANDN U42768 ( .B(n41392), .A(n41393), .Z(n43408) );
  XNOR U42769 ( .A(n43410), .B(n43399), .Z(n41377) );
  NOR U42770 ( .A(n43400), .B(n43411), .Z(n43410) );
  ANDN U42771 ( .B(n36109), .A(n37398), .Z(n43393) );
  XOR U42772 ( .A(n35943), .B(n43412), .Z(n37398) );
  XNOR U42773 ( .A(n41454), .B(n40829), .Z(n35943) );
  XNOR U42774 ( .A(n43413), .B(n43414), .Z(n40829) );
  XNOR U42775 ( .A(n39083), .B(n39297), .Z(n43414) );
  XOR U42776 ( .A(n43415), .B(n43416), .Z(n39297) );
  ANDN U42777 ( .B(n43417), .A(n43418), .Z(n43415) );
  XNOR U42778 ( .A(n43419), .B(n43420), .Z(n39083) );
  ANDN U42779 ( .B(n43421), .A(n43422), .Z(n43419) );
  XOR U42780 ( .A(n39032), .B(n43423), .Z(n43413) );
  XNOR U42781 ( .A(n39041), .B(n37432), .Z(n43423) );
  XNOR U42782 ( .A(n43424), .B(n43425), .Z(n37432) );
  ANDN U42783 ( .B(n43426), .A(n43427), .Z(n43424) );
  XNOR U42784 ( .A(n43428), .B(n43429), .Z(n39041) );
  ANDN U42785 ( .B(n43430), .A(n43431), .Z(n43428) );
  XNOR U42786 ( .A(n43432), .B(n43433), .Z(n39032) );
  ANDN U42787 ( .B(n43434), .A(n43435), .Z(n43432) );
  XOR U42788 ( .A(n43436), .B(n43437), .Z(n41454) );
  XOR U42789 ( .A(n37186), .B(n40466), .Z(n43437) );
  XOR U42790 ( .A(n43438), .B(n42001), .Z(n40466) );
  NOR U42791 ( .A(n42000), .B(n43439), .Z(n43438) );
  XNOR U42792 ( .A(n43440), .B(n41164), .Z(n37186) );
  ANDN U42793 ( .B(n43441), .A(n43442), .Z(n43440) );
  XOR U42794 ( .A(n41158), .B(n43443), .Z(n43436) );
  XOR U42795 ( .A(n37502), .B(n38966), .Z(n43443) );
  XNOR U42796 ( .A(n43444), .B(n41168), .Z(n38966) );
  ANDN U42797 ( .B(n41169), .A(n43445), .Z(n43444) );
  XNOR U42798 ( .A(n43446), .B(n41179), .Z(n37502) );
  NOR U42799 ( .A(n41178), .B(n43447), .Z(n43446) );
  XNOR U42800 ( .A(n43448), .B(n41174), .Z(n41158) );
  ANDN U42801 ( .B(n43449), .A(n43450), .Z(n43448) );
  XOR U42802 ( .A(n43451), .B(n37258), .Z(n36109) );
  XOR U42803 ( .A(n43453), .B(n43454), .Z(n38982) );
  XNOR U42804 ( .A(n38992), .B(n38309), .Z(n43454) );
  XOR U42805 ( .A(n43455), .B(n41699), .Z(n38309) );
  XOR U42806 ( .A(n43456), .B(n43457), .Z(n41699) );
  ANDN U42807 ( .B(n43458), .A(n42901), .Z(n43455) );
  XNOR U42808 ( .A(n43459), .B(n42894), .Z(n38992) );
  AND U42809 ( .A(n42895), .B(n43460), .Z(n43459) );
  XNOR U42810 ( .A(n40432), .B(n43461), .Z(n43453) );
  XOR U42811 ( .A(n39301), .B(n35626), .Z(n43461) );
  XNOR U42812 ( .A(n43462), .B(n41709), .Z(n35626) );
  XOR U42813 ( .A(n43463), .B(n43464), .Z(n41709) );
  ANDN U42814 ( .B(n42891), .A(n43465), .Z(n43462) );
  XOR U42815 ( .A(n43466), .B(n41694), .Z(n39301) );
  XOR U42816 ( .A(n43467), .B(n43468), .Z(n41694) );
  ANDN U42817 ( .B(n42899), .A(n43469), .Z(n43466) );
  XNOR U42818 ( .A(n43470), .B(n41704), .Z(n40432) );
  XOR U42819 ( .A(n43471), .B(n43472), .Z(n41704) );
  XNOR U42820 ( .A(n43474), .B(n39687), .Z(n32610) );
  IV U42821 ( .A(n37395), .Z(n39687) );
  XOR U42822 ( .A(n40955), .B(n37868), .Z(n37395) );
  XNOR U42823 ( .A(n43477), .B(n43384), .Z(n40955) );
  ANDN U42824 ( .B(n43478), .A(n43479), .Z(n43477) );
  ANDN U42825 ( .B(n36105), .A(n37394), .Z(n43474) );
  XOR U42826 ( .A(n38131), .B(n40934), .Z(n37394) );
  XNOR U42827 ( .A(n43480), .B(n43481), .Z(n40934) );
  ANDN U42828 ( .B(n43482), .A(n40864), .Z(n43480) );
  IV U42829 ( .A(n41606), .Z(n38131) );
  XOR U42830 ( .A(n43483), .B(n39180), .Z(n41606) );
  XNOR U42831 ( .A(n43484), .B(n43485), .Z(n39180) );
  XOR U42832 ( .A(n43486), .B(n39246), .Z(n43485) );
  XOR U42833 ( .A(n43487), .B(n43488), .Z(n39246) );
  ANDN U42834 ( .B(n41608), .A(n41609), .Z(n43487) );
  XOR U42835 ( .A(n37953), .B(n43489), .Z(n43484) );
  XOR U42836 ( .A(n38927), .B(n43490), .Z(n43489) );
  XNOR U42837 ( .A(n43491), .B(n41549), .Z(n38927) );
  NOR U42838 ( .A(n40938), .B(n40939), .Z(n43491) );
  XNOR U42839 ( .A(n43492), .B(n40872), .Z(n37953) );
  IV U42840 ( .A(n43493), .Z(n40872) );
  ANDN U42841 ( .B(n40928), .A(n40929), .Z(n43492) );
  XOR U42842 ( .A(n31257), .B(n43495), .Z(n43391) );
  XOR U42843 ( .A(n37389), .B(n31228), .Z(n43495) );
  XNOR U42844 ( .A(n43496), .B(n39705), .Z(n31228) );
  IV U42845 ( .A(n39753), .Z(n39705) );
  XOR U42846 ( .A(n38959), .B(n43497), .Z(n39753) );
  XOR U42847 ( .A(n42905), .B(n43498), .Z(n38959) );
  XOR U42848 ( .A(n43499), .B(n43500), .Z(n42905) );
  XOR U42849 ( .A(n40522), .B(n38392), .Z(n43500) );
  XOR U42850 ( .A(n43501), .B(n39514), .Z(n38392) );
  NOR U42851 ( .A(n43502), .B(n43503), .Z(n43501) );
  XNOR U42852 ( .A(n43504), .B(n39510), .Z(n40522) );
  NOR U42853 ( .A(n43505), .B(n43506), .Z(n43504) );
  XOR U42854 ( .A(n37879), .B(n43507), .Z(n43499) );
  XOR U42855 ( .A(n38170), .B(n43508), .Z(n43507) );
  XNOR U42856 ( .A(n43509), .B(n40364), .Z(n38170) );
  NOR U42857 ( .A(n43510), .B(n43511), .Z(n43509) );
  XNOR U42858 ( .A(n43512), .B(n39501), .Z(n37879) );
  NOR U42859 ( .A(n43513), .B(n43514), .Z(n43512) );
  ANDN U42860 ( .B(n36100), .A(n38223), .Z(n43496) );
  XNOR U42861 ( .A(n42248), .B(n43515), .Z(n38223) );
  XNOR U42862 ( .A(n43516), .B(n43517), .Z(n42248) );
  XOR U42863 ( .A(n42023), .B(n37535), .Z(n36100) );
  XNOR U42864 ( .A(n40339), .B(n42054), .Z(n37535) );
  XNOR U42865 ( .A(n43520), .B(n43521), .Z(n42054) );
  XNOR U42866 ( .A(n37504), .B(n39991), .Z(n43521) );
  XOR U42867 ( .A(n43522), .B(n41824), .Z(n39991) );
  XOR U42868 ( .A(n43523), .B(n43524), .Z(n41823) );
  XNOR U42869 ( .A(n43525), .B(n41827), .Z(n37504) );
  XOR U42870 ( .A(n38101), .B(n43527), .Z(n43520) );
  XOR U42871 ( .A(n41802), .B(n39414), .Z(n43527) );
  XOR U42872 ( .A(n43528), .B(n41834), .Z(n39414) );
  ANDN U42873 ( .B(n41833), .A(n42016), .Z(n43528) );
  XNOR U42874 ( .A(n43529), .B(n43530), .Z(n41833) );
  XOR U42875 ( .A(n43531), .B(n43532), .Z(n41802) );
  XOR U42876 ( .A(n43533), .B(n41838), .Z(n38101) );
  ANDN U42877 ( .B(n41837), .A(n42019), .Z(n43533) );
  XNOR U42878 ( .A(n43534), .B(n43535), .Z(n41837) );
  XNOR U42879 ( .A(n43536), .B(n43537), .Z(n40339) );
  XNOR U42880 ( .A(n37303), .B(n38980), .Z(n43537) );
  XOR U42881 ( .A(n43538), .B(n41808), .Z(n38980) );
  ANDN U42882 ( .B(n40747), .A(n40749), .Z(n43538) );
  XOR U42883 ( .A(n43539), .B(n43540), .Z(n40749) );
  XNOR U42884 ( .A(n43541), .B(n41649), .Z(n40747) );
  XOR U42885 ( .A(n43542), .B(n42885), .Z(n37303) );
  ANDN U42886 ( .B(n40734), .A(n40735), .Z(n43542) );
  XNOR U42887 ( .A(n43543), .B(n43544), .Z(n40735) );
  XOR U42888 ( .A(n43545), .B(n43546), .Z(n40734) );
  XOR U42889 ( .A(n35319), .B(n43547), .Z(n43536) );
  XOR U42890 ( .A(n37793), .B(n37041), .Z(n43547) );
  XNOR U42891 ( .A(n43548), .B(n41818), .Z(n37041) );
  ANDN U42892 ( .B(n40738), .A(n40740), .Z(n43548) );
  XNOR U42893 ( .A(n43549), .B(n43550), .Z(n40740) );
  XNOR U42894 ( .A(n43551), .B(n43552), .Z(n40738) );
  XNOR U42895 ( .A(n43553), .B(n41815), .Z(n37793) );
  XOR U42896 ( .A(n43554), .B(n43555), .Z(n40744) );
  XOR U42897 ( .A(n43556), .B(n43557), .Z(n40743) );
  XOR U42898 ( .A(n43558), .B(n41812), .Z(n35319) );
  XNOR U42899 ( .A(n43559), .B(n43560), .Z(n40752) );
  XOR U42900 ( .A(n43561), .B(n43562), .Z(n40751) );
  XOR U42901 ( .A(n43563), .B(n41828), .Z(n42023) );
  XNOR U42902 ( .A(n43564), .B(n43565), .Z(n41828) );
  ANDN U42903 ( .B(n43526), .A(n43566), .Z(n43563) );
  XNOR U42904 ( .A(n43567), .B(n39697), .Z(n37389) );
  IV U42905 ( .A(n37402), .Z(n39697) );
  XOR U42906 ( .A(n43568), .B(n35311), .Z(n37402) );
  XOR U42907 ( .A(n39887), .B(n43569), .Z(n35311) );
  XOR U42908 ( .A(n43570), .B(n43571), .Z(n39887) );
  XOR U42909 ( .A(n39442), .B(n38089), .Z(n43571) );
  XNOR U42910 ( .A(n43572), .B(n41620), .Z(n38089) );
  XOR U42911 ( .A(n43575), .B(n43576), .Z(n41621) );
  XOR U42912 ( .A(n43577), .B(n43578), .Z(n42173) );
  XNOR U42913 ( .A(n43579), .B(n41469), .Z(n39442) );
  XOR U42914 ( .A(n43580), .B(n43581), .Z(n41469) );
  ANDN U42915 ( .B(n41470), .A(n42181), .Z(n43579) );
  XOR U42916 ( .A(n43582), .B(n43583), .Z(n42181) );
  XOR U42917 ( .A(n43584), .B(n43073), .Z(n41470) );
  XNOR U42918 ( .A(n41023), .B(n43585), .Z(n43570) );
  XOR U42919 ( .A(n37007), .B(n38991), .Z(n43585) );
  XNOR U42920 ( .A(n43586), .B(n41473), .Z(n38991) );
  XOR U42921 ( .A(n43587), .B(n43588), .Z(n41473) );
  ANDN U42922 ( .B(n41474), .A(n42183), .Z(n43586) );
  XOR U42923 ( .A(n43590), .B(n43591), .Z(n41474) );
  XOR U42924 ( .A(n43592), .B(n41464), .Z(n37007) );
  XOR U42925 ( .A(n43593), .B(n43594), .Z(n41464) );
  ANDN U42926 ( .B(n41463), .A(n42178), .Z(n43592) );
  XNOR U42927 ( .A(n43595), .B(n43596), .Z(n42178) );
  XNOR U42928 ( .A(n43599), .B(n41459), .Z(n41023) );
  XOR U42929 ( .A(n43600), .B(n43601), .Z(n41459) );
  ANDN U42930 ( .B(n41460), .A(n42175), .Z(n43599) );
  XNOR U42931 ( .A(n43602), .B(n43603), .Z(n42175) );
  XOR U42932 ( .A(n43604), .B(n43605), .Z(n41460) );
  NOR U42933 ( .A(n37401), .B(n36113), .Z(n43567) );
  XNOR U42934 ( .A(n40252), .B(n36308), .Z(n36113) );
  XNOR U42935 ( .A(n43606), .B(n43607), .Z(n40616) );
  XNOR U42936 ( .A(n39012), .B(n39214), .Z(n43607) );
  XNOR U42937 ( .A(n43608), .B(n43609), .Z(n39214) );
  ANDN U42938 ( .B(n41532), .A(n43610), .Z(n43608) );
  XNOR U42939 ( .A(n43611), .B(n43612), .Z(n39012) );
  ANDN U42940 ( .B(n41527), .A(n41528), .Z(n43611) );
  XOR U42941 ( .A(n39272), .B(n43613), .Z(n43606) );
  XOR U42942 ( .A(n40527), .B(n43614), .Z(n43613) );
  XOR U42943 ( .A(n43615), .B(n43616), .Z(n40527) );
  NOR U42944 ( .A(n41540), .B(n41541), .Z(n43615) );
  XNOR U42945 ( .A(n43617), .B(n43618), .Z(n39272) );
  ANDN U42946 ( .B(n41536), .A(n41537), .Z(n43617) );
  XOR U42947 ( .A(n43620), .B(n42590), .Z(n40252) );
  ANDN U42948 ( .B(n43052), .A(n43621), .Z(n43620) );
  XOR U42949 ( .A(n39936), .B(n42956), .Z(n37401) );
  XNOR U42950 ( .A(n43622), .B(n41990), .Z(n42956) );
  ANDN U42951 ( .B(n43623), .A(n43624), .Z(n43622) );
  XOR U42952 ( .A(n43625), .B(n43626), .Z(n39936) );
  XNOR U42953 ( .A(n43627), .B(n39693), .Z(n31257) );
  IV U42954 ( .A(n37405), .Z(n39693) );
  XOR U42955 ( .A(n43210), .B(n37683), .Z(n37405) );
  XNOR U42956 ( .A(n41063), .B(n43628), .Z(n37683) );
  XOR U42957 ( .A(n43629), .B(n43630), .Z(n41063) );
  XNOR U42958 ( .A(n39662), .B(n39388), .Z(n43630) );
  XOR U42959 ( .A(n43631), .B(n42754), .Z(n39388) );
  NOR U42960 ( .A(n43208), .B(n43207), .Z(n43631) );
  XNOR U42961 ( .A(n43632), .B(n42742), .Z(n39662) );
  ANDN U42962 ( .B(n43204), .A(n43205), .Z(n43632) );
  XOR U42963 ( .A(n40140), .B(n43633), .Z(n43629) );
  XOR U42964 ( .A(n40613), .B(n43634), .Z(n43633) );
  XNOR U42965 ( .A(n43635), .B(n42747), .Z(n40613) );
  ANDN U42966 ( .B(n43212), .A(n43213), .Z(n43635) );
  XNOR U42967 ( .A(n43636), .B(n42738), .Z(n40140) );
  ANDN U42968 ( .B(n43215), .A(n43216), .Z(n43636) );
  XOR U42969 ( .A(n43637), .B(n43638), .Z(n43210) );
  ANDN U42970 ( .B(n43639), .A(n42749), .Z(n43637) );
  ANDN U42971 ( .B(n36096), .A(n37404), .Z(n43627) );
  XNOR U42972 ( .A(n42701), .B(n37005), .Z(n37404) );
  XNOR U42973 ( .A(n41040), .B(n42824), .Z(n37005) );
  XNOR U42974 ( .A(n43640), .B(n43641), .Z(n42824) );
  XNOR U42975 ( .A(n34636), .B(n37842), .Z(n43641) );
  XNOR U42976 ( .A(n43642), .B(n43526), .Z(n37842) );
  ANDN U42977 ( .B(n43566), .A(n41826), .Z(n43642) );
  XNOR U42978 ( .A(n43645), .B(n42019), .Z(n34636) );
  XOR U42979 ( .A(n43646), .B(n43647), .Z(n42019) );
  ANDN U42980 ( .B(n42020), .A(n41836), .Z(n43645) );
  XOR U42981 ( .A(n39864), .B(n43648), .Z(n43640) );
  XOR U42982 ( .A(n40130), .B(n37790), .Z(n43648) );
  XNOR U42983 ( .A(n43649), .B(n42025), .Z(n37790) );
  XOR U42984 ( .A(n42517), .B(n43650), .Z(n42025) );
  ANDN U42985 ( .B(n42026), .A(n41822), .Z(n43649) );
  XNOR U42986 ( .A(n43651), .B(n42809), .Z(n40130) );
  XOR U42987 ( .A(n43590), .B(n43652), .Z(n42809) );
  ANDN U42988 ( .B(n42810), .A(n43653), .Z(n43651) );
  XNOR U42989 ( .A(n43654), .B(n42016), .Z(n39864) );
  XOR U42990 ( .A(n43655), .B(n43656), .Z(n42016) );
  ANDN U42991 ( .B(n42017), .A(n41832), .Z(n43654) );
  XNOR U42992 ( .A(n43657), .B(n43658), .Z(n41040) );
  XOR U42993 ( .A(n39405), .B(n41840), .Z(n43658) );
  XOR U42994 ( .A(n43659), .B(n43660), .Z(n41840) );
  NOR U42995 ( .A(n42705), .B(n42706), .Z(n43659) );
  XNOR U42996 ( .A(n43661), .B(n43662), .Z(n42706) );
  XNOR U42997 ( .A(n43663), .B(n43664), .Z(n39405) );
  ANDN U42998 ( .B(n41853), .A(n42699), .Z(n43663) );
  XOR U42999 ( .A(n43665), .B(n43666), .Z(n41853) );
  XOR U43000 ( .A(n40825), .B(n43667), .Z(n43657) );
  XOR U43001 ( .A(n42011), .B(n39266), .Z(n43667) );
  ANDN U43002 ( .B(n42697), .A(n41857), .Z(n43668) );
  XNOR U43003 ( .A(n43672), .B(n43673), .Z(n42011) );
  ANDN U43004 ( .B(n43674), .A(n42467), .Z(n43672) );
  XNOR U43005 ( .A(n43675), .B(n43676), .Z(n40825) );
  AND U43006 ( .A(n42703), .B(n41849), .Z(n43675) );
  XNOR U43007 ( .A(n42510), .B(n43677), .Z(n41849) );
  XNOR U43008 ( .A(n43678), .B(n43674), .Z(n42701) );
  AND U43009 ( .A(n42467), .B(n42469), .Z(n43678) );
  XNOR U43010 ( .A(n43679), .B(n43680), .Z(n42467) );
  XOR U43011 ( .A(n43681), .B(n35611), .Z(n36096) );
  XOR U43012 ( .A(n43682), .B(n43683), .Z(n33771) );
  XOR U43013 ( .A(n33176), .B(n35394), .Z(n43683) );
  XOR U43014 ( .A(n43684), .B(n34764), .Z(n35394) );
  XNOR U43015 ( .A(n43152), .B(n38242), .Z(n34764) );
  XOR U43016 ( .A(n41659), .B(n43685), .Z(n38242) );
  XOR U43017 ( .A(n43686), .B(n43687), .Z(n41659) );
  XNOR U43018 ( .A(n37913), .B(n43688), .Z(n43687) );
  XOR U43019 ( .A(n43689), .B(n43690), .Z(n37913) );
  XNOR U43020 ( .A(n38453), .B(n43691), .Z(n43686) );
  XOR U43021 ( .A(n39917), .B(n41800), .Z(n43691) );
  XOR U43022 ( .A(n43692), .B(n43693), .Z(n41800) );
  ANDN U43023 ( .B(n43169), .A(n43694), .Z(n43692) );
  XNOR U43024 ( .A(n43695), .B(n43696), .Z(n39917) );
  AND U43025 ( .A(n43165), .B(n43163), .Z(n43695) );
  XNOR U43026 ( .A(n43697), .B(n43698), .Z(n38453) );
  XNOR U43027 ( .A(n43699), .B(n42095), .Z(n43152) );
  AND U43028 ( .A(n38206), .B(n38207), .Z(n43684) );
  XNOR U43029 ( .A(n40686), .B(n35376), .Z(n38207) );
  XNOR U43030 ( .A(n43702), .B(n43703), .Z(n40920) );
  XOR U43031 ( .A(n39544), .B(n36521), .Z(n43703) );
  XOR U43032 ( .A(n43704), .B(n43216), .Z(n36521) );
  XOR U43033 ( .A(n43705), .B(n43706), .Z(n43216) );
  NOR U43034 ( .A(n42736), .B(n42737), .Z(n43704) );
  XNOR U43035 ( .A(n43707), .B(n42526), .Z(n42736) );
  XNOR U43036 ( .A(n43708), .B(n43639), .Z(n39544) );
  XNOR U43037 ( .A(n43709), .B(n43552), .Z(n42749) );
  XOR U43038 ( .A(n39492), .B(n43710), .Z(n43702) );
  XOR U43039 ( .A(n42966), .B(n43200), .Z(n43710) );
  XNOR U43040 ( .A(n43711), .B(n43208), .Z(n43200) );
  XOR U43041 ( .A(n43712), .B(n43713), .Z(n43208) );
  ANDN U43042 ( .B(n42753), .A(n43714), .Z(n43711) );
  XOR U43043 ( .A(n43715), .B(n43716), .Z(n42753) );
  XNOR U43044 ( .A(n43717), .B(n43213), .Z(n42966) );
  XNOR U43045 ( .A(n43718), .B(n43719), .Z(n43213) );
  NOR U43046 ( .A(n42746), .B(n42745), .Z(n43717) );
  XNOR U43047 ( .A(n43720), .B(n42453), .Z(n42745) );
  XNOR U43048 ( .A(n43721), .B(n43205), .Z(n39492) );
  XOR U43049 ( .A(n43722), .B(n43723), .Z(n43205) );
  ANDN U43050 ( .B(n42741), .A(n42740), .Z(n43721) );
  XOR U43051 ( .A(n43724), .B(n42681), .Z(n42740) );
  XNOR U43052 ( .A(n43726), .B(n40023), .Z(n40686) );
  XOR U43053 ( .A(n43728), .B(n37114), .Z(n38206) );
  XNOR U43054 ( .A(n42445), .B(n40374), .Z(n37114) );
  XOR U43055 ( .A(n43729), .B(n43730), .Z(n40374) );
  XNOR U43056 ( .A(n40474), .B(n42123), .Z(n43730) );
  XNOR U43057 ( .A(n43731), .B(n43732), .Z(n42123) );
  ANDN U43058 ( .B(n43733), .A(n43734), .Z(n43731) );
  XNOR U43059 ( .A(n43735), .B(n43736), .Z(n40474) );
  ANDN U43060 ( .B(n42251), .A(n43737), .Z(n43735) );
  XOR U43061 ( .A(n39518), .B(n43738), .Z(n43729) );
  XOR U43062 ( .A(n38534), .B(n36705), .Z(n43738) );
  XOR U43063 ( .A(n43739), .B(n43740), .Z(n36705) );
  ANDN U43064 ( .B(n43517), .A(n43741), .Z(n43739) );
  XNOR U43065 ( .A(n43742), .B(n43743), .Z(n38534) );
  ANDN U43066 ( .B(n43744), .A(n42240), .Z(n43742) );
  XNOR U43067 ( .A(n43745), .B(n43746), .Z(n39518) );
  ANDN U43068 ( .B(n43747), .A(n42244), .Z(n43745) );
  XOR U43069 ( .A(n43748), .B(n43749), .Z(n42445) );
  XOR U43070 ( .A(n38897), .B(n39892), .Z(n43749) );
  XOR U43071 ( .A(n43750), .B(n43751), .Z(n39892) );
  ANDN U43072 ( .B(n43118), .A(n43752), .Z(n43750) );
  XNOR U43073 ( .A(n43753), .B(n42144), .Z(n38897) );
  ANDN U43074 ( .B(n42143), .A(n43122), .Z(n43753) );
  IV U43075 ( .A(n43754), .Z(n42143) );
  XNOR U43076 ( .A(n39623), .B(n43755), .Z(n43748) );
  XOR U43077 ( .A(n39039), .B(n39740), .Z(n43755) );
  XNOR U43078 ( .A(n43756), .B(n42139), .Z(n39740) );
  AND U43079 ( .A(n43127), .B(n42140), .Z(n43756) );
  XOR U43080 ( .A(n43757), .B(n42131), .Z(n39039) );
  NOR U43081 ( .A(n43134), .B(n42130), .Z(n43757) );
  XOR U43082 ( .A(n43758), .B(n42135), .Z(n39623) );
  AND U43083 ( .A(n43130), .B(n42136), .Z(n43758) );
  XOR U43084 ( .A(n43759), .B(n34758), .Z(n33176) );
  XOR U43085 ( .A(n42640), .B(n37884), .Z(n34758) );
  XOR U43086 ( .A(n43760), .B(n41142), .Z(n37884) );
  XNOR U43087 ( .A(n43761), .B(n43762), .Z(n41142) );
  XNOR U43088 ( .A(n39337), .B(n38568), .Z(n43762) );
  XOR U43089 ( .A(n43763), .B(n40688), .Z(n38568) );
  ANDN U43090 ( .B(n40689), .A(n40017), .Z(n43763) );
  XOR U43091 ( .A(n43764), .B(n43765), .Z(n40017) );
  XOR U43092 ( .A(n43766), .B(n43767), .Z(n40689) );
  XNOR U43093 ( .A(n43768), .B(n43727), .Z(n39337) );
  NOR U43094 ( .A(n41144), .B(n40021), .Z(n43768) );
  XOR U43095 ( .A(n43769), .B(n43770), .Z(n40021) );
  XNOR U43096 ( .A(n43771), .B(n42672), .Z(n41144) );
  XNOR U43097 ( .A(n35587), .B(n43772), .Z(n43761) );
  XOR U43098 ( .A(n39979), .B(n40673), .Z(n43772) );
  XOR U43099 ( .A(n43773), .B(n40683), .Z(n40673) );
  ANDN U43100 ( .B(n40684), .A(n40913), .Z(n43773) );
  XNOR U43101 ( .A(n43774), .B(n43775), .Z(n40913) );
  XNOR U43102 ( .A(n43776), .B(n43777), .Z(n40684) );
  XNOR U43103 ( .A(n43778), .B(n40691), .Z(n39979) );
  ANDN U43104 ( .B(n40692), .A(n40203), .Z(n43778) );
  XNOR U43105 ( .A(n42860), .B(n43779), .Z(n40203) );
  XNOR U43106 ( .A(n43780), .B(n43781), .Z(n40692) );
  XNOR U43107 ( .A(n43782), .B(n40679), .Z(n35587) );
  ANDN U43108 ( .B(n40680), .A(n41072), .Z(n43782) );
  XNOR U43109 ( .A(n43783), .B(n43565), .Z(n41072) );
  XOR U43110 ( .A(n43784), .B(n43785), .Z(n40680) );
  XNOR U43111 ( .A(n43786), .B(n43787), .Z(n42640) );
  ANDN U43112 ( .B(n40117), .A(n43788), .Z(n43786) );
  AND U43113 ( .A(n38215), .B(n38214), .Z(n43759) );
  XNOR U43114 ( .A(n43789), .B(n36212), .Z(n38214) );
  XNOR U43115 ( .A(n43791), .B(n43792), .Z(n43498) );
  XNOR U43116 ( .A(n40097), .B(n38932), .Z(n43792) );
  XOR U43117 ( .A(n43793), .B(n42618), .Z(n38932) );
  ANDN U43118 ( .B(n43794), .A(n43795), .Z(n43793) );
  XOR U43119 ( .A(n43796), .B(n42627), .Z(n40097) );
  IV U43120 ( .A(n43797), .Z(n42627) );
  ANDN U43121 ( .B(n43798), .A(n43799), .Z(n43796) );
  XNOR U43122 ( .A(n37079), .B(n43800), .Z(n43791) );
  XOR U43123 ( .A(n38299), .B(n35158), .Z(n43800) );
  XOR U43124 ( .A(n43801), .B(n42632), .Z(n35158) );
  ANDN U43125 ( .B(n43802), .A(n43803), .Z(n43801) );
  XOR U43126 ( .A(n43804), .B(n42622), .Z(n38299) );
  ANDN U43127 ( .B(n43805), .A(n43806), .Z(n43804) );
  XOR U43128 ( .A(n43807), .B(n43808), .Z(n37079) );
  NOR U43129 ( .A(n43809), .B(n43810), .Z(n43807) );
  XNOR U43130 ( .A(n43811), .B(n40569), .Z(n38215) );
  IV U43131 ( .A(n38642), .Z(n40569) );
  XOR U43132 ( .A(n41578), .B(n40429), .Z(n38642) );
  XNOR U43133 ( .A(n43812), .B(n43813), .Z(n40429) );
  XNOR U43134 ( .A(n37780), .B(n37450), .Z(n43813) );
  XNOR U43135 ( .A(n43814), .B(n41385), .Z(n37450) );
  XOR U43136 ( .A(n43815), .B(n43816), .Z(n41385) );
  ANDN U43137 ( .B(n41386), .A(n43817), .Z(n43814) );
  XOR U43138 ( .A(n43818), .B(n41380), .Z(n37780) );
  XOR U43139 ( .A(n43819), .B(n43820), .Z(n41380) );
  ANDN U43140 ( .B(n41381), .A(n43821), .Z(n43818) );
  XNOR U43141 ( .A(n38545), .B(n43822), .Z(n43812) );
  XOR U43142 ( .A(n39944), .B(n41373), .Z(n43822) );
  XNOR U43143 ( .A(n43823), .B(n43400), .Z(n41373) );
  XOR U43144 ( .A(n43824), .B(n43825), .Z(n43400) );
  ANDN U43145 ( .B(n43411), .A(n43826), .Z(n43823) );
  XOR U43146 ( .A(n43827), .B(n41393), .Z(n39944) );
  XOR U43147 ( .A(n43828), .B(n43829), .Z(n41393) );
  ANDN U43148 ( .B(n41394), .A(n43830), .Z(n43827) );
  XOR U43149 ( .A(n43831), .B(n41389), .Z(n38545) );
  XNOR U43150 ( .A(n43832), .B(n43833), .Z(n41389) );
  ANDN U43151 ( .B(n41390), .A(n43834), .Z(n43831) );
  XNOR U43152 ( .A(n43835), .B(n43836), .Z(n41578) );
  XNOR U43153 ( .A(n39020), .B(n36409), .Z(n43836) );
  XOR U43154 ( .A(n43837), .B(n43169), .Z(n36409) );
  XNOR U43155 ( .A(n43838), .B(n41657), .Z(n43169) );
  ANDN U43156 ( .B(n43168), .A(n43839), .Z(n43837) );
  XNOR U43157 ( .A(n43840), .B(n43841), .Z(n39020) );
  ANDN U43158 ( .B(n43182), .A(n43842), .Z(n43840) );
  XNOR U43159 ( .A(n40220), .B(n43843), .Z(n43835) );
  XNOR U43160 ( .A(n41149), .B(n38178), .Z(n43843) );
  XNOR U43161 ( .A(n43844), .B(n43174), .Z(n38178) );
  XNOR U43162 ( .A(n43845), .B(n43846), .Z(n43174) );
  NOR U43163 ( .A(n43847), .B(n43173), .Z(n43844) );
  XOR U43164 ( .A(n43848), .B(n43165), .Z(n41149) );
  XOR U43165 ( .A(n43849), .B(n43088), .Z(n43165) );
  ANDN U43166 ( .B(n43164), .A(n43850), .Z(n43848) );
  XNOR U43167 ( .A(n43851), .B(n43178), .Z(n40220) );
  XOR U43168 ( .A(n43852), .B(n43108), .Z(n43178) );
  ANDN U43169 ( .B(n43853), .A(n43177), .Z(n43851) );
  IV U43170 ( .A(n43854), .Z(n43177) );
  XNOR U43171 ( .A(n34356), .B(n43855), .Z(n43682) );
  XOR U43172 ( .A(n32933), .B(n32401), .Z(n43855) );
  XNOR U43173 ( .A(n43856), .B(n34768), .Z(n32401) );
  XOR U43174 ( .A(n35315), .B(n43857), .Z(n34768) );
  XOR U43175 ( .A(n43858), .B(n41513), .Z(n35315) );
  XNOR U43176 ( .A(n43859), .B(n43860), .Z(n41513) );
  XNOR U43177 ( .A(n37035), .B(n39594), .Z(n43860) );
  XNOR U43178 ( .A(n43861), .B(n40422), .Z(n39594) );
  XNOR U43179 ( .A(n43862), .B(n43863), .Z(n40422) );
  NOR U43180 ( .A(n40838), .B(n40587), .Z(n43861) );
  XNOR U43181 ( .A(n43864), .B(n40413), .Z(n37035) );
  XOR U43182 ( .A(n43865), .B(n43866), .Z(n40413) );
  NOR U43183 ( .A(n40847), .B(n40590), .Z(n43864) );
  XOR U43184 ( .A(n38130), .B(n43867), .Z(n43859) );
  XOR U43185 ( .A(n40581), .B(n36346), .Z(n43867) );
  XNOR U43186 ( .A(n43868), .B(n40426), .Z(n36346) );
  XOR U43187 ( .A(n43869), .B(n41742), .Z(n40426) );
  ANDN U43188 ( .B(n40592), .A(n40842), .Z(n43868) );
  XNOR U43189 ( .A(n43870), .B(n40417), .Z(n40581) );
  XNOR U43190 ( .A(n43871), .B(n43550), .Z(n40417) );
  NOR U43191 ( .A(n40585), .B(n40851), .Z(n43870) );
  XNOR U43192 ( .A(n43872), .B(n40409), .Z(n38130) );
  XNOR U43193 ( .A(n43873), .B(n43321), .Z(n40409) );
  NOR U43194 ( .A(n40594), .B(n40855), .Z(n43872) );
  AND U43195 ( .A(n38234), .B(n38233), .Z(n43856) );
  XNOR U43196 ( .A(n39165), .B(n43874), .Z(n38233) );
  XNOR U43197 ( .A(n41684), .B(n43475), .Z(n39165) );
  XNOR U43198 ( .A(n43875), .B(n43876), .Z(n43475) );
  XOR U43199 ( .A(n39146), .B(n35624), .Z(n43876) );
  XOR U43200 ( .A(n43877), .B(n43354), .Z(n35624) );
  AND U43201 ( .A(n43878), .B(n43355), .Z(n43877) );
  XNOR U43202 ( .A(n43879), .B(n43358), .Z(n39146) );
  XOR U43203 ( .A(n42552), .B(n43881), .Z(n43875) );
  XOR U43204 ( .A(n39243), .B(n37084), .Z(n43881) );
  XNOR U43205 ( .A(n43882), .B(n43366), .Z(n37084) );
  ANDN U43206 ( .B(n42944), .A(n43365), .Z(n43882) );
  XNOR U43207 ( .A(n43883), .B(n43368), .Z(n39243) );
  ANDN U43208 ( .B(n43369), .A(n43884), .Z(n43883) );
  IV U43209 ( .A(n43885), .Z(n43369) );
  XNOR U43210 ( .A(n43886), .B(n43362), .Z(n42552) );
  XOR U43211 ( .A(n43887), .B(n43888), .Z(n41684) );
  XNOR U43212 ( .A(n39837), .B(n41399), .Z(n43888) );
  XOR U43213 ( .A(n43889), .B(n41933), .Z(n41399) );
  XOR U43214 ( .A(n43865), .B(n43890), .Z(n41933) );
  ANDN U43215 ( .B(n43891), .A(n42557), .Z(n43889) );
  IV U43216 ( .A(n43892), .Z(n42557) );
  XNOR U43217 ( .A(n43893), .B(n41938), .Z(n39837) );
  XOR U43218 ( .A(n43894), .B(n43895), .Z(n41938) );
  ANDN U43219 ( .B(n42559), .A(n43896), .Z(n43893) );
  XOR U43220 ( .A(n41230), .B(n43897), .Z(n43887) );
  XOR U43221 ( .A(n39430), .B(n40321), .Z(n43897) );
  XNOR U43222 ( .A(n43898), .B(n41924), .Z(n40321) );
  XOR U43223 ( .A(n43899), .B(n43900), .Z(n41924) );
  ANDN U43224 ( .B(n42564), .A(n43901), .Z(n43898) );
  XOR U43225 ( .A(n43902), .B(n41930), .Z(n39430) );
  XOR U43226 ( .A(n43903), .B(n43904), .Z(n41930) );
  ANDN U43227 ( .B(n43905), .A(n42562), .Z(n43902) );
  IV U43228 ( .A(n43906), .Z(n42562) );
  XNOR U43229 ( .A(n43907), .B(n42567), .Z(n41230) );
  ANDN U43230 ( .B(n43908), .A(n43909), .Z(n43907) );
  XNOR U43231 ( .A(n43910), .B(n37044), .Z(n38234) );
  XOR U43232 ( .A(n42004), .B(n41997), .Z(n37044) );
  XNOR U43233 ( .A(n43911), .B(n43912), .Z(n41997) );
  XNOR U43234 ( .A(n37480), .B(n42168), .Z(n43912) );
  XNOR U43235 ( .A(n43913), .B(n43914), .Z(n42168) );
  NOR U43236 ( .A(n41167), .B(n41168), .Z(n43913) );
  XOR U43237 ( .A(n43915), .B(n43916), .Z(n41168) );
  XOR U43238 ( .A(n43917), .B(n43918), .Z(n37480) );
  ANDN U43239 ( .B(n41163), .A(n41164), .Z(n43917) );
  XNOR U43240 ( .A(n43919), .B(n43920), .Z(n41164) );
  XOR U43241 ( .A(n37618), .B(n43921), .Z(n43911) );
  XOR U43242 ( .A(n41089), .B(n40992), .Z(n43921) );
  XNOR U43243 ( .A(n43922), .B(n43923), .Z(n40992) );
  NOR U43244 ( .A(n41999), .B(n42001), .Z(n43922) );
  XOR U43245 ( .A(n43924), .B(n43925), .Z(n42001) );
  XNOR U43246 ( .A(n43926), .B(n43927), .Z(n41089) );
  NOR U43247 ( .A(n41177), .B(n41179), .Z(n43926) );
  XOR U43248 ( .A(n43928), .B(n43590), .Z(n41179) );
  IV U43249 ( .A(n42214), .Z(n43590) );
  XOR U43250 ( .A(n43929), .B(n43930), .Z(n37618) );
  NOR U43251 ( .A(n41173), .B(n41174), .Z(n43929) );
  XNOR U43252 ( .A(n40856), .B(n43931), .Z(n41174) );
  XOR U43253 ( .A(n43932), .B(n43933), .Z(n42004) );
  XOR U43254 ( .A(n37889), .B(n38675), .Z(n43933) );
  XNOR U43255 ( .A(n43934), .B(n43935), .Z(n38675) );
  NOR U43256 ( .A(n43433), .B(n43936), .Z(n43934) );
  XNOR U43257 ( .A(n43937), .B(n43938), .Z(n37889) );
  ANDN U43258 ( .B(n43425), .A(n43939), .Z(n43937) );
  XOR U43259 ( .A(n38668), .B(n43940), .Z(n43932) );
  XNOR U43260 ( .A(n37836), .B(n43941), .Z(n43940) );
  XOR U43261 ( .A(n43942), .B(n43943), .Z(n37836) );
  NOR U43262 ( .A(n43944), .B(n43429), .Z(n43942) );
  XOR U43263 ( .A(n43945), .B(n43946), .Z(n38668) );
  ANDN U43264 ( .B(n43947), .A(n43948), .Z(n43945) );
  XOR U43265 ( .A(n43949), .B(n36091), .Z(n32933) );
  XOR U43266 ( .A(n37328), .B(n43305), .Z(n36091) );
  XOR U43267 ( .A(n43950), .B(n43951), .Z(n43305) );
  ANDN U43268 ( .B(n40758), .A(n41489), .Z(n43950) );
  XOR U43269 ( .A(n43665), .B(n43952), .Z(n40758) );
  XNOR U43270 ( .A(n39222), .B(n40468), .Z(n37328) );
  XNOR U43271 ( .A(n43953), .B(n43954), .Z(n40468) );
  XNOR U43272 ( .A(n43955), .B(n37423), .Z(n43954) );
  XNOR U43273 ( .A(n43956), .B(n40770), .Z(n37423) );
  ANDN U43274 ( .B(n43301), .A(n41487), .Z(n43956) );
  XOR U43275 ( .A(n43957), .B(n43958), .Z(n41487) );
  XOR U43276 ( .A(n39183), .B(n43959), .Z(n43953) );
  XOR U43277 ( .A(n35934), .B(n38462), .Z(n43959) );
  XNOR U43278 ( .A(n43960), .B(n40760), .Z(n38462) );
  ANDN U43279 ( .B(n41489), .A(n43951), .Z(n43960) );
  XOR U43280 ( .A(n43961), .B(n43962), .Z(n41489) );
  XNOR U43281 ( .A(n43963), .B(n41492), .Z(n35934) );
  XOR U43282 ( .A(n43964), .B(n43965), .Z(n41478) );
  XNOR U43283 ( .A(n43966), .B(n40764), .Z(n39183) );
  ANDN U43284 ( .B(n43296), .A(n41485), .Z(n43966) );
  IV U43285 ( .A(n43297), .Z(n41485) );
  XOR U43286 ( .A(n43967), .B(n43968), .Z(n43297) );
  XOR U43287 ( .A(n43969), .B(n43970), .Z(n39222) );
  XNOR U43288 ( .A(n35511), .B(n38555), .Z(n43970) );
  XNOR U43289 ( .A(n43971), .B(n40456), .Z(n38555) );
  ANDN U43290 ( .B(n43972), .A(n43973), .Z(n43971) );
  XOR U43291 ( .A(n43974), .B(n41185), .Z(n35511) );
  ANDN U43292 ( .B(n43975), .A(n42069), .Z(n43974) );
  XNOR U43293 ( .A(n35801), .B(n43976), .Z(n43969) );
  XNOR U43294 ( .A(n40570), .B(n40135), .Z(n43976) );
  XNOR U43295 ( .A(n43977), .B(n42073), .Z(n40135) );
  AND U43296 ( .A(n43978), .B(n42065), .Z(n43977) );
  XOR U43297 ( .A(n43979), .B(n40453), .Z(n40570) );
  AND U43298 ( .A(n43980), .B(n42060), .Z(n43979) );
  XOR U43299 ( .A(n43981), .B(n40461), .Z(n35801) );
  AND U43300 ( .A(n43982), .B(n43983), .Z(n43981) );
  ANDN U43301 ( .B(n38476), .A(n38915), .Z(n43949) );
  IV U43302 ( .A(n43389), .Z(n38915) );
  XOR U43303 ( .A(n41326), .B(n34617), .Z(n43389) );
  XNOR U43304 ( .A(n43984), .B(n43985), .Z(n40360) );
  XNOR U43305 ( .A(n36398), .B(n37511), .Z(n43985) );
  XOR U43306 ( .A(n43986), .B(n43987), .Z(n37511) );
  NOR U43307 ( .A(n43988), .B(n39505), .Z(n43986) );
  XNOR U43308 ( .A(n43989), .B(n43510), .Z(n36398) );
  NOR U43309 ( .A(n40362), .B(n40363), .Z(n43989) );
  XOR U43310 ( .A(n39840), .B(n43990), .Z(n43984) );
  XOR U43311 ( .A(n39480), .B(n36368), .Z(n43990) );
  XNOR U43312 ( .A(n43991), .B(n43513), .Z(n36368) );
  NOR U43313 ( .A(n39500), .B(n39499), .Z(n43991) );
  XNOR U43314 ( .A(n43992), .B(n43506), .Z(n39480) );
  NOR U43315 ( .A(n39508), .B(n39509), .Z(n43992) );
  XNOR U43316 ( .A(n43993), .B(n43503), .Z(n39840) );
  XNOR U43317 ( .A(n43995), .B(n43996), .Z(n41326) );
  ANDN U43318 ( .B(n43997), .A(n43998), .Z(n43995) );
  XOR U43319 ( .A(n43999), .B(n39528), .Z(n38476) );
  XOR U43320 ( .A(n44000), .B(n34753), .Z(n34356) );
  XNOR U43321 ( .A(n44001), .B(n38775), .Z(n34753) );
  IV U43322 ( .A(n37789), .Z(n38775) );
  XOR U43323 ( .A(n40477), .B(n40465), .Z(n37789) );
  XOR U43324 ( .A(n44002), .B(n44003), .Z(n40465) );
  XNOR U43325 ( .A(n38125), .B(n40139), .Z(n44003) );
  XOR U43326 ( .A(n44004), .B(n40727), .Z(n40139) );
  XOR U43327 ( .A(n44005), .B(n43550), .Z(n40727) );
  ANDN U43328 ( .B(n40728), .A(n44006), .Z(n44004) );
  XOR U43329 ( .A(n44007), .B(n40724), .Z(n38125) );
  XNOR U43330 ( .A(n44008), .B(n44009), .Z(n40724) );
  ANDN U43331 ( .B(n40723), .A(n44010), .Z(n44007) );
  XOR U43332 ( .A(n38167), .B(n44011), .Z(n44002) );
  XNOR U43333 ( .A(n40704), .B(n38420), .Z(n44011) );
  XOR U43334 ( .A(n44012), .B(n40715), .Z(n38420) );
  XOR U43335 ( .A(n44013), .B(n44014), .Z(n40715) );
  ANDN U43336 ( .B(n40714), .A(n44015), .Z(n44012) );
  XNOR U43337 ( .A(n44016), .B(n40711), .Z(n40704) );
  ANDN U43338 ( .B(n44018), .A(n40710), .Z(n44016) );
  XOR U43339 ( .A(n44019), .B(n40720), .Z(n38167) );
  NOR U43340 ( .A(n44020), .B(n44021), .Z(n44019) );
  XOR U43341 ( .A(n44022), .B(n44023), .Z(n40477) );
  XNOR U43342 ( .A(n40055), .B(n39002), .Z(n44023) );
  XNOR U43343 ( .A(n44024), .B(n40306), .Z(n39002) );
  XOR U43344 ( .A(n44025), .B(n44026), .Z(n40306) );
  ANDN U43345 ( .B(n40307), .A(n40161), .Z(n44024) );
  XNOR U43346 ( .A(n44027), .B(n40315), .Z(n40055) );
  XOR U43347 ( .A(n44028), .B(n44029), .Z(n40315) );
  ANDN U43348 ( .B(n40316), .A(n41544), .Z(n44027) );
  XOR U43349 ( .A(n40300), .B(n44030), .Z(n44022) );
  XOR U43350 ( .A(n37220), .B(n39429), .Z(n44030) );
  XNOR U43351 ( .A(n44031), .B(n40319), .Z(n39429) );
  XOR U43352 ( .A(n44032), .B(n44033), .Z(n40319) );
  AND U43353 ( .A(n40398), .B(n40320), .Z(n44031) );
  XNOR U43354 ( .A(n44034), .B(n40312), .Z(n37220) );
  XOR U43355 ( .A(n44035), .B(n44036), .Z(n40312) );
  ANDN U43356 ( .B(n42820), .A(n40311), .Z(n44034) );
  XNOR U43357 ( .A(n44037), .B(n42399), .Z(n40300) );
  XOR U43358 ( .A(n44038), .B(n44039), .Z(n42399) );
  ANDN U43359 ( .B(n42420), .A(n40154), .Z(n44037) );
  AND U43360 ( .A(n38212), .B(n38211), .Z(n44000) );
  XNOR U43361 ( .A(n44040), .B(n36555), .Z(n38211) );
  XNOR U43362 ( .A(n44041), .B(n36219), .Z(n38212) );
  XOR U43363 ( .A(n40520), .B(n40530), .Z(n36219) );
  XOR U43364 ( .A(n44042), .B(n44043), .Z(n40530) );
  XNOR U43365 ( .A(n39090), .B(n37713), .Z(n44043) );
  XOR U43366 ( .A(n44044), .B(n40948), .Z(n37713) );
  ANDN U43367 ( .B(n40949), .A(n43386), .Z(n44044) );
  XOR U43368 ( .A(n44045), .B(n44046), .Z(n39090) );
  ANDN U43369 ( .B(n43373), .A(n42187), .Z(n44045) );
  IV U43370 ( .A(n44047), .Z(n42187) );
  XNOR U43371 ( .A(n39828), .B(n44048), .Z(n44042) );
  XOR U43372 ( .A(n40214), .B(n37029), .Z(n44048) );
  XOR U43373 ( .A(n44049), .B(n40952), .Z(n37029) );
  ANDN U43374 ( .B(n40953), .A(n44050), .Z(n44049) );
  XOR U43375 ( .A(n44051), .B(n40959), .Z(n40214) );
  AND U43376 ( .A(n40960), .B(n43376), .Z(n44051) );
  XOR U43377 ( .A(n44052), .B(n43478), .Z(n39828) );
  ANDN U43378 ( .B(n43479), .A(n43382), .Z(n44052) );
  XNOR U43379 ( .A(n44053), .B(n44054), .Z(n40520) );
  XOR U43380 ( .A(n38551), .B(n40340), .Z(n44054) );
  XOR U43381 ( .A(n44055), .B(n44056), .Z(n40340) );
  ANDN U43382 ( .B(n44057), .A(n42428), .Z(n44055) );
  XNOR U43383 ( .A(n44058), .B(n44059), .Z(n38551) );
  ANDN U43384 ( .B(n44060), .A(n44061), .Z(n44058) );
  XNOR U43385 ( .A(n40942), .B(n44062), .Z(n44053) );
  XOR U43386 ( .A(n38331), .B(n36962), .Z(n44062) );
  XNOR U43387 ( .A(n44063), .B(n44064), .Z(n36962) );
  ANDN U43388 ( .B(n44065), .A(n42433), .Z(n44063) );
  IV U43389 ( .A(n44066), .Z(n42433) );
  XOR U43390 ( .A(n44067), .B(n44068), .Z(n38331) );
  ANDN U43391 ( .B(n44069), .A(n42441), .Z(n44067) );
  IV U43392 ( .A(n44070), .Z(n42441) );
  XNOR U43393 ( .A(n44071), .B(n44072), .Z(n40942) );
  ANDN U43394 ( .B(n44073), .A(n42437), .Z(n44071) );
  XNOR U43395 ( .A(n44074), .B(n28053), .Z(n31293) );
  XNOR U43396 ( .A(n35990), .B(n30514), .Z(n28053) );
  XNOR U43397 ( .A(n32380), .B(n39646), .Z(n30514) );
  XNOR U43398 ( .A(n44075), .B(n44076), .Z(n39646) );
  XOR U43399 ( .A(n34354), .B(n30502), .Z(n44076) );
  XNOR U43400 ( .A(n44077), .B(n35462), .Z(n30502) );
  XOR U43401 ( .A(n43486), .B(n39247), .Z(n35462) );
  IV U43402 ( .A(n37954), .Z(n39247) );
  XNOR U43403 ( .A(n44078), .B(n40876), .Z(n43486) );
  AND U43404 ( .A(n40933), .B(n40932), .Z(n44078) );
  ANDN U43405 ( .B(n35461), .A(n32476), .Z(n44077) );
  XOR U43406 ( .A(n39158), .B(n44079), .Z(n32476) );
  XOR U43407 ( .A(n43140), .B(n44080), .Z(n39158) );
  XOR U43408 ( .A(n44081), .B(n44082), .Z(n43140) );
  XOR U43409 ( .A(n39517), .B(n44083), .Z(n44082) );
  XOR U43410 ( .A(n44084), .B(n44085), .Z(n39517) );
  ANDN U43411 ( .B(n44086), .A(n44087), .Z(n44084) );
  XNOR U43412 ( .A(n39136), .B(n44088), .Z(n44081) );
  XNOR U43413 ( .A(n37419), .B(n33916), .Z(n44088) );
  XOR U43414 ( .A(n44089), .B(n41410), .Z(n33916) );
  NOR U43415 ( .A(n44090), .B(n44091), .Z(n44089) );
  XNOR U43416 ( .A(n44092), .B(n41416), .Z(n37419) );
  ANDN U43417 ( .B(n44093), .A(n44094), .Z(n44092) );
  XOR U43418 ( .A(n44095), .B(n41406), .Z(n39136) );
  ANDN U43419 ( .B(n44096), .A(n44097), .Z(n44095) );
  XNOR U43420 ( .A(n39011), .B(n43614), .Z(n35461) );
  XOR U43421 ( .A(n44098), .B(n44099), .Z(n43614) );
  ANDN U43422 ( .B(n41523), .A(n41524), .Z(n44098) );
  XNOR U43423 ( .A(n44100), .B(n44101), .Z(n42575) );
  XOR U43424 ( .A(n38155), .B(n39742), .Z(n44101) );
  XNOR U43425 ( .A(n44102), .B(n44103), .Z(n39742) );
  ANDN U43426 ( .B(n41540), .A(n44104), .Z(n44102) );
  XOR U43427 ( .A(n44105), .B(n44106), .Z(n41540) );
  XNOR U43428 ( .A(n44107), .B(n44108), .Z(n38155) );
  ANDN U43429 ( .B(n44099), .A(n41523), .Z(n44107) );
  XNOR U43430 ( .A(n44109), .B(n43644), .Z(n41523) );
  XOR U43431 ( .A(n39080), .B(n44110), .Z(n44100) );
  XOR U43432 ( .A(n38845), .B(n37026), .Z(n44110) );
  XNOR U43433 ( .A(n44111), .B(n44112), .Z(n37026) );
  ANDN U43434 ( .B(n43609), .A(n41532), .Z(n44111) );
  XOR U43435 ( .A(n44113), .B(n44114), .Z(n41532) );
  XNOR U43436 ( .A(n44115), .B(n44116), .Z(n38845) );
  NOR U43437 ( .A(n44117), .B(n41536), .Z(n44115) );
  XOR U43438 ( .A(n44118), .B(n44119), .Z(n41536) );
  XOR U43439 ( .A(n44120), .B(n44121), .Z(n39080) );
  NOR U43440 ( .A(n44122), .B(n41527), .Z(n44120) );
  XOR U43441 ( .A(n41598), .B(n44123), .Z(n41527) );
  XNOR U43442 ( .A(n44124), .B(n44125), .Z(n39818) );
  XOR U43443 ( .A(n37542), .B(n40475), .Z(n44125) );
  XOR U43444 ( .A(n44126), .B(n42999), .Z(n40475) );
  XNOR U43445 ( .A(n44128), .B(n43003), .Z(n37542) );
  ANDN U43446 ( .B(n43002), .A(n44129), .Z(n44128) );
  XNOR U43447 ( .A(n40566), .B(n44130), .Z(n44124) );
  XOR U43448 ( .A(n38418), .B(n42967), .Z(n44130) );
  XOR U43449 ( .A(n44131), .B(n42995), .Z(n42967) );
  ANDN U43450 ( .B(n44132), .A(n42994), .Z(n44131) );
  XNOR U43451 ( .A(n44133), .B(n42986), .Z(n38418) );
  ANDN U43452 ( .B(n44134), .A(n44135), .Z(n44133) );
  XNOR U43453 ( .A(n44136), .B(n42990), .Z(n40566) );
  XNOR U43454 ( .A(n44138), .B(n35470), .Z(n34354) );
  XNOR U43455 ( .A(n44139), .B(n38573), .Z(n35470) );
  XOR U43456 ( .A(n42532), .B(n44140), .Z(n38573) );
  XNOR U43457 ( .A(n44141), .B(n44142), .Z(n42532) );
  XNOR U43458 ( .A(n38501), .B(n37845), .Z(n44142) );
  XNOR U43459 ( .A(n44143), .B(n41125), .Z(n37845) );
  NOR U43460 ( .A(n44144), .B(n42270), .Z(n44143) );
  XNOR U43461 ( .A(n44145), .B(n41132), .Z(n38501) );
  NOR U43462 ( .A(n41131), .B(n42262), .Z(n44145) );
  XOR U43463 ( .A(n40247), .B(n44146), .Z(n44141) );
  XNOR U43464 ( .A(n39977), .B(n35788), .Z(n44146) );
  XNOR U43465 ( .A(n44147), .B(n44148), .Z(n35788) );
  NOR U43466 ( .A(n44149), .B(n42258), .Z(n44147) );
  XOR U43467 ( .A(n44150), .B(n43061), .Z(n39977) );
  ANDN U43468 ( .B(n43062), .A(n42273), .Z(n44150) );
  XOR U43469 ( .A(n44151), .B(n41136), .Z(n40247) );
  NOR U43470 ( .A(n42266), .B(n41135), .Z(n44151) );
  ANDN U43471 ( .B(n35469), .A(n34600), .Z(n44138) );
  IV U43472 ( .A(n44152), .Z(n34600) );
  XNOR U43473 ( .A(n35439), .B(n44153), .Z(n44075) );
  XOR U43474 ( .A(n31948), .B(n32387), .Z(n44153) );
  XOR U43475 ( .A(n44154), .B(n35459), .Z(n32387) );
  XOR U43476 ( .A(n44155), .B(n37472), .Z(n35459) );
  XNOR U43477 ( .A(n44156), .B(n44157), .Z(n42050) );
  XNOR U43478 ( .A(n39555), .B(n37916), .Z(n44157) );
  XNOR U43479 ( .A(n44158), .B(n41267), .Z(n37916) );
  XOR U43480 ( .A(n44159), .B(n43925), .Z(n41267) );
  ANDN U43481 ( .B(n41268), .A(n43090), .Z(n44158) );
  IV U43482 ( .A(n44160), .Z(n43090) );
  XNOR U43483 ( .A(n44161), .B(n41261), .Z(n39555) );
  XNOR U43484 ( .A(n42331), .B(n44162), .Z(n41261) );
  IV U43485 ( .A(n44163), .Z(n42331) );
  ANDN U43486 ( .B(n41262), .A(n43076), .Z(n44161) );
  XOR U43487 ( .A(n41038), .B(n44164), .Z(n44156) );
  XOR U43488 ( .A(n41252), .B(n35603), .Z(n44164) );
  XNOR U43489 ( .A(n44165), .B(n41869), .Z(n35603) );
  XOR U43490 ( .A(n44166), .B(n44167), .Z(n41869) );
  ANDN U43491 ( .B(n41868), .A(n43082), .Z(n44165) );
  XNOR U43492 ( .A(n44168), .B(n41257), .Z(n41252) );
  XOR U43493 ( .A(n44169), .B(n42419), .Z(n41257) );
  XNOR U43494 ( .A(n44171), .B(n41272), .Z(n41038) );
  XOR U43495 ( .A(n44172), .B(n44173), .Z(n41272) );
  XNOR U43496 ( .A(n44174), .B(n44175), .Z(n39675) );
  XOR U43497 ( .A(n37475), .B(n37031), .Z(n44175) );
  XOR U43498 ( .A(n44176), .B(n41277), .Z(n37031) );
  XNOR U43499 ( .A(n44177), .B(n44178), .Z(n41277) );
  NOR U43500 ( .A(n41278), .B(n41451), .Z(n44176) );
  XNOR U43501 ( .A(n44179), .B(n44180), .Z(n41451) );
  XOR U43502 ( .A(n44181), .B(n44182), .Z(n41278) );
  XNOR U43503 ( .A(n44183), .B(n41887), .Z(n37475) );
  IV U43504 ( .A(n41281), .Z(n41887) );
  XOR U43505 ( .A(n44184), .B(n43079), .Z(n41281) );
  ANDN U43506 ( .B(n41282), .A(n41438), .Z(n44183) );
  XOR U43507 ( .A(n44185), .B(n44186), .Z(n41438) );
  XOR U43508 ( .A(n44187), .B(n43581), .Z(n41282) );
  XOR U43509 ( .A(n40164), .B(n44188), .Z(n44174) );
  XOR U43510 ( .A(n39287), .B(n37054), .Z(n44188) );
  XNOR U43511 ( .A(n44189), .B(n41286), .Z(n37054) );
  XOR U43512 ( .A(n44190), .B(n44191), .Z(n41286) );
  ANDN U43513 ( .B(n41287), .A(n41448), .Z(n44189) );
  XNOR U43514 ( .A(n44192), .B(n44193), .Z(n41448) );
  XOR U43515 ( .A(n44194), .B(n44195), .Z(n41287) );
  XNOR U43516 ( .A(n44196), .B(n41291), .Z(n39287) );
  XNOR U43517 ( .A(n44197), .B(n43925), .Z(n41291) );
  ANDN U43518 ( .B(n41290), .A(n41445), .Z(n44196) );
  XNOR U43519 ( .A(n44198), .B(n44199), .Z(n41445) );
  XOR U43520 ( .A(n44200), .B(n44201), .Z(n41290) );
  XNOR U43521 ( .A(n44202), .B(n41879), .Z(n40164) );
  XOR U43522 ( .A(n44203), .B(n44204), .Z(n41879) );
  NOR U43523 ( .A(n41441), .B(n41294), .Z(n44202) );
  XNOR U43524 ( .A(n44205), .B(n43825), .Z(n41294) );
  XNOR U43525 ( .A(n44206), .B(n42516), .Z(n41441) );
  IV U43526 ( .A(n44207), .Z(n42516) );
  ANDN U43527 ( .B(n35458), .A(n32472), .Z(n44154) );
  XOR U43528 ( .A(n43380), .B(n37427), .Z(n32472) );
  XOR U43529 ( .A(n41918), .B(n44208), .Z(n37427) );
  XOR U43530 ( .A(n44209), .B(n44210), .Z(n41918) );
  XOR U43531 ( .A(n41572), .B(n39376), .Z(n44210) );
  XOR U43532 ( .A(n44211), .B(n44212), .Z(n39376) );
  NOR U43533 ( .A(n44213), .B(n43358), .Z(n44211) );
  XOR U43534 ( .A(n44214), .B(n44215), .Z(n43358) );
  XOR U43535 ( .A(n44216), .B(n42938), .Z(n41572) );
  NOR U43536 ( .A(n42937), .B(n43368), .Z(n44216) );
  XOR U43537 ( .A(n44217), .B(n44218), .Z(n43368) );
  XOR U43538 ( .A(n44219), .B(n44220), .Z(n42937) );
  XNOR U43539 ( .A(n37348), .B(n44221), .Z(n44209) );
  XNOR U43540 ( .A(n40004), .B(n42928), .Z(n44221) );
  XOR U43541 ( .A(n44222), .B(n42942), .Z(n42928) );
  NOR U43542 ( .A(n43362), .B(n42941), .Z(n44222) );
  XOR U43543 ( .A(n44223), .B(n44224), .Z(n42941) );
  XOR U43544 ( .A(n44225), .B(n44226), .Z(n43362) );
  XNOR U43545 ( .A(n44227), .B(n44228), .Z(n40004) );
  NOR U43546 ( .A(n43353), .B(n43354), .Z(n44227) );
  XNOR U43547 ( .A(n44229), .B(n43574), .Z(n43354) );
  XOR U43548 ( .A(n44230), .B(n42946), .Z(n37348) );
  NOR U43549 ( .A(n43366), .B(n42945), .Z(n44230) );
  XNOR U43550 ( .A(n44231), .B(n44232), .Z(n42945) );
  XNOR U43551 ( .A(n42667), .B(n44233), .Z(n43366) );
  XNOR U43552 ( .A(n44234), .B(n44050), .Z(n43380) );
  XNOR U43553 ( .A(n39848), .B(n44236), .Z(n35458) );
  XNOR U43554 ( .A(n44237), .B(n35466), .Z(n31948) );
  XNOR U43555 ( .A(n44238), .B(n39454), .Z(n35466) );
  ANDN U43556 ( .B(n35467), .A(n32466), .Z(n44237) );
  XOR U43557 ( .A(n41921), .B(n35595), .Z(n32466) );
  IV U43558 ( .A(n37871), .Z(n35595) );
  XOR U43559 ( .A(n42929), .B(n42785), .Z(n37871) );
  XOR U43560 ( .A(n44239), .B(n44240), .Z(n42785) );
  XNOR U43561 ( .A(n44079), .B(n39533), .Z(n44240) );
  XOR U43562 ( .A(n44241), .B(n44090), .Z(n39533) );
  ANDN U43563 ( .B(n44091), .A(n41408), .Z(n44241) );
  XNOR U43564 ( .A(n44242), .B(n44243), .Z(n44079) );
  ANDN U43565 ( .B(n43066), .A(n44244), .Z(n44242) );
  XOR U43566 ( .A(n39159), .B(n44245), .Z(n44239) );
  XOR U43567 ( .A(n39971), .B(n39558), .Z(n44245) );
  XNOR U43568 ( .A(n44246), .B(n44247), .Z(n39558) );
  NOR U43569 ( .A(n44248), .B(n44086), .Z(n44246) );
  XNOR U43570 ( .A(n44249), .B(n44096), .Z(n39971) );
  XNOR U43571 ( .A(n44250), .B(n44093), .Z(n39159) );
  ANDN U43572 ( .B(n44094), .A(n41415), .Z(n44250) );
  XOR U43573 ( .A(n44251), .B(n44252), .Z(n42929) );
  XOR U43574 ( .A(n43139), .B(n36988), .Z(n44252) );
  XNOR U43575 ( .A(n44253), .B(n43901), .Z(n36988) );
  ANDN U43576 ( .B(n41925), .A(n41923), .Z(n44253) );
  XOR U43577 ( .A(n44254), .B(n44255), .Z(n41925) );
  XNOR U43578 ( .A(n44256), .B(n43908), .Z(n43139) );
  ANDN U43579 ( .B(n42566), .A(n44257), .Z(n44256) );
  XOR U43580 ( .A(n37667), .B(n44258), .Z(n44251) );
  XOR U43581 ( .A(n39890), .B(n39420), .Z(n44258) );
  XOR U43582 ( .A(n44259), .B(n43891), .Z(n39420) );
  XOR U43583 ( .A(n44260), .B(n43777), .Z(n41934) );
  NOR U43584 ( .A(n41929), .B(n41928), .Z(n44261) );
  XOR U43585 ( .A(n44262), .B(n44263), .Z(n41929) );
  XNOR U43586 ( .A(n44264), .B(n43896), .Z(n37667) );
  ANDN U43587 ( .B(n41936), .A(n41937), .Z(n44264) );
  XOR U43588 ( .A(n44265), .B(n42163), .Z(n41937) );
  XNOR U43589 ( .A(n44266), .B(n44267), .Z(n41921) );
  NOR U43590 ( .A(n42567), .B(n42566), .Z(n44266) );
  XNOR U43591 ( .A(n42537), .B(n44268), .Z(n42566) );
  XNOR U43592 ( .A(n44269), .B(n44270), .Z(n42567) );
  XOR U43593 ( .A(n44271), .B(n37500), .Z(n35467) );
  IV U43594 ( .A(n38426), .Z(n37500) );
  XOR U43595 ( .A(n41119), .B(n41717), .Z(n38426) );
  XNOR U43596 ( .A(n44272), .B(n44273), .Z(n41717) );
  XOR U43597 ( .A(n39812), .B(n44274), .Z(n44273) );
  XNOR U43598 ( .A(n44275), .B(n42367), .Z(n39812) );
  ANDN U43599 ( .B(n44276), .A(n44277), .Z(n44275) );
  XOR U43600 ( .A(n36554), .B(n44278), .Z(n44272) );
  XOR U43601 ( .A(n44040), .B(n39410), .Z(n44278) );
  XOR U43602 ( .A(n44279), .B(n42379), .Z(n39410) );
  ANDN U43603 ( .B(n44280), .A(n44281), .Z(n44279) );
  XNOR U43604 ( .A(n44282), .B(n42371), .Z(n44040) );
  IV U43605 ( .A(n44283), .Z(n42371) );
  NOR U43606 ( .A(n44284), .B(n44285), .Z(n44282) );
  XNOR U43607 ( .A(n44286), .B(n42384), .Z(n36554) );
  ANDN U43608 ( .B(n44287), .A(n44288), .Z(n44286) );
  XNOR U43609 ( .A(n44289), .B(n44290), .Z(n41119) );
  XOR U43610 ( .A(n38525), .B(n39072), .Z(n44290) );
  XOR U43611 ( .A(n44291), .B(n42291), .Z(n39072) );
  ANDN U43612 ( .B(n44292), .A(n44293), .Z(n44291) );
  XNOR U43613 ( .A(n44294), .B(n42295), .Z(n38525) );
  XOR U43614 ( .A(n39624), .B(n44297), .Z(n44289) );
  XOR U43615 ( .A(n37799), .B(n43040), .Z(n44297) );
  XOR U43616 ( .A(n44298), .B(n44299), .Z(n43040) );
  NOR U43617 ( .A(n44300), .B(n44301), .Z(n44298) );
  XNOR U43618 ( .A(n44302), .B(n42281), .Z(n37799) );
  NOR U43619 ( .A(n44303), .B(n44304), .Z(n44302) );
  XNOR U43620 ( .A(n44305), .B(n42285), .Z(n39624) );
  ANDN U43621 ( .B(n44306), .A(n44307), .Z(n44305) );
  XOR U43622 ( .A(n44308), .B(n36451), .Z(n35439) );
  XOR U43623 ( .A(n38113), .B(n42062), .Z(n36451) );
  XNOR U43624 ( .A(n44309), .B(n43973), .Z(n42062) );
  IV U43625 ( .A(n44310), .Z(n43973) );
  NOR U43626 ( .A(n40457), .B(n40455), .Z(n44309) );
  ANDN U43627 ( .B(n32878), .A(n35987), .Z(n44308) );
  XOR U43628 ( .A(n38320), .B(n44311), .Z(n35987) );
  XOR U43629 ( .A(n44312), .B(n43476), .Z(n38320) );
  XOR U43630 ( .A(n44313), .B(n44314), .Z(n43476) );
  XOR U43631 ( .A(n39261), .B(n43349), .Z(n44314) );
  XOR U43632 ( .A(n44315), .B(n43377), .Z(n43349) );
  NOR U43633 ( .A(n43378), .B(n40959), .Z(n44315) );
  XOR U43634 ( .A(n44316), .B(n44317), .Z(n40959) );
  XOR U43635 ( .A(n44318), .B(n43287), .Z(n43378) );
  XNOR U43636 ( .A(n44319), .B(n43383), .Z(n39261) );
  ANDN U43637 ( .B(n43384), .A(n43478), .Z(n44319) );
  XNOR U43638 ( .A(n44320), .B(n44321), .Z(n43478) );
  XNOR U43639 ( .A(n44322), .B(n44323), .Z(n43384) );
  XOR U43640 ( .A(n36201), .B(n44324), .Z(n44313) );
  XNOR U43641 ( .A(n41757), .B(n40823), .Z(n44324) );
  XNOR U43642 ( .A(n44325), .B(n43374), .Z(n40823) );
  ANDN U43643 ( .B(n42186), .A(n44046), .Z(n44325) );
  IV U43644 ( .A(n42188), .Z(n44046) );
  XOR U43645 ( .A(n44326), .B(n44327), .Z(n42188) );
  XNOR U43646 ( .A(n44328), .B(n44329), .Z(n42186) );
  XNOR U43647 ( .A(n44330), .B(n43387), .Z(n41757) );
  ANDN U43648 ( .B(n40947), .A(n40948), .Z(n44330) );
  XOR U43649 ( .A(n43769), .B(n44331), .Z(n40948) );
  XNOR U43650 ( .A(n44332), .B(n44333), .Z(n40947) );
  XNOR U43651 ( .A(n44334), .B(n44235), .Z(n36201) );
  ANDN U43652 ( .B(n40951), .A(n40952), .Z(n44334) );
  XOR U43653 ( .A(n44335), .B(n44336), .Z(n40952) );
  XNOR U43654 ( .A(n44337), .B(n44338), .Z(n40951) );
  XOR U43655 ( .A(n40657), .B(n44339), .Z(n32878) );
  XOR U43656 ( .A(n44340), .B(n40507), .Z(n40657) );
  XNOR U43657 ( .A(n44341), .B(n44342), .Z(n40507) );
  XNOR U43658 ( .A(n40091), .B(n39809), .Z(n44342) );
  XNOR U43659 ( .A(n44343), .B(n41113), .Z(n39809) );
  NOR U43660 ( .A(n41114), .B(n44344), .Z(n44343) );
  XNOR U43661 ( .A(n44345), .B(n41096), .Z(n40091) );
  ANDN U43662 ( .B(n41097), .A(n44346), .Z(n44345) );
  XOR U43663 ( .A(n39441), .B(n44347), .Z(n44341) );
  XOR U43664 ( .A(n38297), .B(n41090), .Z(n44347) );
  XOR U43665 ( .A(n44348), .B(n41110), .Z(n41090) );
  NOR U43666 ( .A(n44349), .B(n41109), .Z(n44348) );
  XNOR U43667 ( .A(n44350), .B(n41106), .Z(n38297) );
  NOR U43668 ( .A(n41105), .B(n44351), .Z(n44350) );
  XNOR U43669 ( .A(n44352), .B(n41101), .Z(n39441) );
  NOR U43670 ( .A(n41100), .B(n44353), .Z(n44352) );
  XOR U43671 ( .A(n44354), .B(n44355), .Z(n32380) );
  XNOR U43672 ( .A(n31550), .B(n32616), .Z(n44355) );
  XNOR U43673 ( .A(n44356), .B(n38249), .Z(n32616) );
  XOR U43674 ( .A(n36894), .B(n41310), .Z(n38249) );
  XNOR U43675 ( .A(n44357), .B(n44358), .Z(n41310) );
  ANDN U43676 ( .B(n44359), .A(n44360), .Z(n44357) );
  XOR U43677 ( .A(n39355), .B(n43994), .Z(n36894) );
  XNOR U43678 ( .A(n44361), .B(n44362), .Z(n43994) );
  XOR U43679 ( .A(n44363), .B(n37072), .Z(n44362) );
  XOR U43680 ( .A(n44364), .B(n42921), .Z(n37072) );
  NOR U43681 ( .A(n44365), .B(n43996), .Z(n44364) );
  XOR U43682 ( .A(n37335), .B(n44366), .Z(n44361) );
  XNOR U43683 ( .A(n39939), .B(n38663), .Z(n44366) );
  XNOR U43684 ( .A(n44367), .B(n42910), .Z(n38663) );
  ANDN U43685 ( .B(n41319), .A(n41318), .Z(n44367) );
  XOR U43686 ( .A(n44368), .B(n42913), .Z(n39939) );
  ANDN U43687 ( .B(n41322), .A(n41323), .Z(n44368) );
  XOR U43688 ( .A(n44369), .B(n42924), .Z(n37335) );
  ANDN U43689 ( .B(n41334), .A(n41332), .Z(n44369) );
  XNOR U43690 ( .A(n44370), .B(n44371), .Z(n39355) );
  XNOR U43691 ( .A(n36357), .B(n40084), .Z(n44371) );
  XNOR U43692 ( .A(n44372), .B(n44373), .Z(n40084) );
  NOR U43693 ( .A(n44358), .B(n44359), .Z(n44372) );
  XNOR U43694 ( .A(n44374), .B(n44375), .Z(n36357) );
  NOR U43695 ( .A(n41301), .B(n41303), .Z(n44374) );
  XOR U43696 ( .A(n36552), .B(n44376), .Z(n44370) );
  XNOR U43697 ( .A(n37766), .B(n37923), .Z(n44376) );
  XNOR U43698 ( .A(n44377), .B(n44378), .Z(n37923) );
  NOR U43699 ( .A(n41305), .B(n41306), .Z(n44377) );
  IV U43700 ( .A(n44379), .Z(n41305) );
  XNOR U43701 ( .A(n44380), .B(n44381), .Z(n37766) );
  ANDN U43702 ( .B(n41603), .A(n41605), .Z(n44380) );
  XNOR U43703 ( .A(n44382), .B(n44383), .Z(n36552) );
  NOR U43704 ( .A(n44384), .B(n41312), .Z(n44382) );
  NOR U43705 ( .A(n35451), .B(n34584), .Z(n44356) );
  XOR U43706 ( .A(n44385), .B(n34623), .Z(n34584) );
  XNOR U43707 ( .A(n44386), .B(n44387), .Z(n39633) );
  XNOR U43708 ( .A(n37488), .B(n42779), .Z(n44387) );
  XNOR U43709 ( .A(n44388), .B(n43426), .Z(n42779) );
  XOR U43710 ( .A(n44389), .B(n43418), .Z(n37488) );
  ANDN U43711 ( .B(n43946), .A(n43417), .Z(n44389) );
  IV U43712 ( .A(n44390), .Z(n43417) );
  XNOR U43713 ( .A(n37648), .B(n44391), .Z(n44386) );
  XOR U43714 ( .A(n35942), .B(n43412), .Z(n44391) );
  XNOR U43715 ( .A(n44392), .B(n43434), .Z(n43412) );
  ANDN U43716 ( .B(n43435), .A(n43935), .Z(n44392) );
  XNOR U43717 ( .A(n44393), .B(n43421), .Z(n35942) );
  ANDN U43718 ( .B(n43422), .A(n44394), .Z(n44393) );
  XOR U43719 ( .A(n44395), .B(n43430), .Z(n37648) );
  ANDN U43720 ( .B(n43431), .A(n43943), .Z(n44395) );
  XNOR U43721 ( .A(n44396), .B(n44397), .Z(n43569) );
  XNOR U43722 ( .A(n40219), .B(n41453), .Z(n44397) );
  XNOR U43723 ( .A(n44398), .B(n41178), .Z(n41453) );
  XOR U43724 ( .A(n44399), .B(n43280), .Z(n41178) );
  ANDN U43725 ( .B(n43447), .A(n43927), .Z(n44398) );
  XNOR U43726 ( .A(n44400), .B(n43450), .Z(n40219) );
  IV U43727 ( .A(n41175), .Z(n43450) );
  XOR U43728 ( .A(n44401), .B(n44014), .Z(n41175) );
  ANDN U43729 ( .B(n43930), .A(n43449), .Z(n44400) );
  IV U43730 ( .A(n44402), .Z(n43449) );
  XNOR U43731 ( .A(n33930), .B(n44403), .Z(n44396) );
  XOR U43732 ( .A(n38179), .B(n35795), .Z(n44403) );
  XNOR U43733 ( .A(n44404), .B(n42000), .Z(n35795) );
  XOR U43734 ( .A(n44320), .B(n44405), .Z(n42000) );
  IV U43735 ( .A(n43815), .Z(n44320) );
  ANDN U43736 ( .B(n43439), .A(n43923), .Z(n44404) );
  XOR U43737 ( .A(n44406), .B(n41165), .Z(n38179) );
  IV U43738 ( .A(n43442), .Z(n41165) );
  XNOR U43739 ( .A(n42881), .B(n44407), .Z(n43442) );
  ANDN U43740 ( .B(n43918), .A(n43441), .Z(n44406) );
  XOR U43741 ( .A(n44408), .B(n41169), .Z(n33930) );
  XNOR U43742 ( .A(n44409), .B(n44410), .Z(n41169) );
  ANDN U43743 ( .B(n43445), .A(n43914), .Z(n44408) );
  XNOR U43744 ( .A(n42795), .B(n39186), .Z(n35451) );
  XOR U43745 ( .A(n40997), .B(n39642), .Z(n39186) );
  XNOR U43746 ( .A(n44411), .B(n44412), .Z(n39642) );
  XNOR U43747 ( .A(n39797), .B(n38177), .Z(n44412) );
  XNOR U43748 ( .A(n44413), .B(n42478), .Z(n38177) );
  NOR U43749 ( .A(n41895), .B(n41896), .Z(n44413) );
  IV U43750 ( .A(n44414), .Z(n41895) );
  XNOR U43751 ( .A(n44415), .B(n42483), .Z(n39797) );
  NOR U43752 ( .A(n41906), .B(n41904), .Z(n44415) );
  XOR U43753 ( .A(n39225), .B(n44416), .Z(n44411) );
  XOR U43754 ( .A(n39340), .B(n39400), .Z(n44416) );
  XNOR U43755 ( .A(n44417), .B(n42489), .Z(n39400) );
  ANDN U43756 ( .B(n41914), .A(n44418), .Z(n44417) );
  XOR U43757 ( .A(n44419), .B(n42485), .Z(n39340) );
  NOR U43758 ( .A(n41900), .B(n41899), .Z(n44419) );
  XNOR U43759 ( .A(n44420), .B(n42476), .Z(n39225) );
  ANDN U43760 ( .B(n41908), .A(n41910), .Z(n44420) );
  XNOR U43761 ( .A(n44421), .B(n44422), .Z(n40997) );
  XNOR U43762 ( .A(n39516), .B(n44238), .Z(n44422) );
  XOR U43763 ( .A(n44423), .B(n40816), .Z(n44238) );
  ANDN U43764 ( .B(n42802), .A(n42803), .Z(n44423) );
  ANDN U43765 ( .B(n42794), .A(n42793), .Z(n44424) );
  XOR U43766 ( .A(n39453), .B(n44425), .Z(n44421) );
  XOR U43767 ( .A(n42778), .B(n44426), .Z(n44425) );
  XNOR U43768 ( .A(n44427), .B(n44428), .Z(n42778) );
  XOR U43769 ( .A(n44429), .B(n40812), .Z(n39453) );
  NOR U43770 ( .A(n44430), .B(n44431), .Z(n44429) );
  XNOR U43771 ( .A(n44432), .B(n44431), .Z(n42795) );
  AND U43772 ( .A(n40811), .B(n44430), .Z(n44432) );
  XNOR U43773 ( .A(n44433), .B(n38240), .Z(n31550) );
  XOR U43774 ( .A(n44083), .B(n33917), .Z(n38240) );
  IV U43775 ( .A(n37420), .Z(n33917) );
  XOR U43776 ( .A(n44434), .B(n44435), .Z(n42758) );
  XNOR U43777 ( .A(n39796), .B(n44236), .Z(n44435) );
  XNOR U43778 ( .A(n44436), .B(n44437), .Z(n44236) );
  ANDN U43779 ( .B(n44438), .A(n44439), .Z(n44436) );
  XNOR U43780 ( .A(n44440), .B(n44441), .Z(n39796) );
  ANDN U43781 ( .B(n44442), .A(n44443), .Z(n44440) );
  XOR U43782 ( .A(n44444), .B(n44445), .Z(n44434) );
  XOR U43783 ( .A(n36518), .B(n39849), .Z(n44445) );
  NOR U43784 ( .A(n44448), .B(n44449), .Z(n44446) );
  XNOR U43785 ( .A(n44450), .B(n44451), .Z(n36518) );
  ANDN U43786 ( .B(n44452), .A(n44453), .Z(n44450) );
  XNOR U43787 ( .A(n44454), .B(n44455), .Z(n41685) );
  XNOR U43788 ( .A(n38706), .B(n38454), .Z(n44455) );
  XNOR U43789 ( .A(n44456), .B(n43068), .Z(n38454) );
  ANDN U43790 ( .B(n43067), .A(n44243), .Z(n44456) );
  XOR U43791 ( .A(n44457), .B(n44458), .Z(n38706) );
  XOR U43792 ( .A(n44459), .B(n44460), .Z(n44090) );
  XNOR U43793 ( .A(n44461), .B(n44462), .Z(n41410) );
  XOR U43794 ( .A(n37013), .B(n44463), .Z(n44454) );
  XNOR U43795 ( .A(n37508), .B(n35296), .Z(n44463) );
  XOR U43796 ( .A(n44464), .B(n44465), .Z(n35296) );
  ANDN U43797 ( .B(n41406), .A(n44096), .Z(n44464) );
  XOR U43798 ( .A(n44466), .B(n44467), .Z(n44096) );
  XOR U43799 ( .A(n44468), .B(n44469), .Z(n41406) );
  XNOR U43800 ( .A(n44470), .B(n41417), .Z(n37508) );
  ANDN U43801 ( .B(n41416), .A(n44093), .Z(n44470) );
  XOR U43802 ( .A(n44471), .B(n43716), .Z(n44093) );
  XNOR U43803 ( .A(n44472), .B(n44473), .Z(n41416) );
  ANDN U43804 ( .B(n44085), .A(n44247), .Z(n44474) );
  IV U43805 ( .A(n44087), .Z(n44247) );
  XOR U43806 ( .A(n44476), .B(n42659), .Z(n44087) );
  XNOR U43807 ( .A(n44477), .B(n43067), .Z(n44083) );
  XOR U43808 ( .A(n44478), .B(n44479), .Z(n43067) );
  AND U43809 ( .A(n44244), .B(n44243), .Z(n44477) );
  XNOR U43810 ( .A(n44480), .B(n41745), .Z(n44243) );
  ANDN U43811 ( .B(n34596), .A(n34597), .Z(n44433) );
  XOR U43812 ( .A(n39184), .B(n43955), .Z(n34597) );
  XNOR U43813 ( .A(n44481), .B(n40773), .Z(n43955) );
  ANDN U43814 ( .B(n41482), .A(n44482), .Z(n44481) );
  XOR U43815 ( .A(n44483), .B(n44336), .Z(n41482) );
  XNOR U43816 ( .A(n41725), .B(n40571), .Z(n39184) );
  XNOR U43817 ( .A(n44484), .B(n44485), .Z(n40571) );
  XNOR U43818 ( .A(n38612), .B(n38798), .Z(n44485) );
  XNOR U43819 ( .A(n44486), .B(n40452), .Z(n38798) );
  XNOR U43820 ( .A(n44487), .B(n44488), .Z(n40452) );
  ANDN U43821 ( .B(n40453), .A(n43980), .Z(n44486) );
  XOR U43822 ( .A(n44489), .B(n43671), .Z(n40453) );
  XOR U43823 ( .A(n44490), .B(n41186), .Z(n38612) );
  XOR U43824 ( .A(n44491), .B(n44492), .Z(n41186) );
  ANDN U43825 ( .B(n41185), .A(n43975), .Z(n44490) );
  XNOR U43826 ( .A(n44493), .B(n44494), .Z(n41185) );
  XNOR U43827 ( .A(n39702), .B(n44495), .Z(n44484) );
  XNOR U43828 ( .A(n33921), .B(n38920), .Z(n44495) );
  XOR U43829 ( .A(n44496), .B(n42066), .Z(n38920) );
  XOR U43830 ( .A(n44497), .B(n44498), .Z(n42066) );
  ANDN U43831 ( .B(n42073), .A(n43978), .Z(n44496) );
  XOR U43832 ( .A(n44499), .B(n44500), .Z(n42073) );
  XOR U43833 ( .A(n44501), .B(n40457), .Z(n33921) );
  XOR U43834 ( .A(n44502), .B(n44503), .Z(n40457) );
  NOR U43835 ( .A(n40456), .B(n43972), .Z(n44501) );
  XOR U43836 ( .A(n44504), .B(n44505), .Z(n40456) );
  XNOR U43837 ( .A(n44506), .B(n40460), .Z(n39702) );
  ANDN U43838 ( .B(n40461), .A(n43983), .Z(n44506) );
  XNOR U43839 ( .A(n44507), .B(n43303), .Z(n40461) );
  XOR U43840 ( .A(n44508), .B(n44509), .Z(n41725) );
  XOR U43841 ( .A(n37609), .B(n36436), .Z(n44509) );
  XOR U43842 ( .A(n44510), .B(n40759), .Z(n36436) );
  XOR U43843 ( .A(n44511), .B(n44512), .Z(n40759) );
  AND U43844 ( .A(n43951), .B(n40760), .Z(n44510) );
  XOR U43845 ( .A(n44513), .B(n44514), .Z(n40760) );
  XOR U43846 ( .A(n44515), .B(n44516), .Z(n43951) );
  XNOR U43847 ( .A(n44517), .B(n40763), .Z(n37609) );
  XOR U43848 ( .A(n44518), .B(n44519), .Z(n40763) );
  ANDN U43849 ( .B(n40764), .A(n43296), .Z(n44517) );
  XOR U43850 ( .A(n44520), .B(n44521), .Z(n43296) );
  XOR U43851 ( .A(n44522), .B(n44523), .Z(n40764) );
  XOR U43852 ( .A(n40443), .B(n44524), .Z(n44508) );
  XOR U43853 ( .A(n36713), .B(n39669), .Z(n44524) );
  XNOR U43854 ( .A(n44525), .B(n41480), .Z(n39669) );
  XNOR U43855 ( .A(n44526), .B(n43287), .Z(n41480) );
  ANDN U43856 ( .B(n41492), .A(n43310), .Z(n44525) );
  XNOR U43857 ( .A(n44527), .B(n44528), .Z(n43310) );
  XOR U43858 ( .A(n44529), .B(n43540), .Z(n41492) );
  XNOR U43859 ( .A(n44530), .B(n40769), .Z(n36713) );
  XOR U43860 ( .A(n44531), .B(n41657), .Z(n40769) );
  NOR U43861 ( .A(n40770), .B(n43301), .Z(n44530) );
  XNOR U43862 ( .A(n44532), .B(n44533), .Z(n43301) );
  XOR U43863 ( .A(n44536), .B(n40774), .Z(n40443) );
  XOR U43864 ( .A(n44537), .B(n43552), .Z(n40774) );
  ANDN U43865 ( .B(n44482), .A(n40773), .Z(n44536) );
  XOR U43866 ( .A(n44538), .B(n44539), .Z(n40773) );
  IV U43867 ( .A(n43307), .Z(n44482) );
  XOR U43868 ( .A(n44540), .B(n44541), .Z(n43307) );
  XOR U43869 ( .A(n38113), .B(n42058), .Z(n34596) );
  XOR U43870 ( .A(n44542), .B(n43982), .Z(n42058) );
  XOR U43871 ( .A(n44543), .B(n44544), .Z(n40460) );
  XNOR U43872 ( .A(n44545), .B(n44546), .Z(n40661) );
  XOR U43873 ( .A(n39221), .B(n38827), .Z(n44546) );
  XOR U43874 ( .A(n44547), .B(n43983), .Z(n38827) );
  XNOR U43875 ( .A(n44548), .B(n43644), .Z(n43983) );
  NOR U43876 ( .A(n40459), .B(n43982), .Z(n44547) );
  XOR U43877 ( .A(n44551), .B(n42868), .Z(n40459) );
  XNOR U43878 ( .A(n44552), .B(n43980), .Z(n39221) );
  XNOR U43879 ( .A(n44553), .B(n44182), .Z(n43980) );
  NOR U43880 ( .A(n40451), .B(n42060), .Z(n44552) );
  XNOR U43881 ( .A(n44554), .B(n44516), .Z(n42060) );
  IV U43882 ( .A(n42061), .Z(n40451) );
  XOR U43883 ( .A(n44555), .B(n44556), .Z(n42061) );
  XOR U43884 ( .A(n37170), .B(n44557), .Z(n44545) );
  XNOR U43885 ( .A(n35616), .B(n38092), .Z(n44557) );
  XOR U43886 ( .A(n44558), .B(n43975), .Z(n38092) );
  XOR U43887 ( .A(n44559), .B(n43958), .Z(n43975) );
  AND U43888 ( .A(n42069), .B(n41184), .Z(n44558) );
  XNOR U43889 ( .A(n44560), .B(n41883), .Z(n41184) );
  XOR U43890 ( .A(n44561), .B(n43555), .Z(n42069) );
  XNOR U43891 ( .A(n44562), .B(n43978), .Z(n35616) );
  XOR U43892 ( .A(n44563), .B(n44564), .Z(n43978) );
  NOR U43893 ( .A(n42072), .B(n42065), .Z(n44562) );
  XOR U43894 ( .A(n44565), .B(n43965), .Z(n42065) );
  IV U43895 ( .A(n42067), .Z(n42072) );
  XOR U43896 ( .A(n44254), .B(n44566), .Z(n42067) );
  XNOR U43897 ( .A(n44567), .B(n43972), .Z(n37170) );
  XOR U43898 ( .A(n44568), .B(n42450), .Z(n43972) );
  ANDN U43899 ( .B(n40455), .A(n44310), .Z(n44567) );
  XOR U43900 ( .A(n44223), .B(n44569), .Z(n44310) );
  XOR U43901 ( .A(n44570), .B(n44571), .Z(n40455) );
  XOR U43902 ( .A(n44572), .B(n44573), .Z(n43626) );
  XOR U43903 ( .A(n41494), .B(n41961), .Z(n44573) );
  XOR U43904 ( .A(n44574), .B(n41223), .Z(n41961) );
  XOR U43905 ( .A(n44575), .B(n42659), .Z(n41223) );
  ANDN U43906 ( .B(n41990), .A(n44576), .Z(n44574) );
  XOR U43907 ( .A(n42508), .B(n44577), .Z(n41990) );
  XNOR U43908 ( .A(n44578), .B(n41227), .Z(n41494) );
  XOR U43909 ( .A(n44579), .B(n44580), .Z(n41227) );
  AND U43910 ( .A(n41992), .B(n42955), .Z(n44578) );
  XNOR U43911 ( .A(n44581), .B(n44582), .Z(n41992) );
  XOR U43912 ( .A(n39311), .B(n44583), .Z(n44572) );
  XOR U43913 ( .A(n40124), .B(n41862), .Z(n44583) );
  XNOR U43914 ( .A(n44584), .B(n41214), .Z(n41862) );
  XOR U43915 ( .A(n44585), .B(n44586), .Z(n41214) );
  ANDN U43916 ( .B(n42953), .A(n42952), .Z(n44584) );
  IV U43917 ( .A(n41985), .Z(n42952) );
  XOR U43918 ( .A(n44587), .B(n44588), .Z(n41985) );
  XNOR U43919 ( .A(n44589), .B(n41219), .Z(n40124) );
  XNOR U43920 ( .A(n44590), .B(n43468), .Z(n41219) );
  ANDN U43921 ( .B(n41988), .A(n44591), .Z(n44589) );
  XNOR U43922 ( .A(n44592), .B(n44593), .Z(n41988) );
  XNOR U43923 ( .A(n44594), .B(n41982), .Z(n39311) );
  XOR U43924 ( .A(n44595), .B(n44596), .Z(n41983) );
  XOR U43925 ( .A(n29026), .B(n44597), .Z(n44354) );
  XNOR U43926 ( .A(n31015), .B(n32152), .Z(n44597) );
  XNOR U43927 ( .A(n44598), .B(n36593), .Z(n32152) );
  XNOR U43928 ( .A(n44599), .B(n39528), .Z(n36593) );
  IV U43929 ( .A(n40000), .Z(n39528) );
  XOR U43930 ( .A(n42076), .B(n42146), .Z(n40000) );
  XNOR U43931 ( .A(n44600), .B(n44601), .Z(n42146) );
  XOR U43932 ( .A(n43271), .B(n44339), .Z(n44601) );
  XNOR U43933 ( .A(n44602), .B(n41105), .Z(n44339) );
  XOR U43934 ( .A(n44603), .B(n44604), .Z(n41105) );
  AND U43935 ( .A(n44605), .B(n44351), .Z(n44602) );
  XOR U43936 ( .A(n44606), .B(n41114), .Z(n43271) );
  XOR U43937 ( .A(n44607), .B(n44608), .Z(n41114) );
  ANDN U43938 ( .B(n44344), .A(n44609), .Z(n44606) );
  XNOR U43939 ( .A(n41370), .B(n44610), .Z(n44600) );
  XOR U43940 ( .A(n41841), .B(n40658), .Z(n44610) );
  XOR U43941 ( .A(n44611), .B(n41097), .Z(n40658) );
  XNOR U43942 ( .A(n44612), .B(n43920), .Z(n41097) );
  ANDN U43943 ( .B(n44346), .A(n44613), .Z(n44611) );
  XNOR U43944 ( .A(n44614), .B(n41109), .Z(n41841) );
  XOR U43945 ( .A(n44615), .B(n44270), .Z(n41109) );
  ANDN U43946 ( .B(n44349), .A(n44616), .Z(n44614) );
  XNOR U43947 ( .A(n44617), .B(n41100), .Z(n41370) );
  ANDN U43948 ( .B(n44353), .A(n44620), .Z(n44617) );
  XNOR U43949 ( .A(n44621), .B(n44622), .Z(n42076) );
  XNOR U43950 ( .A(n39602), .B(n39487), .Z(n44622) );
  XNOR U43951 ( .A(n44623), .B(n44624), .Z(n39487) );
  ANDN U43952 ( .B(n44625), .A(n44373), .Z(n44623) );
  XOR U43953 ( .A(n44626), .B(n41307), .Z(n39602) );
  IV U43954 ( .A(n44627), .Z(n41307) );
  NOR U43955 ( .A(n44628), .B(n44378), .Z(n44626) );
  XNOR U43956 ( .A(n38943), .B(n44629), .Z(n44621) );
  XOR U43957 ( .A(n35307), .B(n44630), .Z(n44629) );
  XNOR U43958 ( .A(n44631), .B(n41302), .Z(n35307) );
  ANDN U43959 ( .B(n44632), .A(n44375), .Z(n44631) );
  IV U43960 ( .A(n44633), .Z(n44375) );
  XNOR U43961 ( .A(n44634), .B(n41604), .Z(n38943) );
  NOR U43962 ( .A(n44635), .B(n44381), .Z(n44634) );
  ANDN U43963 ( .B(n34588), .A(n35669), .Z(n44598) );
  XOR U43964 ( .A(n44636), .B(n38277), .Z(n35669) );
  XOR U43965 ( .A(n44637), .B(n39328), .Z(n34588) );
  IV U43966 ( .A(n42711), .Z(n39328) );
  XNOR U43967 ( .A(n44638), .B(n44639), .Z(n40223) );
  XNOR U43968 ( .A(n43273), .B(n40270), .Z(n44639) );
  XOR U43969 ( .A(n44640), .B(n41354), .Z(n40270) );
  NOR U43970 ( .A(n44641), .B(n44642), .Z(n44640) );
  XOR U43971 ( .A(n44643), .B(n41345), .Z(n43273) );
  NOR U43972 ( .A(n44644), .B(n44645), .Z(n44643) );
  XOR U43973 ( .A(n38970), .B(n44646), .Z(n44638) );
  XOR U43974 ( .A(n40693), .B(n38720), .Z(n44646) );
  XOR U43975 ( .A(n44647), .B(n41342), .Z(n38720) );
  ANDN U43976 ( .B(n44648), .A(n44649), .Z(n44647) );
  XNOR U43977 ( .A(n44650), .B(n41358), .Z(n40693) );
  NOR U43978 ( .A(n44651), .B(n44652), .Z(n44650) );
  XOR U43979 ( .A(n44653), .B(n41350), .Z(n38970) );
  NOR U43980 ( .A(n44654), .B(n44655), .Z(n44653) );
  XNOR U43981 ( .A(n44657), .B(n35447), .Z(n31015) );
  XNOR U43982 ( .A(n38616), .B(n42933), .Z(n35447) );
  XOR U43983 ( .A(n44658), .B(n43880), .Z(n42933) );
  ANDN U43984 ( .B(n44212), .A(n43357), .Z(n44658) );
  IV U43985 ( .A(n44213), .Z(n43357) );
  XNOR U43986 ( .A(n44659), .B(n44660), .Z(n44213) );
  ANDN U43987 ( .B(n34579), .A(n34580), .Z(n44657) );
  XOR U43988 ( .A(n37314), .B(n43104), .Z(n34580) );
  XNOR U43989 ( .A(n44661), .B(n44662), .Z(n43104) );
  ANDN U43990 ( .B(n40393), .A(n43113), .Z(n44661) );
  XOR U43991 ( .A(n44663), .B(n44664), .Z(n40393) );
  XOR U43992 ( .A(n42592), .B(n42551), .Z(n37314) );
  XNOR U43993 ( .A(n44665), .B(n44666), .Z(n42551) );
  XOR U43994 ( .A(n38141), .B(n44155), .Z(n44666) );
  XOR U43995 ( .A(n44667), .B(n41268), .Z(n44155) );
  XOR U43996 ( .A(n43463), .B(n44668), .Z(n41268) );
  ANDN U43997 ( .B(n43035), .A(n44160), .Z(n44667) );
  XNOR U43998 ( .A(n44669), .B(n43846), .Z(n44160) );
  XOR U43999 ( .A(n43587), .B(n44670), .Z(n43035) );
  XNOR U44000 ( .A(n44671), .B(n41262), .Z(n38141) );
  XOR U44001 ( .A(n44672), .B(n44673), .Z(n41262) );
  ANDN U44002 ( .B(n43076), .A(n43037), .Z(n44671) );
  IV U44003 ( .A(n43077), .Z(n43037) );
  XOR U44004 ( .A(n44674), .B(n43298), .Z(n43077) );
  XOR U44005 ( .A(n44675), .B(n44676), .Z(n43076) );
  XOR U44006 ( .A(n37471), .B(n44677), .Z(n44665) );
  XOR U44007 ( .A(n37881), .B(n42965), .Z(n44677) );
  XNOR U44008 ( .A(n44678), .B(n41258), .Z(n42965) );
  ANDN U44009 ( .B(n43030), .A(n44170), .Z(n44678) );
  IV U44010 ( .A(n43086), .Z(n44170) );
  XOR U44011 ( .A(n44681), .B(n44682), .Z(n43086) );
  XNOR U44012 ( .A(n44683), .B(n44488), .Z(n43030) );
  XNOR U44013 ( .A(n44684), .B(n41868), .Z(n37881) );
  XNOR U44014 ( .A(n44685), .B(n44686), .Z(n41868) );
  XOR U44015 ( .A(n44687), .B(n43543), .Z(n43028) );
  XNOR U44016 ( .A(n44688), .B(n44689), .Z(n43082) );
  XNOR U44017 ( .A(n41271), .B(n44690), .Z(n37471) );
  XNOR U44018 ( .A(n4549), .B(n44691), .Z(n44690) );
  NANDN U44019 ( .A(n43072), .B(n43033), .Z(n44691) );
  XNOR U44020 ( .A(n42319), .B(n44692), .Z(n43033) );
  XOR U44021 ( .A(n44693), .B(n44694), .Z(n43072) );
  XOR U44022 ( .A(n44695), .B(n42337), .Z(n41271) );
  IV U44023 ( .A(n44410), .Z(n42337) );
  XOR U44024 ( .A(n44696), .B(n44697), .Z(n42592) );
  XNOR U44025 ( .A(n38996), .B(n39333), .Z(n44697) );
  XOR U44026 ( .A(n44698), .B(n40390), .Z(n39333) );
  ANDN U44027 ( .B(n43096), .A(n43020), .Z(n44698) );
  IV U44028 ( .A(n43097), .Z(n43020) );
  XOR U44029 ( .A(n44699), .B(n43562), .Z(n43097) );
  XOR U44030 ( .A(n44700), .B(n40395), .Z(n38996) );
  AND U44031 ( .A(n44662), .B(n43113), .Z(n44700) );
  XNOR U44032 ( .A(n44701), .B(n44009), .Z(n43113) );
  XOR U44033 ( .A(n42027), .B(n44702), .Z(n44696) );
  XOR U44034 ( .A(n42048), .B(n39026), .Z(n44702) );
  XNOR U44035 ( .A(n44703), .B(n40385), .Z(n39026) );
  AND U44036 ( .A(n43106), .B(n43015), .Z(n44703) );
  XOR U44037 ( .A(n44704), .B(n44705), .Z(n43015) );
  XNOR U44038 ( .A(n44706), .B(n43039), .Z(n42048) );
  AND U44039 ( .A(n43110), .B(n43022), .Z(n44706) );
  XOR U44040 ( .A(n44707), .B(n44163), .Z(n43022) );
  XNOR U44041 ( .A(n44708), .B(n42573), .Z(n42027) );
  XNOR U44042 ( .A(n44709), .B(n44710), .Z(n43012) );
  XOR U44043 ( .A(n44711), .B(n36420), .Z(n34579) );
  XOR U44044 ( .A(n44712), .B(n35454), .Z(n29026) );
  XOR U44045 ( .A(n39848), .B(n44444), .Z(n35454) );
  XOR U44046 ( .A(n44713), .B(n44714), .Z(n44444) );
  NOR U44047 ( .A(n44715), .B(n44716), .Z(n44713) );
  IV U44048 ( .A(n36519), .Z(n39848) );
  XOR U44049 ( .A(n39632), .B(n38708), .Z(n36519) );
  XNOR U44050 ( .A(n44717), .B(n44718), .Z(n38708) );
  XOR U44051 ( .A(n41182), .B(n39467), .Z(n44718) );
  XOR U44052 ( .A(n44719), .B(n44720), .Z(n39467) );
  ANDN U44053 ( .B(n44441), .A(n44442), .Z(n44719) );
  XNOR U44054 ( .A(n44721), .B(n44722), .Z(n41182) );
  ANDN U44055 ( .B(n44716), .A(n44714), .Z(n44721) );
  XNOR U44056 ( .A(n37724), .B(n44723), .Z(n44717) );
  XOR U44057 ( .A(n42101), .B(n39668), .Z(n44723) );
  XNOR U44058 ( .A(n44724), .B(n44725), .Z(n39668) );
  ANDN U44059 ( .B(n44451), .A(n44452), .Z(n44724) );
  XNOR U44060 ( .A(n44726), .B(n44727), .Z(n42101) );
  NOR U44061 ( .A(n44728), .B(n44438), .Z(n44726) );
  XOR U44062 ( .A(n44729), .B(n44730), .Z(n37724) );
  ANDN U44063 ( .B(n44449), .A(n44447), .Z(n44729) );
  XOR U44064 ( .A(n44731), .B(n44732), .Z(n39632) );
  XNOR U44065 ( .A(n35372), .B(n40828), .Z(n44732) );
  XNOR U44066 ( .A(n44733), .B(n42107), .Z(n40828) );
  ANDN U44067 ( .B(n42108), .A(n42776), .Z(n44733) );
  XNOR U44068 ( .A(n43298), .B(n44734), .Z(n42108) );
  XOR U44069 ( .A(n44735), .B(n44736), .Z(n35372) );
  XNOR U44070 ( .A(n37194), .B(n44737), .Z(n44731) );
  XOR U44071 ( .A(n38940), .B(n37803), .Z(n44737) );
  XNOR U44072 ( .A(n44738), .B(n42121), .Z(n37803) );
  ANDN U44073 ( .B(n42120), .A(n44739), .Z(n44738) );
  XOR U44074 ( .A(n44740), .B(n44741), .Z(n42120) );
  XOR U44075 ( .A(n44742), .B(n42117), .Z(n38940) );
  ANDN U44076 ( .B(n42116), .A(n42773), .Z(n44742) );
  XNOR U44077 ( .A(n44743), .B(n44744), .Z(n42116) );
  XNOR U44078 ( .A(n44745), .B(n42112), .Z(n37194) );
  ANDN U44079 ( .B(n42113), .A(n42763), .Z(n44745) );
  XOR U44080 ( .A(n44746), .B(n44747), .Z(n42113) );
  NOR U44081 ( .A(n34592), .B(n34593), .Z(n44712) );
  XOR U44082 ( .A(n39204), .B(n37939), .Z(n34593) );
  XNOR U44083 ( .A(n39969), .B(n39105), .Z(n37939) );
  XOR U44084 ( .A(n44748), .B(n44749), .Z(n39105) );
  XNOR U44085 ( .A(n38873), .B(n37109), .Z(n44749) );
  XOR U44086 ( .A(n44750), .B(n40604), .Z(n37109) );
  ANDN U44087 ( .B(n40635), .A(n40636), .Z(n44750) );
  XOR U44088 ( .A(n44751), .B(n44523), .Z(n40636) );
  XNOR U44089 ( .A(n44752), .B(n40600), .Z(n38873) );
  ANDN U44090 ( .B(n41596), .A(n44753), .Z(n44752) );
  XNOR U44091 ( .A(n44754), .B(n44755), .Z(n44748) );
  XOR U44092 ( .A(n35088), .B(n39520), .Z(n44755) );
  XNOR U44093 ( .A(n44756), .B(n41600), .Z(n39520) );
  ANDN U44094 ( .B(n39201), .A(n44757), .Z(n44756) );
  XNOR U44095 ( .A(n44758), .B(n44759), .Z(n39201) );
  XNOR U44096 ( .A(n44760), .B(n40611), .Z(n35088) );
  XOR U44097 ( .A(n44761), .B(n44762), .Z(n39208) );
  XOR U44098 ( .A(n44763), .B(n44764), .Z(n39969) );
  XNOR U44099 ( .A(n41799), .B(n44765), .Z(n44764) );
  XNOR U44100 ( .A(n44766), .B(n41556), .Z(n41799) );
  ANDN U44101 ( .B(n40500), .A(n40501), .Z(n44766) );
  XNOR U44102 ( .A(n44767), .B(n44768), .Z(n40501) );
  XNOR U44103 ( .A(n38945), .B(n44769), .Z(n44763) );
  XOR U44104 ( .A(n41140), .B(n39326), .Z(n44769) );
  XNOR U44105 ( .A(n44770), .B(n41563), .Z(n39326) );
  ANDN U44106 ( .B(n40496), .A(n40497), .Z(n44770) );
  XOR U44107 ( .A(n44771), .B(n44494), .Z(n40497) );
  XNOR U44108 ( .A(n44772), .B(n41559), .Z(n41140) );
  ANDN U44109 ( .B(n40487), .A(n40489), .Z(n44772) );
  XOR U44110 ( .A(n44773), .B(n44774), .Z(n40489) );
  XOR U44111 ( .A(n44775), .B(n42167), .Z(n38945) );
  ANDN U44112 ( .B(n40491), .A(n40492), .Z(n44775) );
  XOR U44113 ( .A(n44776), .B(n44777), .Z(n40492) );
  XOR U44114 ( .A(n44778), .B(n44753), .Z(n39204) );
  NOR U44115 ( .A(n40598), .B(n41596), .Z(n44778) );
  XOR U44116 ( .A(n43298), .B(n44779), .Z(n41596) );
  XOR U44117 ( .A(n44780), .B(n44596), .Z(n40598) );
  XNOR U44118 ( .A(n38817), .B(n42655), .Z(n34592) );
  XNOR U44119 ( .A(n44781), .B(n40895), .Z(n42655) );
  AND U44120 ( .A(n41035), .B(n41655), .Z(n44781) );
  XOR U44121 ( .A(n43602), .B(n44782), .Z(n41035) );
  IV U44122 ( .A(n44783), .Z(n43602) );
  XNOR U44123 ( .A(n44784), .B(n35469), .Z(n35990) );
  XOR U44124 ( .A(n44785), .B(n36420), .Z(n35469) );
  XNOR U44125 ( .A(n44786), .B(n44787), .Z(n36420) );
  ANDN U44126 ( .B(n34602), .A(n44152), .Z(n44784) );
  XOR U44127 ( .A(n39325), .B(n44765), .Z(n44152) );
  XNOR U44128 ( .A(n44788), .B(n41566), .Z(n44765) );
  ANDN U44129 ( .B(n40504), .A(n40506), .Z(n44788) );
  XOR U44130 ( .A(n44789), .B(n44790), .Z(n40506) );
  IV U44131 ( .A(n38944), .Z(n39325) );
  XOR U44132 ( .A(n44791), .B(n39356), .Z(n38944) );
  XNOR U44133 ( .A(n44792), .B(n44793), .Z(n39356) );
  XNOR U44134 ( .A(n35081), .B(n38364), .Z(n44793) );
  XNOR U44135 ( .A(n44794), .B(n44795), .Z(n38364) );
  ANDN U44136 ( .B(n41112), .A(n41113), .Z(n44794) );
  XOR U44137 ( .A(n44796), .B(n44797), .Z(n41113) );
  XNOR U44138 ( .A(n44798), .B(n44605), .Z(n35081) );
  ANDN U44139 ( .B(n41104), .A(n41106), .Z(n44798) );
  XOR U44140 ( .A(n44799), .B(n44800), .Z(n41106) );
  XNOR U44141 ( .A(n37689), .B(n44801), .Z(n44792) );
  XOR U44142 ( .A(n44802), .B(n35168), .Z(n44801) );
  XOR U44143 ( .A(n44803), .B(n44616), .Z(n35168) );
  IV U44144 ( .A(n44804), .Z(n44616) );
  AND U44145 ( .A(n41110), .B(n41108), .Z(n44803) );
  XOR U44146 ( .A(n44805), .B(n44806), .Z(n41110) );
  XOR U44147 ( .A(n44807), .B(n44620), .Z(n37689) );
  IV U44148 ( .A(n44808), .Z(n44620) );
  ANDN U44149 ( .B(n41099), .A(n41101), .Z(n44807) );
  XOR U44150 ( .A(n44809), .B(n44810), .Z(n41101) );
  XOR U44151 ( .A(n42715), .B(n40540), .Z(n34602) );
  XNOR U44152 ( .A(n40919), .B(n44811), .Z(n40540) );
  XOR U44153 ( .A(n44812), .B(n44813), .Z(n40919) );
  XNOR U44154 ( .A(n38779), .B(n39793), .Z(n44813) );
  XNOR U44155 ( .A(n44814), .B(n43229), .Z(n39793) );
  NOR U44156 ( .A(n43230), .B(n42727), .Z(n44814) );
  XNOR U44157 ( .A(n44815), .B(n44816), .Z(n43230) );
  XOR U44158 ( .A(n44817), .B(n43234), .Z(n38779) );
  XNOR U44159 ( .A(n38828), .B(n44819), .Z(n44812) );
  XOR U44160 ( .A(n36778), .B(n38983), .Z(n44819) );
  XNOR U44161 ( .A(n44820), .B(n43222), .Z(n38983) );
  NOR U44162 ( .A(n42722), .B(n42724), .Z(n44820) );
  XNOR U44163 ( .A(n44821), .B(n42206), .Z(n42722) );
  XNOR U44164 ( .A(n44822), .B(n44823), .Z(n36778) );
  NOR U44165 ( .A(n42730), .B(n42731), .Z(n44822) );
  XNOR U44166 ( .A(n44824), .B(n43226), .Z(n38828) );
  NOR U44167 ( .A(n42717), .B(n42718), .Z(n44824) );
  XOR U44168 ( .A(n44825), .B(n44263), .Z(n42717) );
  XNOR U44169 ( .A(n44826), .B(n43233), .Z(n42715) );
  XNOR U44170 ( .A(n44827), .B(n43323), .Z(n43233) );
  AND U44171 ( .A(n44818), .B(n44828), .Z(n44826) );
  ANDN U44172 ( .B(n28990), .A(n27610), .Z(n44074) );
  XNOR U44173 ( .A(n38380), .B(n34115), .Z(n27610) );
  XNOR U44174 ( .A(n34221), .B(n38756), .Z(n34115) );
  XOR U44175 ( .A(n44829), .B(n44830), .Z(n38756) );
  XOR U44176 ( .A(n31696), .B(n29915), .Z(n44830) );
  XOR U44177 ( .A(n44831), .B(n40273), .Z(n29915) );
  XOR U44178 ( .A(n39787), .B(n44832), .Z(n40273) );
  IV U44179 ( .A(n37679), .Z(n39787) );
  XOR U44180 ( .A(n43790), .B(n43725), .Z(n37679) );
  XOR U44181 ( .A(n44833), .B(n44834), .Z(n43725) );
  XNOR U44182 ( .A(n37037), .B(n36208), .Z(n44834) );
  XOR U44183 ( .A(n44835), .B(n40914), .Z(n36208) );
  XOR U44184 ( .A(n44836), .B(n44837), .Z(n40914) );
  ANDN U44185 ( .B(n40682), .A(n40683), .Z(n44835) );
  XOR U44186 ( .A(n44838), .B(n44839), .Z(n40683) );
  XOR U44187 ( .A(n44840), .B(n44841), .Z(n40682) );
  XNOR U44188 ( .A(n44842), .B(n41073), .Z(n37037) );
  XOR U44189 ( .A(n43073), .B(n44843), .Z(n41073) );
  ANDN U44190 ( .B(n40679), .A(n41075), .Z(n44842) );
  XOR U44191 ( .A(n44581), .B(n44844), .Z(n41075) );
  IV U44192 ( .A(n44845), .Z(n44581) );
  XOR U44193 ( .A(n44846), .B(n44847), .Z(n40679) );
  XOR U44194 ( .A(n36405), .B(n44848), .Z(n44833) );
  XOR U44195 ( .A(n38808), .B(n38712), .Z(n44848) );
  XNOR U44196 ( .A(n44849), .B(n40022), .Z(n38712) );
  XNOR U44197 ( .A(n44850), .B(n44851), .Z(n40022) );
  ANDN U44198 ( .B(n43727), .A(n40023), .Z(n44849) );
  XOR U44199 ( .A(n43577), .B(n44852), .Z(n40023) );
  XNOR U44200 ( .A(n42537), .B(n44853), .Z(n43727) );
  XNOR U44201 ( .A(n44854), .B(n40019), .Z(n38808) );
  XOR U44202 ( .A(n44855), .B(n44856), .Z(n40019) );
  NOR U44203 ( .A(n40688), .B(n40018), .Z(n44854) );
  XNOR U44204 ( .A(n44857), .B(n43895), .Z(n40018) );
  XOR U44205 ( .A(n44858), .B(n44859), .Z(n40688) );
  XOR U44206 ( .A(n44860), .B(n40205), .Z(n36405) );
  XOR U44207 ( .A(n44861), .B(n44862), .Z(n40205) );
  ANDN U44208 ( .B(n40691), .A(n40204), .Z(n44860) );
  XNOR U44209 ( .A(n44863), .B(n40853), .Z(n40204) );
  XOR U44210 ( .A(n44864), .B(n44865), .Z(n40691) );
  XNOR U44211 ( .A(n44866), .B(n44867), .Z(n43790) );
  XNOR U44212 ( .A(n38584), .B(n39628), .Z(n44867) );
  XOR U44213 ( .A(n44868), .B(n40113), .Z(n39628) );
  XOR U44214 ( .A(n44869), .B(n44870), .Z(n40113) );
  ANDN U44215 ( .B(n40114), .A(n44871), .Z(n44868) );
  XOR U44216 ( .A(n44872), .B(n40702), .Z(n38584) );
  XOR U44217 ( .A(n44873), .B(n44874), .Z(n40702) );
  ANDN U44218 ( .B(n40701), .A(n44875), .Z(n44872) );
  XNOR U44219 ( .A(n38085), .B(n44876), .Z(n44866) );
  XOR U44220 ( .A(n40008), .B(n37182), .Z(n44876) );
  XOR U44221 ( .A(n44877), .B(n42637), .Z(n37182) );
  IV U44222 ( .A(n40103), .Z(n42637) );
  XOR U44223 ( .A(n44878), .B(n41594), .Z(n40103) );
  AND U44224 ( .A(n44879), .B(n40104), .Z(n44877) );
  XOR U44225 ( .A(n44880), .B(n40108), .Z(n40008) );
  XOR U44226 ( .A(n44881), .B(n44882), .Z(n40108) );
  ANDN U44227 ( .B(n44883), .A(n40107), .Z(n44880) );
  XNOR U44228 ( .A(n44884), .B(n40117), .Z(n38085) );
  XOR U44229 ( .A(n44885), .B(n44886), .Z(n40117) );
  ANDN U44230 ( .B(n40118), .A(n44887), .Z(n44884) );
  NOR U44231 ( .A(n35882), .B(n35883), .Z(n44831) );
  XNOR U44232 ( .A(n42408), .B(n36362), .Z(n35883) );
  IV U44233 ( .A(n39014), .Z(n36362) );
  XOR U44234 ( .A(n40149), .B(n40943), .Z(n39014) );
  XNOR U44235 ( .A(n44888), .B(n44889), .Z(n40943) );
  XNOR U44236 ( .A(n39350), .B(n44311), .Z(n44889) );
  XNOR U44237 ( .A(n44890), .B(n42434), .Z(n44311) );
  NOR U44238 ( .A(n44064), .B(n44065), .Z(n44890) );
  XNOR U44239 ( .A(n44891), .B(n44892), .Z(n39350) );
  XOR U44240 ( .A(n39161), .B(n44893), .Z(n44888) );
  XOR U44241 ( .A(n39974), .B(n38321), .Z(n44893) );
  XNOR U44242 ( .A(n44894), .B(n42443), .Z(n38321) );
  XNOR U44243 ( .A(n44895), .B(n44896), .Z(n39974) );
  NOR U44244 ( .A(n44072), .B(n44073), .Z(n44895) );
  XNOR U44245 ( .A(n44897), .B(n42430), .Z(n39161) );
  ANDN U44246 ( .B(n44056), .A(n44057), .Z(n44897) );
  XOR U44247 ( .A(n44898), .B(n44899), .Z(n40149) );
  XNOR U44248 ( .A(n38406), .B(n37846), .Z(n44899) );
  XNOR U44249 ( .A(n44900), .B(n44010), .Z(n37846) );
  XOR U44250 ( .A(n44901), .B(n44494), .Z(n40722) );
  XNOR U44251 ( .A(n44902), .B(n44006), .Z(n38406) );
  NOR U44252 ( .A(n40726), .B(n42782), .Z(n44902) );
  XOR U44253 ( .A(n42546), .B(n44903), .Z(n40726) );
  XOR U44254 ( .A(n44904), .B(n44905), .Z(n44898) );
  XOR U44255 ( .A(n36700), .B(n39322), .Z(n44905) );
  XNOR U44256 ( .A(n44906), .B(n44015), .Z(n39322) );
  IV U44257 ( .A(n44907), .Z(n44015) );
  ANDN U44258 ( .B(n42416), .A(n40713), .Z(n44906) );
  XOR U44259 ( .A(n40856), .B(n44908), .Z(n40713) );
  XNOR U44260 ( .A(n44909), .B(n44021), .Z(n36700) );
  ANDN U44261 ( .B(n44910), .A(n44911), .Z(n44909) );
  XNOR U44262 ( .A(n44912), .B(n44913), .Z(n42408) );
  ANDN U44263 ( .B(n40720), .A(n44910), .Z(n44912) );
  IV U44264 ( .A(n40718), .Z(n44910) );
  XOR U44265 ( .A(n44914), .B(n44915), .Z(n40718) );
  XOR U44266 ( .A(n44459), .B(n44916), .Z(n40720) );
  IV U44267 ( .A(n40330), .Z(n35882) );
  XOR U44268 ( .A(n43634), .B(n39389), .Z(n40330) );
  XNOR U44269 ( .A(n44917), .B(n44918), .Z(n41141) );
  XOR U44270 ( .A(n34639), .B(n39010), .Z(n44918) );
  XOR U44271 ( .A(n44920), .B(n44921), .Z(n42741) );
  ANDN U44272 ( .B(n42742), .A(n43204), .Z(n44919) );
  XOR U44273 ( .A(n44922), .B(n44173), .Z(n43204) );
  XNOR U44274 ( .A(n44923), .B(n44186), .Z(n42742) );
  XNOR U44275 ( .A(n44924), .B(n42751), .Z(n34639) );
  XOR U44276 ( .A(n44925), .B(n43574), .Z(n42751) );
  ANDN U44277 ( .B(n43638), .A(n42750), .Z(n44924) );
  XOR U44278 ( .A(n42712), .B(n44926), .Z(n44917) );
  XNOR U44279 ( .A(n41686), .B(n39854), .Z(n44926) );
  XNOR U44280 ( .A(n44927), .B(n42746), .Z(n39854) );
  XOR U44281 ( .A(n44928), .B(n42153), .Z(n42746) );
  ANDN U44282 ( .B(n42747), .A(n43212), .Z(n44927) );
  XNOR U44283 ( .A(n44929), .B(n44930), .Z(n43212) );
  XNOR U44284 ( .A(n44931), .B(n44932), .Z(n42747) );
  XOR U44285 ( .A(n44933), .B(n43714), .Z(n41686) );
  IV U44286 ( .A(n42755), .Z(n43714) );
  XNOR U44287 ( .A(n44934), .B(n43088), .Z(n42755) );
  ANDN U44288 ( .B(n43207), .A(n42754), .Z(n44933) );
  XNOR U44289 ( .A(n44935), .B(n44936), .Z(n42754) );
  XOR U44290 ( .A(n44937), .B(n44938), .Z(n43207) );
  XNOR U44291 ( .A(n44939), .B(n42737), .Z(n42712) );
  XOR U44292 ( .A(n43559), .B(n44940), .Z(n42737) );
  ANDN U44293 ( .B(n42738), .A(n43215), .Z(n44939) );
  XNOR U44294 ( .A(n44941), .B(n43962), .Z(n43215) );
  XOR U44295 ( .A(n44942), .B(n44943), .Z(n42738) );
  XOR U44296 ( .A(n44946), .B(n42496), .Z(n42750) );
  NOR U44297 ( .A(n43639), .B(n43638), .Z(n44945) );
  XOR U44298 ( .A(n44948), .B(n41745), .Z(n43639) );
  XNOR U44299 ( .A(n44949), .B(n40070), .Z(n31696) );
  XNOR U44300 ( .A(n35583), .B(n44950), .Z(n40070) );
  XNOR U44301 ( .A(n40615), .B(n40512), .Z(n35583) );
  XOR U44302 ( .A(n44951), .B(n44952), .Z(n40512) );
  XOR U44303 ( .A(n40795), .B(n44953), .Z(n44952) );
  XNOR U44304 ( .A(n44954), .B(n42971), .Z(n40795) );
  IV U44305 ( .A(n44955), .Z(n42971) );
  NOR U44306 ( .A(n44956), .B(n41001), .Z(n44954) );
  XOR U44307 ( .A(n36449), .B(n44957), .Z(n44951) );
  XNOR U44308 ( .A(n39617), .B(n37001), .Z(n44957) );
  ANDN U44309 ( .B(n44959), .A(n41005), .Z(n44958) );
  XNOR U44310 ( .A(n44960), .B(n42976), .Z(n39617) );
  IV U44311 ( .A(n44961), .Z(n42976) );
  ANDN U44312 ( .B(n44962), .A(n44963), .Z(n44960) );
  XOR U44313 ( .A(n44964), .B(n42978), .Z(n36449) );
  XOR U44314 ( .A(n44966), .B(n44967), .Z(n40615) );
  XOR U44315 ( .A(n38595), .B(n39816), .Z(n44967) );
  XOR U44316 ( .A(n44968), .B(n42998), .Z(n39816) );
  XNOR U44317 ( .A(n44969), .B(n44970), .Z(n42998) );
  NOR U44318 ( .A(n44127), .B(n44971), .Z(n44968) );
  XOR U44319 ( .A(n44972), .B(n43002), .Z(n38595) );
  XOR U44320 ( .A(n44973), .B(n42340), .Z(n43002) );
  NOR U44321 ( .A(n44974), .B(n44975), .Z(n44972) );
  XNOR U44322 ( .A(n39579), .B(n44976), .Z(n44966) );
  XOR U44323 ( .A(n39047), .B(n37173), .Z(n44976) );
  XOR U44324 ( .A(n44978), .B(n44979), .Z(n42994) );
  NOR U44325 ( .A(n44132), .B(n44980), .Z(n44977) );
  XNOR U44326 ( .A(n44981), .B(n42985), .Z(n39047) );
  IV U44327 ( .A(n44135), .Z(n42985) );
  XOR U44328 ( .A(n44497), .B(n44982), .Z(n44135) );
  NOR U44329 ( .A(n44134), .B(n44983), .Z(n44981) );
  XOR U44330 ( .A(n44984), .B(n42989), .Z(n39579) );
  XOR U44331 ( .A(n44985), .B(n44986), .Z(n42989) );
  NOR U44332 ( .A(n44137), .B(n44987), .Z(n44984) );
  NOR U44333 ( .A(n40071), .B(n37463), .Z(n44949) );
  XOR U44334 ( .A(n44988), .B(n39284), .Z(n37463) );
  IV U44335 ( .A(n38865), .Z(n39284) );
  XOR U44336 ( .A(n41716), .B(n43394), .Z(n38865) );
  XNOR U44337 ( .A(n44989), .B(n44990), .Z(n43394) );
  XNOR U44338 ( .A(n39129), .B(n41915), .Z(n44990) );
  XNOR U44339 ( .A(n44991), .B(n43263), .Z(n41915) );
  IV U44340 ( .A(n44992), .Z(n43263) );
  ANDN U44341 ( .B(n40979), .A(n43262), .Z(n44991) );
  XNOR U44342 ( .A(n44993), .B(n43258), .Z(n39129) );
  ANDN U44343 ( .B(n43259), .A(n44994), .Z(n44993) );
  XNOR U44344 ( .A(n38373), .B(n44995), .Z(n44989) );
  XOR U44345 ( .A(n37165), .B(n43235), .Z(n44995) );
  XOR U44346 ( .A(n44996), .B(n43266), .Z(n43235) );
  NOR U44347 ( .A(n43265), .B(n41361), .Z(n44996) );
  XNOR U44348 ( .A(n44997), .B(n43254), .Z(n37165) );
  ANDN U44349 ( .B(n43255), .A(n40985), .Z(n44997) );
  XNOR U44350 ( .A(n44998), .B(n43269), .Z(n38373) );
  ANDN U44351 ( .B(n43270), .A(n40989), .Z(n44998) );
  XNOR U44352 ( .A(n44999), .B(n45000), .Z(n41716) );
  XNOR U44353 ( .A(n41515), .B(n39598), .Z(n45000) );
  XNOR U44354 ( .A(n45001), .B(n42354), .Z(n39598) );
  XNOR U44355 ( .A(n45002), .B(n44710), .Z(n42354) );
  XNOR U44356 ( .A(n45004), .B(n43008), .Z(n41515) );
  XNOR U44357 ( .A(n45005), .B(n45006), .Z(n43008) );
  ANDN U44358 ( .B(n45007), .A(n43239), .Z(n45004) );
  XNOR U44359 ( .A(n40353), .B(n45008), .Z(n44999) );
  XOR U44360 ( .A(n37317), .B(n39054), .Z(n45008) );
  XNOR U44361 ( .A(n45009), .B(n42350), .Z(n39054) );
  XNOR U44362 ( .A(n45010), .B(n45011), .Z(n42350) );
  XNOR U44363 ( .A(n45013), .B(n42361), .Z(n37317) );
  XNOR U44364 ( .A(n45014), .B(n45015), .Z(n42361) );
  XNOR U44365 ( .A(n45017), .B(n43243), .Z(n40353) );
  XOR U44366 ( .A(n45019), .B(n35579), .Z(n40071) );
  XOR U44367 ( .A(n42784), .B(n45020), .Z(n35579) );
  XOR U44368 ( .A(n45021), .B(n45022), .Z(n42784) );
  XOR U44369 ( .A(n39276), .B(n38456), .Z(n45022) );
  XOR U44370 ( .A(n45023), .B(n44715), .Z(n38456) );
  NOR U44371 ( .A(n44722), .B(n45024), .Z(n45023) );
  XNOR U44372 ( .A(n45025), .B(n44453), .Z(n39276) );
  NOR U44373 ( .A(n45026), .B(n44725), .Z(n45025) );
  XOR U44374 ( .A(n45027), .B(n45028), .Z(n45021) );
  XOR U44375 ( .A(n39218), .B(n45029), .Z(n45028) );
  XNOR U44376 ( .A(n45030), .B(n44448), .Z(n39218) );
  NOR U44377 ( .A(n44730), .B(n45031), .Z(n45030) );
  IV U44378 ( .A(n45032), .Z(n44730) );
  XOR U44379 ( .A(n32905), .B(n45033), .Z(n44829) );
  XOR U44380 ( .A(n34357), .B(n32962), .Z(n45033) );
  XOR U44381 ( .A(n45034), .B(n40064), .Z(n32962) );
  XOR U44382 ( .A(n39962), .B(n39295), .Z(n40064) );
  XOR U44383 ( .A(n44811), .B(n40579), .Z(n39295) );
  XNOR U44384 ( .A(n45035), .B(n45036), .Z(n40579) );
  XNOR U44385 ( .A(n38886), .B(n40521), .Z(n45036) );
  XNOR U44386 ( .A(n45037), .B(n44649), .Z(n40521) );
  ANDN U44387 ( .B(n41340), .A(n41341), .Z(n45037) );
  XNOR U44388 ( .A(n45038), .B(n44641), .Z(n38886) );
  ANDN U44389 ( .B(n41353), .A(n45039), .Z(n45038) );
  XOR U44390 ( .A(n45040), .B(n45041), .Z(n45035) );
  XOR U44391 ( .A(n41082), .B(n38326), .Z(n45041) );
  XNOR U44392 ( .A(n45042), .B(n44652), .Z(n38326) );
  XNOR U44393 ( .A(n45043), .B(n44654), .Z(n41082) );
  XOR U44394 ( .A(n45044), .B(n45045), .Z(n44811) );
  XNOR U44395 ( .A(n34627), .B(n45046), .Z(n45045) );
  XOR U44396 ( .A(n45047), .B(n45048), .Z(n34627) );
  ANDN U44397 ( .B(n45049), .A(n45050), .Z(n45047) );
  XNOR U44398 ( .A(n39382), .B(n45051), .Z(n45044) );
  XOR U44399 ( .A(n39920), .B(n40663), .Z(n45051) );
  XNOR U44400 ( .A(n45052), .B(n45053), .Z(n40663) );
  ANDN U44401 ( .B(n39953), .A(n39954), .Z(n45052) );
  XOR U44402 ( .A(n45054), .B(n45055), .Z(n39920) );
  ANDN U44403 ( .B(n39957), .A(n39958), .Z(n45054) );
  XNOR U44404 ( .A(n45056), .B(n45057), .Z(n39382) );
  ANDN U44405 ( .B(n39965), .A(n45058), .Z(n45056) );
  XNOR U44406 ( .A(n45059), .B(n45049), .Z(n39962) );
  ANDN U44407 ( .B(n45060), .A(n45061), .Z(n45059) );
  ANDN U44408 ( .B(n35876), .A(n35877), .Z(n45034) );
  XOR U44409 ( .A(n43490), .B(n37954), .Z(n35877) );
  XOR U44410 ( .A(n45062), .B(n41579), .Z(n37954) );
  XNOR U44411 ( .A(n45063), .B(n45064), .Z(n41579) );
  XNOR U44412 ( .A(n39734), .B(n38831), .Z(n45064) );
  XOR U44413 ( .A(n45065), .B(n43147), .Z(n38831) );
  NOR U44414 ( .A(n42098), .B(n43146), .Z(n45065) );
  XOR U44415 ( .A(n45066), .B(n43150), .Z(n39734) );
  ANDN U44416 ( .B(n42084), .A(n43149), .Z(n45066) );
  XOR U44417 ( .A(n37311), .B(n45067), .Z(n45063) );
  XOR U44418 ( .A(n35525), .B(n43142), .Z(n45067) );
  XNOR U44419 ( .A(n45068), .B(n43701), .Z(n43142) );
  ANDN U44420 ( .B(n45069), .A(n43700), .Z(n45068) );
  XNOR U44421 ( .A(n45070), .B(n43159), .Z(n35525) );
  ANDN U44422 ( .B(n42088), .A(n43158), .Z(n45070) );
  XNOR U44423 ( .A(n45071), .B(n43155), .Z(n37311) );
  ANDN U44424 ( .B(n45072), .A(n45073), .Z(n45071) );
  XNOR U44425 ( .A(n45074), .B(n40866), .Z(n43490) );
  IV U44426 ( .A(n45075), .Z(n40866) );
  ANDN U44427 ( .B(n43481), .A(n43482), .Z(n45074) );
  XOR U44428 ( .A(n42287), .B(n37523), .Z(n35876) );
  XOR U44429 ( .A(n40371), .B(n41147), .Z(n37523) );
  XNOR U44430 ( .A(n45076), .B(n45077), .Z(n41147) );
  XOR U44431 ( .A(n38683), .B(n38919), .Z(n45077) );
  XNOR U44432 ( .A(n45078), .B(n41131), .Z(n38919) );
  AND U44433 ( .A(n42263), .B(n42262), .Z(n45078) );
  XOR U44434 ( .A(n45081), .B(n45082), .Z(n42262) );
  XNOR U44435 ( .A(n45083), .B(n41126), .Z(n38683) );
  IV U44436 ( .A(n44144), .Z(n41126) );
  XOR U44437 ( .A(n45084), .B(n45085), .Z(n44144) );
  AND U44438 ( .A(n42270), .B(n42271), .Z(n45083) );
  XOR U44439 ( .A(n45086), .B(n43713), .Z(n42270) );
  XOR U44440 ( .A(n42530), .B(n45087), .Z(n45076) );
  XOR U44441 ( .A(n41576), .B(n39273), .Z(n45087) );
  XNOR U44442 ( .A(n45088), .B(n43062), .Z(n39273) );
  XNOR U44443 ( .A(n45089), .B(n44837), .Z(n43062) );
  XNOR U44444 ( .A(n45090), .B(n45091), .Z(n42273) );
  XOR U44445 ( .A(n45092), .B(n41135), .Z(n41576) );
  AND U44446 ( .A(n42266), .B(n42267), .Z(n45092) );
  XNOR U44447 ( .A(n45094), .B(n42526), .Z(n42266) );
  XNOR U44448 ( .A(n45095), .B(n45096), .Z(n42530) );
  ANDN U44449 ( .B(n42258), .A(n42260), .Z(n45095) );
  XNOR U44450 ( .A(n45097), .B(n42340), .Z(n42258) );
  XOR U44451 ( .A(n45098), .B(n45099), .Z(n40371) );
  XOR U44452 ( .A(n38572), .B(n40575), .Z(n45099) );
  XOR U44453 ( .A(n45100), .B(n44304), .Z(n40575) );
  NOR U44454 ( .A(n45101), .B(n42280), .Z(n45100) );
  XOR U44455 ( .A(n45102), .B(n44306), .Z(n38572) );
  ANDN U44456 ( .B(n42283), .A(n42284), .Z(n45102) );
  XOR U44457 ( .A(n38837), .B(n45103), .Z(n45098) );
  XOR U44458 ( .A(n44139), .B(n38791), .Z(n45103) );
  XOR U44459 ( .A(n45104), .B(n44295), .Z(n38791) );
  AND U44460 ( .A(n42294), .B(n42293), .Z(n45104) );
  XOR U44461 ( .A(n45105), .B(n44301), .Z(n44139) );
  ANDN U44462 ( .B(n45106), .A(n45107), .Z(n45105) );
  XNOR U44463 ( .A(n45108), .B(n44293), .Z(n38837) );
  XNOR U44464 ( .A(n45109), .B(n45110), .Z(n42287) );
  ANDN U44465 ( .B(n44299), .A(n45106), .Z(n45109) );
  XOR U44466 ( .A(n45111), .B(n40324), .Z(n34357) );
  IV U44467 ( .A(n40068), .Z(n40324) );
  XNOR U44468 ( .A(n43941), .B(n37837), .Z(n40068) );
  XOR U44469 ( .A(n42169), .B(n40210), .Z(n37837) );
  XNOR U44470 ( .A(n45112), .B(n45113), .Z(n40210) );
  XOR U44471 ( .A(n38156), .B(n40186), .Z(n45113) );
  XOR U44472 ( .A(n45114), .B(n43431), .Z(n40186) );
  XNOR U44473 ( .A(n44688), .B(n45115), .Z(n43431) );
  XOR U44474 ( .A(n45116), .B(n45117), .Z(n43943) );
  IV U44475 ( .A(n45118), .Z(n43944) );
  XNOR U44476 ( .A(n45119), .B(n44390), .Z(n38156) );
  XOR U44477 ( .A(n45120), .B(n45121), .Z(n44390) );
  NOR U44478 ( .A(n43946), .B(n43947), .Z(n45119) );
  XOR U44479 ( .A(n45122), .B(n45123), .Z(n43946) );
  XOR U44480 ( .A(n44385), .B(n45124), .Z(n45112) );
  XOR U44481 ( .A(n39402), .B(n34622), .Z(n45124) );
  XNOR U44482 ( .A(n45125), .B(n43427), .Z(n34622) );
  XOR U44483 ( .A(n45126), .B(n45127), .Z(n43427) );
  NOR U44484 ( .A(n45128), .B(n43938), .Z(n45125) );
  XOR U44485 ( .A(n44704), .B(n45129), .Z(n43938) );
  XNOR U44486 ( .A(n45130), .B(n43435), .Z(n39402) );
  XNOR U44487 ( .A(n44864), .B(n45132), .Z(n43935) );
  XNOR U44488 ( .A(n45133), .B(n43422), .Z(n44385) );
  XOR U44489 ( .A(n45134), .B(n45135), .Z(n43422) );
  XOR U44490 ( .A(n45137), .B(n45138), .Z(n42169) );
  XNOR U44491 ( .A(n35310), .B(n41710), .Z(n45138) );
  XOR U44492 ( .A(n45139), .B(n43447), .Z(n41710) );
  XNOR U44493 ( .A(n42312), .B(n45140), .Z(n43447) );
  XOR U44494 ( .A(n43346), .B(n45141), .Z(n43927) );
  XNOR U44495 ( .A(n45142), .B(n44789), .Z(n41177) );
  XOR U44496 ( .A(n45143), .B(n44402), .Z(n35310) );
  XOR U44497 ( .A(n45144), .B(n45145), .Z(n44402) );
  ANDN U44498 ( .B(n41173), .A(n43930), .Z(n45143) );
  XOR U44499 ( .A(n45146), .B(n44659), .Z(n43930) );
  XOR U44500 ( .A(n45147), .B(n45148), .Z(n41173) );
  XOR U44501 ( .A(n40900), .B(n45149), .Z(n45137) );
  XNOR U44502 ( .A(n43568), .B(n39656), .Z(n45149) );
  XNOR U44503 ( .A(n45150), .B(n43439), .Z(n39656) );
  XNOR U44504 ( .A(n45151), .B(n45152), .Z(n43439) );
  XOR U44505 ( .A(n45153), .B(n42673), .Z(n43923) );
  IV U44506 ( .A(n45154), .Z(n42673) );
  XNOR U44507 ( .A(n45155), .B(n42510), .Z(n41999) );
  XOR U44508 ( .A(n45156), .B(n43445), .Z(n43568) );
  XOR U44509 ( .A(n45157), .B(n43784), .Z(n43445) );
  AND U44510 ( .A(n43914), .B(n41167), .Z(n45156) );
  XOR U44511 ( .A(n45158), .B(n45159), .Z(n41167) );
  XNOR U44512 ( .A(n45160), .B(n42319), .Z(n43914) );
  XOR U44513 ( .A(n45161), .B(n43441), .Z(n40900) );
  XNOR U44514 ( .A(n45162), .B(n44869), .Z(n43441) );
  NOR U44515 ( .A(n41163), .B(n43918), .Z(n45161) );
  XNOR U44516 ( .A(n45163), .B(n43769), .Z(n43918) );
  XOR U44517 ( .A(n45164), .B(n44535), .Z(n41163) );
  XNOR U44518 ( .A(n45165), .B(n44394), .Z(n43941) );
  XNOR U44519 ( .A(n45166), .B(n45167), .Z(n44394) );
  NOR U44520 ( .A(n45136), .B(n43420), .Z(n45165) );
  ANDN U44521 ( .B(n38759), .A(n37973), .Z(n45111) );
  XNOR U44522 ( .A(n45169), .B(n45170), .Z(n42055) );
  XNOR U44523 ( .A(n39634), .B(n39084), .Z(n45170) );
  XOR U44524 ( .A(n45171), .B(n41850), .Z(n39084) );
  XOR U44525 ( .A(n45172), .B(n45173), .Z(n41850) );
  ANDN U44526 ( .B(n41851), .A(n43676), .Z(n45171) );
  XOR U44527 ( .A(n45174), .B(n41858), .Z(n39634) );
  XOR U44528 ( .A(n45175), .B(n43920), .Z(n41858) );
  XNOR U44529 ( .A(n37847), .B(n45176), .Z(n45169) );
  XOR U44530 ( .A(n38274), .B(n38560), .Z(n45176) );
  XNOR U44531 ( .A(n45177), .B(n42469), .Z(n38560) );
  XNOR U44532 ( .A(n45178), .B(n43329), .Z(n42469) );
  ANDN U44533 ( .B(n42468), .A(n43673), .Z(n45177) );
  XNOR U44534 ( .A(n45179), .B(n42707), .Z(n38274) );
  XNOR U44535 ( .A(n44869), .B(n45180), .Z(n42707) );
  ANDN U44536 ( .B(n42709), .A(n43660), .Z(n45179) );
  XOR U44537 ( .A(n45181), .B(n41854), .Z(n37847) );
  XOR U44538 ( .A(n45182), .B(n44550), .Z(n41854) );
  ANDN U44539 ( .B(n41855), .A(n43664), .Z(n45181) );
  IV U44540 ( .A(n45183), .Z(n43664) );
  XOR U44541 ( .A(n45184), .B(n45185), .Z(n38449) );
  XNOR U44542 ( .A(n37019), .B(n38923), .Z(n45185) );
  XOR U44543 ( .A(n45186), .B(n42228), .Z(n38923) );
  ANDN U44544 ( .B(n42229), .A(n41054), .Z(n45186) );
  IV U44545 ( .A(n45187), .Z(n41054) );
  XOR U44546 ( .A(n45188), .B(n41957), .Z(n37019) );
  ANDN U44547 ( .B(n45189), .A(n45190), .Z(n45188) );
  XNOR U44548 ( .A(n38494), .B(n45191), .Z(n45184) );
  XOR U44549 ( .A(n41842), .B(n40651), .Z(n45191) );
  XOR U44550 ( .A(n45192), .B(n41954), .Z(n40651) );
  XNOR U44551 ( .A(n45193), .B(n41950), .Z(n41842) );
  XOR U44552 ( .A(n45195), .B(n45196), .Z(n38494) );
  NOR U44553 ( .A(n42007), .B(n41050), .Z(n45195) );
  XNOR U44554 ( .A(n42092), .B(n38667), .Z(n38759) );
  IV U44555 ( .A(n39025), .Z(n38667) );
  XOR U44556 ( .A(n43483), .B(n41570), .Z(n39025) );
  XOR U44557 ( .A(n45197), .B(n45198), .Z(n41570) );
  XNOR U44558 ( .A(n40568), .B(n43811), .Z(n45198) );
  XNOR U44559 ( .A(n45199), .B(n43854), .Z(n43811) );
  XOR U44560 ( .A(n44585), .B(n45200), .Z(n43854) );
  NOR U44561 ( .A(n43853), .B(n43690), .Z(n45199) );
  XNOR U44562 ( .A(n45201), .B(n43164), .Z(n40568) );
  XOR U44563 ( .A(n45202), .B(n45203), .Z(n43164) );
  XNOR U44564 ( .A(n38641), .B(n45204), .Z(n45197) );
  XOR U44565 ( .A(n39426), .B(n39170), .Z(n45204) );
  XNOR U44566 ( .A(n45205), .B(n43182), .Z(n39170) );
  XOR U44567 ( .A(n45206), .B(n42691), .Z(n43182) );
  XNOR U44568 ( .A(n45208), .B(n43168), .Z(n39426) );
  XOR U44569 ( .A(n45209), .B(n43335), .Z(n43168) );
  ANDN U44570 ( .B(n43839), .A(n43693), .Z(n45208) );
  XNOR U44571 ( .A(n45210), .B(n43173), .Z(n38641) );
  XOR U44572 ( .A(n45211), .B(n44571), .Z(n43173) );
  XOR U44573 ( .A(n45212), .B(n45213), .Z(n43483) );
  XNOR U44574 ( .A(n41577), .B(n39665), .Z(n45213) );
  XOR U44575 ( .A(n45214), .B(n43158), .Z(n39665) );
  XOR U44576 ( .A(n45215), .B(n45216), .Z(n43158) );
  NOR U44577 ( .A(n42089), .B(n42088), .Z(n45214) );
  XOR U44578 ( .A(n42540), .B(n45217), .Z(n42088) );
  XOR U44579 ( .A(n45218), .B(n43146), .Z(n41577) );
  XOR U44580 ( .A(n45219), .B(n43329), .Z(n43146) );
  ANDN U44581 ( .B(n42098), .A(n42099), .Z(n45218) );
  XOR U44582 ( .A(n45220), .B(n45221), .Z(n42098) );
  XOR U44583 ( .A(n39488), .B(n45222), .Z(n45212) );
  XNOR U44584 ( .A(n40038), .B(n38962), .Z(n45222) );
  XNOR U44585 ( .A(n45223), .B(n43156), .Z(n38962) );
  IV U44586 ( .A(n45073), .Z(n43156) );
  XNOR U44587 ( .A(n45224), .B(n44182), .Z(n45073) );
  NOR U44588 ( .A(n45225), .B(n45072), .Z(n45223) );
  XNOR U44589 ( .A(n45226), .B(n43149), .Z(n40038) );
  XNOR U44590 ( .A(n45227), .B(n43323), .Z(n43149) );
  ANDN U44591 ( .B(n42086), .A(n42084), .Z(n45226) );
  XOR U44592 ( .A(n45228), .B(n45229), .Z(n42084) );
  XOR U44593 ( .A(n45230), .B(n43700), .Z(n39488) );
  XOR U44594 ( .A(n45231), .B(n45232), .Z(n43700) );
  ANDN U44595 ( .B(n42094), .A(n42096), .Z(n45230) );
  IV U44596 ( .A(n45069), .Z(n42094) );
  XNOR U44597 ( .A(n45233), .B(n42453), .Z(n45069) );
  XNOR U44598 ( .A(n45234), .B(n45072), .Z(n42092) );
  XNOR U44599 ( .A(n45235), .B(n45236), .Z(n45072) );
  ANDN U44600 ( .B(n45225), .A(n43154), .Z(n45234) );
  XOR U44601 ( .A(n45237), .B(n40062), .Z(n32905) );
  XOR U44602 ( .A(n37782), .B(n42426), .Z(n40062) );
  XNOR U44603 ( .A(n45238), .B(n44061), .Z(n42426) );
  IV U44604 ( .A(n45239), .Z(n44061) );
  NOR U44605 ( .A(n45240), .B(n44892), .Z(n45238) );
  IV U44606 ( .A(n35799), .Z(n37782) );
  XOR U44607 ( .A(n40705), .B(n44208), .Z(n35799) );
  XNOR U44608 ( .A(n45241), .B(n45242), .Z(n44208) );
  XNOR U44609 ( .A(n38939), .B(n39859), .Z(n45242) );
  XNOR U44610 ( .A(n45243), .B(n44047), .Z(n39859) );
  XOR U44611 ( .A(n45244), .B(n45245), .Z(n44047) );
  ANDN U44612 ( .B(n43374), .A(n43373), .Z(n45243) );
  XNOR U44613 ( .A(n45246), .B(n45247), .Z(n43373) );
  XNOR U44614 ( .A(n45248), .B(n45249), .Z(n43374) );
  XNOR U44615 ( .A(n45250), .B(n40960), .Z(n38939) );
  XOR U44616 ( .A(n44783), .B(n45251), .Z(n40960) );
  NOR U44617 ( .A(n43377), .B(n43376), .Z(n45250) );
  XNOR U44618 ( .A(n45252), .B(n45253), .Z(n43376) );
  XNOR U44619 ( .A(n45254), .B(n45255), .Z(n43377) );
  XOR U44620 ( .A(n40528), .B(n45256), .Z(n45241) );
  XOR U44621 ( .A(n40516), .B(n37801), .Z(n45256) );
  XNOR U44622 ( .A(n45257), .B(n40953), .Z(n37801) );
  XNOR U44623 ( .A(n44680), .B(n45258), .Z(n40953) );
  ANDN U44624 ( .B(n44050), .A(n44235), .Z(n45257) );
  XNOR U44625 ( .A(n45259), .B(n45260), .Z(n44235) );
  XOR U44626 ( .A(n45261), .B(n43962), .Z(n44050) );
  XNOR U44627 ( .A(n45262), .B(n43479), .Z(n40516) );
  XOR U44628 ( .A(n45263), .B(n44837), .Z(n43479) );
  ANDN U44629 ( .B(n43382), .A(n43383), .Z(n45262) );
  XOR U44630 ( .A(n45264), .B(n44839), .Z(n43383) );
  XNOR U44631 ( .A(n41652), .B(n45265), .Z(n43382) );
  XNOR U44632 ( .A(n45266), .B(n40949), .Z(n40528) );
  XNOR U44633 ( .A(n45267), .B(n45268), .Z(n40949) );
  ANDN U44634 ( .B(n43386), .A(n43387), .Z(n45266) );
  XOR U44635 ( .A(n45269), .B(n44167), .Z(n43387) );
  XOR U44636 ( .A(n45270), .B(n44479), .Z(n43386) );
  XOR U44637 ( .A(n45271), .B(n45272), .Z(n40705) );
  XOR U44638 ( .A(n36218), .B(n39253), .Z(n45272) );
  XOR U44639 ( .A(n45273), .B(n44073), .Z(n39253) );
  XOR U44640 ( .A(n45274), .B(n45275), .Z(n44073) );
  ANDN U44641 ( .B(n42437), .A(n42439), .Z(n45273) );
  XOR U44642 ( .A(n45276), .B(n43895), .Z(n42437) );
  XNOR U44643 ( .A(n45277), .B(n44057), .Z(n36218) );
  XOR U44644 ( .A(n45278), .B(n42877), .Z(n44057) );
  ANDN U44645 ( .B(n42428), .A(n42429), .Z(n45277) );
  XOR U44646 ( .A(n45279), .B(n45280), .Z(n42428) );
  XOR U44647 ( .A(n37083), .B(n45281), .Z(n45271) );
  XOR U44648 ( .A(n44041), .B(n37433), .Z(n45281) );
  XNOR U44649 ( .A(n45282), .B(n44065), .Z(n37433) );
  XOR U44650 ( .A(n44316), .B(n45283), .Z(n44065) );
  ANDN U44651 ( .B(n42435), .A(n44066), .Z(n45282) );
  XOR U44652 ( .A(n45284), .B(n44528), .Z(n44066) );
  XNOR U44653 ( .A(n45285), .B(n44069), .Z(n44041) );
  XOR U44654 ( .A(n45244), .B(n45286), .Z(n44069) );
  NOR U44655 ( .A(n44070), .B(n42442), .Z(n45285) );
  XOR U44656 ( .A(n45287), .B(n45117), .Z(n44070) );
  XNOR U44657 ( .A(n45288), .B(n44060), .Z(n37083) );
  XOR U44658 ( .A(n45289), .B(n43327), .Z(n44060) );
  ANDN U44659 ( .B(n45240), .A(n45239), .Z(n45288) );
  XOR U44660 ( .A(n45290), .B(n44106), .Z(n45239) );
  NOR U44661 ( .A(n35886), .B(n35888), .Z(n45237) );
  XNOR U44662 ( .A(n45291), .B(n45292), .Z(n35888) );
  XNOR U44663 ( .A(n42601), .B(n35932), .Z(n35886) );
  XOR U44664 ( .A(n40578), .B(n42049), .Z(n35932) );
  XOR U44665 ( .A(n45293), .B(n45294), .Z(n42049) );
  XOR U44666 ( .A(n36793), .B(n38084), .Z(n45294) );
  XOR U44667 ( .A(n45295), .B(n40384), .Z(n38084) );
  XNOR U44668 ( .A(n45296), .B(n45006), .Z(n40384) );
  ANDN U44669 ( .B(n40385), .A(n43106), .Z(n45295) );
  XOR U44670 ( .A(n45297), .B(n44845), .Z(n43106) );
  XOR U44671 ( .A(n42685), .B(n45298), .Z(n40385) );
  IV U44672 ( .A(n45159), .Z(n42685) );
  XOR U44673 ( .A(n45299), .B(n40394), .Z(n36793) );
  XOR U44674 ( .A(n45300), .B(n45301), .Z(n40394) );
  ANDN U44675 ( .B(n40395), .A(n44662), .Z(n45299) );
  XOR U44676 ( .A(n45302), .B(n45303), .Z(n44662) );
  XOR U44677 ( .A(n45304), .B(n43774), .Z(n40395) );
  XNOR U44678 ( .A(n40377), .B(n45305), .Z(n45293) );
  XOR U44679 ( .A(n37686), .B(n39058), .Z(n45305) );
  XNOR U44680 ( .A(n45306), .B(n43024), .Z(n39058) );
  XOR U44681 ( .A(n45307), .B(n45308), .Z(n43024) );
  ANDN U44682 ( .B(n43039), .A(n43110), .Z(n45306) );
  XNOR U44683 ( .A(n45309), .B(n44680), .Z(n43110) );
  XOR U44684 ( .A(n45310), .B(n45311), .Z(n43039) );
  XOR U44685 ( .A(n45312), .B(n40391), .Z(n37686) );
  XOR U44686 ( .A(n45154), .B(n45313), .Z(n40391) );
  ANDN U44687 ( .B(n40390), .A(n43096), .Z(n45312) );
  XNOR U44688 ( .A(n44688), .B(n45314), .Z(n43096) );
  XNOR U44689 ( .A(n45315), .B(n45316), .Z(n40390) );
  XNOR U44690 ( .A(n45317), .B(n42572), .Z(n40377) );
  XNOR U44691 ( .A(n45318), .B(n41742), .Z(n42572) );
  ANDN U44692 ( .B(n42573), .A(n43100), .Z(n45317) );
  XOR U44693 ( .A(n45319), .B(n45320), .Z(n43100) );
  XOR U44694 ( .A(n45321), .B(n45322), .Z(n42573) );
  XOR U44695 ( .A(n45323), .B(n45324), .Z(n40578) );
  XOR U44696 ( .A(n38351), .B(n38664), .Z(n45324) );
  XNOR U44697 ( .A(n45325), .B(n40228), .Z(n38664) );
  ANDN U44698 ( .B(n42596), .A(n42597), .Z(n45325) );
  XOR U44699 ( .A(n41888), .B(n45326), .Z(n42597) );
  XOR U44700 ( .A(n40232), .B(n45327), .Z(n38351) );
  XNOR U44701 ( .A(n11417), .B(n45328), .Z(n45327) );
  OR U44702 ( .A(n42599), .B(n42600), .Z(n45328) );
  XNOR U44703 ( .A(n44743), .B(n45329), .Z(n42600) );
  XOR U44704 ( .A(n38536), .B(n45330), .Z(n45323) );
  XOR U44705 ( .A(n39832), .B(n39120), .Z(n45330) );
  XNOR U44706 ( .A(n45331), .B(n40237), .Z(n39120) );
  ANDN U44707 ( .B(n45332), .A(n43289), .Z(n45331) );
  XNOR U44708 ( .A(n45333), .B(n40245), .Z(n39832) );
  ANDN U44709 ( .B(n42604), .A(n42605), .Z(n45333) );
  XOR U44710 ( .A(n45334), .B(n43594), .Z(n42605) );
  XNOR U44711 ( .A(n45335), .B(n40241), .Z(n38536) );
  ANDN U44712 ( .B(n42608), .A(n42609), .Z(n45335) );
  XOR U44713 ( .A(n45336), .B(n43323), .Z(n42609) );
  XNOR U44714 ( .A(n45337), .B(n45332), .Z(n42601) );
  XOR U44715 ( .A(n45338), .B(n45339), .Z(n40236) );
  XOR U44716 ( .A(n42881), .B(n45340), .Z(n43289) );
  XOR U44717 ( .A(n45341), .B(n45342), .Z(n34221) );
  XOR U44718 ( .A(n40043), .B(n30794), .Z(n45342) );
  XOR U44719 ( .A(n45343), .B(n38721), .Z(n30794) );
  XNOR U44720 ( .A(n44426), .B(n39454), .Z(n38721) );
  XNOR U44721 ( .A(n45344), .B(n45345), .Z(n39799) );
  XNOR U44722 ( .A(n42471), .B(n38884), .Z(n45345) );
  XNOR U44723 ( .A(n45346), .B(n42486), .Z(n38884) );
  ANDN U44724 ( .B(n41899), .A(n42485), .Z(n45346) );
  XOR U44725 ( .A(n45347), .B(n44180), .Z(n42485) );
  IV U44726 ( .A(n43319), .Z(n44180) );
  XNOR U44727 ( .A(n45348), .B(n45349), .Z(n41899) );
  XNOR U44728 ( .A(n45350), .B(n42482), .Z(n42471) );
  AND U44729 ( .A(n42483), .B(n41904), .Z(n45350) );
  XOR U44730 ( .A(n45351), .B(n45352), .Z(n41904) );
  XOR U44731 ( .A(n45353), .B(n45354), .Z(n42483) );
  XOR U44732 ( .A(n41180), .B(n45355), .Z(n45344) );
  XNOR U44733 ( .A(n37210), .B(n41611), .Z(n45355) );
  XNOR U44734 ( .A(n45356), .B(n42479), .Z(n41611) );
  ANDN U44735 ( .B(n42478), .A(n44414), .Z(n45356) );
  XOR U44736 ( .A(n45357), .B(n45358), .Z(n44414) );
  XOR U44737 ( .A(n42319), .B(n45359), .Z(n42478) );
  XOR U44738 ( .A(n45360), .B(n42475), .Z(n37210) );
  ANDN U44739 ( .B(n42476), .A(n41908), .Z(n45360) );
  XOR U44740 ( .A(n45303), .B(n45361), .Z(n41908) );
  XOR U44741 ( .A(n45362), .B(n43088), .Z(n42476) );
  XNOR U44742 ( .A(n45363), .B(n45364), .Z(n41180) );
  ANDN U44743 ( .B(n42489), .A(n41912), .Z(n45363) );
  IV U44744 ( .A(n44418), .Z(n41912) );
  XOR U44745 ( .A(n45365), .B(n43781), .Z(n44418) );
  XOR U44746 ( .A(n45366), .B(n42461), .Z(n42489) );
  XNOR U44747 ( .A(n45367), .B(n45368), .Z(n40534) );
  XNOR U44748 ( .A(n38995), .B(n40800), .Z(n45368) );
  XOR U44749 ( .A(n45369), .B(n40817), .Z(n40800) );
  NOR U44750 ( .A(n42802), .B(n40816), .Z(n45369) );
  XNOR U44751 ( .A(n45372), .B(n43535), .Z(n42802) );
  IV U44752 ( .A(n45358), .Z(n43535) );
  XOR U44753 ( .A(n45373), .B(n40813), .Z(n38995) );
  ANDN U44754 ( .B(n44431), .A(n40812), .Z(n45373) );
  XOR U44755 ( .A(n45374), .B(n45352), .Z(n40812) );
  IV U44756 ( .A(n44469), .Z(n45352) );
  XOR U44757 ( .A(n44743), .B(n45375), .Z(n44431) );
  XOR U44758 ( .A(n37839), .B(n45376), .Z(n45367) );
  XOR U44759 ( .A(n36556), .B(n38081), .Z(n45376) );
  XOR U44760 ( .A(n45377), .B(n45378), .Z(n38081) );
  ANDN U44761 ( .B(n44428), .A(n42798), .Z(n45377) );
  XOR U44762 ( .A(n45379), .B(n45249), .Z(n42798) );
  XNOR U44763 ( .A(n45380), .B(n40820), .Z(n36556) );
  ANDN U44764 ( .B(n40821), .A(n45381), .Z(n45380) );
  XNOR U44765 ( .A(n45382), .B(n40808), .Z(n37839) );
  ANDN U44766 ( .B(n42793), .A(n40807), .Z(n45382) );
  XOR U44767 ( .A(n45383), .B(n44336), .Z(n40807) );
  XOR U44768 ( .A(n45384), .B(n43319), .Z(n42793) );
  XNOR U44769 ( .A(n45385), .B(n40821), .Z(n44426) );
  XNOR U44770 ( .A(n45386), .B(n45387), .Z(n40821) );
  ANDN U44771 ( .B(n42791), .A(n42790), .Z(n45385) );
  IV U44772 ( .A(n45381), .Z(n42790) );
  XOR U44773 ( .A(n45388), .B(n45389), .Z(n45381) );
  ANDN U44774 ( .B(n38382), .A(n38002), .Z(n45343) );
  XOR U44775 ( .A(n44904), .B(n36701), .Z(n38002) );
  XOR U44776 ( .A(n44312), .B(n42818), .Z(n36701) );
  XNOR U44777 ( .A(n45390), .B(n45391), .Z(n42818) );
  XNOR U44778 ( .A(n39296), .B(n38949), .Z(n45391) );
  XOR U44779 ( .A(n45392), .B(n40714), .Z(n38949) );
  XOR U44780 ( .A(n45393), .B(n42166), .Z(n40714) );
  NOR U44781 ( .A(n44907), .B(n42416), .Z(n45392) );
  XOR U44782 ( .A(n45394), .B(n45395), .Z(n42416) );
  XNOR U44783 ( .A(n45396), .B(n45397), .Z(n44907) );
  XOR U44784 ( .A(n45399), .B(n44193), .Z(n40723) );
  ANDN U44785 ( .B(n44010), .A(n42410), .Z(n45398) );
  XOR U44786 ( .A(n45400), .B(n45401), .Z(n42410) );
  XOR U44787 ( .A(n45402), .B(n45403), .Z(n44010) );
  XNOR U44788 ( .A(n40463), .B(n45404), .Z(n45390) );
  XOR U44789 ( .A(n39825), .B(n38307), .Z(n45404) );
  XNOR U44790 ( .A(n45405), .B(n44020), .Z(n38307) );
  IV U44791 ( .A(n40719), .Z(n44020) );
  XOR U44792 ( .A(n45406), .B(n44106), .Z(n40719) );
  ANDN U44793 ( .B(n44021), .A(n44913), .Z(n45405) );
  IV U44794 ( .A(n44911), .Z(n44913) );
  XOR U44795 ( .A(n45407), .B(n42522), .Z(n44911) );
  XOR U44796 ( .A(n45274), .B(n45408), .Z(n44021) );
  XNOR U44797 ( .A(n45410), .B(n44191), .Z(n40710) );
  ANDN U44798 ( .B(n42414), .A(n44018), .Z(n45409) );
  XOR U44799 ( .A(n45411), .B(n40728), .Z(n40463) );
  XNOR U44800 ( .A(n45412), .B(n43719), .Z(n40728) );
  XNOR U44801 ( .A(n45413), .B(n42309), .Z(n44006) );
  XOR U44802 ( .A(n45414), .B(n45415), .Z(n42782) );
  XOR U44803 ( .A(n45416), .B(n45417), .Z(n44312) );
  XNOR U44804 ( .A(n38403), .B(n38730), .Z(n45417) );
  XNOR U44805 ( .A(n45418), .B(n42439), .Z(n38730) );
  XOR U44806 ( .A(n45419), .B(n44201), .Z(n42439) );
  ANDN U44807 ( .B(n44072), .A(n42438), .Z(n45418) );
  IV U44808 ( .A(n44896), .Z(n42438) );
  XNOR U44809 ( .A(n45420), .B(n42325), .Z(n44896) );
  XOR U44810 ( .A(n44680), .B(n45421), .Z(n44072) );
  XNOR U44811 ( .A(n45422), .B(n42429), .Z(n38403) );
  XNOR U44812 ( .A(n45423), .B(n44009), .Z(n42429) );
  ANDN U44813 ( .B(n42430), .A(n44056), .Z(n45422) );
  XNOR U44814 ( .A(n45424), .B(n45425), .Z(n44056) );
  XNOR U44815 ( .A(n45426), .B(n40853), .Z(n42430) );
  XNOR U44816 ( .A(n38782), .B(n45429), .Z(n45416) );
  XOR U44817 ( .A(n37263), .B(n42422), .Z(n45429) );
  XOR U44818 ( .A(n45430), .B(n42435), .Z(n42422) );
  XNOR U44819 ( .A(n45431), .B(n42166), .Z(n42435) );
  AND U44820 ( .A(n42434), .B(n44064), .Z(n45430) );
  XNOR U44821 ( .A(n43722), .B(n45432), .Z(n44064) );
  XOR U44822 ( .A(n45433), .B(n44619), .Z(n42434) );
  XOR U44823 ( .A(n45434), .B(n45240), .Z(n37263) );
  XOR U44824 ( .A(n42214), .B(n45435), .Z(n45240) );
  XOR U44825 ( .A(n45436), .B(n45437), .Z(n42214) );
  ANDN U44826 ( .B(n44892), .A(n44059), .Z(n45434) );
  XNOR U44827 ( .A(n41874), .B(n45438), .Z(n44059) );
  XOR U44828 ( .A(n45439), .B(n45440), .Z(n44892) );
  XOR U44829 ( .A(n45441), .B(n42442), .Z(n38782) );
  XOR U44830 ( .A(n45442), .B(n45443), .Z(n42442) );
  ANDN U44831 ( .B(n42443), .A(n44068), .Z(n45441) );
  XOR U44832 ( .A(n42689), .B(n45444), .Z(n44068) );
  XNOR U44833 ( .A(n43595), .B(n45445), .Z(n42443) );
  XOR U44834 ( .A(n45447), .B(n45448), .Z(n44018) );
  NOR U44835 ( .A(n40709), .B(n42414), .Z(n45446) );
  XNOR U44836 ( .A(n42510), .B(n45449), .Z(n42414) );
  XOR U44837 ( .A(n45450), .B(n45451), .Z(n42510) );
  XOR U44838 ( .A(n45452), .B(n45453), .Z(n40709) );
  XOR U44839 ( .A(n42355), .B(n38149), .Z(n38382) );
  IV U44840 ( .A(n39399), .Z(n38149) );
  XNOR U44841 ( .A(n40370), .B(n40974), .Z(n39399) );
  XNOR U44842 ( .A(n45454), .B(n45455), .Z(n40974) );
  XOR U44843 ( .A(n38951), .B(n39805), .Z(n45455) );
  XNOR U44844 ( .A(n45456), .B(n45018), .Z(n39805) );
  ANDN U44845 ( .B(n45457), .A(n43241), .Z(n45456) );
  XNOR U44846 ( .A(n45458), .B(n45007), .Z(n38951) );
  ANDN U44847 ( .B(n43006), .A(n43007), .Z(n45458) );
  XOR U44848 ( .A(n45459), .B(n44841), .Z(n43007) );
  XNOR U44849 ( .A(n41993), .B(n45460), .Z(n45454) );
  XNOR U44850 ( .A(n39884), .B(n39844), .Z(n45460) );
  XNOR U44851 ( .A(n45461), .B(n45003), .Z(n39844) );
  NOR U44852 ( .A(n42352), .B(n42353), .Z(n45461) );
  XOR U44853 ( .A(n45462), .B(n45463), .Z(n42353) );
  XNOR U44854 ( .A(n45464), .B(n45016), .Z(n39884) );
  ANDN U44855 ( .B(n42359), .A(n42360), .Z(n45464) );
  XNOR U44856 ( .A(n45465), .B(n45466), .Z(n42360) );
  XNOR U44857 ( .A(n45467), .B(n45012), .Z(n41993) );
  NOR U44858 ( .A(n42348), .B(n42349), .Z(n45467) );
  XOR U44859 ( .A(n45468), .B(n43846), .Z(n42349) );
  XOR U44860 ( .A(n45469), .B(n45470), .Z(n40370) );
  XNOR U44861 ( .A(n40967), .B(n38099), .Z(n45470) );
  XNOR U44862 ( .A(n45471), .B(n44287), .Z(n38099) );
  ANDN U44863 ( .B(n42382), .A(n42383), .Z(n45471) );
  ANDN U44864 ( .B(n42378), .A(n42380), .Z(n45472) );
  XOR U44865 ( .A(n45473), .B(n45474), .Z(n45469) );
  XOR U44866 ( .A(n39861), .B(n38563), .Z(n45474) );
  XOR U44867 ( .A(n45475), .B(n45476), .Z(n38563) );
  XOR U44868 ( .A(n45477), .B(n45478), .Z(n39861) );
  ANDN U44869 ( .B(n42365), .A(n42366), .Z(n45477) );
  XNOR U44870 ( .A(n45479), .B(n45457), .Z(n42355) );
  AND U44871 ( .A(n43241), .B(n43243), .Z(n45479) );
  XOR U44872 ( .A(n40843), .B(n45480), .Z(n43243) );
  XNOR U44873 ( .A(n45481), .B(n45482), .Z(n43241) );
  XOR U44874 ( .A(n45483), .B(n38704), .Z(n40043) );
  XNOR U44875 ( .A(n42127), .B(n38027), .Z(n38704) );
  XNOR U44876 ( .A(n44787), .B(n39076), .Z(n38027) );
  XNOR U44877 ( .A(n45484), .B(n45485), .Z(n39076) );
  XNOR U44878 ( .A(n42047), .B(n45486), .Z(n45485) );
  XOR U44879 ( .A(n45487), .B(n41239), .Z(n42047) );
  NOR U44880 ( .A(n39902), .B(n39901), .Z(n45487) );
  XNOR U44881 ( .A(n45488), .B(n42157), .Z(n39902) );
  XOR U44882 ( .A(n41152), .B(n45489), .Z(n45484) );
  XOR U44883 ( .A(n40968), .B(n39931), .Z(n45489) );
  XNOR U44884 ( .A(n45490), .B(n41247), .Z(n39931) );
  NOR U44885 ( .A(n39897), .B(n39898), .Z(n45490) );
  XNOR U44886 ( .A(n45491), .B(n45492), .Z(n39898) );
  XNOR U44887 ( .A(n45493), .B(n41243), .Z(n40968) );
  ANDN U44888 ( .B(n39916), .A(n39914), .Z(n45493) );
  XOR U44889 ( .A(n45494), .B(n44039), .Z(n39916) );
  XNOR U44890 ( .A(n45495), .B(n41237), .Z(n41152) );
  NOR U44891 ( .A(n42459), .B(n39910), .Z(n45495) );
  IV U44892 ( .A(n39911), .Z(n42459) );
  XNOR U44893 ( .A(n45496), .B(n45497), .Z(n39911) );
  XOR U44894 ( .A(n45498), .B(n45499), .Z(n44787) );
  XNOR U44895 ( .A(n39358), .B(n39427), .Z(n45499) );
  XNOR U44896 ( .A(n45500), .B(n43131), .Z(n39427) );
  NOR U44897 ( .A(n43132), .B(n42135), .Z(n45500) );
  XOR U44898 ( .A(n45501), .B(n43656), .Z(n42135) );
  XOR U44899 ( .A(n44254), .B(n45502), .Z(n43132) );
  IV U44900 ( .A(n43576), .Z(n44254) );
  XNOR U44901 ( .A(n45503), .B(n43123), .Z(n39358) );
  ANDN U44902 ( .B(n42144), .A(n43124), .Z(n45503) );
  XOR U44903 ( .A(n45504), .B(n45505), .Z(n43124) );
  XOR U44904 ( .A(n45506), .B(n44472), .Z(n42144) );
  XNOR U44905 ( .A(n36392), .B(n45507), .Z(n45498) );
  XOR U44906 ( .A(n38111), .B(n43114), .Z(n45507) );
  XNOR U44907 ( .A(n45508), .B(n43135), .Z(n43114) );
  AND U44908 ( .A(n42129), .B(n42131), .Z(n45508) );
  XOR U44909 ( .A(n44659), .B(n45509), .Z(n42131) );
  XOR U44910 ( .A(n45510), .B(n45453), .Z(n42129) );
  XOR U44911 ( .A(n45511), .B(n43128), .Z(n38111) );
  NOR U44912 ( .A(n42139), .B(n42138), .Z(n45511) );
  XNOR U44913 ( .A(n42456), .B(n45512), .Z(n42138) );
  IV U44914 ( .A(n45315), .Z(n42456) );
  XOR U44915 ( .A(n45513), .B(n45514), .Z(n42139) );
  XNOR U44916 ( .A(n45515), .B(n43120), .Z(n36392) );
  ANDN U44917 ( .B(n43119), .A(n45516), .Z(n45515) );
  XNOR U44918 ( .A(n45517), .B(n43119), .Z(n42127) );
  XOR U44919 ( .A(n45518), .B(n45519), .Z(n43119) );
  ANDN U44920 ( .B(n43752), .A(n43751), .Z(n45517) );
  IV U44921 ( .A(n45516), .Z(n43751) );
  XOR U44922 ( .A(n45520), .B(n42153), .Z(n45516) );
  ANDN U44923 ( .B(n40053), .A(n38006), .Z(n45483) );
  XOR U44924 ( .A(n31660), .B(n45521), .Z(n45341) );
  XNOR U44925 ( .A(n31749), .B(n36038), .Z(n45521) );
  XNOR U44926 ( .A(n45522), .B(n38713), .Z(n36038) );
  IV U44927 ( .A(n40056), .Z(n38713) );
  XOR U44928 ( .A(n45291), .B(n45523), .Z(n40056) );
  IV U44929 ( .A(n38339), .Z(n45291) );
  XNOR U44930 ( .A(n43452), .B(n42124), .Z(n38339) );
  XNOR U44931 ( .A(n45524), .B(n45525), .Z(n42124) );
  XOR U44932 ( .A(n36419), .B(n38954), .Z(n45525) );
  XOR U44933 ( .A(n45526), .B(n42246), .Z(n38954) );
  ANDN U44934 ( .B(n43746), .A(n43747), .Z(n45526) );
  XNOR U44935 ( .A(n45527), .B(n42253), .Z(n36419) );
  ANDN U44936 ( .B(n43736), .A(n45528), .Z(n45527) );
  XOR U44937 ( .A(n44711), .B(n45529), .Z(n45524) );
  XOR U44938 ( .A(n40623), .B(n44785), .Z(n45529) );
  XOR U44939 ( .A(n45530), .B(n43518), .Z(n44785) );
  ANDN U44940 ( .B(n43741), .A(n43740), .Z(n45530) );
  XNOR U44941 ( .A(n45531), .B(n45532), .Z(n40623) );
  ANDN U44942 ( .B(n43732), .A(n43733), .Z(n45531) );
  XOR U44943 ( .A(n45533), .B(n42241), .Z(n44711) );
  ANDN U44944 ( .B(n43743), .A(n43744), .Z(n45533) );
  XNOR U44945 ( .A(n45534), .B(n45535), .Z(n43452) );
  XNOR U44946 ( .A(n43494), .B(n45536), .Z(n45535) );
  XNOR U44947 ( .A(n45537), .B(n39726), .Z(n43494) );
  ANDN U44948 ( .B(n45538), .A(n45539), .Z(n45537) );
  XOR U44949 ( .A(n37010), .B(n45540), .Z(n45534) );
  XNOR U44950 ( .A(n43390), .B(n38857), .Z(n45540) );
  XOR U44951 ( .A(n45541), .B(n45542), .Z(n38857) );
  ANDN U44952 ( .B(n45543), .A(n45544), .Z(n45541) );
  XNOR U44953 ( .A(n45545), .B(n39731), .Z(n43390) );
  ANDN U44954 ( .B(n45546), .A(n45547), .Z(n45545) );
  XNOR U44955 ( .A(n45548), .B(n39721), .Z(n37010) );
  ANDN U44956 ( .B(n45549), .A(n45550), .Z(n45548) );
  ANDN U44957 ( .B(n37998), .A(n38387), .Z(n45522) );
  XOR U44958 ( .A(n34633), .B(n42031), .Z(n38387) );
  XNOR U44959 ( .A(n45551), .B(n45552), .Z(n42031) );
  ANDN U44960 ( .B(n41766), .A(n41767), .Z(n45551) );
  XNOR U44961 ( .A(n45553), .B(n45554), .Z(n41767) );
  XNOR U44962 ( .A(n41943), .B(n43184), .Z(n34633) );
  XNOR U44963 ( .A(n45555), .B(n45556), .Z(n43184) );
  XNOR U44964 ( .A(n38139), .B(n37520), .Z(n45556) );
  XNOR U44965 ( .A(n45557), .B(n42874), .Z(n37520) );
  ANDN U44966 ( .B(n42038), .A(n41779), .Z(n45557) );
  XOR U44967 ( .A(n45154), .B(n45558), .Z(n41779) );
  XNOR U44968 ( .A(n45559), .B(n42883), .Z(n38139) );
  ANDN U44969 ( .B(n42033), .A(n41762), .Z(n45559) );
  XNOR U44970 ( .A(n40840), .B(n45560), .Z(n41762) );
  XNOR U44971 ( .A(n38116), .B(n45561), .Z(n45555) );
  XNOR U44972 ( .A(n37908), .B(n39416), .Z(n45561) );
  XNOR U44973 ( .A(n45562), .B(n42869), .Z(n39416) );
  ANDN U44974 ( .B(n42036), .A(n41771), .Z(n45562) );
  XNOR U44975 ( .A(n45563), .B(n42496), .Z(n41771) );
  XOR U44976 ( .A(n45564), .B(n42878), .Z(n37908) );
  ANDN U44977 ( .B(n42040), .A(n41775), .Z(n45564) );
  XOR U44978 ( .A(n45565), .B(n45566), .Z(n41775) );
  XOR U44979 ( .A(n45567), .B(n42865), .Z(n38116) );
  ANDN U44980 ( .B(n45552), .A(n41766), .Z(n45567) );
  XOR U44981 ( .A(n45568), .B(n45569), .Z(n41766) );
  XOR U44982 ( .A(n45570), .B(n45571), .Z(n41943) );
  XNOR U44983 ( .A(n45572), .B(n39277), .Z(n45571) );
  XNOR U44984 ( .A(n45573), .B(n42853), .Z(n39277) );
  ANDN U44985 ( .B(n41617), .A(n41615), .Z(n45573) );
  XNOR U44986 ( .A(n45574), .B(n45575), .Z(n41617) );
  XOR U44987 ( .A(n39813), .B(n45576), .Z(n45570) );
  XOR U44988 ( .A(n39390), .B(n39521), .Z(n45576) );
  XNOR U44989 ( .A(n45577), .B(n42861), .Z(n39521) );
  ANDN U44990 ( .B(n39575), .A(n39573), .Z(n45577) );
  XOR U44991 ( .A(n45578), .B(n41874), .Z(n39575) );
  XNOR U44992 ( .A(n45579), .B(n42844), .Z(n39390) );
  NOR U44993 ( .A(n40121), .B(n40120), .Z(n45579) );
  XOR U44994 ( .A(n45580), .B(n45565), .Z(n40121) );
  XNOR U44995 ( .A(n45581), .B(n42857), .Z(n39813) );
  NOR U44996 ( .A(n41790), .B(n41941), .Z(n45581) );
  XNOR U44997 ( .A(n45582), .B(n45583), .Z(n41790) );
  XOR U44998 ( .A(n42624), .B(n33927), .Z(n37998) );
  XNOR U44999 ( .A(n40359), .B(n43760), .Z(n33927) );
  XNOR U45000 ( .A(n45584), .B(n45585), .Z(n43760) );
  XNOR U45001 ( .A(n39476), .B(n38519), .Z(n45585) );
  XNOR U45002 ( .A(n45586), .B(n44875), .Z(n38519) );
  NOR U45003 ( .A(n40700), .B(n42639), .Z(n45586) );
  XOR U45004 ( .A(n45587), .B(n45588), .Z(n40700) );
  XNOR U45005 ( .A(n45589), .B(n45590), .Z(n39476) );
  NOR U45006 ( .A(n40106), .B(n42645), .Z(n45589) );
  XOR U45007 ( .A(n45591), .B(n45592), .Z(n40106) );
  XOR U45008 ( .A(n40350), .B(n45593), .Z(n45584) );
  XOR U45009 ( .A(n39928), .B(n37795), .Z(n45593) );
  XNOR U45010 ( .A(n45594), .B(n44887), .Z(n37795) );
  IV U45011 ( .A(n45595), .Z(n44887) );
  ANDN U45012 ( .B(n43787), .A(n40116), .Z(n45594) );
  IV U45013 ( .A(n43788), .Z(n40116) );
  XOR U45014 ( .A(n45596), .B(n45597), .Z(n43788) );
  XNOR U45015 ( .A(n45598), .B(n44871), .Z(n39928) );
  NOR U45016 ( .A(n45599), .B(n40112), .Z(n45598) );
  XOR U45017 ( .A(n45600), .B(n44167), .Z(n40112) );
  IV U45018 ( .A(n41878), .Z(n44167) );
  XNOR U45019 ( .A(n44879), .B(n45601), .Z(n40350) );
  XOR U45020 ( .A(n45602), .B(n4407), .Z(n45601) );
  NANDN U45021 ( .A(rc_i[0]), .B(n31711), .Z(n4407) );
  ANDN U45022 ( .B(n42636), .A(n40102), .Z(n45602) );
  XNOR U45023 ( .A(n42689), .B(n45603), .Z(n40102) );
  XOR U45024 ( .A(n45604), .B(n45605), .Z(n40359) );
  XNOR U45025 ( .A(n39282), .B(n45606), .Z(n45605) );
  NOR U45026 ( .A(n42620), .B(n42621), .Z(n45607) );
  XOR U45027 ( .A(n38182), .B(n45608), .Z(n45604) );
  XOR U45028 ( .A(n41719), .B(n39271), .Z(n45608) );
  NOR U45029 ( .A(n42617), .B(n42616), .Z(n45609) );
  XNOR U45030 ( .A(n45610), .B(n43810), .Z(n41719) );
  NOR U45031 ( .A(n45611), .B(n45612), .Z(n45610) );
  XOR U45032 ( .A(n45613), .B(n43798), .Z(n38182) );
  ANDN U45033 ( .B(n42628), .A(n42626), .Z(n45613) );
  XNOR U45034 ( .A(n45614), .B(n45611), .Z(n42624) );
  ANDN U45035 ( .B(n45612), .A(n43808), .Z(n45614) );
  XOR U45036 ( .A(n45615), .B(n38709), .Z(n31749) );
  XNOR U45037 ( .A(n39930), .B(n45486), .Z(n38709) );
  XOR U45038 ( .A(n45616), .B(n41250), .Z(n45486) );
  NOR U45039 ( .A(n39907), .B(n39906), .Z(n45616) );
  XNOR U45040 ( .A(n45617), .B(n42329), .Z(n39907) );
  XNOR U45041 ( .A(n42817), .B(n43136), .Z(n39930) );
  XNOR U45042 ( .A(n45618), .B(n45619), .Z(n43136) );
  XOR U45043 ( .A(n40269), .B(n39814), .Z(n45619) );
  XNOR U45044 ( .A(n45620), .B(n41244), .Z(n39814) );
  XNOR U45045 ( .A(n45621), .B(n45622), .Z(n41244) );
  XOR U45046 ( .A(n45623), .B(n43594), .Z(n41243) );
  XOR U45047 ( .A(n41733), .B(n45624), .Z(n39914) );
  XOR U45048 ( .A(n45625), .B(n41251), .Z(n40269) );
  XOR U45049 ( .A(n45626), .B(n45627), .Z(n41251) );
  ANDN U45050 ( .B(n39906), .A(n41250), .Z(n45625) );
  XOR U45051 ( .A(n45628), .B(n45629), .Z(n41250) );
  XNOR U45052 ( .A(n45630), .B(n45631), .Z(n39906) );
  XNOR U45053 ( .A(n39946), .B(n45632), .Z(n45618) );
  XOR U45054 ( .A(n39306), .B(n40476), .Z(n45632) );
  XNOR U45055 ( .A(n45633), .B(n41236), .Z(n40476) );
  XOR U45056 ( .A(n45634), .B(n45635), .Z(n41236) );
  XOR U45057 ( .A(n45636), .B(n42160), .Z(n41237) );
  XOR U45058 ( .A(n45637), .B(n42318), .Z(n39910) );
  IV U45059 ( .A(n42301), .Z(n42318) );
  XNOR U45060 ( .A(n45638), .B(n41246), .Z(n39306) );
  XNOR U45061 ( .A(n43091), .B(n45639), .Z(n41246) );
  XOR U45062 ( .A(n40843), .B(n45640), .Z(n39897) );
  IV U45063 ( .A(n43583), .Z(n40843) );
  XNOR U45064 ( .A(n45641), .B(n44604), .Z(n41247) );
  XNOR U45065 ( .A(n45642), .B(n41240), .Z(n39946) );
  XOR U45066 ( .A(n45643), .B(n42852), .Z(n41240) );
  IV U45067 ( .A(n45644), .Z(n42852) );
  ANDN U45068 ( .B(n39901), .A(n41239), .Z(n45642) );
  XNOR U45069 ( .A(n45645), .B(n45646), .Z(n41239) );
  XOR U45070 ( .A(n45647), .B(n45260), .Z(n39901) );
  XOR U45071 ( .A(n45648), .B(n45649), .Z(n42817) );
  XOR U45072 ( .A(n38774), .B(n39137), .Z(n45649) );
  XOR U45073 ( .A(n45650), .B(n40316), .Z(n39137) );
  XNOR U45074 ( .A(n41639), .B(n45651), .Z(n40316) );
  XOR U45075 ( .A(n45652), .B(n44263), .Z(n41544) );
  XOR U45076 ( .A(n45653), .B(n45448), .Z(n41545) );
  XNOR U45077 ( .A(n45654), .B(n40320), .Z(n38774) );
  XOR U45078 ( .A(n45655), .B(n45656), .Z(n40320) );
  ANDN U45079 ( .B(n40399), .A(n40398), .Z(n45654) );
  XNOR U45080 ( .A(n45658), .B(n43846), .Z(n40399) );
  XNOR U45081 ( .A(n44001), .B(n45659), .Z(n45648) );
  XOR U45082 ( .A(n39093), .B(n37788), .Z(n45659) );
  XOR U45083 ( .A(n45660), .B(n42420), .Z(n37788) );
  XNOR U45084 ( .A(n44163), .B(n45661), .Z(n42420) );
  ANDN U45085 ( .B(n40154), .A(n40155), .Z(n45660) );
  XOR U45086 ( .A(n45662), .B(n44859), .Z(n40155) );
  XNOR U45087 ( .A(n45665), .B(n40311), .Z(n39093) );
  ANDN U45088 ( .B(n42393), .A(n42820), .Z(n45665) );
  XOR U45089 ( .A(n45667), .B(n45167), .Z(n42820) );
  XOR U45090 ( .A(n45668), .B(n45669), .Z(n42393) );
  XOR U45091 ( .A(n45670), .B(n40307), .Z(n44001) );
  XNOR U45092 ( .A(n45671), .B(n44336), .Z(n40307) );
  XOR U45093 ( .A(n45672), .B(n45673), .Z(n40161) );
  XOR U45094 ( .A(n43091), .B(n45674), .Z(n40163) );
  ANDN U45095 ( .B(n38390), .A(n37989), .Z(n45615) );
  XNOR U45096 ( .A(n43048), .B(n38900), .Z(n35611) );
  XNOR U45097 ( .A(n45676), .B(n45677), .Z(n38900) );
  XOR U45098 ( .A(n36969), .B(n39925), .Z(n45677) );
  XOR U45099 ( .A(n45678), .B(n44987), .Z(n39925) );
  XNOR U45100 ( .A(n44316), .B(n45679), .Z(n42990) );
  XNOR U45101 ( .A(n45680), .B(n44971), .Z(n36969) );
  ANDN U45102 ( .B(n42999), .A(n45681), .Z(n45680) );
  XNOR U45103 ( .A(n42846), .B(n45682), .Z(n42999) );
  XOR U45104 ( .A(n39667), .B(n45683), .Z(n45676) );
  XOR U45105 ( .A(n45684), .B(n37615), .Z(n45683) );
  XNOR U45106 ( .A(n45685), .B(n44975), .Z(n37615) );
  ANDN U45107 ( .B(n43003), .A(n45686), .Z(n45685) );
  XOR U45108 ( .A(n45687), .B(n45688), .Z(n43003) );
  XNOR U45109 ( .A(n45689), .B(n44983), .Z(n39667) );
  XNOR U45110 ( .A(n45690), .B(n43865), .Z(n42986) );
  XOR U45111 ( .A(n45691), .B(n45692), .Z(n43048) );
  XNOR U45112 ( .A(n38421), .B(n39850), .Z(n45692) );
  XOR U45113 ( .A(n45693), .B(n41524), .Z(n39850) );
  XOR U45114 ( .A(n45694), .B(n41740), .Z(n41524) );
  ANDN U45115 ( .B(n41525), .A(n44108), .Z(n45693) );
  IV U45116 ( .A(n45695), .Z(n44108) );
  XOR U45117 ( .A(n45696), .B(n41528), .Z(n38421) );
  XNOR U45118 ( .A(n45697), .B(n45698), .Z(n41528) );
  AND U45119 ( .A(n44121), .B(n41529), .Z(n45696) );
  XOR U45120 ( .A(n39615), .B(n45699), .Z(n45691) );
  XOR U45121 ( .A(n41518), .B(n39540), .Z(n45699) );
  XNOR U45122 ( .A(n45700), .B(n41541), .Z(n39540) );
  XOR U45123 ( .A(n45701), .B(n44218), .Z(n41541) );
  XNOR U45124 ( .A(n45702), .B(n41537), .Z(n41518) );
  XOR U45125 ( .A(n45703), .B(n44759), .Z(n41537) );
  AND U45126 ( .A(n41538), .B(n44116), .Z(n45702) );
  XNOR U45127 ( .A(n45704), .B(n43610), .Z(n39615) );
  IV U45128 ( .A(n41533), .Z(n43610) );
  XOR U45129 ( .A(n45705), .B(n44533), .Z(n41533) );
  AND U45130 ( .A(n44112), .B(n41534), .Z(n45704) );
  XOR U45131 ( .A(n38616), .B(n42932), .Z(n38390) );
  XOR U45132 ( .A(n45706), .B(n43878), .Z(n42932) );
  XOR U45133 ( .A(n45707), .B(n44327), .Z(n43353) );
  IV U45134 ( .A(n44503), .Z(n44327) );
  XOR U45135 ( .A(n43141), .B(n40216), .Z(n38616) );
  XOR U45136 ( .A(n45708), .B(n45709), .Z(n40216) );
  XNOR U45137 ( .A(n39164), .B(n37787), .Z(n45709) );
  XOR U45138 ( .A(n45710), .B(n43885), .Z(n37787) );
  XOR U45139 ( .A(n45711), .B(n41594), .Z(n43885) );
  ANDN U45140 ( .B(n42938), .A(n42936), .Z(n45710) );
  IV U45141 ( .A(n43884), .Z(n42936) );
  XOR U45142 ( .A(n45712), .B(n44114), .Z(n43884) );
  XOR U45143 ( .A(n44704), .B(n45713), .Z(n42938) );
  XNOR U45144 ( .A(n45714), .B(n43359), .Z(n39164) );
  XOR U45145 ( .A(n45715), .B(n41878), .Z(n43359) );
  XNOR U45146 ( .A(n45716), .B(n45717), .Z(n41878) );
  NOR U45147 ( .A(n43880), .B(n44212), .Z(n45714) );
  XNOR U45148 ( .A(n45718), .B(n45656), .Z(n44212) );
  XOR U45149 ( .A(n43874), .B(n45720), .Z(n45708) );
  XOR U45150 ( .A(n38751), .B(n38645), .Z(n45720) );
  XNOR U45151 ( .A(n45721), .B(n43355), .Z(n38645) );
  XOR U45152 ( .A(n44535), .B(n45722), .Z(n43355) );
  NOR U45153 ( .A(n44228), .B(n43878), .Z(n45721) );
  XNOR U45154 ( .A(n45723), .B(n45724), .Z(n43878) );
  XOR U45155 ( .A(n42537), .B(n45725), .Z(n44228) );
  IV U45156 ( .A(n41735), .Z(n42537) );
  XOR U45157 ( .A(n45728), .B(n43365), .Z(n38751) );
  XOR U45158 ( .A(n44935), .B(n45729), .Z(n43365) );
  NOR U45159 ( .A(n42946), .B(n42944), .Z(n45728) );
  XOR U45160 ( .A(n45730), .B(n44608), .Z(n42944) );
  XOR U45161 ( .A(n45731), .B(n43713), .Z(n42946) );
  XNOR U45162 ( .A(n45732), .B(n43363), .Z(n43874) );
  XOR U45163 ( .A(n45733), .B(n45734), .Z(n43363) );
  NOR U45164 ( .A(n42942), .B(n42940), .Z(n45732) );
  XOR U45165 ( .A(n45735), .B(n44747), .Z(n42940) );
  XOR U45166 ( .A(n43311), .B(n45736), .Z(n42942) );
  XNOR U45167 ( .A(n45737), .B(n45738), .Z(n43141) );
  XNOR U45168 ( .A(n38439), .B(n40696), .Z(n45738) );
  XNOR U45169 ( .A(n45739), .B(n42568), .Z(n40696) );
  IV U45170 ( .A(n43909), .Z(n42568) );
  XOR U45171 ( .A(n45740), .B(n45453), .Z(n43909) );
  ANDN U45172 ( .B(n44257), .A(n43908), .Z(n45739) );
  XNOR U45173 ( .A(n45741), .B(n43594), .Z(n43908) );
  IV U45174 ( .A(n44267), .Z(n44257) );
  XNOR U45175 ( .A(n45742), .B(n42325), .Z(n44267) );
  XNOR U45176 ( .A(n45743), .B(n42559), .Z(n38439) );
  XOR U45177 ( .A(n45744), .B(n45588), .Z(n42559) );
  ANDN U45178 ( .B(n43896), .A(n41936), .Z(n45743) );
  XOR U45179 ( .A(n45745), .B(n44220), .Z(n41936) );
  XOR U45180 ( .A(n43083), .B(n45746), .Z(n43896) );
  XNOR U45181 ( .A(n41683), .B(n45747), .Z(n45737) );
  XOR U45182 ( .A(n39069), .B(n38819), .Z(n45747) );
  XOR U45183 ( .A(n45748), .B(n42564), .Z(n38819) );
  XOR U45184 ( .A(n45749), .B(n41745), .Z(n42564) );
  XNOR U45185 ( .A(n45750), .B(n45751), .Z(n41745) );
  AND U45186 ( .A(n43901), .B(n41923), .Z(n45748) );
  XNOR U45187 ( .A(n45752), .B(n45753), .Z(n41923) );
  XOR U45188 ( .A(n45754), .B(n44593), .Z(n43901) );
  XOR U45189 ( .A(n45755), .B(n43906), .Z(n39069) );
  XOR U45190 ( .A(n45756), .B(n45216), .Z(n43906) );
  ANDN U45191 ( .B(n41928), .A(n43905), .Z(n45755) );
  XOR U45192 ( .A(n45757), .B(n43716), .Z(n43905) );
  XNOR U45193 ( .A(n45758), .B(n45759), .Z(n41928) );
  XOR U45194 ( .A(n45760), .B(n43892), .Z(n41683) );
  XOR U45195 ( .A(n45761), .B(n44410), .Z(n43892) );
  ANDN U45196 ( .B(n41932), .A(n43891), .Z(n45760) );
  XNOR U45197 ( .A(n45762), .B(n44469), .Z(n43891) );
  XOR U45198 ( .A(n45763), .B(n45764), .Z(n41932) );
  XOR U45199 ( .A(n44953), .B(n37002), .Z(n38716) );
  XOR U45200 ( .A(n39817), .B(n45766), .Z(n37002) );
  XOR U45201 ( .A(n45767), .B(n45768), .Z(n39817) );
  XNOR U45202 ( .A(n42786), .B(n38971), .Z(n45768) );
  XOR U45203 ( .A(n45769), .B(n41003), .Z(n38971) );
  XOR U45204 ( .A(n45770), .B(n45279), .Z(n41003) );
  ANDN U45205 ( .B(n44956), .A(n44955), .Z(n45769) );
  XOR U45206 ( .A(n45771), .B(n43079), .Z(n44955) );
  XNOR U45207 ( .A(n45772), .B(n41006), .Z(n42786) );
  XOR U45208 ( .A(n44461), .B(n45773), .Z(n41006) );
  NOR U45209 ( .A(n42973), .B(n44959), .Z(n45772) );
  XNOR U45210 ( .A(n45774), .B(n43722), .Z(n42973) );
  XNOR U45211 ( .A(n39481), .B(n45775), .Z(n45767) );
  XOR U45212 ( .A(n39921), .B(n39672), .Z(n45775) );
  XOR U45213 ( .A(n45776), .B(n41016), .Z(n39672) );
  XOR U45214 ( .A(n45777), .B(n45778), .Z(n41016) );
  ANDN U45215 ( .B(n44963), .A(n44961), .Z(n45776) );
  XOR U45216 ( .A(n45779), .B(n45554), .Z(n44961) );
  XOR U45217 ( .A(n45780), .B(n41012), .Z(n39921) );
  XOR U45218 ( .A(n45781), .B(n45782), .Z(n41012) );
  ANDN U45219 ( .B(n42980), .A(n45783), .Z(n45780) );
  XNOR U45220 ( .A(n45784), .B(n41020), .Z(n39481) );
  NOR U45221 ( .A(n44965), .B(n42978), .Z(n45784) );
  XNOR U45222 ( .A(n45786), .B(n45787), .Z(n42978) );
  XOR U45223 ( .A(n45788), .B(n42980), .Z(n44953) );
  XOR U45224 ( .A(n45789), .B(n45790), .Z(n42980) );
  ANDN U45225 ( .B(n45783), .A(n41010), .Z(n45788) );
  ANDN U45226 ( .B(n38385), .A(n37993), .Z(n45765) );
  XOR U45227 ( .A(n42104), .B(n36547), .Z(n37993) );
  XOR U45228 ( .A(n39298), .B(n45020), .Z(n36547) );
  XNOR U45229 ( .A(n45791), .B(n45792), .Z(n45020) );
  XOR U45230 ( .A(n36453), .B(n38272), .Z(n45792) );
  XNOR U45231 ( .A(n45793), .B(n45794), .Z(n38272) );
  ANDN U45232 ( .B(n42121), .A(n42119), .Z(n45793) );
  XOR U45233 ( .A(n43577), .B(n45795), .Z(n42121) );
  XNOR U45234 ( .A(n45796), .B(n45797), .Z(n36453) );
  ANDN U45235 ( .B(n45798), .A(n44736), .Z(n45796) );
  XOR U45236 ( .A(n42003), .B(n45799), .Z(n45791) );
  XNOR U45237 ( .A(n38657), .B(n35770), .Z(n45799) );
  XNOR U45238 ( .A(n45800), .B(n42774), .Z(n35770) );
  ANDN U45239 ( .B(n42115), .A(n42117), .Z(n45800) );
  XNOR U45240 ( .A(n43819), .B(n45801), .Z(n42117) );
  XNOR U45241 ( .A(n45802), .B(n42762), .Z(n38657) );
  ANDN U45242 ( .B(n42112), .A(n42111), .Z(n45802) );
  XNOR U45243 ( .A(n42872), .B(n45803), .Z(n42112) );
  XNOR U45244 ( .A(n45804), .B(n42777), .Z(n42003) );
  AND U45245 ( .A(n42106), .B(n42107), .Z(n45804) );
  XOR U45246 ( .A(n45805), .B(n43781), .Z(n42107) );
  XOR U45247 ( .A(n45806), .B(n45807), .Z(n39298) );
  XOR U45248 ( .A(n37670), .B(n40036), .Z(n45807) );
  XOR U45249 ( .A(n45808), .B(n43936), .Z(n40036) );
  XOR U45250 ( .A(n45809), .B(n42526), .Z(n43936) );
  ANDN U45251 ( .B(n43433), .A(n43434), .Z(n45808) );
  XOR U45252 ( .A(n45810), .B(n40856), .Z(n43434) );
  XNOR U45253 ( .A(n45811), .B(n44182), .Z(n43433) );
  XNOR U45254 ( .A(n45812), .B(n45136), .Z(n37670) );
  XNOR U45255 ( .A(n45813), .B(n45814), .Z(n45136) );
  ANDN U45256 ( .B(n43420), .A(n43421), .Z(n45812) );
  XNOR U45257 ( .A(n44497), .B(n45815), .Z(n43421) );
  XOR U45258 ( .A(n44337), .B(n45816), .Z(n43420) );
  XOR U45259 ( .A(n40941), .B(n45817), .Z(n45806) );
  XNOR U45260 ( .A(n43910), .B(n37043), .Z(n45817) );
  XOR U45261 ( .A(n45818), .B(n45118), .Z(n37043) );
  XOR U45262 ( .A(n45819), .B(n41649), .Z(n45118) );
  ANDN U45263 ( .B(n43429), .A(n43430), .Z(n45818) );
  XNOR U45264 ( .A(n45820), .B(n45821), .Z(n43430) );
  XOR U45265 ( .A(n42881), .B(n45822), .Z(n43429) );
  XNOR U45266 ( .A(n45823), .B(n45128), .Z(n43910) );
  IV U45267 ( .A(n43939), .Z(n45128) );
  XOR U45268 ( .A(n45824), .B(n44886), .Z(n43939) );
  IV U45269 ( .A(n44841), .Z(n44886) );
  NOR U45270 ( .A(n43425), .B(n43426), .Z(n45823) );
  XOR U45271 ( .A(n45825), .B(n43706), .Z(n43426) );
  XNOR U45272 ( .A(n45826), .B(n45006), .Z(n43425) );
  XNOR U45273 ( .A(n45827), .B(n43947), .Z(n40941) );
  XNOR U45274 ( .A(n45828), .B(n45829), .Z(n43947) );
  ANDN U45275 ( .B(n43418), .A(n43416), .Z(n45827) );
  IV U45276 ( .A(n43948), .Z(n43416) );
  XOR U45277 ( .A(n45830), .B(n43895), .Z(n43948) );
  XOR U45278 ( .A(n45831), .B(n45268), .Z(n43418) );
  XNOR U45279 ( .A(n45832), .B(n45798), .Z(n42104) );
  ANDN U45280 ( .B(n44736), .A(n42765), .Z(n45832) );
  XNOR U45281 ( .A(n45833), .B(n42877), .Z(n42765) );
  XOR U45282 ( .A(n45834), .B(n45753), .Z(n44736) );
  XOR U45283 ( .A(n44630), .B(n35308), .Z(n38385) );
  XNOR U45284 ( .A(n44340), .B(n40336), .Z(n35308) );
  XNOR U45285 ( .A(n45835), .B(n45836), .Z(n40336) );
  XNOR U45286 ( .A(n39421), .B(n38620), .Z(n45836) );
  XOR U45287 ( .A(n45838), .B(n45371), .Z(n41323) );
  ANDN U45288 ( .B(n41324), .A(n45839), .Z(n45837) );
  XOR U45289 ( .A(n45840), .B(n44232), .Z(n41324) );
  XNOR U45290 ( .A(n45841), .B(n45842), .Z(n39421) );
  NOR U45291 ( .A(n41329), .B(n42917), .Z(n45841) );
  IV U45292 ( .A(n42916), .Z(n41329) );
  XNOR U45293 ( .A(n45843), .B(n45443), .Z(n42916) );
  XOR U45294 ( .A(n39493), .B(n45844), .Z(n45835) );
  XOR U45295 ( .A(n38967), .B(n39439), .Z(n45844) );
  XNOR U45296 ( .A(n45845), .B(n44365), .Z(n39439) );
  IV U45297 ( .A(n43998), .Z(n44365) );
  XOR U45298 ( .A(n45723), .B(n45846), .Z(n43998) );
  ANDN U45299 ( .B(n42922), .A(n43997), .Z(n45845) );
  IV U45300 ( .A(n42920), .Z(n43997) );
  XOR U45301 ( .A(n45847), .B(n45673), .Z(n42920) );
  XOR U45302 ( .A(n45848), .B(n41334), .Z(n38967) );
  NOR U45303 ( .A(n42925), .B(n41333), .Z(n45848) );
  XOR U45304 ( .A(n41874), .B(n45850), .Z(n41333) );
  XOR U45305 ( .A(n45852), .B(n45853), .Z(n41319) );
  ANDN U45306 ( .B(n41320), .A(n42909), .Z(n45851) );
  XOR U45307 ( .A(n45854), .B(n45497), .Z(n41320) );
  XOR U45308 ( .A(n45855), .B(n45856), .Z(n44340) );
  XOR U45309 ( .A(n41297), .B(n38523), .Z(n45856) );
  XOR U45310 ( .A(n45857), .B(n41306), .Z(n38523) );
  XOR U45311 ( .A(n45858), .B(n45859), .Z(n41306) );
  ANDN U45312 ( .B(n44628), .A(n44627), .Z(n45857) );
  XOR U45313 ( .A(n45860), .B(n45861), .Z(n44627) );
  XNOR U45314 ( .A(n45862), .B(n44359), .Z(n41297) );
  XNOR U45315 ( .A(n45863), .B(n42526), .Z(n44359) );
  XNOR U45316 ( .A(n45726), .B(n45864), .Z(n42526) );
  XOR U45317 ( .A(n45865), .B(n45866), .Z(n45726) );
  XNOR U45318 ( .A(n43299), .B(n45867), .Z(n45866) );
  XNOR U45319 ( .A(n45868), .B(n45869), .Z(n43299) );
  ANDN U45320 ( .B(n45870), .A(n45871), .Z(n45868) );
  XOR U45321 ( .A(n44734), .B(n45872), .Z(n45865) );
  XOR U45322 ( .A(n44674), .B(n44779), .Z(n45872) );
  XNOR U45323 ( .A(n45873), .B(n45874), .Z(n44779) );
  XNOR U45324 ( .A(n45877), .B(n45878), .Z(n44674) );
  NOR U45325 ( .A(n45879), .B(n45880), .Z(n45877) );
  XNOR U45326 ( .A(n45881), .B(n45882), .Z(n44734) );
  NOR U45327 ( .A(n45883), .B(n45884), .Z(n45881) );
  ANDN U45328 ( .B(n44360), .A(n44625), .Z(n45862) );
  IV U45329 ( .A(n44624), .Z(n44360) );
  XOR U45330 ( .A(n45885), .B(n43833), .Z(n44624) );
  XOR U45331 ( .A(n38862), .B(n45886), .Z(n45855) );
  XOR U45332 ( .A(n39831), .B(n39752), .Z(n45886) );
  XNOR U45333 ( .A(n45887), .B(n41303), .Z(n39752) );
  XNOR U45334 ( .A(n43600), .B(n45888), .Z(n41303) );
  NOR U45335 ( .A(n44632), .B(n41302), .Z(n45887) );
  XNOR U45336 ( .A(n45889), .B(n45890), .Z(n41302) );
  XNOR U45337 ( .A(n45891), .B(n41605), .Z(n39831) );
  XOR U45338 ( .A(n45892), .B(n45453), .Z(n41605) );
  XOR U45339 ( .A(n45893), .B(n45894), .Z(n45453) );
  ANDN U45340 ( .B(n44635), .A(n41604), .Z(n45891) );
  XOR U45341 ( .A(n45895), .B(n42550), .Z(n41604) );
  XNOR U45342 ( .A(n45896), .B(n44384), .Z(n38862) );
  IV U45343 ( .A(n41314), .Z(n44384) );
  XOR U45344 ( .A(n45897), .B(n45898), .Z(n41314) );
  NOR U45345 ( .A(n41313), .B(n45899), .Z(n45896) );
  XNOR U45346 ( .A(n45900), .B(n41313), .Z(n44630) );
  XNOR U45347 ( .A(n45901), .B(n45902), .Z(n41313) );
  ANDN U45348 ( .B(n45899), .A(n44383), .Z(n45900) );
  XOR U45349 ( .A(n45903), .B(n40053), .Z(n38380) );
  XOR U45350 ( .A(n34626), .B(n45046), .Z(n40053) );
  XNOR U45351 ( .A(n45904), .B(n45905), .Z(n45046) );
  ANDN U45352 ( .B(n40077), .A(n40078), .Z(n45904) );
  XOR U45353 ( .A(n45906), .B(n39795), .Z(n34626) );
  XNOR U45354 ( .A(n45907), .B(n45908), .Z(n39795) );
  XNOR U45355 ( .A(n39327), .B(n44637), .Z(n45908) );
  XOR U45356 ( .A(n45909), .B(n45910), .Z(n44637) );
  NOR U45357 ( .A(n45905), .B(n40077), .Z(n45909) );
  XOR U45358 ( .A(n45911), .B(n45912), .Z(n40077) );
  XOR U45359 ( .A(n45913), .B(n45914), .Z(n39327) );
  ANDN U45360 ( .B(n45058), .A(n45057), .Z(n45913) );
  IV U45361 ( .A(n39964), .Z(n45058) );
  XOR U45362 ( .A(n45915), .B(n45916), .Z(n39964) );
  XNOR U45363 ( .A(n42710), .B(n45917), .Z(n45907) );
  XOR U45364 ( .A(n40437), .B(n43063), .Z(n45917) );
  XNOR U45365 ( .A(n45918), .B(n45919), .Z(n43063) );
  XNOR U45366 ( .A(n4687), .B(n45920), .Z(n45919) );
  OR U45367 ( .A(n39953), .B(n45053), .Z(n45920) );
  XOR U45368 ( .A(n45921), .B(n45922), .Z(n39953) );
  XOR U45369 ( .A(n45923), .B(n45924), .Z(n40437) );
  XOR U45370 ( .A(n45926), .B(n45927), .Z(n42710) );
  XOR U45371 ( .A(n45928), .B(n44500), .Z(n39957) );
  ANDN U45372 ( .B(n38006), .A(n38703), .Z(n45903) );
  IV U45373 ( .A(n38008), .Z(n38703) );
  XNOR U45374 ( .A(n44274), .B(n36555), .Z(n38008) );
  XOR U45375 ( .A(n43042), .B(n41516), .Z(n36555) );
  XNOR U45376 ( .A(n45929), .B(n45930), .Z(n41516) );
  XNOR U45377 ( .A(n37324), .B(n40515), .Z(n45930) );
  XNOR U45378 ( .A(n45931), .B(n42366), .Z(n40515) );
  XOR U45379 ( .A(n45932), .B(n44492), .Z(n42366) );
  AND U45380 ( .A(n42367), .B(n44277), .Z(n45931) );
  XOR U45381 ( .A(n45933), .B(n43524), .Z(n42367) );
  XNOR U45382 ( .A(n45934), .B(n42380), .Z(n37324) );
  XNOR U45383 ( .A(n45935), .B(n42402), .Z(n42380) );
  ANDN U45384 ( .B(n44281), .A(n42379), .Z(n45934) );
  XOR U45385 ( .A(n45936), .B(n41657), .Z(n42379) );
  XNOR U45386 ( .A(n45937), .B(n45938), .Z(n41657) );
  XNOR U45387 ( .A(n39663), .B(n45939), .Z(n45929) );
  XNOR U45388 ( .A(n40624), .B(n40007), .Z(n45939) );
  XOR U45389 ( .A(n45940), .B(n42383), .Z(n40007) );
  XOR U45390 ( .A(n45310), .B(n45941), .Z(n42383) );
  AND U45391 ( .A(n42384), .B(n44288), .Z(n45940) );
  XOR U45392 ( .A(n45942), .B(n45644), .Z(n42384) );
  XNOR U45393 ( .A(n45943), .B(n42370), .Z(n40624) );
  ANDN U45394 ( .B(n44285), .A(n44283), .Z(n45943) );
  XOR U45395 ( .A(n45944), .B(n45945), .Z(n44283) );
  XNOR U45396 ( .A(n45946), .B(n42375), .Z(n39663) );
  XOR U45397 ( .A(n45947), .B(n42501), .Z(n42375) );
  ANDN U45398 ( .B(n42376), .A(n45948), .Z(n45946) );
  XNOR U45399 ( .A(n45949), .B(n45950), .Z(n43042) );
  XNOR U45400 ( .A(n38261), .B(n38499), .Z(n45950) );
  XOR U45401 ( .A(n45951), .B(n42294), .Z(n38499) );
  XOR U45402 ( .A(n45952), .B(n45953), .Z(n42294) );
  ANDN U45403 ( .B(n42295), .A(n44296), .Z(n45951) );
  XNOR U45404 ( .A(n45954), .B(n43327), .Z(n42295) );
  XNOR U45405 ( .A(n45955), .B(n42280), .Z(n38261) );
  XNOR U45406 ( .A(n45956), .B(n45091), .Z(n42280) );
  ANDN U45407 ( .B(n42281), .A(n45957), .Z(n45955) );
  XOR U45408 ( .A(n45958), .B(n44839), .Z(n42281) );
  XNOR U45409 ( .A(n42254), .B(n45959), .Z(n45949) );
  XNOR U45410 ( .A(n41718), .B(n38603), .Z(n45959) );
  XNOR U45411 ( .A(n45960), .B(n42284), .Z(n38603) );
  XNOR U45412 ( .A(n45961), .B(n45443), .Z(n42284) );
  ANDN U45413 ( .B(n42285), .A(n45962), .Z(n45960) );
  XNOR U45414 ( .A(n45963), .B(n42681), .Z(n42285) );
  XNOR U45415 ( .A(n45964), .B(n45106), .Z(n41718) );
  XOR U45416 ( .A(n44579), .B(n45965), .Z(n45106) );
  NOR U45417 ( .A(n45966), .B(n44299), .Z(n45964) );
  XOR U45418 ( .A(n45967), .B(n43781), .Z(n44299) );
  IV U45419 ( .A(n45968), .Z(n43781) );
  XNOR U45420 ( .A(n45969), .B(n42290), .Z(n42254) );
  XOR U45421 ( .A(n42689), .B(n45970), .Z(n42290) );
  ANDN U45422 ( .B(n42291), .A(n44292), .Z(n45969) );
  XNOR U45423 ( .A(n45971), .B(n45172), .Z(n42291) );
  XOR U45424 ( .A(n45972), .B(n42376), .Z(n44274) );
  XNOR U45425 ( .A(n45973), .B(n45974), .Z(n42376) );
  ANDN U45426 ( .B(n45948), .A(n45476), .Z(n45972) );
  IV U45427 ( .A(n45975), .Z(n45476) );
  XOR U45428 ( .A(n45976), .B(n38037), .Z(n38006) );
  XNOR U45429 ( .A(n45977), .B(n44944), .Z(n38037) );
  XOR U45430 ( .A(n45978), .B(n45979), .Z(n44944) );
  XNOR U45431 ( .A(n35305), .B(n38377), .Z(n45979) );
  XNOR U45432 ( .A(n45980), .B(n44818), .Z(n38377) );
  XOR U45433 ( .A(n45981), .B(n45982), .Z(n44818) );
  NOR U45434 ( .A(n43232), .B(n44828), .Z(n45980) );
  XNOR U45435 ( .A(n45983), .B(n42731), .Z(n35305) );
  XOR U45436 ( .A(n45984), .B(n43303), .Z(n42731) );
  NOR U45437 ( .A(n45985), .B(n42732), .Z(n45983) );
  XNOR U45438 ( .A(n39948), .B(n45986), .Z(n45978) );
  XNOR U45439 ( .A(n39385), .B(n39365), .Z(n45986) );
  XNOR U45440 ( .A(n45987), .B(n42727), .Z(n39365) );
  XNOR U45441 ( .A(n45988), .B(n43574), .Z(n42727) );
  NOR U45442 ( .A(n43228), .B(n42728), .Z(n45987) );
  XOR U45443 ( .A(n45989), .B(n42718), .Z(n39385) );
  XNOR U45444 ( .A(n45990), .B(n42681), .Z(n42718) );
  ANDN U45445 ( .B(n42719), .A(n43225), .Z(n45989) );
  XOR U45446 ( .A(n45991), .B(n42724), .Z(n39948) );
  XOR U45447 ( .A(n45992), .B(n45993), .Z(n42724) );
  NOR U45448 ( .A(n43221), .B(n42723), .Z(n45991) );
  XOR U45449 ( .A(n35651), .B(n31632), .Z(n28990) );
  XNOR U45450 ( .A(n45994), .B(n45995), .Z(n38225) );
  XOR U45451 ( .A(n32830), .B(n29272), .Z(n45995) );
  XNOR U45452 ( .A(n45996), .B(n35426), .Z(n29272) );
  XOR U45453 ( .A(n42585), .B(n38640), .Z(n35426) );
  XOR U45454 ( .A(n39743), .B(n41148), .Z(n38640) );
  XNOR U45455 ( .A(n45997), .B(n45998), .Z(n41148) );
  XOR U45456 ( .A(n43047), .B(n38508), .Z(n45998) );
  XOR U45457 ( .A(n45999), .B(n41497), .Z(n38508) );
  XOR U45458 ( .A(n43665), .B(n46000), .Z(n41497) );
  AND U45459 ( .A(n42580), .B(n42579), .Z(n45999) );
  XNOR U45460 ( .A(n46001), .B(n42550), .Z(n42579) );
  XNOR U45461 ( .A(n46002), .B(n40264), .Z(n43047) );
  XOR U45462 ( .A(n46003), .B(n42342), .Z(n40264) );
  ANDN U45463 ( .B(n46004), .A(n43055), .Z(n46002) );
  XNOR U45464 ( .A(n37345), .B(n46005), .Z(n45997) );
  XNOR U45465 ( .A(n41754), .B(n40695), .Z(n46005) );
  XOR U45466 ( .A(n46006), .B(n40261), .Z(n40695) );
  XOR U45467 ( .A(n46008), .B(n44596), .Z(n42582) );
  XNOR U45468 ( .A(n46009), .B(n40257), .Z(n41754) );
  XOR U45469 ( .A(n46010), .B(n44523), .Z(n40257) );
  ANDN U45470 ( .B(n42816), .A(n42815), .Z(n46009) );
  XOR U45471 ( .A(n45386), .B(n46011), .Z(n42815) );
  XNOR U45472 ( .A(n46012), .B(n43053), .Z(n37345) );
  IV U45473 ( .A(n43621), .Z(n43053) );
  XOR U45474 ( .A(n46013), .B(n45448), .Z(n43621) );
  IV U45475 ( .A(n46014), .Z(n45448) );
  ANDN U45476 ( .B(n42588), .A(n42589), .Z(n46012) );
  XOR U45477 ( .A(n46015), .B(n44503), .Z(n42588) );
  XOR U45478 ( .A(n46016), .B(n46017), .Z(n39743) );
  XOR U45479 ( .A(n37712), .B(n37048), .Z(n46017) );
  XOR U45480 ( .A(n46018), .B(n41538), .Z(n37048) );
  XOR U45481 ( .A(n46019), .B(n44777), .Z(n41538) );
  NOR U45482 ( .A(n43618), .B(n44116), .Z(n46018) );
  XNOR U45483 ( .A(n42846), .B(n46020), .Z(n44116) );
  IV U45484 ( .A(n46021), .Z(n42846) );
  IV U45485 ( .A(n44117), .Z(n43618) );
  XOR U45486 ( .A(n46022), .B(n46023), .Z(n44117) );
  XNOR U45487 ( .A(n46024), .B(n41525), .Z(n37712) );
  XOR U45488 ( .A(n46025), .B(n42419), .Z(n41525) );
  NOR U45489 ( .A(n45695), .B(n44099), .Z(n46024) );
  XNOR U45490 ( .A(n46026), .B(n46027), .Z(n44099) );
  XNOR U45491 ( .A(n46028), .B(n43108), .Z(n45695) );
  XOR U45492 ( .A(n35610), .B(n46029), .Z(n46016) );
  XOR U45493 ( .A(n45675), .B(n43681), .Z(n46029) );
  XNOR U45494 ( .A(n46030), .B(n41542), .Z(n43681) );
  XOR U45495 ( .A(n46031), .B(n46032), .Z(n41542) );
  NOR U45496 ( .A(n43616), .B(n44103), .Z(n46030) );
  XNOR U45497 ( .A(n46033), .B(n43916), .Z(n44103) );
  IV U45498 ( .A(n44104), .Z(n43616) );
  XNOR U45499 ( .A(n46035), .B(n41529), .Z(n45675) );
  XNOR U45500 ( .A(n42667), .B(n46036), .Z(n41529) );
  NOR U45501 ( .A(n43612), .B(n44121), .Z(n46035) );
  XOR U45502 ( .A(n46037), .B(n45597), .Z(n44121) );
  IV U45503 ( .A(n44263), .Z(n45597) );
  XOR U45504 ( .A(n46038), .B(n45938), .Z(n44263) );
  XNOR U45505 ( .A(n46039), .B(n46040), .Z(n45938) );
  XNOR U45506 ( .A(n46041), .B(n46042), .Z(n46040) );
  XOR U45507 ( .A(n46043), .B(n46044), .Z(n46039) );
  XOR U45508 ( .A(n45433), .B(n44618), .Z(n46044) );
  XNOR U45509 ( .A(n46045), .B(n46046), .Z(n44618) );
  ANDN U45510 ( .B(n46047), .A(n46048), .Z(n46045) );
  XNOR U45511 ( .A(n46049), .B(n46050), .Z(n45433) );
  ANDN U45512 ( .B(n46051), .A(n46052), .Z(n46049) );
  IV U45513 ( .A(n44122), .Z(n43612) );
  XOR U45514 ( .A(n46053), .B(n46054), .Z(n44122) );
  XNOR U45515 ( .A(n46055), .B(n41534), .Z(n35610) );
  XNOR U45516 ( .A(n46056), .B(n46057), .Z(n41534) );
  NOR U45517 ( .A(n43609), .B(n44112), .Z(n46055) );
  XNOR U45518 ( .A(n46058), .B(n46059), .Z(n44112) );
  XNOR U45519 ( .A(n46060), .B(n40849), .Z(n43609) );
  XOR U45520 ( .A(n46061), .B(n43055), .Z(n42585) );
  XOR U45521 ( .A(n46062), .B(n43337), .Z(n43055) );
  NOR U45522 ( .A(n46004), .B(n40263), .Z(n46061) );
  ANDN U45523 ( .B(n34204), .A(n38228), .Z(n45996) );
  IV U45524 ( .A(n35427), .Z(n38228) );
  XOR U45525 ( .A(n43219), .B(n37000), .Z(n35427) );
  XNOR U45526 ( .A(n43628), .B(n44656), .Z(n37000) );
  XOR U45527 ( .A(n46063), .B(n46064), .Z(n44656) );
  XNOR U45528 ( .A(n38753), .B(n37866), .Z(n46064) );
  XOR U45529 ( .A(n46065), .B(n39966), .Z(n37866) );
  ANDN U45530 ( .B(n45057), .A(n46066), .Z(n46065) );
  XOR U45531 ( .A(n46067), .B(n46068), .Z(n45057) );
  XNOR U45532 ( .A(n46069), .B(n40079), .Z(n38753) );
  XOR U45533 ( .A(n46070), .B(n46071), .Z(n45905) );
  XOR U45534 ( .A(n46072), .B(n46073), .Z(n46063) );
  XNOR U45535 ( .A(n39119), .B(n35939), .Z(n46073) );
  XNOR U45536 ( .A(n46074), .B(n39959), .Z(n35939) );
  ANDN U45537 ( .B(n45927), .A(n45055), .Z(n46074) );
  XOR U45538 ( .A(n42668), .B(n46075), .Z(n45055) );
  XNOR U45539 ( .A(n46076), .B(n45060), .Z(n39119) );
  NOR U45540 ( .A(n45048), .B(n45924), .Z(n46076) );
  XOR U45541 ( .A(n46077), .B(n44564), .Z(n45048) );
  XNOR U45542 ( .A(n46078), .B(n46079), .Z(n43628) );
  XNOR U45543 ( .A(n39843), .B(n38465), .Z(n46079) );
  XOR U45544 ( .A(n46080), .B(n42719), .Z(n38465) );
  XOR U45545 ( .A(n46081), .B(n45216), .Z(n42719) );
  AND U45546 ( .A(n43226), .B(n43225), .Z(n46080) );
  XNOR U45547 ( .A(n46082), .B(n45902), .Z(n43225) );
  XOR U45548 ( .A(n46083), .B(n44207), .Z(n43226) );
  XNOR U45549 ( .A(n46084), .B(n42723), .Z(n39843) );
  XOR U45550 ( .A(n46085), .B(n46086), .Z(n42723) );
  AND U45551 ( .A(n43222), .B(n43221), .Z(n46084) );
  XOR U45552 ( .A(n46087), .B(n43555), .Z(n43221) );
  IV U45553 ( .A(n43472), .Z(n43555) );
  XOR U45554 ( .A(n46088), .B(n46068), .Z(n43222) );
  IV U45555 ( .A(n45753), .Z(n46068) );
  XOR U45556 ( .A(n38036), .B(n46089), .Z(n46078) );
  XOR U45557 ( .A(n39458), .B(n45976), .Z(n46089) );
  XOR U45558 ( .A(n46090), .B(n42732), .Z(n45976) );
  XOR U45559 ( .A(n45159), .B(n46091), .Z(n42732) );
  AND U45560 ( .A(n44823), .B(n45985), .Z(n46090) );
  XOR U45561 ( .A(n46092), .B(n44828), .Z(n39458) );
  XNOR U45562 ( .A(n46093), .B(n45249), .Z(n44828) );
  ANDN U45563 ( .B(n43232), .A(n43234), .Z(n46092) );
  XOR U45564 ( .A(n46094), .B(n44777), .Z(n43234) );
  XOR U45565 ( .A(n46095), .B(n45091), .Z(n43232) );
  XOR U45566 ( .A(n46096), .B(n42728), .Z(n38036) );
  XOR U45567 ( .A(n46097), .B(n42877), .Z(n42728) );
  XNOR U45568 ( .A(n46098), .B(n43846), .Z(n43228) );
  XNOR U45569 ( .A(n46099), .B(n46100), .Z(n43846) );
  XOR U45570 ( .A(n46101), .B(n44806), .Z(n43229) );
  XNOR U45571 ( .A(n46102), .B(n45985), .Z(n43219) );
  XOR U45572 ( .A(n46103), .B(n46104), .Z(n45985) );
  ANDN U45573 ( .B(n42730), .A(n44823), .Z(n46102) );
  XOR U45574 ( .A(n46105), .B(n44119), .Z(n44823) );
  XOR U45575 ( .A(n46106), .B(n46107), .Z(n42730) );
  XNOR U45576 ( .A(n45684), .B(n36970), .Z(n34204) );
  XOR U45577 ( .A(n40533), .B(n41519), .Z(n36970) );
  XNOR U45578 ( .A(n46108), .B(n46109), .Z(n41519) );
  XOR U45579 ( .A(n35623), .B(n39130), .Z(n46109) );
  XOR U45580 ( .A(n46110), .B(n44132), .Z(n39130) );
  XNOR U45581 ( .A(n46111), .B(n44816), .Z(n44132) );
  ANDN U45582 ( .B(n44980), .A(n42993), .Z(n46110) );
  XNOR U45583 ( .A(n46112), .B(n44127), .Z(n35623) );
  XNOR U45584 ( .A(n46113), .B(n42309), .Z(n44127) );
  ANDN U45585 ( .B(n44971), .A(n42997), .Z(n46112) );
  IV U45586 ( .A(n45681), .Z(n42997) );
  XNOR U45587 ( .A(n45786), .B(n46114), .Z(n45681) );
  XNOR U45588 ( .A(n44693), .B(n46115), .Z(n44971) );
  XNOR U45589 ( .A(n44950), .B(n46116), .Z(n46108) );
  XOR U45590 ( .A(n39749), .B(n35584), .Z(n46116) );
  XNOR U45591 ( .A(n46117), .B(n44134), .Z(n35584) );
  XOR U45592 ( .A(n46118), .B(n44328), .Z(n44134) );
  IV U45593 ( .A(n44225), .Z(n44328) );
  ANDN U45594 ( .B(n44983), .A(n42984), .Z(n46117) );
  XNOR U45595 ( .A(n46119), .B(n46120), .Z(n42984) );
  XOR U45596 ( .A(n46121), .B(n45922), .Z(n44983) );
  XNOR U45597 ( .A(n46122), .B(n44137), .Z(n39749) );
  XNOR U45598 ( .A(n45565), .B(n46123), .Z(n44137) );
  ANDN U45599 ( .B(n44987), .A(n42988), .Z(n46122) );
  XOR U45600 ( .A(n46124), .B(n44199), .Z(n42988) );
  XOR U45601 ( .A(n43583), .B(n46125), .Z(n44987) );
  XOR U45602 ( .A(n46126), .B(n46127), .Z(n43583) );
  XNOR U45603 ( .A(n46128), .B(n44974), .Z(n44950) );
  IV U45604 ( .A(n44129), .Z(n44974) );
  XOR U45605 ( .A(n46129), .B(n43530), .Z(n44129) );
  IV U45606 ( .A(n45759), .Z(n43530) );
  ANDN U45607 ( .B(n44975), .A(n43001), .Z(n46128) );
  IV U45608 ( .A(n45686), .Z(n43001) );
  XOR U45609 ( .A(n46130), .B(n43108), .Z(n45686) );
  XNOR U45610 ( .A(n46131), .B(n45894), .Z(n43108) );
  XNOR U45611 ( .A(n46132), .B(n46133), .Z(n45894) );
  XNOR U45612 ( .A(n44187), .B(n46134), .Z(n46133) );
  XOR U45613 ( .A(n46135), .B(n46136), .Z(n44187) );
  ANDN U45614 ( .B(n46137), .A(n46138), .Z(n46135) );
  XOR U45615 ( .A(n46139), .B(n46140), .Z(n46132) );
  XOR U45616 ( .A(n43580), .B(n42493), .Z(n46140) );
  XNOR U45617 ( .A(n46141), .B(n46142), .Z(n42493) );
  XNOR U45618 ( .A(n46145), .B(n46146), .Z(n43580) );
  AND U45619 ( .A(n46147), .B(n46148), .Z(n46145) );
  XOR U45620 ( .A(n44847), .B(n46149), .Z(n44975) );
  XOR U45621 ( .A(n46150), .B(n46151), .Z(n40533) );
  XOR U45622 ( .A(n39586), .B(n37645), .Z(n46151) );
  XOR U45623 ( .A(n46152), .B(n44965), .Z(n37645) );
  XOR U45624 ( .A(n46153), .B(n42503), .Z(n44965) );
  ANDN U45625 ( .B(n41018), .A(n41019), .Z(n46152) );
  XNOR U45626 ( .A(n45148), .B(n46154), .Z(n41019) );
  XNOR U45627 ( .A(n46155), .B(n45466), .Z(n41018) );
  XNOR U45628 ( .A(n46156), .B(n45783), .Z(n39586) );
  XOR U45629 ( .A(n46157), .B(n46158), .Z(n45783) );
  ANDN U45630 ( .B(n41010), .A(n41011), .Z(n46156) );
  XNOR U45631 ( .A(n44472), .B(n46159), .Z(n41011) );
  XOR U45632 ( .A(n44225), .B(n46160), .Z(n41010) );
  XOR U45633 ( .A(n40511), .B(n46161), .Z(n46150) );
  XOR U45634 ( .A(n38679), .B(n39079), .Z(n46161) );
  XNOR U45635 ( .A(n46162), .B(n44963), .Z(n39079) );
  XOR U45636 ( .A(n46163), .B(n44767), .Z(n44963) );
  NOR U45637 ( .A(n44962), .B(n41015), .Z(n46162) );
  XNOR U45638 ( .A(n46164), .B(n46165), .Z(n41015) );
  IV U45639 ( .A(n41014), .Z(n44962) );
  XOR U45640 ( .A(n46166), .B(n46167), .Z(n41014) );
  XNOR U45641 ( .A(n46168), .B(n44956), .Z(n38679) );
  XOR U45642 ( .A(n46169), .B(n44743), .Z(n44956) );
  ANDN U45643 ( .B(n41001), .A(n41002), .Z(n46168) );
  XOR U45644 ( .A(n46170), .B(n43671), .Z(n41002) );
  XNOR U45645 ( .A(n46171), .B(n46172), .Z(n41001) );
  XNOR U45646 ( .A(n46173), .B(n44959), .Z(n40511) );
  XOR U45647 ( .A(n45322), .B(n46174), .Z(n44959) );
  IV U45648 ( .A(n44693), .Z(n45322) );
  XOR U45649 ( .A(n46175), .B(n45898), .Z(n41005) );
  IV U45650 ( .A(n46176), .Z(n45898) );
  XOR U45651 ( .A(n46177), .B(n46178), .Z(n41007) );
  XNOR U45652 ( .A(n46179), .B(n44980), .Z(n45684) );
  XNOR U45653 ( .A(n46171), .B(n46180), .Z(n44980) );
  IV U45654 ( .A(n46181), .Z(n46171) );
  ANDN U45655 ( .B(n42993), .A(n42995), .Z(n46179) );
  XOR U45656 ( .A(n46182), .B(n46183), .Z(n42995) );
  XOR U45657 ( .A(n46184), .B(n46185), .Z(n42993) );
  XOR U45658 ( .A(n43508), .B(n37880), .Z(n35423) );
  IV U45659 ( .A(n38171), .Z(n37880) );
  XNOR U45660 ( .A(n40335), .B(n40098), .Z(n38171) );
  XNOR U45661 ( .A(n46187), .B(n46188), .Z(n40098) );
  XOR U45662 ( .A(n40143), .B(n42612), .Z(n46188) );
  XOR U45663 ( .A(n46189), .B(n42617), .Z(n42612) );
  XOR U45664 ( .A(n46190), .B(n43280), .Z(n42617) );
  IV U45665 ( .A(n43706), .Z(n43280) );
  XOR U45666 ( .A(n46191), .B(n46192), .Z(n43706) );
  AND U45667 ( .A(n43795), .B(n42618), .Z(n46189) );
  XNOR U45668 ( .A(n46193), .B(n46194), .Z(n42618) );
  XOR U45669 ( .A(n46195), .B(n42628), .Z(n40143) );
  XOR U45670 ( .A(n46196), .B(n45395), .Z(n42628) );
  ANDN U45671 ( .B(n43799), .A(n43797), .Z(n46195) );
  XOR U45672 ( .A(n46197), .B(n46198), .Z(n43797) );
  XOR U45673 ( .A(n39448), .B(n46199), .Z(n46187) );
  XOR U45674 ( .A(n40995), .B(n39937), .Z(n46199) );
  XNOR U45675 ( .A(n46200), .B(n42631), .Z(n39937) );
  ANDN U45676 ( .B(n42632), .A(n43802), .Z(n46200) );
  XNOR U45677 ( .A(n46201), .B(n45121), .Z(n42632) );
  XNOR U45678 ( .A(n46202), .B(n42621), .Z(n40995) );
  XOR U45679 ( .A(n46203), .B(n42306), .Z(n42621) );
  XOR U45680 ( .A(n45252), .B(n46204), .Z(n42622) );
  IV U45681 ( .A(n46205), .Z(n43806) );
  XNOR U45682 ( .A(n46206), .B(n45612), .Z(n39448) );
  XNOR U45683 ( .A(n46207), .B(n46208), .Z(n45612) );
  XOR U45684 ( .A(n44163), .B(n46209), .Z(n43808) );
  XNOR U45685 ( .A(n46210), .B(n46211), .Z(n44163) );
  XOR U45686 ( .A(n46212), .B(n46213), .Z(n40335) );
  XNOR U45687 ( .A(n38023), .B(n38850), .Z(n46213) );
  XNOR U45688 ( .A(n46214), .B(n39500), .Z(n38850) );
  XOR U45689 ( .A(n42872), .B(n46215), .Z(n39500) );
  IV U45690 ( .A(n44663), .Z(n42872) );
  AND U45691 ( .A(n39501), .B(n43514), .Z(n46214) );
  XNOR U45692 ( .A(n46216), .B(n42404), .Z(n39501) );
  IV U45693 ( .A(n45252), .Z(n42404) );
  XNOR U45694 ( .A(n46217), .B(n39509), .Z(n38023) );
  XNOR U45695 ( .A(n45151), .B(n46218), .Z(n39509) );
  XOR U45696 ( .A(n42517), .B(n46219), .Z(n39510) );
  XNOR U45697 ( .A(n39289), .B(n46220), .Z(n46212) );
  XNOR U45698 ( .A(n35515), .B(n38671), .Z(n46220) );
  XNOR U45699 ( .A(n46221), .B(n40363), .Z(n38671) );
  XOR U45700 ( .A(n46222), .B(n42166), .Z(n40363) );
  AND U45701 ( .A(n40364), .B(n43511), .Z(n46221) );
  XOR U45702 ( .A(n46223), .B(n42683), .Z(n40364) );
  XOR U45703 ( .A(n46224), .B(n39513), .Z(n35515) );
  XOR U45704 ( .A(n43865), .B(n46225), .Z(n39513) );
  ANDN U45705 ( .B(n39514), .A(n46226), .Z(n46224) );
  XOR U45706 ( .A(n45014), .B(n46227), .Z(n39514) );
  XOR U45707 ( .A(n46228), .B(n39505), .Z(n39289) );
  XNOR U45708 ( .A(n46229), .B(n46198), .Z(n39505) );
  XNOR U45709 ( .A(n46231), .B(n39506), .Z(n43508) );
  XOR U45710 ( .A(n45348), .B(n46232), .Z(n39506) );
  ANDN U45711 ( .B(n43987), .A(n46230), .Z(n46231) );
  ANDN U45712 ( .B(n34200), .A(n46233), .Z(n46186) );
  IV U45713 ( .A(n35424), .Z(n46233) );
  XOR U45714 ( .A(n45473), .B(n38564), .Z(n35424) );
  XOR U45715 ( .A(n41994), .B(n44140), .Z(n38564) );
  XNOR U45716 ( .A(n46234), .B(n46235), .Z(n44140) );
  XNOR U45717 ( .A(n40622), .B(n38143), .Z(n46235) );
  XOR U45718 ( .A(n46236), .B(n44307), .Z(n38143) );
  IV U45719 ( .A(n45962), .Z(n44307) );
  XOR U45720 ( .A(n46139), .B(n42494), .Z(n45962) );
  XNOR U45721 ( .A(n46237), .B(n46238), .Z(n46139) );
  ANDN U45722 ( .B(n46239), .A(n46240), .Z(n46237) );
  NOR U45723 ( .A(n44306), .B(n42283), .Z(n46236) );
  XOR U45724 ( .A(n46241), .B(n45397), .Z(n42283) );
  XNOR U45725 ( .A(n45565), .B(n46242), .Z(n44306) );
  XNOR U45726 ( .A(n46243), .B(n44292), .Z(n40622) );
  XOR U45727 ( .A(n46244), .B(n44915), .Z(n44292) );
  XOR U45728 ( .A(n42395), .B(n46245), .Z(n42289) );
  XOR U45729 ( .A(n46246), .B(n43083), .Z(n44293) );
  XOR U45730 ( .A(n41021), .B(n46247), .Z(n46234) );
  XOR U45731 ( .A(n41118), .B(n40436), .Z(n46247) );
  XNOR U45732 ( .A(n46248), .B(n45966), .Z(n40436) );
  IV U45733 ( .A(n44300), .Z(n45966) );
  XOR U45734 ( .A(n46249), .B(n45203), .Z(n44300) );
  ANDN U45735 ( .B(n44301), .A(n45110), .Z(n46248) );
  IV U45736 ( .A(n45107), .Z(n45110) );
  XNOR U45737 ( .A(n46250), .B(n42306), .Z(n45107) );
  XNOR U45738 ( .A(n46251), .B(n42327), .Z(n44301) );
  XNOR U45739 ( .A(n46252), .B(n45957), .Z(n41118) );
  IV U45740 ( .A(n44303), .Z(n45957) );
  XOR U45741 ( .A(n46253), .B(n41883), .Z(n44303) );
  ANDN U45742 ( .B(n44304), .A(n42279), .Z(n46252) );
  IV U45743 ( .A(n45101), .Z(n42279) );
  XNOR U45744 ( .A(n46254), .B(n46166), .Z(n45101) );
  XOR U45745 ( .A(n44845), .B(n46255), .Z(n44304) );
  XNOR U45746 ( .A(n46256), .B(n44296), .Z(n41021) );
  XOR U45747 ( .A(n46257), .B(n45644), .Z(n44296) );
  ANDN U45748 ( .B(n44295), .A(n42293), .Z(n46256) );
  XNOR U45749 ( .A(n46258), .B(n43965), .Z(n42293) );
  XOR U45750 ( .A(n46259), .B(n45274), .Z(n44295) );
  IV U45751 ( .A(n43330), .Z(n45274) );
  XOR U45752 ( .A(n46260), .B(n46261), .Z(n41994) );
  XNOR U45753 ( .A(n44271), .B(n37499), .Z(n46261) );
  XOR U45754 ( .A(n46262), .B(n44281), .Z(n37499) );
  XOR U45755 ( .A(n44461), .B(n46263), .Z(n44281) );
  NOR U45756 ( .A(n44280), .B(n42378), .Z(n46262) );
  XNOR U45757 ( .A(n45504), .B(n46264), .Z(n42378) );
  XNOR U45758 ( .A(n46265), .B(n44191), .Z(n44280) );
  XOR U45759 ( .A(n46266), .B(n44277), .Z(n44271) );
  XNOR U45760 ( .A(n46267), .B(n42681), .Z(n44277) );
  XNOR U45761 ( .A(n46268), .B(n46269), .Z(n42681) );
  NOR U45762 ( .A(n44276), .B(n42365), .Z(n46266) );
  XOR U45763 ( .A(n46270), .B(n44673), .Z(n42365) );
  IV U45764 ( .A(n45478), .Z(n44276) );
  XOR U45765 ( .A(n42689), .B(n46271), .Z(n45478) );
  XOR U45766 ( .A(n46272), .B(n46273), .Z(n42689) );
  XNOR U45767 ( .A(n38425), .B(n46274), .Z(n46260) );
  XNOR U45768 ( .A(n40832), .B(n40298), .Z(n46274) );
  XOR U45769 ( .A(n46275), .B(n44288), .Z(n40298) );
  XOR U45770 ( .A(n46276), .B(n45463), .Z(n44288) );
  IV U45771 ( .A(n44014), .Z(n45463) );
  NOR U45772 ( .A(n44287), .B(n42382), .Z(n46275) );
  XOR U45773 ( .A(n45789), .B(n46277), .Z(n42382) );
  XOR U45774 ( .A(n46278), .B(n45386), .Z(n44287) );
  XOR U45775 ( .A(n46279), .B(n45948), .Z(n40832) );
  XOR U45776 ( .A(n46280), .B(n41883), .Z(n45948) );
  NOR U45777 ( .A(n45975), .B(n42374), .Z(n46279) );
  XOR U45778 ( .A(n46281), .B(n46282), .Z(n42374) );
  XOR U45779 ( .A(n46283), .B(n44882), .Z(n45975) );
  XNOR U45780 ( .A(n46284), .B(n44285), .Z(n38425) );
  XOR U45781 ( .A(n46285), .B(n45395), .Z(n44285) );
  IV U45782 ( .A(n46286), .Z(n45395) );
  ANDN U45783 ( .B(n44284), .A(n42369), .Z(n46284) );
  XNOR U45784 ( .A(n46287), .B(n44284), .Z(n45473) );
  XOR U45785 ( .A(n43784), .B(n46288), .Z(n44284) );
  ANDN U45786 ( .B(n42369), .A(n42370), .Z(n46287) );
  XOR U45787 ( .A(n46289), .B(n46032), .Z(n42370) );
  XOR U45788 ( .A(n42319), .B(n46290), .Z(n42369) );
  XNOR U45789 ( .A(n46291), .B(n46292), .Z(n42319) );
  XNOR U45790 ( .A(n42249), .B(n39213), .Z(n34200) );
  IV U45791 ( .A(n43515), .Z(n39213) );
  XOR U45792 ( .A(n41232), .B(n40641), .Z(n43515) );
  XOR U45793 ( .A(n46293), .B(n46294), .Z(n40641) );
  XOR U45794 ( .A(n39885), .B(n37113), .Z(n46294) );
  XOR U45795 ( .A(n46295), .B(n43744), .Z(n37113) );
  XOR U45796 ( .A(n46296), .B(n45656), .Z(n43744) );
  ANDN U45797 ( .B(n42240), .A(n42242), .Z(n46295) );
  XNOR U45798 ( .A(n44337), .B(n46297), .Z(n42240) );
  XNOR U45799 ( .A(n46298), .B(n43747), .Z(n39885) );
  XOR U45800 ( .A(n46166), .B(n46299), .Z(n43747) );
  XOR U45801 ( .A(n46300), .B(n43765), .Z(n42244) );
  XOR U45802 ( .A(n43728), .B(n46301), .Z(n46293) );
  XOR U45803 ( .A(n42947), .B(n38993), .Z(n46301) );
  XNOR U45804 ( .A(n46302), .B(n43733), .Z(n38993) );
  XOR U45805 ( .A(n44535), .B(n46303), .Z(n43733) );
  NOR U45806 ( .A(n46304), .B(n46305), .Z(n46302) );
  XOR U45807 ( .A(n46307), .B(n45339), .Z(n43741) );
  NOR U45808 ( .A(n43519), .B(n43517), .Z(n46306) );
  XOR U45809 ( .A(n46308), .B(n46120), .Z(n43517) );
  XNOR U45810 ( .A(n46309), .B(n45528), .Z(n43728) );
  IV U45811 ( .A(n43737), .Z(n45528) );
  XOR U45812 ( .A(n46310), .B(n45011), .Z(n43737) );
  NOR U45813 ( .A(n42252), .B(n42251), .Z(n46309) );
  XOR U45814 ( .A(n46311), .B(n45764), .Z(n42251) );
  IV U45815 ( .A(n46312), .Z(n42252) );
  XOR U45816 ( .A(n46313), .B(n46314), .Z(n41232) );
  XNOR U45817 ( .A(n37149), .B(n39866), .Z(n46314) );
  XNOR U45818 ( .A(n46315), .B(n42140), .Z(n39866) );
  XOR U45819 ( .A(n46316), .B(n43916), .Z(n42140) );
  NOR U45820 ( .A(n43128), .B(n43127), .Z(n46315) );
  XOR U45821 ( .A(n46317), .B(n44837), .Z(n43127) );
  XOR U45822 ( .A(n46318), .B(n45644), .Z(n43128) );
  XOR U45823 ( .A(n46319), .B(n46192), .Z(n45644) );
  XNOR U45824 ( .A(n46320), .B(n46321), .Z(n46192) );
  XNOR U45825 ( .A(n46015), .B(n45707), .Z(n46321) );
  XOR U45826 ( .A(n46322), .B(n46323), .Z(n45707) );
  ANDN U45827 ( .B(n46324), .A(n46325), .Z(n46322) );
  XOR U45828 ( .A(n46326), .B(n46327), .Z(n46015) );
  ANDN U45829 ( .B(n46328), .A(n46329), .Z(n46326) );
  XNOR U45830 ( .A(n46330), .B(n46331), .Z(n46320) );
  XOR U45831 ( .A(n44502), .B(n44326), .Z(n46331) );
  XOR U45832 ( .A(n46332), .B(n46333), .Z(n44326) );
  ANDN U45833 ( .B(n46334), .A(n46335), .Z(n46332) );
  XNOR U45834 ( .A(n46336), .B(n46337), .Z(n44502) );
  ANDN U45835 ( .B(n46338), .A(n46339), .Z(n46336) );
  XNOR U45836 ( .A(n46340), .B(n42136), .Z(n37149) );
  ANDN U45837 ( .B(n43131), .A(n43130), .Z(n46340) );
  XOR U45838 ( .A(n46342), .B(n46343), .Z(n43130) );
  XOR U45839 ( .A(n46344), .B(n44604), .Z(n43131) );
  IV U45840 ( .A(n42210), .Z(n44604) );
  XOR U45841 ( .A(n42444), .B(n46345), .Z(n46313) );
  XNOR U45842 ( .A(n39762), .B(n37505), .Z(n46345) );
  XOR U45843 ( .A(n46346), .B(n42130), .Z(n37505) );
  XOR U45844 ( .A(n46347), .B(n42309), .Z(n42130) );
  AND U45845 ( .A(n43135), .B(n43134), .Z(n46346) );
  XOR U45846 ( .A(n46350), .B(n45629), .Z(n43134) );
  XOR U45847 ( .A(n46351), .B(n45339), .Z(n43135) );
  XNOR U45848 ( .A(n46352), .B(n43754), .Z(n39762) );
  XOR U45849 ( .A(n46353), .B(n45425), .Z(n43754) );
  IV U45850 ( .A(n44774), .Z(n45425) );
  AND U45851 ( .A(n43122), .B(n43123), .Z(n46352) );
  XNOR U45852 ( .A(n46354), .B(n43767), .Z(n43123) );
  XOR U45853 ( .A(n46355), .B(n44550), .Z(n43122) );
  XOR U45854 ( .A(n46356), .B(n43752), .Z(n42444) );
  XOR U45855 ( .A(n46357), .B(n45371), .Z(n43752) );
  ANDN U45856 ( .B(n43120), .A(n43118), .Z(n46356) );
  XOR U45857 ( .A(n46358), .B(n42498), .Z(n43118) );
  XOR U45858 ( .A(n43311), .B(n46359), .Z(n43120) );
  XNOR U45859 ( .A(n46360), .B(n43734), .Z(n42249) );
  IV U45860 ( .A(n46304), .Z(n43734) );
  XOR U45861 ( .A(n46361), .B(n43680), .Z(n46304) );
  ANDN U45862 ( .B(n46305), .A(n45532), .Z(n46360) );
  XNOR U45863 ( .A(n32599), .B(n46362), .Z(n45994) );
  XOR U45864 ( .A(n35399), .B(n31640), .Z(n46362) );
  XNOR U45865 ( .A(n46363), .B(n35431), .Z(n31640) );
  XOR U45866 ( .A(n45536), .B(n37011), .Z(n35431) );
  XOR U45867 ( .A(n44786), .B(n40434), .Z(n37011) );
  XNOR U45868 ( .A(n46364), .B(n46365), .Z(n40434) );
  XNOR U45869 ( .A(n38930), .B(n38557), .Z(n46365) );
  XNOR U45870 ( .A(n46366), .B(n39730), .Z(n38557) );
  IV U45871 ( .A(n46367), .Z(n39730) );
  ANDN U45872 ( .B(n39731), .A(n45546), .Z(n46366) );
  XOR U45873 ( .A(n46368), .B(n40849), .Z(n39731) );
  IV U45874 ( .A(n43457), .Z(n40849) );
  XOR U45875 ( .A(n46369), .B(n39720), .Z(n38930) );
  XOR U45876 ( .A(n46370), .B(n44218), .Z(n39721) );
  IV U45877 ( .A(n44593), .Z(n44218) );
  XNOR U45878 ( .A(n46348), .B(n46371), .Z(n44593) );
  XNOR U45879 ( .A(n46372), .B(n46373), .Z(n46348) );
  XOR U45880 ( .A(n45447), .B(n46013), .Z(n46373) );
  XOR U45881 ( .A(n46374), .B(n46375), .Z(n46013) );
  NOR U45882 ( .A(n46376), .B(n46377), .Z(n46374) );
  XNOR U45883 ( .A(n46378), .B(n46379), .Z(n45447) );
  ANDN U45884 ( .B(n46380), .A(n46381), .Z(n46378) );
  XOR U45885 ( .A(n46382), .B(n46383), .Z(n46372) );
  XOR U45886 ( .A(n45653), .B(n46384), .Z(n46383) );
  XNOR U45887 ( .A(n46385), .B(n46386), .Z(n45653) );
  ANDN U45888 ( .B(n46387), .A(n46388), .Z(n46385) );
  XNOR U45889 ( .A(n38647), .B(n46389), .Z(n46364) );
  XOR U45890 ( .A(n37205), .B(n39710), .Z(n46389) );
  XOR U45891 ( .A(n46390), .B(n39727), .Z(n39710) );
  ANDN U45892 ( .B(n39726), .A(n45538), .Z(n46390) );
  XOR U45893 ( .A(n46391), .B(n44862), .Z(n39726) );
  XOR U45894 ( .A(n46392), .B(n46393), .Z(n37205) );
  ANDN U45895 ( .B(n45544), .A(n39716), .Z(n46392) );
  IV U45896 ( .A(n45542), .Z(n39716) );
  XOR U45897 ( .A(n46394), .B(n42223), .Z(n45542) );
  IV U45898 ( .A(n46395), .Z(n45544) );
  XNOR U45899 ( .A(n46396), .B(n40645), .Z(n38647) );
  XOR U45900 ( .A(n46398), .B(n46399), .Z(n44786) );
  XNOR U45901 ( .A(n39403), .B(n41139), .Z(n46399) );
  XNOR U45902 ( .A(n46400), .B(n46312), .Z(n41139) );
  XOR U45903 ( .A(n46401), .B(n43550), .Z(n46312) );
  ANDN U45904 ( .B(n42253), .A(n43736), .Z(n46400) );
  XOR U45905 ( .A(n44874), .B(n46402), .Z(n43736) );
  IV U45906 ( .A(n46403), .Z(n44874) );
  XOR U45907 ( .A(n46404), .B(n46405), .Z(n42253) );
  XOR U45908 ( .A(n46406), .B(n42242), .Z(n39403) );
  XOR U45909 ( .A(n46407), .B(n42419), .Z(n42242) );
  NOR U45910 ( .A(n43743), .B(n42241), .Z(n46406) );
  XOR U45911 ( .A(n46410), .B(n42153), .Z(n42241) );
  IV U45912 ( .A(n46107), .Z(n42153) );
  XOR U45913 ( .A(n46411), .B(n46412), .Z(n46107) );
  XNOR U45914 ( .A(n46413), .B(n46414), .Z(n43743) );
  XNOR U45915 ( .A(n39268), .B(n46415), .Z(n46398) );
  XOR U45916 ( .A(n40272), .B(n42235), .Z(n46415) );
  XOR U45917 ( .A(n46416), .B(n43519), .Z(n42235) );
  XOR U45918 ( .A(n46417), .B(n45127), .Z(n43519) );
  ANDN U45919 ( .B(n43740), .A(n43518), .Z(n46416) );
  XOR U45920 ( .A(n46418), .B(n45443), .Z(n43518) );
  XOR U45921 ( .A(n45504), .B(n46419), .Z(n43740) );
  XNOR U45922 ( .A(n46420), .B(n42245), .Z(n40272) );
  XOR U45923 ( .A(n46421), .B(n46422), .Z(n42245) );
  ANDN U45924 ( .B(n42246), .A(n43746), .Z(n46420) );
  XOR U45925 ( .A(n46423), .B(n41731), .Z(n43746) );
  XOR U45926 ( .A(n46424), .B(n45358), .Z(n42246) );
  XOR U45927 ( .A(n46425), .B(n46305), .Z(n39268) );
  XNOR U45928 ( .A(n46426), .B(n44469), .Z(n46305) );
  XOR U45929 ( .A(n46429), .B(n42503), .Z(n43732) );
  XOR U45930 ( .A(n46430), .B(n44467), .Z(n45532) );
  XNOR U45931 ( .A(n46431), .B(n40644), .Z(n45536) );
  XNOR U45932 ( .A(n46432), .B(n42877), .Z(n40644) );
  XNOR U45933 ( .A(n46433), .B(n46434), .Z(n42877) );
  AND U45934 ( .A(n46435), .B(n46397), .Z(n46431) );
  XOR U45935 ( .A(n41701), .B(n38446), .Z(n35432) );
  IV U45936 ( .A(n37640), .Z(n38446) );
  XNOR U45937 ( .A(n40730), .B(n40640), .Z(n37640) );
  XNOR U45938 ( .A(n46436), .B(n46437), .Z(n40640) );
  XOR U45939 ( .A(n39459), .B(n35631), .Z(n46437) );
  XNOR U45940 ( .A(n46438), .B(n45539), .Z(n35631) );
  IV U45941 ( .A(n46439), .Z(n45539) );
  ANDN U45942 ( .B(n39725), .A(n39727), .Z(n46438) );
  XOR U45943 ( .A(n46440), .B(n43524), .Z(n39727) );
  IV U45944 ( .A(n46183), .Z(n43524) );
  XOR U45945 ( .A(n46441), .B(n45550), .Z(n39459) );
  ANDN U45946 ( .B(n39719), .A(n39720), .Z(n46441) );
  XOR U45947 ( .A(n46442), .B(n46443), .Z(n39720) );
  XNOR U45948 ( .A(n36432), .B(n46444), .Z(n46436) );
  XOR U45949 ( .A(n40372), .B(n39152), .Z(n46444) );
  XNOR U45950 ( .A(n46445), .B(n45547), .Z(n39152) );
  ANDN U45951 ( .B(n39729), .A(n46367), .Z(n46445) );
  XOR U45952 ( .A(n46446), .B(n46447), .Z(n46367) );
  XOR U45953 ( .A(n46448), .B(n45543), .Z(n40372) );
  ANDN U45954 ( .B(n39715), .A(n46393), .Z(n46448) );
  IV U45955 ( .A(n39717), .Z(n46393) );
  XOR U45956 ( .A(n46449), .B(n43335), .Z(n39717) );
  IV U45957 ( .A(n45268), .Z(n43335) );
  XNOR U45958 ( .A(n46450), .B(n46451), .Z(n45268) );
  XNOR U45959 ( .A(n46452), .B(n46435), .Z(n36432) );
  XOR U45960 ( .A(n46453), .B(n45260), .Z(n40645) );
  XOR U45961 ( .A(n46454), .B(n46455), .Z(n40730) );
  XOR U45962 ( .A(n38910), .B(n46456), .Z(n46455) );
  XNOR U45963 ( .A(n46457), .B(n43465), .Z(n38910) );
  IV U45964 ( .A(n46458), .Z(n43465) );
  ANDN U45965 ( .B(n41707), .A(n42890), .Z(n46457) );
  IV U45966 ( .A(n41708), .Z(n42890) );
  XOR U45967 ( .A(n46181), .B(n46459), .Z(n41708) );
  XNOR U45968 ( .A(n37622), .B(n46460), .Z(n46454) );
  XOR U45969 ( .A(n38495), .B(n36315), .Z(n46460) );
  XNOR U45970 ( .A(n46461), .B(n43458), .Z(n36315) );
  ANDN U45971 ( .B(n41697), .A(n41698), .Z(n46461) );
  XOR U45972 ( .A(n46462), .B(n45734), .Z(n41698) );
  XOR U45973 ( .A(n46463), .B(n43469), .Z(n38495) );
  ANDN U45974 ( .B(n41693), .A(n42898), .Z(n46463) );
  IV U45975 ( .A(n41695), .Z(n42898) );
  XOR U45976 ( .A(n46464), .B(n44797), .Z(n41695) );
  XNOR U45977 ( .A(n46465), .B(n43460), .Z(n37622) );
  AND U45978 ( .A(n42893), .B(n46466), .Z(n46465) );
  XNOR U45979 ( .A(n46467), .B(n46466), .Z(n41701) );
  NOR U45980 ( .A(n42893), .B(n42894), .Z(n46467) );
  XNOR U45981 ( .A(n45151), .B(n46468), .Z(n42894) );
  XNOR U45982 ( .A(n46469), .B(n44178), .Z(n42893) );
  IV U45983 ( .A(n42496), .Z(n44178) );
  XOR U45984 ( .A(n46470), .B(n46371), .Z(n42496) );
  XNOR U45985 ( .A(n46471), .B(n46472), .Z(n46371) );
  XNOR U45986 ( .A(n46473), .B(n45925), .Z(n46472) );
  XNOR U45987 ( .A(n46474), .B(n46475), .Z(n45925) );
  XOR U45988 ( .A(n43074), .B(n46478), .Z(n46471) );
  XOR U45989 ( .A(n43584), .B(n44843), .Z(n46478) );
  XNOR U45990 ( .A(n46479), .B(n46480), .Z(n44843) );
  NOR U45991 ( .A(n46481), .B(n46482), .Z(n46479) );
  XNOR U45992 ( .A(n46483), .B(n46484), .Z(n43584) );
  XNOR U45993 ( .A(n46487), .B(n46488), .Z(n43074) );
  XOR U45994 ( .A(n38181), .B(n45606), .Z(n34208) );
  XNOR U45995 ( .A(n46491), .B(n43803), .Z(n45606) );
  NOR U45996 ( .A(n42630), .B(n42631), .Z(n46491) );
  XOR U45997 ( .A(n46492), .B(n43671), .Z(n42631) );
  XNOR U45998 ( .A(n40352), .B(n39842), .Z(n38181) );
  XNOR U45999 ( .A(n46493), .B(n46494), .Z(n39842) );
  XOR U46000 ( .A(n43789), .B(n36211), .Z(n46494) );
  XOR U46001 ( .A(n46495), .B(n43799), .Z(n36211) );
  XOR U46002 ( .A(n46496), .B(n44014), .Z(n43799) );
  XOR U46003 ( .A(n46497), .B(n46498), .Z(n44014) );
  ANDN U46004 ( .B(n42626), .A(n43798), .Z(n46495) );
  XOR U46005 ( .A(n46499), .B(n44809), .Z(n43798) );
  IV U46006 ( .A(n45244), .Z(n44809) );
  XOR U46007 ( .A(n46500), .B(n46501), .Z(n42626) );
  XNOR U46008 ( .A(n46502), .B(n43809), .Z(n43789) );
  XOR U46009 ( .A(n46503), .B(n45902), .Z(n43809) );
  AND U46010 ( .A(n45611), .B(n43810), .Z(n46502) );
  XOR U46011 ( .A(n46504), .B(n44762), .Z(n43810) );
  XOR U46012 ( .A(n46505), .B(n46506), .Z(n45611) );
  XNOR U46013 ( .A(n37708), .B(n46507), .Z(n46493) );
  XNOR U46014 ( .A(n40509), .B(n39375), .Z(n46507) );
  XOR U46015 ( .A(n46508), .B(n46205), .Z(n39375) );
  XOR U46016 ( .A(n46509), .B(n46510), .Z(n46205) );
  ANDN U46017 ( .B(n42620), .A(n43805), .Z(n46508) );
  XOR U46018 ( .A(n46511), .B(n46512), .Z(n43805) );
  XNOR U46019 ( .A(n46514), .B(n43802), .Z(n40509) );
  XNOR U46020 ( .A(n44680), .B(n46515), .Z(n43802) );
  XNOR U46021 ( .A(n46516), .B(n46517), .Z(n44680) );
  AND U46022 ( .A(n42630), .B(n43803), .Z(n46514) );
  XOR U46023 ( .A(n45828), .B(n46518), .Z(n43803) );
  XOR U46024 ( .A(n46519), .B(n44747), .Z(n42630) );
  XNOR U46025 ( .A(n46520), .B(n43795), .Z(n37708) );
  XOR U46026 ( .A(n46521), .B(n45491), .Z(n43795) );
  IV U46027 ( .A(n44935), .Z(n45491) );
  ANDN U46028 ( .B(n42616), .A(n43794), .Z(n46520) );
  XNOR U46029 ( .A(n46522), .B(n43819), .Z(n43794) );
  XNOR U46030 ( .A(n42504), .B(n46523), .Z(n42616) );
  XOR U46031 ( .A(n46524), .B(n46525), .Z(n40352) );
  XNOR U46032 ( .A(n37680), .B(n39332), .Z(n46525) );
  XNOR U46033 ( .A(n46526), .B(n40701), .Z(n39332) );
  XOR U46034 ( .A(n46527), .B(n46528), .Z(n40701) );
  AND U46035 ( .A(n42639), .B(n44875), .Z(n46526) );
  XNOR U46036 ( .A(n46529), .B(n43565), .Z(n44875) );
  XOR U46037 ( .A(n46530), .B(n44747), .Z(n42639) );
  IV U46038 ( .A(n45403), .Z(n44747) );
  XNOR U46039 ( .A(n46533), .B(n40114), .Z(n37680) );
  XOR U46040 ( .A(n46534), .B(n43895), .Z(n40114) );
  XOR U46041 ( .A(n46535), .B(n46536), .Z(n43895) );
  ANDN U46042 ( .B(n44871), .A(n42643), .Z(n46533) );
  IV U46043 ( .A(n45599), .Z(n42643) );
  XNOR U46044 ( .A(n46537), .B(n43920), .Z(n45599) );
  XOR U46045 ( .A(n46538), .B(n43102), .Z(n44871) );
  XNOR U46046 ( .A(n44832), .B(n46539), .Z(n46524) );
  XOR U46047 ( .A(n39788), .B(n40822), .Z(n46539) );
  XOR U46048 ( .A(n46540), .B(n40104), .Z(n40822) );
  XNOR U46049 ( .A(n44767), .B(n46541), .Z(n40104) );
  NOR U46050 ( .A(n42636), .B(n44879), .Z(n46540) );
  XNOR U46051 ( .A(n46542), .B(n45443), .Z(n44879) );
  XOR U46052 ( .A(n43819), .B(n46545), .Z(n42636) );
  XOR U46053 ( .A(n46546), .B(n40118), .Z(n39788) );
  XOR U46054 ( .A(n46547), .B(n42306), .Z(n40118) );
  NOR U46055 ( .A(n45595), .B(n43787), .Z(n46546) );
  XNOR U46056 ( .A(n46548), .B(n44492), .Z(n43787) );
  XOR U46057 ( .A(n45159), .B(n46549), .Z(n45595) );
  XOR U46058 ( .A(n46550), .B(n46551), .Z(n45159) );
  XNOR U46059 ( .A(n46552), .B(n40107), .Z(n44832) );
  ANDN U46060 ( .B(n42645), .A(n44883), .Z(n46552) );
  IV U46061 ( .A(n45590), .Z(n44883) );
  XOR U46062 ( .A(n46554), .B(n42219), .Z(n45590) );
  XNOR U46063 ( .A(n42546), .B(n46555), .Z(n42645) );
  IV U46064 ( .A(n44686), .Z(n42546) );
  XNOR U46065 ( .A(n46556), .B(n39590), .Z(n35399) );
  XOR U46066 ( .A(n45029), .B(n39219), .Z(n39590) );
  XNOR U46067 ( .A(n46557), .B(n44443), .Z(n45029) );
  NOR U46068 ( .A(n46558), .B(n44720), .Z(n46557) );
  AND U46069 ( .A(n35640), .B(n34195), .Z(n46556) );
  XOR U46070 ( .A(n41830), .B(n38486), .Z(n34195) );
  XNOR U46071 ( .A(n46559), .B(n46560), .Z(n42693) );
  XNOR U46072 ( .A(n42823), .B(n39089), .Z(n46560) );
  XNOR U46073 ( .A(n46561), .B(n42810), .Z(n39089) );
  XOR U46074 ( .A(n46562), .B(n42340), .Z(n42810) );
  AND U46075 ( .A(n43532), .B(n43653), .Z(n46561) );
  XNOR U46076 ( .A(n46563), .B(n42017), .Z(n42823) );
  XOR U46077 ( .A(n46564), .B(n43540), .Z(n42017) );
  AND U46078 ( .A(n41832), .B(n41834), .Z(n46563) );
  XOR U46079 ( .A(n45697), .B(n46565), .Z(n41834) );
  XNOR U46080 ( .A(n46566), .B(n43552), .Z(n41832) );
  XOR U46081 ( .A(n41117), .B(n46567), .Z(n46559) );
  XOR U46082 ( .A(n40141), .B(n35324), .Z(n46567) );
  XNOR U46083 ( .A(n46568), .B(n43566), .Z(n35324) );
  XOR U46084 ( .A(n46569), .B(n42157), .Z(n43566) );
  ANDN U46085 ( .B(n41826), .A(n41827), .Z(n46568) );
  XOR U46086 ( .A(n46570), .B(n43662), .Z(n41827) );
  IV U46087 ( .A(n46571), .Z(n43662) );
  XNOR U46088 ( .A(n46572), .B(n46573), .Z(n41826) );
  XNOR U46089 ( .A(n46574), .B(n42026), .Z(n40141) );
  XNOR U46090 ( .A(n46575), .B(n42672), .Z(n42026) );
  XOR U46091 ( .A(n46576), .B(n45664), .Z(n41822) );
  XOR U46092 ( .A(n46577), .B(n42450), .Z(n41824) );
  IV U46093 ( .A(n45588), .Z(n42450) );
  XOR U46094 ( .A(n46578), .B(n46579), .Z(n45588) );
  XNOR U46095 ( .A(n46580), .B(n42020), .Z(n41117) );
  XNOR U46096 ( .A(n43577), .B(n46581), .Z(n42020) );
  AND U46097 ( .A(n41836), .B(n41838), .Z(n46580) );
  XOR U46098 ( .A(n43330), .B(n46582), .Z(n41838) );
  XOR U46099 ( .A(n46583), .B(n46584), .Z(n43330) );
  XNOR U46100 ( .A(n46585), .B(n43329), .Z(n41836) );
  XOR U46101 ( .A(n46586), .B(n46587), .Z(n42886) );
  XNOR U46102 ( .A(n38490), .B(n38832), .Z(n46587) );
  XOR U46103 ( .A(n46588), .B(n40739), .Z(n38832) );
  ANDN U46104 ( .B(n41818), .A(n42828), .Z(n46588) );
  IV U46105 ( .A(n41817), .Z(n42828) );
  XOR U46106 ( .A(n46166), .B(n46590), .Z(n41817) );
  XNOR U46107 ( .A(n46591), .B(n42219), .Z(n41818) );
  XNOR U46108 ( .A(n46592), .B(n40753), .Z(n38490) );
  XNOR U46109 ( .A(n42517), .B(n46593), .Z(n40753) );
  IV U46110 ( .A(n46207), .Z(n42517) );
  XOR U46111 ( .A(n46594), .B(n46595), .Z(n46207) );
  XOR U46112 ( .A(n46596), .B(n44856), .Z(n41811) );
  XOR U46113 ( .A(n46021), .B(n46597), .Z(n41812) );
  XOR U46114 ( .A(n39073), .B(n46598), .Z(n46586) );
  XOR U46115 ( .A(n37514), .B(n41688), .Z(n46598) );
  XOR U46116 ( .A(n46599), .B(n40736), .Z(n41688) );
  XOR U46117 ( .A(n46600), .B(n46601), .Z(n40736) );
  AND U46118 ( .A(n42885), .B(n42832), .Z(n46599) );
  XNOR U46119 ( .A(n46056), .B(n46602), .Z(n42832) );
  IV U46120 ( .A(n44316), .Z(n46056) );
  XNOR U46121 ( .A(n46470), .B(n46603), .Z(n44316) );
  XOR U46122 ( .A(n46604), .B(n46605), .Z(n46470) );
  XOR U46123 ( .A(n44771), .B(n44214), .Z(n46605) );
  XOR U46124 ( .A(n46606), .B(n46607), .Z(n44214) );
  NOR U46125 ( .A(n46608), .B(n46609), .Z(n46606) );
  XNOR U46126 ( .A(n46610), .B(n46611), .Z(n44771) );
  XOR U46127 ( .A(n44901), .B(n46614), .Z(n46604) );
  XNOR U46128 ( .A(n44493), .B(n46615), .Z(n46614) );
  XOR U46129 ( .A(n46616), .B(n46617), .Z(n44493) );
  ANDN U46130 ( .B(n46618), .A(n46619), .Z(n46616) );
  XNOR U46131 ( .A(n46620), .B(n46621), .Z(n44901) );
  XOR U46132 ( .A(n44783), .B(n46624), .Z(n42885) );
  XOR U46133 ( .A(n46625), .B(n40745), .Z(n37514) );
  IV U46134 ( .A(n42834), .Z(n40745) );
  XNOR U46135 ( .A(n46626), .B(n42340), .Z(n42834) );
  XOR U46136 ( .A(n45716), .B(n46627), .Z(n42340) );
  XOR U46137 ( .A(n46628), .B(n46629), .Z(n45716) );
  XNOR U46138 ( .A(n46630), .B(n46631), .Z(n46629) );
  XOR U46139 ( .A(n46632), .B(n46633), .Z(n46628) );
  XOR U46140 ( .A(n46634), .B(n46635), .Z(n46633) );
  AND U46141 ( .A(n41814), .B(n41815), .Z(n46625) );
  XNOR U46142 ( .A(n46636), .B(n42160), .Z(n41815) );
  XOR U46143 ( .A(n46637), .B(n46638), .Z(n41814) );
  XOR U46144 ( .A(n46639), .B(n40748), .Z(n39073) );
  XNOR U46145 ( .A(n46640), .B(n44333), .Z(n40748) );
  IV U46146 ( .A(n44528), .Z(n44333) );
  ANDN U46147 ( .B(n41808), .A(n41807), .Z(n46639) );
  IV U46148 ( .A(n42836), .Z(n41807) );
  XOR U46149 ( .A(n44850), .B(n46642), .Z(n41808) );
  XNOR U46150 ( .A(n46643), .B(n43653), .Z(n41830) );
  XOR U46151 ( .A(n46644), .B(n45308), .Z(n43653) );
  NOR U46152 ( .A(n42808), .B(n43532), .Z(n46643) );
  XOR U46153 ( .A(n43598), .B(n46645), .Z(n43532) );
  XOR U46154 ( .A(n46646), .B(n44106), .Z(n42808) );
  XOR U46155 ( .A(n41043), .B(n36537), .Z(n35640) );
  XOR U46156 ( .A(n42012), .B(n40442), .Z(n36537) );
  XNOR U46157 ( .A(n46647), .B(n46648), .Z(n40442) );
  XOR U46158 ( .A(n45168), .B(n42464), .Z(n46648) );
  XNOR U46159 ( .A(n46649), .B(n45190), .Z(n42464) );
  IV U46160 ( .A(n41958), .Z(n45190) );
  XOR U46161 ( .A(n46650), .B(n45858), .Z(n41958) );
  NOR U46162 ( .A(n45189), .B(n41059), .Z(n46649) );
  IV U46163 ( .A(n41058), .Z(n45189) );
  XOR U46164 ( .A(n45828), .B(n46651), .Z(n41058) );
  XNOR U46165 ( .A(n46652), .B(n42229), .Z(n45168) );
  XNOR U46166 ( .A(n46653), .B(n42223), .Z(n42229) );
  ANDN U46167 ( .B(n41056), .A(n45187), .Z(n46652) );
  XOR U46168 ( .A(n46654), .B(n44195), .Z(n45187) );
  XOR U46169 ( .A(n37676), .B(n46655), .Z(n46647) );
  XOR U46170 ( .A(n39819), .B(n35928), .Z(n46655) );
  XNOR U46171 ( .A(n46656), .B(n41955), .Z(n35928) );
  XOR U46172 ( .A(n46657), .B(n44032), .Z(n41955) );
  ANDN U46173 ( .B(n41045), .A(n41046), .Z(n46656) );
  XNOR U46174 ( .A(n45386), .B(n46658), .Z(n41045) );
  XOR U46175 ( .A(n46659), .B(n42007), .Z(n39819) );
  XOR U46176 ( .A(n46660), .B(n44579), .Z(n42007) );
  AND U46177 ( .A(n41052), .B(n41050), .Z(n46659) );
  XOR U46178 ( .A(n46661), .B(n46405), .Z(n41050) );
  XNOR U46179 ( .A(n46662), .B(n41949), .Z(n37676) );
  XOR U46180 ( .A(n46663), .B(n44969), .Z(n41949) );
  IV U46181 ( .A(n43967), .Z(n44969) );
  ANDN U46182 ( .B(n45194), .A(n46664), .Z(n46662) );
  XOR U46183 ( .A(n46665), .B(n46666), .Z(n42012) );
  XNOR U46184 ( .A(n37509), .B(n39006), .Z(n46666) );
  XOR U46185 ( .A(n46667), .B(n42709), .Z(n39006) );
  XNOR U46186 ( .A(n42329), .B(n46668), .Z(n42709) );
  XOR U46187 ( .A(n46669), .B(n44119), .Z(n42705) );
  XOR U46188 ( .A(n46510), .B(n46670), .Z(n43660) );
  IV U46189 ( .A(n43311), .Z(n46510) );
  XNOR U46190 ( .A(n46671), .B(n46672), .Z(n43311) );
  XOR U46191 ( .A(n46673), .B(n41855), .Z(n37509) );
  XOR U46192 ( .A(n46674), .B(n45203), .Z(n41855) );
  ANDN U46193 ( .B(n42699), .A(n45183), .Z(n46673) );
  XOR U46194 ( .A(n46675), .B(n46676), .Z(n45183) );
  XNOR U46195 ( .A(n46677), .B(n42306), .Z(n42699) );
  XOR U46196 ( .A(n46678), .B(n46679), .Z(n42306) );
  XOR U46197 ( .A(n42053), .B(n46680), .Z(n46665) );
  XNOR U46198 ( .A(n40342), .B(n38842), .Z(n46680) );
  XNOR U46199 ( .A(n46681), .B(n41851), .Z(n38842) );
  XOR U46200 ( .A(n46682), .B(n43594), .Z(n41851) );
  XNOR U46201 ( .A(n46683), .B(n46684), .Z(n43594) );
  ANDN U46202 ( .B(n43676), .A(n42703), .Z(n46681) );
  XOR U46203 ( .A(n46382), .B(n46014), .Z(n42703) );
  XNOR U46204 ( .A(n46685), .B(n46686), .Z(n46382) );
  NOR U46205 ( .A(n46687), .B(n46688), .Z(n46685) );
  XOR U46206 ( .A(n42508), .B(n46689), .Z(n43676) );
  IV U46207 ( .A(n45148), .Z(n42508) );
  XNOR U46208 ( .A(n46690), .B(n46691), .Z(n45148) );
  XOR U46209 ( .A(n46692), .B(n42468), .Z(n40342) );
  XOR U46210 ( .A(n46693), .B(n42672), .Z(n42468) );
  XOR U46211 ( .A(n46694), .B(n46695), .Z(n42672) );
  ANDN U46212 ( .B(n43673), .A(n43674), .Z(n46692) );
  XNOR U46213 ( .A(n42667), .B(n46696), .Z(n43674) );
  XNOR U46214 ( .A(n45386), .B(n46697), .Z(n43673) );
  XNOR U46215 ( .A(n46698), .B(n46699), .Z(n45386) );
  XNOR U46216 ( .A(n46700), .B(n41859), .Z(n42053) );
  XOR U46217 ( .A(n46701), .B(n46702), .Z(n41859) );
  NOR U46218 ( .A(n43669), .B(n42697), .Z(n46700) );
  XNOR U46219 ( .A(n46703), .B(n45554), .Z(n42697) );
  XOR U46220 ( .A(n46704), .B(n42402), .Z(n43669) );
  IV U46221 ( .A(n44193), .Z(n42402) );
  XOR U46222 ( .A(n46705), .B(n46706), .Z(n44193) );
  XNOR U46223 ( .A(n46707), .B(n45194), .Z(n41043) );
  XNOR U46224 ( .A(n46708), .B(n45121), .Z(n45194) );
  ANDN U46225 ( .B(n46664), .A(n41948), .Z(n46707) );
  XOR U46226 ( .A(n46709), .B(n35434), .Z(n32599) );
  XOR U46227 ( .A(n43187), .B(n37630), .Z(n35434) );
  XOR U46228 ( .A(n43625), .B(n39418), .Z(n37630) );
  XNOR U46229 ( .A(n46710), .B(n46711), .Z(n39418) );
  XOR U46230 ( .A(n41418), .B(n38317), .Z(n46711) );
  XOR U46231 ( .A(n46712), .B(n41780), .Z(n38317) );
  XOR U46232 ( .A(n46713), .B(n46032), .Z(n41780) );
  NOR U46233 ( .A(n42038), .B(n42874), .Z(n46712) );
  XNOR U46234 ( .A(n46714), .B(n45397), .Z(n42874) );
  XOR U46235 ( .A(n46715), .B(n46601), .Z(n42038) );
  XNOR U46236 ( .A(n46716), .B(n42879), .Z(n41418) );
  XOR U46237 ( .A(n46717), .B(n46158), .Z(n42879) );
  NOR U46238 ( .A(n42040), .B(n42878), .Z(n46716) );
  XOR U46239 ( .A(n45504), .B(n46718), .Z(n42878) );
  XNOR U46240 ( .A(n44472), .B(n46719), .Z(n42040) );
  XOR U46241 ( .A(n38876), .B(n46720), .Z(n46710) );
  XOR U46242 ( .A(n38157), .B(n42838), .Z(n46720) );
  XNOR U46243 ( .A(n46721), .B(n41764), .Z(n42838) );
  XNOR U46244 ( .A(n46722), .B(n45339), .Z(n41764) );
  NOR U46245 ( .A(n42033), .B(n42883), .Z(n46721) );
  XOR U46246 ( .A(n46723), .B(n43644), .Z(n42883) );
  XOR U46247 ( .A(n46724), .B(n45982), .Z(n42033) );
  IV U46248 ( .A(n42550), .Z(n45982) );
  XNOR U46249 ( .A(n46725), .B(n46726), .Z(n42550) );
  XNOR U46250 ( .A(n46727), .B(n41768), .Z(n38157) );
  XOR U46251 ( .A(n43463), .B(n46728), .Z(n41768) );
  XOR U46252 ( .A(n45583), .B(n46729), .Z(n45552) );
  XOR U46253 ( .A(n46730), .B(n45203), .Z(n42865) );
  XNOR U46254 ( .A(n46731), .B(n46732), .Z(n45203) );
  XNOR U46255 ( .A(n46733), .B(n41772), .Z(n38876) );
  XOR U46256 ( .A(n46734), .B(n44759), .Z(n41772) );
  IV U46257 ( .A(n46735), .Z(n44759) );
  NOR U46258 ( .A(n42869), .B(n42036), .Z(n46733) );
  XNOR U46259 ( .A(n46736), .B(n44539), .Z(n42036) );
  IV U46260 ( .A(n44673), .Z(n44539) );
  XOR U46261 ( .A(n46737), .B(n45861), .Z(n42869) );
  XOR U46262 ( .A(n46738), .B(n46739), .Z(n43625) );
  XOR U46263 ( .A(n40003), .B(n38441), .Z(n46739) );
  XOR U46264 ( .A(n46740), .B(n41207), .Z(n38441) );
  XNOR U46265 ( .A(n46741), .B(n46032), .Z(n41207) );
  ANDN U46266 ( .B(n43194), .A(n43193), .Z(n46740) );
  XNOR U46267 ( .A(n46742), .B(n43719), .Z(n43193) );
  XNOR U46268 ( .A(n46743), .B(n41197), .Z(n40003) );
  XNOR U46269 ( .A(n46744), .B(n46745), .Z(n41197) );
  NOR U46270 ( .A(n43198), .B(n41965), .Z(n46743) );
  XOR U46271 ( .A(n46746), .B(n45123), .Z(n41965) );
  XOR U46272 ( .A(n35633), .B(n46747), .Z(n46738) );
  XOR U46273 ( .A(n40347), .B(n39546), .Z(n46747) );
  XNOR U46274 ( .A(n46748), .B(n41973), .Z(n39546) );
  XOR U46275 ( .A(n44675), .B(n46749), .Z(n41973) );
  ANDN U46276 ( .B(n43190), .A(n43189), .Z(n46748) );
  XOR U46277 ( .A(n43600), .B(n46750), .Z(n43189) );
  XOR U46278 ( .A(n42881), .B(n46752), .Z(n41192) );
  XNOR U46279 ( .A(n46753), .B(n46754), .Z(n42881) );
  NOR U46280 ( .A(n46755), .B(n41977), .Z(n46751) );
  XOR U46281 ( .A(n46756), .B(n45569), .Z(n41977) );
  IV U46282 ( .A(n43196), .Z(n46755) );
  XNOR U46283 ( .A(n46757), .B(n41202), .Z(n35633) );
  XNOR U46284 ( .A(n46631), .B(n46758), .Z(n41202) );
  XNOR U46285 ( .A(n46759), .B(n45875), .Z(n46631) );
  ANDN U46286 ( .B(n46760), .A(n46761), .Z(n46759) );
  ANDN U46287 ( .B(n46762), .A(n46763), .Z(n46757) );
  XNOR U46288 ( .A(n46764), .B(n41967), .Z(n43187) );
  IV U46289 ( .A(n46763), .Z(n41967) );
  XOR U46290 ( .A(n46181), .B(n46765), .Z(n46763) );
  NOR U46291 ( .A(n46762), .B(n41201), .Z(n46764) );
  AND U46292 ( .A(n35435), .B(n34191), .Z(n46709) );
  XNOR U46293 ( .A(n37110), .B(n44754), .Z(n34191) );
  XNOR U46294 ( .A(n46766), .B(n40608), .Z(n44754) );
  ANDN U46295 ( .B(n39195), .A(n39197), .Z(n46766) );
  XOR U46296 ( .A(n46767), .B(n44774), .Z(n39197) );
  XNOR U46297 ( .A(n44791), .B(n43858), .Z(n37110) );
  XNOR U46298 ( .A(n46768), .B(n46769), .Z(n43858) );
  XOR U46299 ( .A(n38785), .B(n37850), .Z(n46769) );
  XOR U46300 ( .A(n46770), .B(n41591), .Z(n37850) );
  XNOR U46301 ( .A(n46771), .B(n43550), .Z(n41591) );
  XNOR U46302 ( .A(n46772), .B(n46269), .Z(n43550) );
  XNOR U46303 ( .A(n46773), .B(n46774), .Z(n46269) );
  XNOR U46304 ( .A(n46114), .B(n46775), .Z(n46774) );
  XNOR U46305 ( .A(n46776), .B(n46777), .Z(n46114) );
  ANDN U46306 ( .B(n46778), .A(n46779), .Z(n46776) );
  XNOR U46307 ( .A(n46780), .B(n46781), .Z(n46773) );
  XOR U46308 ( .A(n45787), .B(n46782), .Z(n46781) );
  XOR U46309 ( .A(n46783), .B(n46784), .Z(n45787) );
  ANDN U46310 ( .B(n46785), .A(n46786), .Z(n46783) );
  NOR U46311 ( .A(n39199), .B(n41600), .Z(n46770) );
  XNOR U46312 ( .A(n46787), .B(n44550), .Z(n41600) );
  IV U46313 ( .A(n44757), .Z(n39199) );
  XOR U46314 ( .A(n43899), .B(n46788), .Z(n44757) );
  XNOR U46315 ( .A(n46789), .B(n40599), .Z(n38785) );
  XNOR U46316 ( .A(n46790), .B(n44921), .Z(n40599) );
  ANDN U46317 ( .B(n44753), .A(n40600), .Z(n46789) );
  XOR U46318 ( .A(n46791), .B(n45669), .Z(n40600) );
  XNOR U46319 ( .A(n45789), .B(n46792), .Z(n44753) );
  IV U46320 ( .A(n41639), .Z(n45789) );
  XOR U46321 ( .A(n46793), .B(n46794), .Z(n41639) );
  XOR U46322 ( .A(n39209), .B(n46795), .Z(n46768) );
  XOR U46323 ( .A(n39234), .B(n35330), .Z(n46795) );
  XNOR U46324 ( .A(n46796), .B(n40612), .Z(n35330) );
  XOR U46325 ( .A(n40856), .B(n46797), .Z(n40612) );
  XNOR U46326 ( .A(n46798), .B(n46799), .Z(n40856) );
  NOR U46327 ( .A(n39206), .B(n40611), .Z(n46796) );
  XOR U46328 ( .A(n46800), .B(n41644), .Z(n40611) );
  IV U46329 ( .A(n45734), .Z(n41644) );
  XNOR U46330 ( .A(n46801), .B(n46120), .Z(n39206) );
  XNOR U46331 ( .A(n46802), .B(n40609), .Z(n39234) );
  XNOR U46332 ( .A(n46803), .B(n44336), .Z(n40609) );
  XNOR U46333 ( .A(n46551), .B(n46804), .Z(n44336) );
  XOR U46334 ( .A(n46805), .B(n46806), .Z(n46551) );
  XOR U46335 ( .A(n44946), .B(n44177), .Z(n46806) );
  XNOR U46336 ( .A(n46807), .B(n46808), .Z(n44177) );
  ANDN U46337 ( .B(n46809), .A(n46810), .Z(n46807) );
  XOR U46338 ( .A(n46811), .B(n46812), .Z(n44946) );
  ANDN U46339 ( .B(n46482), .A(n46813), .Z(n46811) );
  XNOR U46340 ( .A(n45563), .B(n46814), .Z(n46805) );
  XOR U46341 ( .A(n42495), .B(n46469), .Z(n46814) );
  XOR U46342 ( .A(n46815), .B(n46490), .Z(n46469) );
  ANDN U46343 ( .B(n46489), .A(n46816), .Z(n46815) );
  XOR U46344 ( .A(n46817), .B(n46477), .Z(n42495) );
  AND U46345 ( .A(n46818), .B(n46476), .Z(n46817) );
  XOR U46346 ( .A(n46819), .B(n46486), .Z(n45563) );
  ANDN U46347 ( .B(n46485), .A(n46820), .Z(n46819) );
  NOR U46348 ( .A(n39195), .B(n40608), .Z(n46802) );
  XOR U46349 ( .A(n46821), .B(n44943), .Z(n40608) );
  XNOR U46350 ( .A(n46822), .B(n43962), .Z(n39195) );
  IV U46351 ( .A(n41747), .Z(n43962) );
  XNOR U46352 ( .A(n46825), .B(n40603), .Z(n39209) );
  XOR U46353 ( .A(n46826), .B(n46185), .Z(n40603) );
  ANDN U46354 ( .B(n40604), .A(n40635), .Z(n46825) );
  XNOR U46355 ( .A(n43595), .B(n46827), .Z(n40635) );
  IV U46356 ( .A(n44789), .Z(n43595) );
  XNOR U46357 ( .A(n46828), .B(n46829), .Z(n44789) );
  XOR U46358 ( .A(n46830), .B(n43656), .Z(n40604) );
  IV U46359 ( .A(n43833), .Z(n43656) );
  XNOR U46360 ( .A(n46679), .B(n46831), .Z(n43833) );
  XNOR U46361 ( .A(n46832), .B(n46833), .Z(n46679) );
  XOR U46362 ( .A(n46165), .B(n46834), .Z(n46833) );
  XNOR U46363 ( .A(n46835), .B(n46836), .Z(n46165) );
  ANDN U46364 ( .B(n46837), .A(n46838), .Z(n46835) );
  XOR U46365 ( .A(n46839), .B(n46840), .Z(n46832) );
  XNOR U46366 ( .A(n46841), .B(n45890), .Z(n46840) );
  XNOR U46367 ( .A(n46842), .B(n46843), .Z(n45890) );
  ANDN U46368 ( .B(n46844), .A(n46845), .Z(n46842) );
  XOR U46369 ( .A(n46846), .B(n46847), .Z(n44791) );
  XNOR U46370 ( .A(n39371), .B(n40793), .Z(n46847) );
  XNOR U46371 ( .A(n46848), .B(n41564), .Z(n40793) );
  XNOR U46372 ( .A(n46849), .B(n43303), .Z(n41564) );
  XOR U46373 ( .A(n46850), .B(n45864), .Z(n43303) );
  XNOR U46374 ( .A(n46851), .B(n46852), .Z(n45864) );
  XNOR U46375 ( .A(n46565), .B(n45698), .Z(n46852) );
  XNOR U46376 ( .A(n46853), .B(n46854), .Z(n45698) );
  ANDN U46377 ( .B(n46855), .A(n46856), .Z(n46853) );
  XOR U46378 ( .A(n46857), .B(n46858), .Z(n46565) );
  ANDN U46379 ( .B(n46859), .A(n46860), .Z(n46857) );
  XOR U46380 ( .A(n45173), .B(n46861), .Z(n46851) );
  XNOR U46381 ( .A(n45971), .B(n46862), .Z(n46861) );
  XNOR U46382 ( .A(n46863), .B(n46864), .Z(n45971) );
  ANDN U46383 ( .B(n46865), .A(n46866), .Z(n46863) );
  XOR U46384 ( .A(n46867), .B(n46868), .Z(n45173) );
  ANDN U46385 ( .B(n46869), .A(n46870), .Z(n46867) );
  ANDN U46386 ( .B(n41563), .A(n40496), .Z(n46848) );
  XOR U46387 ( .A(n44845), .B(n46871), .Z(n40496) );
  XOR U46388 ( .A(n46872), .B(n46873), .Z(n44845) );
  XNOR U46389 ( .A(n46874), .B(n45260), .Z(n41563) );
  XNOR U46390 ( .A(n46875), .B(n41558), .Z(n39371) );
  XOR U46391 ( .A(n46876), .B(n45121), .Z(n41558) );
  IV U46392 ( .A(n46877), .Z(n45121) );
  ANDN U46393 ( .B(n41559), .A(n40487), .Z(n46875) );
  XNOR U46394 ( .A(n45688), .B(n46878), .Z(n40487) );
  XOR U46395 ( .A(n45583), .B(n46879), .Z(n41559) );
  XNOR U46396 ( .A(n38543), .B(n46880), .Z(n46846) );
  XOR U46397 ( .A(n41550), .B(n39142), .Z(n46880) );
  XNOR U46398 ( .A(n46881), .B(n41567), .Z(n39142) );
  XNOR U46399 ( .A(n46882), .B(n42503), .Z(n41567) );
  IV U46400 ( .A(n45514), .Z(n42503) );
  ANDN U46401 ( .B(n41566), .A(n40504), .Z(n46881) );
  XOR U46402 ( .A(n46885), .B(n42223), .Z(n40504) );
  IV U46403 ( .A(n46886), .Z(n42223) );
  XOR U46404 ( .A(n46887), .B(n44882), .Z(n41566) );
  XNOR U46405 ( .A(n46888), .B(n42150), .Z(n41550) );
  XNOR U46406 ( .A(n46889), .B(n44915), .Z(n42150) );
  ANDN U46407 ( .B(n42167), .A(n40491), .Z(n46888) );
  XNOR U46408 ( .A(n46890), .B(n46735), .Z(n40491) );
  XNOR U46409 ( .A(n46891), .B(n44182), .Z(n42167) );
  XNOR U46410 ( .A(n46892), .B(n46627), .Z(n44182) );
  XNOR U46411 ( .A(n46893), .B(n46894), .Z(n46627) );
  XNOR U46412 ( .A(n42684), .B(n46895), .Z(n46894) );
  XNOR U46413 ( .A(n46896), .B(n46897), .Z(n42684) );
  ANDN U46414 ( .B(n46898), .A(n46899), .Z(n46896) );
  XOR U46415 ( .A(n46900), .B(n46901), .Z(n46893) );
  XOR U46416 ( .A(n46223), .B(n46023), .Z(n46901) );
  XNOR U46417 ( .A(n46902), .B(n46903), .Z(n46023) );
  ANDN U46418 ( .B(n46904), .A(n46905), .Z(n46902) );
  XNOR U46419 ( .A(n46906), .B(n46907), .Z(n46223) );
  ANDN U46420 ( .B(n46908), .A(n46909), .Z(n46906) );
  XOR U46421 ( .A(n46910), .B(n41555), .Z(n38543) );
  XOR U46422 ( .A(n41652), .B(n46911), .Z(n41555) );
  ANDN U46423 ( .B(n41556), .A(n40500), .Z(n46910) );
  XOR U46424 ( .A(n46912), .B(n44232), .Z(n40500) );
  IV U46425 ( .A(n43777), .Z(n44232) );
  XOR U46426 ( .A(n46913), .B(n46914), .Z(n43777) );
  XOR U46427 ( .A(n46915), .B(n41598), .Z(n41556) );
  XOR U46428 ( .A(n40804), .B(n38343), .Z(n35435) );
  IV U46429 ( .A(n39259), .Z(n38343) );
  XNOR U46430 ( .A(n40277), .B(n45766), .Z(n39259) );
  XNOR U46431 ( .A(n46916), .B(n46917), .Z(n45766) );
  XNOR U46432 ( .A(n39853), .B(n41890), .Z(n46917) );
  XOR U46433 ( .A(n46918), .B(n44430), .Z(n41890) );
  XOR U46434 ( .A(n46919), .B(n42210), .Z(n44430) );
  ANDN U46435 ( .B(n40813), .A(n40811), .Z(n46918) );
  XNOR U46436 ( .A(n46922), .B(n44882), .Z(n40811) );
  XOR U46437 ( .A(n43598), .B(n46923), .Z(n40813) );
  XNOR U46438 ( .A(n46924), .B(n42791), .Z(n39853) );
  XOR U46439 ( .A(n46925), .B(n44533), .Z(n42791) );
  ANDN U46440 ( .B(n40819), .A(n40820), .Z(n46924) );
  XOR U46441 ( .A(n46926), .B(n45646), .Z(n40820) );
  XOR U46442 ( .A(n46927), .B(n44220), .Z(n40819) );
  XOR U46443 ( .A(n39348), .B(n46928), .Z(n46916) );
  XNOR U46444 ( .A(n41371), .B(n39112), .Z(n46928) );
  XNOR U46445 ( .A(n46929), .B(n42803), .Z(n39112) );
  XNOR U46446 ( .A(n43774), .B(n46930), .Z(n42803) );
  IV U46447 ( .A(n45228), .Z(n43774) );
  ANDN U46448 ( .B(n40817), .A(n40815), .Z(n46929) );
  XNOR U46449 ( .A(n46931), .B(n46932), .Z(n40815) );
  XOR U46450 ( .A(n46675), .B(n46933), .Z(n40817) );
  XNOR U46451 ( .A(n46934), .B(n42794), .Z(n41371) );
  XNOR U46452 ( .A(n46935), .B(n45006), .Z(n42794) );
  ANDN U46453 ( .B(n40806), .A(n40808), .Z(n46934) );
  XOR U46454 ( .A(n46936), .B(n43647), .Z(n40808) );
  IV U46455 ( .A(n43102), .Z(n43647) );
  XNOR U46456 ( .A(n46937), .B(n45554), .Z(n40806) );
  XNOR U46457 ( .A(n46938), .B(n42800), .Z(n39348) );
  XNOR U46458 ( .A(n46939), .B(n43079), .Z(n42800) );
  IV U46459 ( .A(n46940), .Z(n43079) );
  ANDN U46460 ( .B(n45378), .A(n42799), .Z(n46938) );
  XOR U46461 ( .A(n46941), .B(n46942), .Z(n40277) );
  XNOR U46462 ( .A(n39068), .B(n37691), .Z(n46942) );
  XNOR U46463 ( .A(n46943), .B(n41896), .Z(n37691) );
  XOR U46464 ( .A(n44675), .B(n46944), .Z(n41896) );
  IV U46465 ( .A(n44850), .Z(n44675) );
  XNOR U46466 ( .A(n46945), .B(n46946), .Z(n44850) );
  NOR U46467 ( .A(n42479), .B(n41897), .Z(n46943) );
  XOR U46468 ( .A(n46615), .B(n44215), .Z(n41897) );
  IV U46469 ( .A(n44494), .Z(n44215) );
  XNOR U46470 ( .A(n46947), .B(n46948), .Z(n44494) );
  XNOR U46471 ( .A(n46949), .B(n46950), .Z(n46615) );
  XOR U46472 ( .A(n46953), .B(n44519), .Z(n42479) );
  IV U46473 ( .A(n42501), .Z(n44519) );
  XNOR U46474 ( .A(n46954), .B(n46535), .Z(n42501) );
  XOR U46475 ( .A(n46955), .B(n46956), .Z(n46535) );
  XNOR U46476 ( .A(n44586), .B(n46878), .Z(n46956) );
  XOR U46477 ( .A(n46957), .B(n46958), .Z(n46878) );
  XOR U46478 ( .A(n46961), .B(n46962), .Z(n44586) );
  XOR U46479 ( .A(n45200), .B(n46965), .Z(n46955) );
  XOR U46480 ( .A(n45687), .B(n46966), .Z(n46965) );
  XOR U46481 ( .A(n46967), .B(n46968), .Z(n45687) );
  XOR U46482 ( .A(n46971), .B(n46972), .Z(n45200) );
  NOR U46483 ( .A(n46973), .B(n46974), .Z(n46971) );
  XNOR U46484 ( .A(n46975), .B(n41900), .Z(n39068) );
  XNOR U46485 ( .A(n46976), .B(n46120), .Z(n41900) );
  NOR U46486 ( .A(n41901), .B(n42486), .Z(n46975) );
  XOR U46487 ( .A(n45911), .B(n46977), .Z(n42486) );
  IV U46488 ( .A(n44704), .Z(n45911) );
  XOR U46489 ( .A(n46978), .B(n46824), .Z(n44704) );
  XOR U46490 ( .A(n46979), .B(n46980), .Z(n46824) );
  XOR U46491 ( .A(n44701), .B(n45423), .Z(n46980) );
  XOR U46492 ( .A(n46981), .B(n46982), .Z(n45423) );
  XNOR U46493 ( .A(n46985), .B(n46986), .Z(n44701) );
  ANDN U46494 ( .B(n46987), .A(n46988), .Z(n46985) );
  XOR U46495 ( .A(n46989), .B(n46990), .Z(n46979) );
  XOR U46496 ( .A(n46991), .B(n44008), .Z(n46990) );
  XNOR U46497 ( .A(n46992), .B(n46993), .Z(n44008) );
  NOR U46498 ( .A(n46994), .B(n46995), .Z(n46992) );
  XNOR U46499 ( .A(n45080), .B(n46996), .Z(n41901) );
  XOR U46500 ( .A(n38769), .B(n46997), .Z(n46941) );
  XOR U46501 ( .A(n41751), .B(n37852), .Z(n46997) );
  XNOR U46502 ( .A(n46998), .B(n41906), .Z(n37852) );
  XNOR U46503 ( .A(n44032), .B(n46999), .Z(n41906) );
  NOR U46504 ( .A(n42482), .B(n41905), .Z(n46998) );
  XOR U46505 ( .A(n45697), .B(n46862), .Z(n41905) );
  XNOR U46506 ( .A(n47000), .B(n47001), .Z(n46862) );
  ANDN U46507 ( .B(n47002), .A(n47003), .Z(n47000) );
  IV U46508 ( .A(n45172), .Z(n45697) );
  XOR U46509 ( .A(n46517), .B(n47004), .Z(n45172) );
  XOR U46510 ( .A(n47005), .B(n47006), .Z(n46517) );
  XNOR U46511 ( .A(n44615), .B(n44269), .Z(n47006) );
  XNOR U46512 ( .A(n47007), .B(n47008), .Z(n44269) );
  ANDN U46513 ( .B(n46854), .A(n46855), .Z(n47007) );
  XNOR U46514 ( .A(n47009), .B(n47010), .Z(n44615) );
  ANDN U46515 ( .B(n47001), .A(n47002), .Z(n47009) );
  XOR U46516 ( .A(n44563), .B(n47011), .Z(n47005) );
  XOR U46517 ( .A(n46077), .B(n47012), .Z(n47011) );
  XNOR U46518 ( .A(n47013), .B(n47014), .Z(n46077) );
  NOR U46519 ( .A(n46859), .B(n46858), .Z(n47013) );
  XNOR U46520 ( .A(n47015), .B(n47016), .Z(n44563) );
  NOR U46521 ( .A(n46865), .B(n46864), .Z(n47015) );
  XOR U46522 ( .A(n46042), .B(n44619), .Z(n42482) );
  XNOR U46523 ( .A(n47017), .B(n47018), .Z(n46042) );
  ANDN U46524 ( .B(n47019), .A(n47020), .Z(n47017) );
  XNOR U46525 ( .A(n47021), .B(n41910), .Z(n41751) );
  XOR U46526 ( .A(n47022), .B(n46571), .Z(n41910) );
  NOR U46527 ( .A(n41909), .B(n42475), .Z(n47021) );
  XNOR U46528 ( .A(n47023), .B(n42498), .Z(n42475) );
  XOR U46529 ( .A(n45630), .B(n47024), .Z(n41909) );
  XOR U46530 ( .A(n47025), .B(n41914), .Z(n38769) );
  XOR U46531 ( .A(n47026), .B(n42654), .Z(n41914) );
  NOR U46532 ( .A(n45364), .B(n41913), .Z(n47025) );
  XNOR U46533 ( .A(n47027), .B(n42513), .Z(n41913) );
  IV U46534 ( .A(n42488), .Z(n45364) );
  XNOR U46535 ( .A(n47028), .B(n45006), .Z(n42488) );
  XNOR U46536 ( .A(n47029), .B(n47030), .Z(n45006) );
  XOR U46537 ( .A(n47031), .B(n42799), .Z(n40804) );
  XOR U46538 ( .A(n47032), .B(n47033), .Z(n42799) );
  NOR U46539 ( .A(n45378), .B(n44428), .Z(n47031) );
  XOR U46540 ( .A(n45953), .B(n47034), .Z(n44428) );
  XOR U46541 ( .A(n47035), .B(n43457), .Z(n45378) );
  XNOR U46542 ( .A(n47036), .B(n47037), .Z(n45751) );
  XNOR U46543 ( .A(n46215), .B(n45803), .Z(n47037) );
  XOR U46544 ( .A(n47038), .B(n47039), .Z(n45803) );
  ANDN U46545 ( .B(n47040), .A(n47041), .Z(n47038) );
  XNOR U46546 ( .A(n47042), .B(n47043), .Z(n46215) );
  ANDN U46547 ( .B(n47044), .A(n47045), .Z(n47042) );
  XOR U46548 ( .A(n42873), .B(n47046), .Z(n47036) );
  XOR U46549 ( .A(n47047), .B(n44664), .Z(n47046) );
  XNOR U46550 ( .A(n47048), .B(n47049), .Z(n44664) );
  ANDN U46551 ( .B(n47050), .A(n47051), .Z(n47048) );
  XOR U46552 ( .A(n47052), .B(n47053), .Z(n42873) );
  ANDN U46553 ( .B(n47054), .A(n47055), .Z(n47052) );
  XNOR U46554 ( .A(n47057), .B(n47058), .Z(n33147) );
  XNOR U46555 ( .A(n32295), .B(n31027), .Z(n47058) );
  XNOR U46556 ( .A(n47059), .B(n33756), .Z(n31027) );
  XNOR U46557 ( .A(n42298), .B(n37797), .Z(n33756) );
  XOR U46558 ( .A(n41663), .B(n39106), .Z(n37797) );
  XNOR U46559 ( .A(n47060), .B(n47061), .Z(n39106) );
  XOR U46560 ( .A(n37087), .B(n40034), .Z(n47061) );
  XNOR U46561 ( .A(n47062), .B(n40587), .Z(n40034) );
  XOR U46562 ( .A(n47064), .B(n45664), .Z(n40838) );
  XOR U46563 ( .A(n47065), .B(n44512), .Z(n40420) );
  XNOR U46564 ( .A(n47066), .B(n40592), .Z(n37087) );
  XNOR U46565 ( .A(n47067), .B(n44544), .Z(n40592) );
  XNOR U46566 ( .A(n47068), .B(n43565), .Z(n40842) );
  XNOR U46567 ( .A(n47069), .B(n42461), .Z(n40424) );
  XOR U46568 ( .A(n35316), .B(n47070), .Z(n47060) );
  XOR U46569 ( .A(n43857), .B(n42230), .Z(n47070) );
  XNOR U46570 ( .A(n47071), .B(n40585), .Z(n42230) );
  XOR U46571 ( .A(n47072), .B(n44541), .Z(n40585) );
  ANDN U46572 ( .B(n40851), .A(n40416), .Z(n47071) );
  XOR U46573 ( .A(n47073), .B(n46528), .Z(n40416) );
  XNOR U46574 ( .A(n41733), .B(n47074), .Z(n40851) );
  IV U46575 ( .A(n45279), .Z(n41733) );
  XOR U46576 ( .A(n47075), .B(n47076), .Z(n46191) );
  XNOR U46577 ( .A(n46944), .B(n44851), .Z(n47076) );
  XOR U46578 ( .A(n47077), .B(n47078), .Z(n44851) );
  ANDN U46579 ( .B(n47079), .A(n46379), .Z(n47077) );
  XNOR U46580 ( .A(n47080), .B(n47081), .Z(n46944) );
  ANDN U46581 ( .B(n47082), .A(n46686), .Z(n47080) );
  XOR U46582 ( .A(n46642), .B(n47083), .Z(n47075) );
  XOR U46583 ( .A(n44676), .B(n46749), .Z(n47083) );
  XNOR U46584 ( .A(n47084), .B(n47085), .Z(n46749) );
  ANDN U46585 ( .B(n47086), .A(n46386), .Z(n47084) );
  XNOR U46586 ( .A(n47087), .B(n47088), .Z(n44676) );
  ANDN U46587 ( .B(n47089), .A(n46375), .Z(n47087) );
  XNOR U46588 ( .A(n47090), .B(n47091), .Z(n46642) );
  ANDN U46589 ( .B(n47092), .A(n47093), .Z(n47090) );
  XNOR U46590 ( .A(n47095), .B(n40594), .Z(n43857) );
  XOR U46591 ( .A(n45244), .B(n47096), .Z(n40594) );
  XOR U46592 ( .A(n47097), .B(n47098), .Z(n45244) );
  ANDN U46593 ( .B(n40855), .A(n40858), .Z(n47095) );
  XOR U46594 ( .A(n42683), .B(n46900), .Z(n40855) );
  XNOR U46595 ( .A(n47100), .B(n47101), .Z(n46900) );
  ANDN U46596 ( .B(n47102), .A(n47103), .Z(n47100) );
  XNOR U46597 ( .A(n40590), .B(n47104), .Z(n35316) );
  XNOR U46598 ( .A(n11417), .B(n47105), .Z(n47104) );
  XNOR U46599 ( .A(n44783), .B(n47106), .Z(n40411) );
  XOR U46600 ( .A(n47107), .B(n47108), .Z(n44783) );
  XOR U46601 ( .A(n47109), .B(n45135), .Z(n40847) );
  XOR U46602 ( .A(n47110), .B(n42654), .Z(n40590) );
  IV U46603 ( .A(n46601), .Z(n42654) );
  XNOR U46604 ( .A(n47111), .B(n47112), .Z(n46531) );
  XOR U46605 ( .A(n47113), .B(n44321), .Z(n47112) );
  XNOR U46606 ( .A(n47114), .B(n46959), .Z(n44321) );
  ANDN U46607 ( .B(n47115), .A(n47116), .Z(n47114) );
  XOR U46608 ( .A(n44405), .B(n47117), .Z(n47111) );
  XNOR U46609 ( .A(n47118), .B(n43816), .Z(n47117) );
  XOR U46610 ( .A(n47119), .B(n47120), .Z(n43816) );
  AND U46611 ( .A(n47121), .B(n47122), .Z(n47119) );
  XNOR U46612 ( .A(n47123), .B(n46969), .Z(n44405) );
  AND U46613 ( .A(n47124), .B(n47125), .Z(n47123) );
  XOR U46614 ( .A(n47127), .B(n47128), .Z(n41663) );
  XOR U46615 ( .A(n37927), .B(n41499), .Z(n47128) );
  XOR U46616 ( .A(n47129), .B(n40565), .Z(n41499) );
  XNOR U46617 ( .A(n44686), .B(n47130), .Z(n40565) );
  AND U46618 ( .A(n42217), .B(n41508), .Z(n47129) );
  XOR U46619 ( .A(n47133), .B(n45664), .Z(n41508) );
  XNOR U46620 ( .A(n43342), .B(n47134), .Z(n42217) );
  XNOR U46621 ( .A(n47135), .B(n40557), .Z(n37927) );
  XNOR U46622 ( .A(n47136), .B(n46745), .Z(n40557) );
  IV U46623 ( .A(n44479), .Z(n46745) );
  ANDN U46624 ( .B(n41510), .A(n42204), .Z(n47135) );
  XOR U46625 ( .A(n38410), .B(n47137), .Z(n47127) );
  XOR U46626 ( .A(n40365), .B(n39659), .Z(n47137) );
  XNOR U46627 ( .A(n47138), .B(n40561), .Z(n39659) );
  XOR U46628 ( .A(n47139), .B(n43916), .Z(n40561) );
  ANDN U46629 ( .B(n42304), .A(n41512), .Z(n47138) );
  XOR U46630 ( .A(n47140), .B(n47141), .Z(n41512) );
  IV U46631 ( .A(n42208), .Z(n42304) );
  XOR U46632 ( .A(n47142), .B(n42327), .Z(n42208) );
  IV U46633 ( .A(n44516), .Z(n42327) );
  XNOR U46634 ( .A(n47143), .B(n47144), .Z(n44516) );
  XNOR U46635 ( .A(n47145), .B(n40548), .Z(n40365) );
  XOR U46636 ( .A(n47146), .B(n45135), .Z(n40548) );
  ANDN U46637 ( .B(n41503), .A(n42221), .Z(n47145) );
  IV U46638 ( .A(n42311), .Z(n42221) );
  XNOR U46639 ( .A(n47147), .B(n42166), .Z(n42311) );
  XOR U46640 ( .A(n47148), .B(n47149), .Z(n42166) );
  XNOR U46641 ( .A(n46134), .B(n42494), .Z(n41503) );
  IV U46642 ( .A(n43581), .Z(n42494) );
  XOR U46643 ( .A(n47152), .B(n47153), .Z(n46134) );
  ANDN U46644 ( .B(n47154), .A(n47155), .Z(n47152) );
  XOR U46645 ( .A(n47156), .B(n40551), .Z(n38410) );
  XOR U46646 ( .A(n47157), .B(n46178), .Z(n40551) );
  ANDN U46647 ( .B(n42213), .A(n41505), .Z(n47156) );
  XNOR U46648 ( .A(n47158), .B(n44114), .Z(n41505) );
  XOR U46649 ( .A(n43598), .B(n47159), .Z(n42213) );
  XOR U46650 ( .A(n47160), .B(n41510), .Z(n42298) );
  XOR U46651 ( .A(n47161), .B(n47162), .Z(n41510) );
  ANDN U46652 ( .B(n42204), .A(n40555), .Z(n47160) );
  XNOR U46653 ( .A(n42329), .B(n47163), .Z(n40555) );
  XOR U46654 ( .A(n47164), .B(n43321), .Z(n42204) );
  ANDN U46655 ( .B(n33757), .A(n38849), .Z(n47059) );
  IV U46656 ( .A(n35649), .Z(n38849) );
  XOR U46657 ( .A(n46456), .B(n37623), .Z(n35649) );
  XOR U46658 ( .A(n40338), .B(n40373), .Z(n37623) );
  XNOR U46659 ( .A(n47165), .B(n47166), .Z(n40373) );
  XNOR U46660 ( .A(n45523), .B(n45292), .Z(n47166) );
  XNOR U46661 ( .A(n47167), .B(n45546), .Z(n45292) );
  XOR U46662 ( .A(n45080), .B(n47168), .Z(n45546) );
  ANDN U46663 ( .B(n45547), .A(n39729), .Z(n47167) );
  XNOR U46664 ( .A(n47169), .B(n45011), .Z(n39729) );
  XOR U46665 ( .A(n47170), .B(n46286), .Z(n45547) );
  XNOR U46666 ( .A(n47171), .B(n45538), .Z(n45523) );
  XOR U46667 ( .A(n47172), .B(n44816), .Z(n45538) );
  NOR U46668 ( .A(n46439), .B(n39725), .Z(n47171) );
  XOR U46669 ( .A(n41874), .B(n47173), .Z(n39725) );
  XOR U46670 ( .A(n47174), .B(n47175), .Z(n46798) );
  XNOR U46671 ( .A(n45795), .B(n44852), .Z(n47175) );
  XNOR U46672 ( .A(n47176), .B(n47177), .Z(n44852) );
  ANDN U46673 ( .B(n47178), .A(n47179), .Z(n47176) );
  XNOR U46674 ( .A(n47180), .B(n47181), .Z(n45795) );
  ANDN U46675 ( .B(n47182), .A(n47183), .Z(n47180) );
  XOR U46676 ( .A(n47184), .B(n47185), .Z(n47174) );
  XOR U46677 ( .A(n43578), .B(n46581), .Z(n47185) );
  XNOR U46678 ( .A(n47186), .B(n47187), .Z(n46581) );
  ANDN U46679 ( .B(n47188), .A(n47189), .Z(n47186) );
  XNOR U46680 ( .A(n47190), .B(n47191), .Z(n43578) );
  ANDN U46681 ( .B(n47192), .A(n47193), .Z(n47190) );
  XOR U46682 ( .A(n47194), .B(n47195), .Z(n47108) );
  XNOR U46683 ( .A(n47196), .B(n46736), .Z(n47195) );
  XNOR U46684 ( .A(n47197), .B(n47198), .Z(n46736) );
  NOR U46685 ( .A(n47199), .B(n47200), .Z(n47197) );
  XOR U46686 ( .A(n46270), .B(n47201), .Z(n47194) );
  XOR U46687 ( .A(n44538), .B(n44672), .Z(n47201) );
  XNOR U46688 ( .A(n47202), .B(n47203), .Z(n44672) );
  ANDN U46689 ( .B(n47204), .A(n47205), .Z(n47202) );
  XNOR U46690 ( .A(n47206), .B(n47207), .Z(n44538) );
  NOR U46691 ( .A(n47208), .B(n47209), .Z(n47206) );
  XNOR U46692 ( .A(n47210), .B(n47211), .Z(n46270) );
  NOR U46693 ( .A(n47212), .B(n47213), .Z(n47210) );
  XNOR U46694 ( .A(n47214), .B(n45554), .Z(n46439) );
  XOR U46695 ( .A(n46099), .B(n47215), .Z(n45554) );
  XOR U46696 ( .A(n47216), .B(n47217), .Z(n46099) );
  XOR U46697 ( .A(n47218), .B(n44660), .Z(n47217) );
  XNOR U46698 ( .A(n47219), .B(n47220), .Z(n44660) );
  ANDN U46699 ( .B(n47221), .A(n47222), .Z(n47219) );
  XNOR U46700 ( .A(n45509), .B(n47223), .Z(n47216) );
  XOR U46701 ( .A(n45146), .B(n47224), .Z(n47223) );
  XNOR U46702 ( .A(n47225), .B(n47226), .Z(n45146) );
  ANDN U46703 ( .B(n47227), .A(n47228), .Z(n47225) );
  XOR U46704 ( .A(n47229), .B(n47230), .Z(n45509) );
  AND U46705 ( .A(n47231), .B(n47232), .Z(n47229) );
  XOR U46706 ( .A(n38340), .B(n47233), .Z(n47165) );
  XOR U46707 ( .A(n42009), .B(n39629), .Z(n47233) );
  XNOR U46708 ( .A(n47234), .B(n45549), .Z(n39629) );
  XOR U46709 ( .A(n47235), .B(n45664), .Z(n45549) );
  ANDN U46710 ( .B(n45550), .A(n39719), .Z(n47234) );
  XOR U46711 ( .A(n46512), .B(n47238), .Z(n39719) );
  IV U46712 ( .A(n42668), .Z(n46512) );
  XNOR U46713 ( .A(n47239), .B(n42206), .Z(n45550) );
  XNOR U46714 ( .A(n47240), .B(n46397), .Z(n42009) );
  XOR U46715 ( .A(n45303), .B(n47241), .Z(n46397) );
  NOR U46716 ( .A(n40643), .B(n46435), .Z(n47240) );
  XOR U46717 ( .A(n47242), .B(n44943), .Z(n46435) );
  IV U46718 ( .A(n43765), .Z(n44943) );
  XNOR U46719 ( .A(n47246), .B(n46395), .Z(n38340) );
  XOR U46720 ( .A(n47247), .B(n44220), .Z(n46395) );
  XNOR U46721 ( .A(n47248), .B(n47249), .Z(n44220) );
  NOR U46722 ( .A(n39715), .B(n45543), .Z(n47246) );
  XNOR U46723 ( .A(n47250), .B(n42163), .Z(n45543) );
  XNOR U46724 ( .A(n47251), .B(n46120), .Z(n39715) );
  XOR U46725 ( .A(n47254), .B(n47255), .Z(n40338) );
  XOR U46726 ( .A(n43451), .B(n40573), .Z(n47255) );
  XNOR U46727 ( .A(n47256), .B(n42903), .Z(n40573) );
  XOR U46728 ( .A(n47257), .B(n44774), .Z(n42903) );
  ANDN U46729 ( .B(n41703), .A(n43473), .Z(n47256) );
  XNOR U46730 ( .A(n47260), .B(n42891), .Z(n43451) );
  XNOR U46731 ( .A(n47261), .B(n44119), .Z(n42891) );
  NOR U46732 ( .A(n46458), .B(n41707), .Z(n47260) );
  XOR U46733 ( .A(n47262), .B(n44777), .Z(n41707) );
  IV U46734 ( .A(n44932), .Z(n44777) );
  XOR U46735 ( .A(n47264), .B(n47265), .Z(n46794) );
  XNOR U46736 ( .A(n45217), .B(n47266), .Z(n47265) );
  XOR U46737 ( .A(n47267), .B(n47268), .Z(n45217) );
  ANDN U46738 ( .B(n47269), .A(n47270), .Z(n47267) );
  XNOR U46739 ( .A(n43333), .B(n47271), .Z(n47264) );
  XOR U46740 ( .A(n43589), .B(n42541), .Z(n47271) );
  XNOR U46741 ( .A(n47272), .B(n47273), .Z(n42541) );
  ANDN U46742 ( .B(n47274), .A(n47275), .Z(n47272) );
  XNOR U46743 ( .A(n47276), .B(n47277), .Z(n43589) );
  NOR U46744 ( .A(n47278), .B(n47279), .Z(n47276) );
  XNOR U46745 ( .A(n47280), .B(n47281), .Z(n43333) );
  AND U46746 ( .A(n47282), .B(n47283), .Z(n47280) );
  XOR U46747 ( .A(n47284), .B(n42219), .Z(n46458) );
  XNOR U46748 ( .A(n47285), .B(n47286), .Z(n45937) );
  XNOR U46749 ( .A(n46422), .B(n47287), .Z(n47286) );
  XNOR U46750 ( .A(n47288), .B(n47289), .Z(n46422) );
  ANDN U46751 ( .B(n47290), .A(n47291), .Z(n47288) );
  XOR U46752 ( .A(n47292), .B(n47293), .Z(n47285) );
  XOR U46753 ( .A(n45777), .B(n47294), .Z(n47293) );
  XNOR U46754 ( .A(n47295), .B(n47296), .Z(n45777) );
  ANDN U46755 ( .B(n47297), .A(n47298), .Z(n47295) );
  XNOR U46756 ( .A(n47299), .B(n47300), .Z(n46127) );
  XOR U46757 ( .A(n44836), .B(n45263), .Z(n47300) );
  XNOR U46758 ( .A(n47301), .B(n47282), .Z(n45263) );
  ANDN U46759 ( .B(n47302), .A(n47303), .Z(n47301) );
  XNOR U46760 ( .A(n47304), .B(n47279), .Z(n44836) );
  AND U46761 ( .A(n47305), .B(n47306), .Z(n47304) );
  XOR U46762 ( .A(n47307), .B(n47308), .Z(n47299) );
  XOR U46763 ( .A(n45089), .B(n46317), .Z(n47308) );
  XNOR U46764 ( .A(n47309), .B(n47310), .Z(n46317) );
  ANDN U46765 ( .B(n47311), .A(n47312), .Z(n47309) );
  XNOR U46766 ( .A(n47313), .B(n47275), .Z(n45089) );
  ANDN U46767 ( .B(n47314), .A(n47315), .Z(n47313) );
  XOR U46768 ( .A(n37257), .B(n47316), .Z(n47254) );
  XOR U46769 ( .A(n40664), .B(n41137), .Z(n47316) );
  XOR U46770 ( .A(n47317), .B(n42901), .Z(n41137) );
  XNOR U46771 ( .A(n47318), .B(n44201), .Z(n42901) );
  NOR U46772 ( .A(n43458), .B(n41697), .Z(n47317) );
  XOR U46773 ( .A(n44225), .B(n47319), .Z(n41697) );
  XNOR U46774 ( .A(n47320), .B(n47321), .Z(n44225) );
  XOR U46775 ( .A(n47322), .B(n41585), .Z(n43458) );
  IV U46776 ( .A(n42524), .Z(n41585) );
  XNOR U46777 ( .A(n47323), .B(n42899), .Z(n40664) );
  XOR U46778 ( .A(n47324), .B(n45221), .Z(n42899) );
  XNOR U46779 ( .A(n45953), .B(n47325), .Z(n41693) );
  XOR U46780 ( .A(n47326), .B(n43546), .Z(n43469) );
  IV U46781 ( .A(n46178), .Z(n43546) );
  XNOR U46782 ( .A(n47327), .B(n42895), .Z(n37257) );
  XOR U46783 ( .A(n47328), .B(n43557), .Z(n42895) );
  IV U46784 ( .A(n44571), .Z(n43557) );
  NOR U46785 ( .A(n46466), .B(n43460), .Z(n47327) );
  XNOR U46786 ( .A(n46330), .B(n44503), .Z(n43460) );
  XOR U46787 ( .A(n46946), .B(n46409), .Z(n44503) );
  XNOR U46788 ( .A(n47329), .B(n47330), .Z(n46409) );
  XNOR U46789 ( .A(n42396), .B(n47331), .Z(n47330) );
  XNOR U46790 ( .A(n47332), .B(n47333), .Z(n42396) );
  ANDN U46791 ( .B(n46333), .A(n46334), .Z(n47332) );
  XOR U46792 ( .A(n42463), .B(n47334), .Z(n47329) );
  XOR U46793 ( .A(n47335), .B(n46245), .Z(n47334) );
  XNOR U46794 ( .A(n47336), .B(n47337), .Z(n46245) );
  NOR U46795 ( .A(n46337), .B(n46338), .Z(n47336) );
  XNOR U46796 ( .A(n47338), .B(n47339), .Z(n42463) );
  XNOR U46797 ( .A(n47340), .B(n47341), .Z(n46946) );
  XNOR U46798 ( .A(n46091), .B(n46549), .Z(n47341) );
  XNOR U46799 ( .A(n47342), .B(n46381), .Z(n46549) );
  NOR U46800 ( .A(n47078), .B(n47079), .Z(n47342) );
  IV U46801 ( .A(n47343), .Z(n47078) );
  XNOR U46802 ( .A(n47344), .B(n46688), .Z(n46091) );
  ANDN U46803 ( .B(n47081), .A(n47082), .Z(n47344) );
  XOR U46804 ( .A(n45298), .B(n47345), .Z(n47340) );
  XOR U46805 ( .A(n45158), .B(n42686), .Z(n47345) );
  XNOR U46806 ( .A(n47346), .B(n46377), .Z(n42686) );
  XNOR U46807 ( .A(n47347), .B(n46388), .Z(n45158) );
  ANDN U46808 ( .B(n47085), .A(n47086), .Z(n47347) );
  XOR U46809 ( .A(n47348), .B(n47349), .Z(n45298) );
  XNOR U46810 ( .A(n47350), .B(n47351), .Z(n46330) );
  ANDN U46811 ( .B(n47352), .A(n47353), .Z(n47350) );
  XNOR U46812 ( .A(n42329), .B(n47354), .Z(n46466) );
  XNOR U46813 ( .A(n47357), .B(n43473), .Z(n46456) );
  XOR U46814 ( .A(n47358), .B(n43719), .Z(n43473) );
  NOR U46815 ( .A(n41703), .B(n41705), .Z(n47357) );
  XOR U46816 ( .A(n47359), .B(n46528), .Z(n41705) );
  IV U46817 ( .A(n44862), .Z(n46528) );
  XNOR U46818 ( .A(n46793), .B(n47360), .Z(n44862) );
  XOR U46819 ( .A(n47361), .B(n47362), .Z(n46793) );
  XOR U46820 ( .A(n44936), .B(n45729), .Z(n47362) );
  XNOR U46821 ( .A(n47363), .B(n47364), .Z(n45729) );
  ANDN U46822 ( .B(n47365), .A(n47366), .Z(n47363) );
  XOR U46823 ( .A(n47367), .B(n47368), .Z(n44936) );
  ANDN U46824 ( .B(n47369), .A(n47370), .Z(n47367) );
  XNOR U46825 ( .A(n45492), .B(n47371), .Z(n47361) );
  XOR U46826 ( .A(n46521), .B(n47372), .Z(n47371) );
  XNOR U46827 ( .A(n47373), .B(n47374), .Z(n46521) );
  ANDN U46828 ( .B(n47375), .A(n47289), .Z(n47373) );
  XNOR U46829 ( .A(n47376), .B(n47377), .Z(n45492) );
  ANDN U46830 ( .B(n47378), .A(n47296), .Z(n47376) );
  XOR U46831 ( .A(n47379), .B(n46932), .Z(n41703) );
  IV U46832 ( .A(n45519), .Z(n46932) );
  XOR U46833 ( .A(n41801), .B(n43688), .Z(n33757) );
  XNOR U46834 ( .A(n47380), .B(n45207), .Z(n43688) );
  ANDN U46835 ( .B(n43180), .A(n43841), .Z(n47380) );
  IV U46836 ( .A(n43181), .Z(n43841) );
  XOR U46837 ( .A(n47381), .B(n46447), .Z(n43181) );
  IV U46838 ( .A(n46414), .Z(n46447) );
  XNOR U46839 ( .A(n42647), .B(n42080), .Z(n41801) );
  XNOR U46840 ( .A(n47382), .B(n47383), .Z(n42080) );
  XNOR U46841 ( .A(n39868), .B(n38894), .Z(n47383) );
  XNOR U46842 ( .A(n47384), .B(n43842), .Z(n38894) );
  XOR U46843 ( .A(n47385), .B(n45117), .Z(n43842) );
  XOR U46844 ( .A(n46403), .B(n47386), .Z(n45207) );
  XOR U46845 ( .A(n47387), .B(n47388), .Z(n43180) );
  XNOR U46846 ( .A(n47389), .B(n43850), .Z(n39868) );
  XOR U46847 ( .A(n47390), .B(n46198), .Z(n43850) );
  NOR U46848 ( .A(n43696), .B(n43163), .Z(n47389) );
  XOR U46849 ( .A(n47391), .B(n44520), .Z(n43163) );
  XOR U46850 ( .A(n47392), .B(n46343), .Z(n43696) );
  IV U46851 ( .A(n43829), .Z(n46343) );
  XOR U46852 ( .A(n39691), .B(n47393), .Z(n47382) );
  XNOR U46853 ( .A(n41568), .B(n40638), .Z(n47393) );
  XNOR U46854 ( .A(n47394), .B(n43839), .Z(n40638) );
  XNOR U46855 ( .A(n47395), .B(n43680), .Z(n43839) );
  XOR U46856 ( .A(n47396), .B(n47397), .Z(n43693) );
  IV U46857 ( .A(n43167), .Z(n43694) );
  XOR U46858 ( .A(n47398), .B(n45922), .Z(n43167) );
  XNOR U46859 ( .A(n47400), .B(n44488), .Z(n43853) );
  ANDN U46860 ( .B(n43690), .A(n43176), .Z(n47399) );
  XNOR U46861 ( .A(n43346), .B(n47401), .Z(n43176) );
  XOR U46862 ( .A(n47402), .B(n45247), .Z(n43690) );
  XNOR U46863 ( .A(n47403), .B(n43847), .Z(n39691) );
  XOR U46864 ( .A(n47404), .B(n44467), .Z(n43847) );
  NOR U46865 ( .A(n43698), .B(n43172), .Z(n47403) );
  XOR U46866 ( .A(n47405), .B(n45080), .Z(n43172) );
  XNOR U46867 ( .A(n47406), .B(n47407), .Z(n43698) );
  XOR U46868 ( .A(n47408), .B(n47409), .Z(n42647) );
  XNOR U46869 ( .A(n44636), .B(n38816), .Z(n47409) );
  XOR U46870 ( .A(n47410), .B(n43821), .Z(n38816) );
  ANDN U46871 ( .B(n43402), .A(n41379), .Z(n47410) );
  XOR U46872 ( .A(n42860), .B(n47411), .Z(n41379) );
  XOR U46873 ( .A(n47412), .B(n43834), .Z(n44636) );
  ANDN U46874 ( .B(n43405), .A(n41388), .Z(n47412) );
  XOR U46875 ( .A(n44535), .B(n47413), .Z(n41388) );
  XOR U46876 ( .A(n46131), .B(n47414), .Z(n44535) );
  XOR U46877 ( .A(n47415), .B(n47416), .Z(n46131) );
  XOR U46878 ( .A(n47417), .B(n46157), .Z(n47416) );
  XOR U46879 ( .A(n47418), .B(n47419), .Z(n46157) );
  ANDN U46880 ( .B(n47420), .A(n47421), .Z(n47418) );
  XOR U46881 ( .A(n43336), .B(n47422), .Z(n47415) );
  XOR U46882 ( .A(n46062), .B(n46717), .Z(n47422) );
  XOR U46883 ( .A(n47423), .B(n47424), .Z(n46717) );
  ANDN U46884 ( .B(n47425), .A(n47426), .Z(n47423) );
  XOR U46885 ( .A(n47427), .B(n47428), .Z(n46062) );
  ANDN U46886 ( .B(n47429), .A(n47430), .Z(n47427) );
  XNOR U46887 ( .A(n47431), .B(n47432), .Z(n43336) );
  ANDN U46888 ( .B(n47433), .A(n47434), .Z(n47431) );
  XNOR U46889 ( .A(n38276), .B(n47435), .Z(n47408) );
  XOR U46890 ( .A(n39474), .B(n47436), .Z(n47435) );
  XOR U46891 ( .A(n47437), .B(n43826), .Z(n39474) );
  ANDN U46892 ( .B(n43398), .A(n43399), .Z(n47437) );
  XOR U46893 ( .A(n47438), .B(n46176), .Z(n43399) );
  XOR U46894 ( .A(n47439), .B(n43830), .Z(n38276) );
  IV U46895 ( .A(n47440), .Z(n43830) );
  ANDN U46896 ( .B(n43409), .A(n41392), .Z(n47439) );
  XNOR U46897 ( .A(n47441), .B(n43468), .Z(n41392) );
  IV U46898 ( .A(n46443), .Z(n43468) );
  XNOR U46899 ( .A(n47442), .B(n33747), .Z(n32295) );
  XOR U46900 ( .A(n45027), .B(n39219), .Z(n33747) );
  XNOR U46901 ( .A(n47443), .B(n47444), .Z(n42005) );
  XOR U46902 ( .A(n38907), .B(n39285), .Z(n47444) );
  XNOR U46903 ( .A(n47445), .B(n42763), .Z(n39285) );
  XNOR U46904 ( .A(n47446), .B(n44201), .Z(n42763) );
  ANDN U46905 ( .B(n42111), .A(n42762), .Z(n47445) );
  XOR U46906 ( .A(n47447), .B(n47448), .Z(n42762) );
  XNOR U46907 ( .A(n47449), .B(n44500), .Z(n42111) );
  IV U46908 ( .A(n47450), .Z(n44500) );
  XOR U46909 ( .A(n47451), .B(n42776), .Z(n38907) );
  XOR U46910 ( .A(n47452), .B(n45135), .Z(n42776) );
  XOR U46911 ( .A(n47453), .B(n47454), .Z(n45135) );
  ANDN U46912 ( .B(n42777), .A(n42106), .Z(n47451) );
  XOR U46913 ( .A(n47455), .B(n47456), .Z(n42106) );
  XOR U46914 ( .A(n44032), .B(n47457), .Z(n42777) );
  IV U46915 ( .A(n45820), .Z(n44032) );
  XNOR U46916 ( .A(n47458), .B(n47459), .Z(n45820) );
  XNOR U46917 ( .A(n40209), .B(n47460), .Z(n47443) );
  XNOR U46918 ( .A(n38965), .B(n38892), .Z(n47460) );
  XNOR U46919 ( .A(n47461), .B(n44739), .Z(n38892) );
  IV U46920 ( .A(n42771), .Z(n44739) );
  XOR U46921 ( .A(n47462), .B(n45646), .Z(n42771) );
  ANDN U46922 ( .B(n42119), .A(n42770), .Z(n47461) );
  IV U46923 ( .A(n45794), .Z(n42770) );
  XOR U46924 ( .A(n47463), .B(n42691), .Z(n45794) );
  XNOR U46925 ( .A(n47464), .B(n45397), .Z(n42119) );
  XOR U46926 ( .A(n47465), .B(n42766), .Z(n38965) );
  XNOR U46927 ( .A(n47466), .B(n44533), .Z(n42766) );
  IV U46928 ( .A(n45575), .Z(n44533) );
  XNOR U46929 ( .A(n47467), .B(n47468), .Z(n45575) );
  NOR U46930 ( .A(n45797), .B(n45798), .Z(n47465) );
  XNOR U46931 ( .A(n47469), .B(n45497), .Z(n45798) );
  IV U46932 ( .A(n42767), .Z(n45797) );
  XOR U46933 ( .A(n47470), .B(n42301), .Z(n42767) );
  XOR U46934 ( .A(n47471), .B(n42773), .Z(n40209) );
  XNOR U46935 ( .A(n44864), .B(n47472), .Z(n42773) );
  ANDN U46936 ( .B(n42774), .A(n42115), .Z(n47471) );
  XOR U46937 ( .A(n47473), .B(n45249), .Z(n42115) );
  XOR U46938 ( .A(n45080), .B(n47474), .Z(n42774) );
  XNOR U46939 ( .A(n47477), .B(n47478), .Z(n44080) );
  XNOR U46940 ( .A(n37864), .B(n36966), .Z(n47478) );
  XNOR U46941 ( .A(n47479), .B(n44438), .Z(n36966) );
  XOR U46942 ( .A(n47480), .B(n44882), .Z(n44438) );
  XOR U46943 ( .A(n46516), .B(n45428), .Z(n44882) );
  XOR U46944 ( .A(n47481), .B(n47482), .Z(n45428) );
  XNOR U46945 ( .A(n47483), .B(n45482), .Z(n47482) );
  XOR U46946 ( .A(n47484), .B(n46987), .Z(n45482) );
  AND U46947 ( .A(n47485), .B(n47486), .Z(n47484) );
  XOR U46948 ( .A(n45782), .B(n47487), .Z(n47481) );
  XOR U46949 ( .A(n47488), .B(n47489), .Z(n47487) );
  XNOR U46950 ( .A(n47490), .B(n46995), .Z(n45782) );
  NOR U46951 ( .A(n47491), .B(n47492), .Z(n47490) );
  XOR U46952 ( .A(n47493), .B(n47494), .Z(n46516) );
  XNOR U46953 ( .A(n45326), .B(n41889), .Z(n47494) );
  XNOR U46954 ( .A(n47495), .B(n47496), .Z(n41889) );
  XNOR U46955 ( .A(n47499), .B(n47500), .Z(n45326) );
  NOR U46956 ( .A(n47501), .B(n47502), .Z(n47499) );
  XOR U46957 ( .A(n47503), .B(n47504), .Z(n47493) );
  XOR U46958 ( .A(n42679), .B(n47141), .Z(n47504) );
  XNOR U46959 ( .A(n47505), .B(n47506), .Z(n47141) );
  XNOR U46960 ( .A(n47509), .B(n47510), .Z(n42679) );
  ANDN U46961 ( .B(n47511), .A(n47512), .Z(n47509) );
  AND U46962 ( .A(n44439), .B(n47513), .Z(n47479) );
  XNOR U46963 ( .A(n47514), .B(n44452), .Z(n37864) );
  XNOR U46964 ( .A(n47515), .B(n43574), .Z(n44452) );
  XNOR U46965 ( .A(n47516), .B(n47517), .Z(n43574) );
  AND U46966 ( .A(n45026), .B(n44453), .Z(n47514) );
  XNOR U46967 ( .A(n47518), .B(n43719), .Z(n44453) );
  XOR U46968 ( .A(n42757), .B(n47521), .Z(n47477) );
  XOR U46969 ( .A(n35164), .B(n38164), .Z(n47521) );
  XOR U46970 ( .A(n47522), .B(n44716), .Z(n38164) );
  XOR U46971 ( .A(n47523), .B(n45569), .Z(n44716) );
  AND U46972 ( .A(n44715), .B(n45024), .Z(n47522) );
  XNOR U46973 ( .A(n45252), .B(n47524), .Z(n44715) );
  XOR U46974 ( .A(n47525), .B(n47526), .Z(n45252) );
  XOR U46975 ( .A(n47527), .B(n44449), .Z(n35164) );
  XNOR U46976 ( .A(n47528), .B(n47529), .Z(n44449) );
  AND U46977 ( .A(n45031), .B(n44448), .Z(n47527) );
  XOR U46978 ( .A(n45786), .B(n46782), .Z(n44448) );
  XNOR U46979 ( .A(n47530), .B(n47531), .Z(n46782) );
  ANDN U46980 ( .B(n47532), .A(n47533), .Z(n47530) );
  XNOR U46981 ( .A(n47534), .B(n44442), .Z(n42757) );
  XNOR U46982 ( .A(n47535), .B(n43920), .Z(n44442) );
  XNOR U46983 ( .A(n47536), .B(n47537), .Z(n43920) );
  AND U46984 ( .A(n46558), .B(n44443), .Z(n47534) );
  XNOR U46985 ( .A(n47538), .B(n47450), .Z(n44443) );
  XNOR U46986 ( .A(n47539), .B(n44439), .Z(n45027) );
  XOR U46987 ( .A(n47540), .B(n41742), .Z(n44439) );
  NOR U46988 ( .A(n47513), .B(n44727), .Z(n47539) );
  ANDN U46989 ( .B(n37586), .A(n37585), .Z(n47442) );
  IV U46990 ( .A(n33748), .Z(n37585) );
  XOR U46991 ( .A(n46072), .B(n35940), .Z(n33748) );
  XOR U46992 ( .A(n47541), .B(n47542), .Z(n45977) );
  XOR U46993 ( .A(n39618), .B(n38776), .Z(n47542) );
  XOR U46994 ( .A(n47543), .B(n39958), .Z(n38776) );
  XOR U46995 ( .A(n47544), .B(n45221), .Z(n39958) );
  ANDN U46996 ( .B(n39959), .A(n45927), .Z(n47543) );
  XOR U46997 ( .A(n47545), .B(n46405), .Z(n45927) );
  IV U46998 ( .A(n44512), .Z(n46405) );
  XNOR U46999 ( .A(n47249), .B(n47546), .Z(n44512) );
  XNOR U47000 ( .A(n47547), .B(n47548), .Z(n47249) );
  XNOR U47001 ( .A(n47549), .B(n44478), .Z(n47548) );
  XOR U47002 ( .A(n47550), .B(n47551), .Z(n44478) );
  ANDN U47003 ( .B(n47552), .A(n47553), .Z(n47550) );
  XNOR U47004 ( .A(n45270), .B(n47554), .Z(n47547) );
  XOR U47005 ( .A(n46744), .B(n47136), .Z(n47554) );
  XOR U47006 ( .A(n47555), .B(n47556), .Z(n47136) );
  ANDN U47007 ( .B(n47557), .A(n47558), .Z(n47555) );
  XOR U47008 ( .A(n47559), .B(n47560), .Z(n46744) );
  ANDN U47009 ( .B(n47561), .A(n47562), .Z(n47559) );
  XOR U47010 ( .A(n47563), .B(n47564), .Z(n45270) );
  AND U47011 ( .A(n47565), .B(n47566), .Z(n47563) );
  XOR U47012 ( .A(n47567), .B(n45814), .Z(n39959) );
  XNOR U47013 ( .A(n47568), .B(n45050), .Z(n39618) );
  IV U47014 ( .A(n45061), .Z(n45050) );
  XOR U47015 ( .A(n46022), .B(n46895), .Z(n45061) );
  XNOR U47016 ( .A(n47569), .B(n47570), .Z(n46895) );
  ANDN U47017 ( .B(n47571), .A(n47572), .Z(n47569) );
  IV U47018 ( .A(n42683), .Z(n46022) );
  XNOR U47019 ( .A(n47573), .B(n47574), .Z(n42683) );
  ANDN U47020 ( .B(n45924), .A(n45060), .Z(n47568) );
  XOR U47021 ( .A(n47575), .B(n46183), .Z(n45060) );
  XNOR U47022 ( .A(n47576), .B(n47577), .Z(n46183) );
  XNOR U47023 ( .A(n47578), .B(n45629), .Z(n45924) );
  IV U47024 ( .A(n44806), .Z(n45629) );
  XOR U47025 ( .A(n47579), .B(n47580), .Z(n44806) );
  XNOR U47026 ( .A(n39187), .B(n47581), .Z(n47541) );
  XNOR U47027 ( .A(n39245), .B(n38861), .Z(n47581) );
  XOR U47028 ( .A(n47582), .B(n39954), .Z(n38861) );
  XOR U47029 ( .A(n47583), .B(n47456), .Z(n39954) );
  XNOR U47030 ( .A(n47585), .B(n44191), .Z(n39965) );
  ANDN U47031 ( .B(n39966), .A(n45914), .Z(n47584) );
  IV U47032 ( .A(n46066), .Z(n45914) );
  XOR U47033 ( .A(n46421), .B(n47287), .Z(n46066) );
  XNOR U47034 ( .A(n47586), .B(n47370), .Z(n47287) );
  ANDN U47035 ( .B(n47587), .A(n47588), .Z(n47586) );
  XOR U47036 ( .A(n47589), .B(n47590), .Z(n39966) );
  XOR U47037 ( .A(n47591), .B(n40078), .Z(n39187) );
  XNOR U47038 ( .A(n47592), .B(n45085), .Z(n40078) );
  ANDN U47039 ( .B(n40079), .A(n45910), .Z(n47591) );
  XNOR U47040 ( .A(n45300), .B(n47593), .Z(n45910) );
  IV U47041 ( .A(n44520), .Z(n45300) );
  XOR U47042 ( .A(n47594), .B(n44816), .Z(n40079) );
  XNOR U47043 ( .A(n47595), .B(n47596), .Z(n43274) );
  XOR U47044 ( .A(n38469), .B(n41335), .Z(n47596) );
  XNOR U47045 ( .A(n47597), .B(n41355), .Z(n41335) );
  IV U47046 ( .A(n45039), .Z(n41355) );
  XOR U47047 ( .A(n47598), .B(n44488), .Z(n45039) );
  ANDN U47048 ( .B(n44642), .A(n41354), .Z(n47597) );
  XOR U47049 ( .A(n43967), .B(n47599), .Z(n41354) );
  XNOR U47050 ( .A(n47600), .B(n47601), .Z(n38469) );
  ANDN U47051 ( .B(n44645), .A(n41345), .Z(n47600) );
  XOR U47052 ( .A(n47602), .B(n47603), .Z(n41345) );
  XOR U47053 ( .A(n40647), .B(n47604), .Z(n47595) );
  XNOR U47054 ( .A(n39529), .B(n37060), .Z(n47604) );
  XNOR U47055 ( .A(n47605), .B(n41341), .Z(n37060) );
  XOR U47056 ( .A(n47606), .B(n44550), .Z(n41341) );
  XNOR U47057 ( .A(n47607), .B(n46427), .Z(n44550) );
  XNOR U47058 ( .A(n47608), .B(n47609), .Z(n46427) );
  XNOR U47059 ( .A(n47610), .B(n45846), .Z(n47609) );
  XNOR U47060 ( .A(n47611), .B(n47612), .Z(n45846) );
  ANDN U47061 ( .B(n47613), .A(n47614), .Z(n47611) );
  XNOR U47062 ( .A(n45724), .B(n47615), .Z(n47608) );
  XOR U47063 ( .A(n40839), .B(n45560), .Z(n47615) );
  XNOR U47064 ( .A(n47616), .B(n47617), .Z(n45560) );
  ANDN U47065 ( .B(n47618), .A(n47619), .Z(n47616) );
  XNOR U47066 ( .A(n47620), .B(n47621), .Z(n40839) );
  ANDN U47067 ( .B(n47622), .A(n47623), .Z(n47620) );
  XNOR U47068 ( .A(n47624), .B(n47625), .Z(n45724) );
  ANDN U47069 ( .B(n41342), .A(n44648), .Z(n47605) );
  XNOR U47070 ( .A(n46403), .B(n47628), .Z(n41342) );
  XNOR U47071 ( .A(n47629), .B(n41359), .Z(n39529) );
  XOR U47072 ( .A(n47630), .B(n45371), .Z(n41359) );
  ANDN U47073 ( .B(n44651), .A(n41358), .Z(n47629) );
  XOR U47074 ( .A(n47631), .B(n47632), .Z(n41358) );
  XNOR U47075 ( .A(n47633), .B(n41351), .Z(n40647) );
  XOR U47076 ( .A(n47634), .B(n44039), .Z(n41351) );
  IV U47077 ( .A(n47590), .Z(n44039) );
  ANDN U47078 ( .B(n44655), .A(n41350), .Z(n47633) );
  XOR U47079 ( .A(n46632), .B(n46758), .Z(n41350) );
  XNOR U47080 ( .A(n47635), .B(n47636), .Z(n46632) );
  AND U47081 ( .A(n47637), .B(n47638), .Z(n47635) );
  XNOR U47082 ( .A(n47639), .B(n39955), .Z(n46072) );
  XNOR U47083 ( .A(n47640), .B(n47641), .Z(n39955) );
  ANDN U47084 ( .B(n45053), .A(n45918), .Z(n47639) );
  XOR U47085 ( .A(n44459), .B(n47642), .Z(n45918) );
  IV U47086 ( .A(n44847), .Z(n44459) );
  XOR U47087 ( .A(n46210), .B(n47643), .Z(n44847) );
  XOR U47088 ( .A(n47644), .B(n47645), .Z(n46210) );
  XOR U47089 ( .A(n47578), .B(n45628), .Z(n47645) );
  XOR U47090 ( .A(n47646), .B(n47647), .Z(n45628) );
  ANDN U47091 ( .B(n47648), .A(n47649), .Z(n47646) );
  XNOR U47092 ( .A(n47650), .B(n47651), .Z(n47578) );
  AND U47093 ( .A(n47652), .B(n47653), .Z(n47650) );
  XOR U47094 ( .A(n44805), .B(n47654), .Z(n47644) );
  XOR U47095 ( .A(n46101), .B(n46350), .Z(n47654) );
  XNOR U47096 ( .A(n47655), .B(n47656), .Z(n46350) );
  ANDN U47097 ( .B(n47657), .A(n47658), .Z(n47655) );
  XNOR U47098 ( .A(n47659), .B(n47660), .Z(n46101) );
  ANDN U47099 ( .B(n47661), .A(n47662), .Z(n47659) );
  XNOR U47100 ( .A(n47663), .B(n47664), .Z(n44805) );
  XNOR U47101 ( .A(n47667), .B(n45091), .Z(n45053) );
  XNOR U47102 ( .A(n38126), .B(n41210), .Z(n37586) );
  XOR U47103 ( .A(n47668), .B(n42961), .Z(n41210) );
  NOR U47104 ( .A(n41981), .B(n41982), .Z(n47668) );
  XOR U47105 ( .A(n45014), .B(n47669), .Z(n41982) );
  IV U47106 ( .A(n38985), .Z(n38126) );
  XOR U47107 ( .A(n42028), .B(n39704), .Z(n38985) );
  XOR U47108 ( .A(n47670), .B(n47671), .Z(n39704) );
  XOR U47109 ( .A(n38628), .B(n37933), .Z(n47671) );
  XOR U47110 ( .A(n47672), .B(n43624), .Z(n37933) );
  IV U47111 ( .A(n44576), .Z(n43624) );
  XOR U47112 ( .A(n47673), .B(n44741), .Z(n44576) );
  ANDN U47113 ( .B(n41222), .A(n43623), .Z(n47672) );
  IV U47114 ( .A(n41221), .Z(n43623) );
  XOR U47115 ( .A(n46635), .B(n47674), .Z(n41221) );
  XNOR U47116 ( .A(n47675), .B(n45871), .Z(n46635) );
  AND U47117 ( .A(n47676), .B(n47677), .Z(n47675) );
  XNOR U47118 ( .A(n47678), .B(n47679), .Z(n41222) );
  XNOR U47119 ( .A(n47680), .B(n42953), .Z(n38628) );
  XOR U47120 ( .A(n47681), .B(n43102), .Z(n42953) );
  ANDN U47121 ( .B(n41213), .A(n41212), .Z(n47680) );
  XOR U47122 ( .A(n43346), .B(n47684), .Z(n41212) );
  XOR U47123 ( .A(n47685), .B(n44544), .Z(n41213) );
  XOR U47124 ( .A(n42948), .B(n47686), .Z(n47670) );
  XNOR U47125 ( .A(n41797), .B(n37721), .Z(n47686) );
  XNOR U47126 ( .A(n47687), .B(n42962), .Z(n37721) );
  XOR U47127 ( .A(n47012), .B(n44270), .Z(n42962) );
  IV U47128 ( .A(n44564), .Z(n44270) );
  XOR U47129 ( .A(n47688), .B(n47689), .Z(n44564) );
  XNOR U47130 ( .A(n47690), .B(n47691), .Z(n47012) );
  NOR U47131 ( .A(n46869), .B(n46868), .Z(n47690) );
  ANDN U47132 ( .B(n41981), .A(n42961), .Z(n47687) );
  XOR U47133 ( .A(n46021), .B(n47692), .Z(n42961) );
  XNOR U47134 ( .A(n47693), .B(n47694), .Z(n46021) );
  XNOR U47135 ( .A(n47695), .B(n42157), .Z(n41981) );
  XOR U47136 ( .A(n47696), .B(n42955), .Z(n41797) );
  XOR U47137 ( .A(n47697), .B(n42325), .Z(n42955) );
  ANDN U47138 ( .B(n41226), .A(n41225), .Z(n47696) );
  XOR U47139 ( .A(n47698), .B(n47450), .Z(n41225) );
  XNOR U47140 ( .A(n46883), .B(n47699), .Z(n47450) );
  XNOR U47141 ( .A(n47700), .B(n47701), .Z(n46883) );
  XOR U47142 ( .A(n44204), .B(n45180), .Z(n47701) );
  XNOR U47143 ( .A(n47702), .B(n47703), .Z(n45180) );
  ANDN U47144 ( .B(n47704), .A(n47705), .Z(n47702) );
  XOR U47145 ( .A(n47706), .B(n47707), .Z(n44204) );
  ANDN U47146 ( .B(n47708), .A(n47709), .Z(n47706) );
  XOR U47147 ( .A(n47710), .B(n47711), .Z(n47700) );
  XOR U47148 ( .A(n45162), .B(n44870), .Z(n47711) );
  XNOR U47149 ( .A(n47712), .B(n47713), .Z(n44870) );
  ANDN U47150 ( .B(n47714), .A(n47715), .Z(n47712) );
  XNOR U47151 ( .A(n47716), .B(n47717), .Z(n45162) );
  ANDN U47152 ( .B(n47718), .A(n47719), .Z(n47716) );
  XNOR U47153 ( .A(n47720), .B(n45221), .Z(n41226) );
  XNOR U47154 ( .A(n47721), .B(n46731), .Z(n45221) );
  XOR U47155 ( .A(n47722), .B(n47723), .Z(n46731) );
  XOR U47156 ( .A(n46701), .B(n47724), .Z(n47723) );
  XNOR U47157 ( .A(n47725), .B(n47726), .Z(n46701) );
  XNOR U47158 ( .A(n44194), .B(n47729), .Z(n47722) );
  XNOR U47159 ( .A(n46654), .B(n47730), .Z(n47729) );
  XNOR U47160 ( .A(n47731), .B(n47732), .Z(n46654) );
  AND U47161 ( .A(n47733), .B(n47734), .Z(n47731) );
  XOR U47162 ( .A(n47735), .B(n47736), .Z(n44194) );
  AND U47163 ( .A(n47737), .B(n47738), .Z(n47735) );
  XNOR U47164 ( .A(n47739), .B(n44591), .Z(n42948) );
  IV U47165 ( .A(n42959), .Z(n44591) );
  XNOR U47166 ( .A(n47740), .B(n47407), .Z(n42959) );
  ANDN U47167 ( .B(n41217), .A(n41218), .Z(n47739) );
  XOR U47168 ( .A(n43083), .B(n47741), .Z(n41218) );
  XOR U47169 ( .A(n46772), .B(n47030), .Z(n43083) );
  XNOR U47170 ( .A(n47742), .B(n47743), .Z(n47030) );
  XOR U47171 ( .A(n45235), .B(n47744), .Z(n47743) );
  XNOR U47172 ( .A(n47745), .B(n47746), .Z(n45235) );
  AND U47173 ( .A(n47747), .B(n47748), .Z(n47745) );
  XOR U47174 ( .A(n47749), .B(n47750), .Z(n47742) );
  XOR U47175 ( .A(n47751), .B(n46053), .Z(n47750) );
  XNOR U47176 ( .A(n47752), .B(n47753), .Z(n46053) );
  AND U47177 ( .A(n47754), .B(n47755), .Z(n47752) );
  XOR U47178 ( .A(n47756), .B(n47757), .Z(n46772) );
  XOR U47179 ( .A(n45831), .B(n46449), .Z(n47757) );
  XNOR U47180 ( .A(n47758), .B(n47759), .Z(n46449) );
  AND U47181 ( .A(n47760), .B(n47761), .Z(n47758) );
  XNOR U47182 ( .A(n47762), .B(n47763), .Z(n45831) );
  AND U47183 ( .A(n47764), .B(n47765), .Z(n47762) );
  XOR U47184 ( .A(n45267), .B(n47766), .Z(n47756) );
  XNOR U47185 ( .A(n45209), .B(n43334), .Z(n47766) );
  XOR U47186 ( .A(n47767), .B(n47768), .Z(n43334) );
  ANDN U47187 ( .B(n47769), .A(n47770), .Z(n47767) );
  XNOR U47188 ( .A(n47771), .B(n47772), .Z(n45209) );
  ANDN U47189 ( .B(n47773), .A(n47774), .Z(n47771) );
  XNOR U47190 ( .A(n47775), .B(n47776), .Z(n45267) );
  ANDN U47191 ( .B(n47777), .A(n47778), .Z(n47775) );
  XOR U47192 ( .A(n47779), .B(n44859), .Z(n41217) );
  XOR U47193 ( .A(n47780), .B(n47781), .Z(n42028) );
  XNOR U47194 ( .A(n38694), .B(n39228), .Z(n47781) );
  XNOR U47195 ( .A(n47782), .B(n43196), .Z(n39228) );
  XNOR U47196 ( .A(n47783), .B(n47407), .Z(n43196) );
  ANDN U47197 ( .B(n41191), .A(n41976), .Z(n47782) );
  IV U47198 ( .A(n41193), .Z(n41976) );
  XOR U47199 ( .A(n43598), .B(n47784), .Z(n41193) );
  XNOR U47200 ( .A(n47525), .B(n47785), .Z(n43598) );
  XOR U47201 ( .A(n47786), .B(n47787), .Z(n47525) );
  XOR U47202 ( .A(n45116), .B(n45287), .Z(n47787) );
  XOR U47203 ( .A(n47788), .B(n47789), .Z(n45287) );
  NOR U47204 ( .A(n47790), .B(n47791), .Z(n47788) );
  XNOR U47205 ( .A(n47792), .B(n47793), .Z(n45116) );
  NOR U47206 ( .A(n47794), .B(n47795), .Z(n47792) );
  XOR U47207 ( .A(n47385), .B(n47796), .Z(n47786) );
  XOR U47208 ( .A(n47797), .B(n42842), .Z(n47796) );
  XNOR U47209 ( .A(n47798), .B(n47799), .Z(n42842) );
  NOR U47210 ( .A(n47800), .B(n47801), .Z(n47798) );
  XNOR U47211 ( .A(n47802), .B(n47803), .Z(n47385) );
  NOR U47212 ( .A(n47804), .B(n47805), .Z(n47802) );
  XNOR U47213 ( .A(n47806), .B(n42822), .Z(n41191) );
  XNOR U47214 ( .A(n47807), .B(n43194), .Z(n38694) );
  XNOR U47215 ( .A(n47808), .B(n44199), .Z(n43194) );
  IV U47216 ( .A(n47809), .Z(n44199) );
  AND U47217 ( .A(n41205), .B(n41206), .Z(n47807) );
  XOR U47218 ( .A(n47810), .B(n45764), .Z(n41206) );
  IV U47219 ( .A(n44986), .Z(n45764) );
  XNOR U47220 ( .A(n47811), .B(n45011), .Z(n41205) );
  XNOR U47221 ( .A(n39175), .B(n47812), .Z(n47780) );
  XOR U47222 ( .A(n38655), .B(n43183), .Z(n47812) );
  XOR U47223 ( .A(n47813), .B(n43198), .Z(n43183) );
  XOR U47224 ( .A(n47814), .B(n46414), .Z(n43198) );
  ANDN U47225 ( .B(n41195), .A(n41196), .Z(n47813) );
  XNOR U47226 ( .A(n47815), .B(n44173), .Z(n41196) );
  XOR U47227 ( .A(n43665), .B(n47816), .Z(n41195) );
  XNOR U47228 ( .A(n46828), .B(n47817), .Z(n43665) );
  XOR U47229 ( .A(n47818), .B(n47819), .Z(n46828) );
  XNOR U47230 ( .A(n47820), .B(n43828), .Z(n47819) );
  XOR U47231 ( .A(n47821), .B(n47822), .Z(n43828) );
  XOR U47232 ( .A(n47825), .B(n47826), .Z(n47818) );
  XOR U47233 ( .A(n46342), .B(n47392), .Z(n47826) );
  XOR U47234 ( .A(n47827), .B(n47828), .Z(n47392) );
  XNOR U47235 ( .A(n47831), .B(n47832), .Z(n46342) );
  XNOR U47236 ( .A(n47835), .B(n46762), .Z(n38655) );
  XNOR U47237 ( .A(n47836), .B(n43562), .Z(n46762) );
  AND U47238 ( .A(n41201), .B(n41203), .Z(n47835) );
  XNOR U47239 ( .A(n47837), .B(n46735), .Z(n41203) );
  XNOR U47240 ( .A(n47838), .B(n47839), .Z(n46735) );
  XOR U47241 ( .A(n47840), .B(n46282), .Z(n41201) );
  XNOR U47242 ( .A(n47841), .B(n43190), .Z(n39175) );
  XNOR U47243 ( .A(n47842), .B(n44596), .Z(n43190) );
  IV U47244 ( .A(n43863), .Z(n44596) );
  XNOR U47245 ( .A(n47843), .B(n47844), .Z(n43863) );
  AND U47246 ( .A(n42043), .B(n41972), .Z(n47841) );
  XNOR U47247 ( .A(n47845), .B(n44710), .Z(n41972) );
  XOR U47248 ( .A(n47846), .B(n46176), .Z(n42043) );
  XOR U47249 ( .A(n32979), .B(n47847), .Z(n47057) );
  XNOR U47250 ( .A(n33700), .B(n31931), .Z(n47847) );
  XOR U47251 ( .A(n47848), .B(n33760), .Z(n31931) );
  XOR U47252 ( .A(n44802), .B(n35082), .Z(n33760) );
  XOR U47253 ( .A(n40085), .B(n41551), .Z(n35082) );
  XNOR U47254 ( .A(n47849), .B(n47850), .Z(n41551) );
  XOR U47255 ( .A(n39527), .B(n44599), .Z(n47850) );
  XOR U47256 ( .A(n47851), .B(n44351), .Z(n44599) );
  XNOR U47257 ( .A(n47852), .B(n45968), .Z(n44351) );
  XNOR U47258 ( .A(n45717), .B(n46823), .Z(n45968) );
  XNOR U47259 ( .A(n47853), .B(n47854), .Z(n46823) );
  XNOR U47260 ( .A(n46697), .B(n46011), .Z(n47854) );
  XNOR U47261 ( .A(n47855), .B(n47856), .Z(n46011) );
  ANDN U47262 ( .B(n47857), .A(n47500), .Z(n47855) );
  XNOR U47263 ( .A(n47858), .B(n47859), .Z(n46697) );
  ANDN U47264 ( .B(n47860), .A(n47510), .Z(n47858) );
  XOR U47265 ( .A(n46658), .B(n47861), .Z(n47853) );
  XOR U47266 ( .A(n46278), .B(n45387), .Z(n47861) );
  XNOR U47267 ( .A(n47862), .B(n47863), .Z(n45387) );
  ANDN U47268 ( .B(n47864), .A(n47865), .Z(n47862) );
  XNOR U47269 ( .A(n47866), .B(n47867), .Z(n46278) );
  ANDN U47270 ( .B(n47868), .A(n47496), .Z(n47866) );
  XNOR U47271 ( .A(n47869), .B(n47870), .Z(n46658) );
  ANDN U47272 ( .B(n47871), .A(n47506), .Z(n47869) );
  XNOR U47273 ( .A(n47872), .B(n47873), .Z(n45717) );
  XNOR U47274 ( .A(n41741), .B(n47874), .Z(n47873) );
  XOR U47275 ( .A(n47875), .B(n46866), .Z(n41741) );
  IV U47276 ( .A(n47876), .Z(n46866) );
  ANDN U47277 ( .B(n47877), .A(n47016), .Z(n47875) );
  XOR U47278 ( .A(n45318), .B(n47878), .Z(n47872) );
  XOR U47279 ( .A(n43869), .B(n47540), .Z(n47878) );
  XNOR U47280 ( .A(n47879), .B(n47003), .Z(n47540) );
  ANDN U47281 ( .B(n47880), .A(n47010), .Z(n47879) );
  IV U47282 ( .A(n47881), .Z(n47010) );
  XNOR U47283 ( .A(n47882), .B(n46870), .Z(n43869) );
  ANDN U47284 ( .B(n47883), .A(n47691), .Z(n47882) );
  XNOR U47285 ( .A(n47884), .B(n46856), .Z(n45318) );
  ANDN U47286 ( .B(n47885), .A(n47008), .Z(n47884) );
  NOR U47287 ( .A(n41104), .B(n44605), .Z(n47851) );
  XNOR U47288 ( .A(n47886), .B(n43680), .Z(n44605) );
  XOR U47289 ( .A(n47887), .B(n47517), .Z(n43680) );
  XNOR U47290 ( .A(n47888), .B(n47889), .Z(n47517) );
  XNOR U47291 ( .A(n46263), .B(n44462), .Z(n47889) );
  XOR U47292 ( .A(n47890), .B(n47891), .Z(n44462) );
  ANDN U47293 ( .B(n47892), .A(n47893), .Z(n47890) );
  XNOR U47294 ( .A(n47894), .B(n47895), .Z(n46263) );
  NOR U47295 ( .A(n47896), .B(n47897), .Z(n47894) );
  XOR U47296 ( .A(n47898), .B(n47899), .Z(n47888) );
  XOR U47297 ( .A(n45773), .B(n46638), .Z(n47899) );
  XNOR U47298 ( .A(n47900), .B(n47901), .Z(n46638) );
  NOR U47299 ( .A(n47902), .B(n47903), .Z(n47900) );
  XNOR U47300 ( .A(n47904), .B(n47905), .Z(n45773) );
  NOR U47301 ( .A(n47906), .B(n47907), .Z(n47904) );
  XOR U47302 ( .A(n41652), .B(n47908), .Z(n41104) );
  IV U47303 ( .A(n43605), .Z(n41652) );
  XNOR U47304 ( .A(n47909), .B(n46671), .Z(n43605) );
  XOR U47305 ( .A(n47910), .B(n47911), .Z(n46671) );
  XNOR U47306 ( .A(n47912), .B(n45993), .Z(n47911) );
  XOR U47307 ( .A(n47913), .B(n47914), .Z(n45993) );
  AND U47308 ( .A(n47915), .B(n47916), .Z(n47913) );
  XNOR U47309 ( .A(n46218), .B(n47917), .Z(n47910) );
  XOR U47310 ( .A(n45152), .B(n46468), .Z(n47917) );
  XNOR U47311 ( .A(n47918), .B(n47919), .Z(n46468) );
  AND U47312 ( .A(n47822), .B(n47920), .Z(n47918) );
  XNOR U47313 ( .A(n47921), .B(n47922), .Z(n45152) );
  AND U47314 ( .A(n47923), .B(n47924), .Z(n47921) );
  XOR U47315 ( .A(n47925), .B(n47926), .Z(n46218) );
  ANDN U47316 ( .B(n47927), .A(n47832), .Z(n47925) );
  XNOR U47317 ( .A(n47928), .B(n44349), .Z(n39527) );
  XOR U47318 ( .A(n47929), .B(n47930), .Z(n44349) );
  NOR U47319 ( .A(n44804), .B(n41108), .Z(n47928) );
  XNOR U47320 ( .A(n47931), .B(n42325), .Z(n41108) );
  XOR U47321 ( .A(n47458), .B(n47932), .Z(n42325) );
  XOR U47322 ( .A(n47933), .B(n47934), .Z(n47458) );
  XOR U47323 ( .A(n47247), .B(n44219), .Z(n47934) );
  XOR U47324 ( .A(n47935), .B(n47561), .Z(n44219) );
  AND U47325 ( .A(n47936), .B(n47562), .Z(n47935) );
  XNOR U47326 ( .A(n47937), .B(n47566), .Z(n47247) );
  NOR U47327 ( .A(n47565), .B(n47938), .Z(n47937) );
  XOR U47328 ( .A(n46927), .B(n47939), .Z(n47933) );
  XOR U47329 ( .A(n45785), .B(n45745), .Z(n47939) );
  XNOR U47330 ( .A(n47940), .B(n47552), .Z(n45745) );
  XNOR U47331 ( .A(n47942), .B(n47557), .Z(n45785) );
  ANDN U47332 ( .B(n47558), .A(n47943), .Z(n47942) );
  XNOR U47333 ( .A(n47944), .B(n47945), .Z(n46927) );
  XNOR U47334 ( .A(n47948), .B(n44173), .Z(n44804) );
  XOR U47335 ( .A(n43999), .B(n47949), .Z(n47849) );
  XOR U47336 ( .A(n39999), .B(n40966), .Z(n47949) );
  XNOR U47337 ( .A(n47950), .B(n44346), .Z(n40966) );
  XNOR U47338 ( .A(n45889), .B(n46834), .Z(n44346) );
  XOR U47339 ( .A(n47951), .B(n47952), .Z(n46834) );
  ANDN U47340 ( .B(n47953), .A(n47954), .Z(n47951) );
  IV U47341 ( .A(n46164), .Z(n45889) );
  ANDN U47342 ( .B(n44613), .A(n41095), .Z(n47950) );
  XNOR U47343 ( .A(n47955), .B(n44344), .Z(n39999) );
  XOR U47344 ( .A(n44585), .B(n46966), .Z(n44344) );
  XNOR U47345 ( .A(n47956), .B(n47957), .Z(n46966) );
  NOR U47346 ( .A(n47958), .B(n47120), .Z(n47956) );
  IV U47347 ( .A(n45688), .Z(n44585) );
  XOR U47348 ( .A(n47785), .B(n47959), .Z(n45688) );
  XNOR U47349 ( .A(n47960), .B(n47961), .Z(n47785) );
  XOR U47350 ( .A(n44554), .B(n42326), .Z(n47961) );
  XOR U47351 ( .A(n47962), .B(n47121), .Z(n42326) );
  ANDN U47352 ( .B(n47958), .A(n47963), .Z(n47962) );
  XNOR U47353 ( .A(n47964), .B(n47124), .Z(n44554) );
  NOR U47354 ( .A(n46970), .B(n46968), .Z(n47964) );
  XNOR U47355 ( .A(n46251), .B(n47965), .Z(n47960) );
  XOR U47356 ( .A(n47142), .B(n44515), .Z(n47965) );
  XNOR U47357 ( .A(n47966), .B(n47967), .Z(n44515) );
  XNOR U47358 ( .A(n47968), .B(n47116), .Z(n47142) );
  NOR U47359 ( .A(n46960), .B(n46958), .Z(n47968) );
  XNOR U47360 ( .A(n47969), .B(n47970), .Z(n46251) );
  NOR U47361 ( .A(n46964), .B(n46962), .Z(n47969) );
  NOR U47362 ( .A(n44795), .B(n41112), .Z(n47955) );
  XOR U47363 ( .A(n45228), .B(n47971), .Z(n41112) );
  XNOR U47364 ( .A(n47972), .B(n46753), .Z(n45228) );
  XOR U47365 ( .A(n47973), .B(n47974), .Z(n46753) );
  XNOR U47366 ( .A(n47669), .B(n45015), .Z(n47974) );
  XNOR U47367 ( .A(n47975), .B(n47976), .Z(n45015) );
  ANDN U47368 ( .B(n47977), .A(n47978), .Z(n47975) );
  XNOR U47369 ( .A(n47979), .B(n47980), .Z(n47669) );
  ANDN U47370 ( .B(n47981), .A(n47982), .Z(n47979) );
  XOR U47371 ( .A(n47983), .B(n47984), .Z(n47973) );
  XOR U47372 ( .A(n47985), .B(n46227), .Z(n47984) );
  XNOR U47373 ( .A(n47986), .B(n47987), .Z(n46227) );
  NOR U47374 ( .A(n47988), .B(n47989), .Z(n47986) );
  IV U47375 ( .A(n44609), .Z(n44795) );
  XOR U47376 ( .A(n47990), .B(n43716), .Z(n44609) );
  IV U47377 ( .A(n47991), .Z(n43716) );
  XNOR U47378 ( .A(n47992), .B(n44353), .Z(n43999) );
  XOR U47379 ( .A(n43346), .B(n47993), .Z(n44353) );
  XOR U47380 ( .A(n47994), .B(n47995), .Z(n43346) );
  NOR U47381 ( .A(n44808), .B(n41099), .Z(n47992) );
  XNOR U47382 ( .A(n47996), .B(n44816), .Z(n41099) );
  XOR U47383 ( .A(n46543), .B(n47997), .Z(n44816) );
  XNOR U47384 ( .A(n47998), .B(n47999), .Z(n46543) );
  XOR U47385 ( .A(n46554), .B(n47284), .Z(n47999) );
  XOR U47386 ( .A(n48000), .B(n47302), .Z(n47284) );
  AND U47387 ( .A(n47281), .B(n47303), .Z(n48000) );
  XNOR U47388 ( .A(n48001), .B(n47306), .Z(n46554) );
  ANDN U47389 ( .B(n48002), .A(n47305), .Z(n48001) );
  XOR U47390 ( .A(n42218), .B(n48003), .Z(n47998) );
  XOR U47391 ( .A(n46513), .B(n46591), .Z(n48003) );
  XNOR U47392 ( .A(n48004), .B(n47311), .Z(n46591) );
  ANDN U47393 ( .B(n47312), .A(n48005), .Z(n48004) );
  XNOR U47394 ( .A(n48006), .B(n47314), .Z(n46513) );
  ANDN U47395 ( .B(n47315), .A(n47273), .Z(n48006) );
  XOR U47396 ( .A(n48007), .B(n48008), .Z(n42218) );
  ANDN U47397 ( .B(n47268), .A(n48009), .Z(n48007) );
  XOR U47398 ( .A(n44978), .B(n48010), .Z(n44808) );
  IV U47399 ( .A(n45583), .Z(n44978) );
  XOR U47400 ( .A(n48011), .B(n48012), .Z(n45583) );
  XOR U47401 ( .A(n48013), .B(n48014), .Z(n40085) );
  XOR U47402 ( .A(n39335), .B(n35609), .Z(n48014) );
  XNOR U47403 ( .A(n48015), .B(n44628), .Z(n35609) );
  XOR U47404 ( .A(n48016), .B(n47930), .Z(n44628) );
  IV U47405 ( .A(n45656), .Z(n47930) );
  XOR U47406 ( .A(n47467), .B(n48017), .Z(n45656) );
  XOR U47407 ( .A(n48018), .B(n48019), .Z(n47467) );
  XNOR U47408 ( .A(n42658), .B(n45634), .Z(n48019) );
  XNOR U47409 ( .A(n48020), .B(n46144), .Z(n45634) );
  NOR U47410 ( .A(n48021), .B(n48022), .Z(n48020) );
  XOR U47411 ( .A(n48023), .B(n47155), .Z(n42658) );
  NOR U47412 ( .A(n48024), .B(n48025), .Z(n48023) );
  XNOR U47413 ( .A(n44476), .B(n48026), .Z(n48018) );
  XNOR U47414 ( .A(n48027), .B(n44575), .Z(n48026) );
  XNOR U47415 ( .A(n48028), .B(n46138), .Z(n44575) );
  NOR U47416 ( .A(n48029), .B(n48030), .Z(n48028) );
  XOR U47417 ( .A(n48031), .B(n46240), .Z(n44476) );
  NOR U47418 ( .A(n48032), .B(n48033), .Z(n48031) );
  ANDN U47419 ( .B(n44378), .A(n44379), .Z(n48015) );
  XNOR U47420 ( .A(n43577), .B(n47184), .Z(n44379) );
  XNOR U47421 ( .A(n48034), .B(n48035), .Z(n47184) );
  ANDN U47422 ( .B(n48036), .A(n48037), .Z(n48034) );
  XNOR U47423 ( .A(n48038), .B(n48039), .Z(n43577) );
  XOR U47424 ( .A(n43463), .B(n48040), .Z(n44378) );
  XNOR U47425 ( .A(n45436), .B(n47453), .Z(n43463) );
  XOR U47426 ( .A(n48041), .B(n48042), .Z(n47453) );
  XOR U47427 ( .A(n43919), .B(n46537), .Z(n48042) );
  XOR U47428 ( .A(n48043), .B(n47213), .Z(n46537) );
  ANDN U47429 ( .B(n48044), .A(n48045), .Z(n48043) );
  XNOR U47430 ( .A(n48046), .B(n47205), .Z(n43919) );
  ANDN U47431 ( .B(n48047), .A(n48048), .Z(n48046) );
  XOR U47432 ( .A(n47535), .B(n48049), .Z(n48041) );
  XNOR U47433 ( .A(n45175), .B(n44612), .Z(n48049) );
  XNOR U47434 ( .A(n48050), .B(n47200), .Z(n44612) );
  ANDN U47435 ( .B(n48051), .A(n48052), .Z(n48050) );
  XNOR U47436 ( .A(n48053), .B(n48054), .Z(n45175) );
  ANDN U47437 ( .B(n48055), .A(n48056), .Z(n48053) );
  XNOR U47438 ( .A(n48057), .B(n47209), .Z(n47535) );
  ANDN U47439 ( .B(n48058), .A(n48059), .Z(n48057) );
  XOR U47440 ( .A(n48060), .B(n48061), .Z(n45436) );
  XNOR U47441 ( .A(n43340), .B(n44709), .Z(n48061) );
  XNOR U47442 ( .A(n48062), .B(n48063), .Z(n44709) );
  ANDN U47443 ( .B(n48064), .A(n48065), .Z(n48062) );
  XNOR U47444 ( .A(n48066), .B(n48067), .Z(n43340) );
  ANDN U47445 ( .B(n48068), .A(n48069), .Z(n48066) );
  XOR U47446 ( .A(n48070), .B(n48071), .Z(n48060) );
  XOR U47447 ( .A(n47845), .B(n45002), .Z(n48071) );
  XNOR U47448 ( .A(n48072), .B(n48073), .Z(n45002) );
  ANDN U47449 ( .B(n48074), .A(n48075), .Z(n48072) );
  XNOR U47450 ( .A(n48076), .B(n48077), .Z(n47845) );
  ANDN U47451 ( .B(n48078), .A(n48079), .Z(n48076) );
  XNOR U47452 ( .A(n48080), .B(n44632), .Z(n39335) );
  XOR U47453 ( .A(n45778), .B(n47294), .Z(n44632) );
  XNOR U47454 ( .A(n48081), .B(n47366), .Z(n47294) );
  ANDN U47455 ( .B(n48082), .A(n48083), .Z(n48081) );
  ANDN U47456 ( .B(n41301), .A(n44633), .Z(n48080) );
  XOR U47457 ( .A(n48084), .B(n41594), .Z(n44633) );
  IV U47458 ( .A(n44323), .Z(n41594) );
  XOR U47459 ( .A(n47577), .B(n48085), .Z(n44323) );
  XNOR U47460 ( .A(n48086), .B(n48087), .Z(n47577) );
  XOR U47461 ( .A(n48088), .B(n47815), .Z(n48087) );
  XOR U47462 ( .A(n48089), .B(n48090), .Z(n47815) );
  ANDN U47463 ( .B(n48091), .A(n48092), .Z(n48089) );
  XOR U47464 ( .A(n44922), .B(n48093), .Z(n48086) );
  XOR U47465 ( .A(n44172), .B(n47948), .Z(n48093) );
  XNOR U47466 ( .A(n48094), .B(n48095), .Z(n47948) );
  ANDN U47467 ( .B(n48096), .A(n48097), .Z(n48094) );
  XNOR U47468 ( .A(n48098), .B(n48099), .Z(n44172) );
  ANDN U47469 ( .B(n48100), .A(n48101), .Z(n48098) );
  XNOR U47470 ( .A(n48102), .B(n48103), .Z(n44922) );
  ANDN U47471 ( .B(n48104), .A(n48105), .Z(n48102) );
  XOR U47472 ( .A(n48106), .B(n42342), .Z(n41301) );
  IV U47473 ( .A(n45247), .Z(n42342) );
  XNOR U47474 ( .A(n48108), .B(n48109), .Z(n47580) );
  XNOR U47475 ( .A(n48110), .B(n48111), .Z(n48109) );
  XNOR U47476 ( .A(n43723), .B(n48112), .Z(n48108) );
  XOR U47477 ( .A(n45774), .B(n45432), .Z(n48112) );
  XNOR U47478 ( .A(n48113), .B(n48114), .Z(n45432) );
  ANDN U47479 ( .B(n47656), .A(n47657), .Z(n48113) );
  XOR U47480 ( .A(n48115), .B(n48116), .Z(n45774) );
  ANDN U47481 ( .B(n47660), .A(n48117), .Z(n48115) );
  XOR U47482 ( .A(n48118), .B(n48119), .Z(n43723) );
  ANDN U47483 ( .B(n47664), .A(n47666), .Z(n48118) );
  XNOR U47484 ( .A(n41939), .B(n48120), .Z(n48013) );
  XOR U47485 ( .A(n42074), .B(n35092), .Z(n48120) );
  XNOR U47486 ( .A(n48121), .B(n44625), .Z(n35092) );
  XOR U47487 ( .A(n48122), .B(n48123), .Z(n44625) );
  AND U47488 ( .A(n44373), .B(n44358), .Z(n48121) );
  XOR U47489 ( .A(n48124), .B(n44029), .Z(n44358) );
  IV U47490 ( .A(n42461), .Z(n44029) );
  XOR U47491 ( .A(n46732), .B(n46754), .Z(n42461) );
  XNOR U47492 ( .A(n48125), .B(n48126), .Z(n46754) );
  XNOR U47493 ( .A(n48127), .B(n43551), .Z(n48126) );
  XOR U47494 ( .A(n48128), .B(n48129), .Z(n43551) );
  AND U47495 ( .A(n48130), .B(n48131), .Z(n48128) );
  XOR U47496 ( .A(n44537), .B(n48132), .Z(n48125) );
  XOR U47497 ( .A(n43709), .B(n46566), .Z(n48132) );
  XNOR U47498 ( .A(n48133), .B(n48134), .Z(n46566) );
  ANDN U47499 ( .B(n48135), .A(n48136), .Z(n48133) );
  XNOR U47500 ( .A(n48137), .B(n48138), .Z(n43709) );
  ANDN U47501 ( .B(n48139), .A(n48140), .Z(n48137) );
  XOR U47502 ( .A(n48141), .B(n48142), .Z(n44537) );
  ANDN U47503 ( .B(n48143), .A(n48144), .Z(n48141) );
  XOR U47504 ( .A(n48145), .B(n48146), .Z(n46732) );
  XNOR U47505 ( .A(n48147), .B(n43343), .Z(n48146) );
  XOR U47506 ( .A(n48148), .B(n48149), .Z(n43343) );
  ANDN U47507 ( .B(n48150), .A(n48151), .Z(n48148) );
  XNOR U47508 ( .A(n47134), .B(n48152), .Z(n48145) );
  XOR U47509 ( .A(n48153), .B(n47641), .Z(n48152) );
  XNOR U47510 ( .A(n48154), .B(n48155), .Z(n47641) );
  ANDN U47511 ( .B(n48156), .A(n48157), .Z(n48154) );
  XOR U47512 ( .A(n48158), .B(n48159), .Z(n47134) );
  ANDN U47513 ( .B(n48160), .A(n48161), .Z(n48158) );
  XOR U47514 ( .A(n47820), .B(n43829), .Z(n44373) );
  XOR U47515 ( .A(n48162), .B(n47923), .Z(n47820) );
  ANDN U47516 ( .B(n48163), .A(n48164), .Z(n48162) );
  XOR U47517 ( .A(n48165), .B(n44635), .Z(n42074) );
  XNOR U47518 ( .A(n47549), .B(n44479), .Z(n44635) );
  XOR U47519 ( .A(n48167), .B(n48168), .Z(n45451) );
  XOR U47520 ( .A(n45374), .B(n46426), .Z(n48168) );
  XOR U47521 ( .A(n48169), .B(n47626), .Z(n46426) );
  ANDN U47522 ( .B(n48170), .A(n47627), .Z(n48169) );
  XOR U47523 ( .A(n48171), .B(n47623), .Z(n45374) );
  NOR U47524 ( .A(n48172), .B(n47622), .Z(n48171) );
  XOR U47525 ( .A(n44468), .B(n48173), .Z(n48167) );
  XOR U47526 ( .A(n45351), .B(n45762), .Z(n48173) );
  XOR U47527 ( .A(n48174), .B(n47619), .Z(n45762) );
  ANDN U47528 ( .B(n48175), .A(n47618), .Z(n48174) );
  XNOR U47529 ( .A(n48176), .B(n48177), .Z(n45351) );
  NOR U47530 ( .A(n48178), .B(n47613), .Z(n48176) );
  XNOR U47531 ( .A(n48179), .B(n48180), .Z(n44468) );
  NOR U47532 ( .A(n48181), .B(n48182), .Z(n48179) );
  XOR U47533 ( .A(n48183), .B(n48184), .Z(n47549) );
  ANDN U47534 ( .B(n47945), .A(n47947), .Z(n48183) );
  ANDN U47535 ( .B(n44381), .A(n41603), .Z(n48165) );
  XOR U47536 ( .A(n46634), .B(n47674), .Z(n41603) );
  XNOR U47537 ( .A(n48185), .B(n45884), .Z(n46634) );
  ANDN U47538 ( .B(n48186), .A(n48187), .Z(n48185) );
  XOR U47539 ( .A(n48188), .B(n47590), .Z(n44381) );
  XNOR U47540 ( .A(n48189), .B(n48190), .Z(n47590) );
  XOR U47541 ( .A(n48191), .B(n45899), .Z(n41939) );
  XNOR U47542 ( .A(n48192), .B(n43088), .Z(n45899) );
  XOR U47543 ( .A(n48195), .B(n46286), .Z(n44383) );
  XOR U47544 ( .A(n48196), .B(n47263), .Z(n46286) );
  XNOR U47545 ( .A(n48197), .B(n48198), .Z(n47263) );
  XNOR U47546 ( .A(n43650), .B(n46208), .Z(n48198) );
  XOR U47547 ( .A(n48199), .B(n48200), .Z(n46208) );
  NOR U47548 ( .A(n48201), .B(n48202), .Z(n48199) );
  XNOR U47549 ( .A(n48203), .B(n48204), .Z(n43650) );
  NOR U47550 ( .A(n48205), .B(n48206), .Z(n48203) );
  XNOR U47551 ( .A(n46593), .B(n48207), .Z(n48197) );
  XOR U47552 ( .A(n46219), .B(n42518), .Z(n48207) );
  XOR U47553 ( .A(n48208), .B(n48209), .Z(n42518) );
  ANDN U47554 ( .B(n48210), .A(n48211), .Z(n48208) );
  XOR U47555 ( .A(n48212), .B(n48213), .Z(n46219) );
  ANDN U47556 ( .B(n48214), .A(n48215), .Z(n48212) );
  XNOR U47557 ( .A(n48216), .B(n48217), .Z(n46593) );
  ANDN U47558 ( .B(n48218), .A(n48219), .Z(n48216) );
  XNOR U47559 ( .A(n48220), .B(n45853), .Z(n41312) );
  XOR U47560 ( .A(n48221), .B(n44613), .Z(n44802) );
  XOR U47561 ( .A(n48222), .B(n46176), .Z(n44613) );
  XNOR U47562 ( .A(n48223), .B(n48224), .Z(n47126) );
  XNOR U47563 ( .A(n48225), .B(n47161), .Z(n48224) );
  XOR U47564 ( .A(n48226), .B(n48227), .Z(n47161) );
  NOR U47565 ( .A(n48228), .B(n48229), .Z(n48226) );
  XNOR U47566 ( .A(n47685), .B(n48230), .Z(n48223) );
  XOR U47567 ( .A(n44543), .B(n47067), .Z(n48230) );
  XNOR U47568 ( .A(n48231), .B(n48232), .Z(n47067) );
  XOR U47569 ( .A(n48235), .B(n48236), .Z(n44543) );
  ANDN U47570 ( .B(n48237), .A(n48238), .Z(n48235) );
  XOR U47571 ( .A(n48239), .B(n48240), .Z(n47685) );
  ANDN U47572 ( .B(n48241), .A(n48242), .Z(n48239) );
  ANDN U47573 ( .B(n41095), .A(n41096), .Z(n48221) );
  XOR U47574 ( .A(n48244), .B(n43562), .Z(n41096) );
  XOR U47575 ( .A(n45450), .B(n48245), .Z(n43562) );
  XOR U47576 ( .A(n48246), .B(n48247), .Z(n45450) );
  XOR U47577 ( .A(n44205), .B(n48248), .Z(n48247) );
  XNOR U47578 ( .A(n48249), .B(n48250), .Z(n44205) );
  ANDN U47579 ( .B(n48251), .A(n48252), .Z(n48249) );
  XNOR U47580 ( .A(n43824), .B(n48253), .Z(n48246) );
  XOR U47581 ( .A(n44587), .B(n48254), .Z(n48253) );
  XOR U47582 ( .A(n48255), .B(n48256), .Z(n44587) );
  AND U47583 ( .A(n48257), .B(n48258), .Z(n48255) );
  XNOR U47584 ( .A(n48259), .B(n48260), .Z(n43824) );
  AND U47585 ( .A(n48261), .B(n48262), .Z(n48259) );
  XNOR U47586 ( .A(n48263), .B(n45260), .Z(n41095) );
  XOR U47587 ( .A(n48264), .B(n48265), .Z(n45260) );
  AND U47588 ( .A(n33761), .B(n35654), .Z(n47848) );
  XNOR U47589 ( .A(n41127), .B(n39344), .Z(n35654) );
  IV U47590 ( .A(n38253), .Z(n39344) );
  XOR U47591 ( .A(n43041), .B(n43619), .Z(n38253) );
  XNOR U47592 ( .A(n48266), .B(n48267), .Z(n43619) );
  XNOR U47593 ( .A(n37685), .B(n42574), .Z(n48267) );
  XNOR U47594 ( .A(n48268), .B(n42583), .Z(n42574) );
  XNOR U47595 ( .A(n48269), .B(n44856), .Z(n42583) );
  IV U47596 ( .A(n44921), .Z(n44856) );
  XOR U47597 ( .A(n46126), .B(n48270), .Z(n44921) );
  XOR U47598 ( .A(n48271), .B(n48272), .Z(n46126) );
  XOR U47599 ( .A(n44159), .B(n48273), .Z(n48272) );
  XNOR U47600 ( .A(n48274), .B(n48215), .Z(n44159) );
  AND U47601 ( .A(n48275), .B(n48276), .Z(n48274) );
  XOR U47602 ( .A(n43924), .B(n48277), .Z(n48271) );
  XNOR U47603 ( .A(n48278), .B(n44197), .Z(n48277) );
  XOR U47604 ( .A(n48279), .B(n48219), .Z(n44197) );
  ANDN U47605 ( .B(n48280), .A(n48281), .Z(n48279) );
  XNOR U47606 ( .A(n48282), .B(n48202), .Z(n43924) );
  AND U47607 ( .A(n48283), .B(n48284), .Z(n48282) );
  ANDN U47608 ( .B(n40259), .A(n40260), .Z(n48268) );
  XNOR U47609 ( .A(n42312), .B(n48285), .Z(n40260) );
  IV U47610 ( .A(n46103), .Z(n42312) );
  XNOR U47611 ( .A(n48286), .B(n43644), .Z(n40259) );
  XOR U47612 ( .A(n47909), .B(n48287), .Z(n43644) );
  XOR U47613 ( .A(n48288), .B(n48289), .Z(n47909) );
  XOR U47614 ( .A(n45854), .B(n48290), .Z(n48289) );
  XNOR U47615 ( .A(n48291), .B(n48292), .Z(n45854) );
  XOR U47616 ( .A(n47469), .B(n48295), .Z(n48288) );
  XOR U47617 ( .A(n45496), .B(n48296), .Z(n48295) );
  XNOR U47618 ( .A(n48297), .B(n48298), .Z(n45496) );
  ANDN U47619 ( .B(n48299), .A(n48300), .Z(n48297) );
  XOR U47620 ( .A(n48301), .B(n48302), .Z(n47469) );
  NOR U47621 ( .A(n48303), .B(n48304), .Z(n48301) );
  XNOR U47622 ( .A(n48305), .B(n42580), .Z(n37685) );
  XOR U47623 ( .A(n45626), .B(n48306), .Z(n42580) );
  IV U47624 ( .A(n45303), .Z(n45626) );
  XNOR U47625 ( .A(n48307), .B(n48308), .Z(n45303) );
  ANDN U47626 ( .B(n41496), .A(n41498), .Z(n48305) );
  XOR U47627 ( .A(n48309), .B(n46059), .Z(n41498) );
  IV U47628 ( .A(n45216), .Z(n46059) );
  XNOR U47629 ( .A(n48310), .B(n48311), .Z(n45216) );
  XOR U47630 ( .A(n47744), .B(n46054), .Z(n41496) );
  XOR U47631 ( .A(n48312), .B(n48313), .Z(n47744) );
  AND U47632 ( .A(n48314), .B(n48315), .Z(n48312) );
  XNOR U47633 ( .A(n37702), .B(n48316), .Z(n48266) );
  XOR U47634 ( .A(n36512), .B(n38922), .Z(n48316) );
  XOR U47635 ( .A(n48317), .B(n42589), .Z(n38922) );
  XOR U47636 ( .A(n48318), .B(n47407), .Z(n42589) );
  ANDN U47637 ( .B(n42590), .A(n43052), .Z(n48317) );
  XOR U47638 ( .A(n45310), .B(n48319), .Z(n43052) );
  IV U47639 ( .A(n44223), .Z(n45310) );
  XOR U47640 ( .A(n48321), .B(n48322), .Z(n47236) );
  XOR U47641 ( .A(n48323), .B(n47446), .Z(n48322) );
  XOR U47642 ( .A(n48324), .B(n46786), .Z(n47446) );
  ANDN U47643 ( .B(n48325), .A(n48326), .Z(n48324) );
  XOR U47644 ( .A(n44200), .B(n48327), .Z(n48321) );
  XOR U47645 ( .A(n45419), .B(n47318), .Z(n48327) );
  XNOR U47646 ( .A(n48328), .B(n46779), .Z(n47318) );
  ANDN U47647 ( .B(n48329), .A(n48330), .Z(n48328) );
  XNOR U47648 ( .A(n48331), .B(n48332), .Z(n45419) );
  ANDN U47649 ( .B(n48333), .A(n48334), .Z(n48331) );
  XNOR U47650 ( .A(n48335), .B(n48336), .Z(n44200) );
  ANDN U47651 ( .B(n48337), .A(n48338), .Z(n48335) );
  XOR U47652 ( .A(n48339), .B(n45127), .Z(n42590) );
  XNOR U47653 ( .A(n48340), .B(n42816), .Z(n36512) );
  XOR U47654 ( .A(n43815), .B(n47113), .Z(n42816) );
  XOR U47655 ( .A(n48341), .B(n46974), .Z(n47113) );
  ANDN U47656 ( .B(n48342), .A(n47967), .Z(n48341) );
  ANDN U47657 ( .B(n40255), .A(n40256), .Z(n48340) );
  XOR U47658 ( .A(n48343), .B(n47603), .Z(n40256) );
  XOR U47659 ( .A(n44935), .B(n47372), .Z(n40255) );
  XOR U47660 ( .A(n48344), .B(n48345), .Z(n47372) );
  ANDN U47661 ( .B(n48346), .A(n48347), .Z(n48344) );
  XOR U47662 ( .A(n48348), .B(n48349), .Z(n44935) );
  XNOR U47663 ( .A(n48350), .B(n46004), .Z(n37702) );
  XOR U47664 ( .A(n48351), .B(n44106), .Z(n46004) );
  XNOR U47665 ( .A(n46945), .B(n48352), .Z(n44106) );
  XOR U47666 ( .A(n48353), .B(n48354), .Z(n46945) );
  XOR U47667 ( .A(n46803), .B(n44335), .Z(n48354) );
  XOR U47668 ( .A(n48355), .B(n46482), .Z(n44335) );
  XOR U47669 ( .A(round_reg[1578]), .B(n48356), .Z(n46482) );
  ANDN U47670 ( .B(n46813), .A(n48357), .Z(n48355) );
  XNOR U47671 ( .A(n48358), .B(n46809), .Z(n46803) );
  ANDN U47672 ( .B(n46810), .A(n48359), .Z(n48358) );
  XOR U47673 ( .A(n45671), .B(n48360), .Z(n48353) );
  XOR U47674 ( .A(n44483), .B(n45383), .Z(n48360) );
  XNOR U47675 ( .A(n48361), .B(n46489), .Z(n45383) );
  XOR U47676 ( .A(round_reg[1295]), .B(n48362), .Z(n46489) );
  ANDN U47677 ( .B(n46816), .A(n48363), .Z(n48361) );
  XNOR U47678 ( .A(n48364), .B(n46485), .Z(n44483) );
  XOR U47679 ( .A(round_reg[1452]), .B(n48365), .Z(n46485) );
  ANDN U47680 ( .B(n46820), .A(n48366), .Z(n48364) );
  XNOR U47681 ( .A(n48367), .B(n46476), .Z(n45671) );
  XNOR U47682 ( .A(round_reg[1513]), .B(n48368), .Z(n46476) );
  NOR U47683 ( .A(n46818), .B(n48369), .Z(n48367) );
  ANDN U47684 ( .B(n40263), .A(n40265), .Z(n48350) );
  XOR U47685 ( .A(n48370), .B(n46178), .Z(n40265) );
  XOR U47686 ( .A(n47994), .B(n45727), .Z(n46178) );
  XOR U47687 ( .A(n48371), .B(n48372), .Z(n45727) );
  XOR U47688 ( .A(n47523), .B(n45568), .Z(n48372) );
  XOR U47689 ( .A(n48373), .B(n48374), .Z(n45568) );
  ANDN U47690 ( .B(n48375), .A(n46907), .Z(n48373) );
  XNOR U47691 ( .A(n48376), .B(n48377), .Z(n47523) );
  ANDN U47692 ( .B(n48378), .A(n46897), .Z(n48376) );
  XOR U47693 ( .A(n48379), .B(n48380), .Z(n48371) );
  XOR U47694 ( .A(n48381), .B(n46756), .Z(n48380) );
  XNOR U47695 ( .A(n48382), .B(n48383), .Z(n46756) );
  ANDN U47696 ( .B(n48384), .A(n46903), .Z(n48382) );
  XOR U47697 ( .A(n48385), .B(n48386), .Z(n47994) );
  XNOR U47698 ( .A(n48387), .B(n48388), .Z(n48386) );
  XOR U47699 ( .A(n46826), .B(n48389), .Z(n48385) );
  XOR U47700 ( .A(n46500), .B(n46184), .Z(n48389) );
  XNOR U47701 ( .A(n48390), .B(n47055), .Z(n46184) );
  ANDN U47702 ( .B(n48391), .A(n48392), .Z(n48390) );
  XNOR U47703 ( .A(n48393), .B(n48394), .Z(n46500) );
  ANDN U47704 ( .B(n48395), .A(n48396), .Z(n48393) );
  XNOR U47705 ( .A(n48397), .B(n47051), .Z(n46826) );
  NOR U47706 ( .A(n48398), .B(n48399), .Z(n48397) );
  XOR U47707 ( .A(n48400), .B(n48401), .Z(n40263) );
  XOR U47708 ( .A(n48402), .B(n48403), .Z(n43041) );
  XNOR U47709 ( .A(n35523), .B(n40970), .Z(n48403) );
  XNOR U47710 ( .A(n48404), .B(n42271), .Z(n40970) );
  XNOR U47711 ( .A(n41749), .B(n48405), .Z(n42271) );
  IV U47712 ( .A(n44579), .Z(n41749) );
  XOR U47713 ( .A(n48406), .B(n46799), .Z(n44579) );
  XNOR U47714 ( .A(n48407), .B(n48408), .Z(n46799) );
  XOR U47715 ( .A(n46430), .B(n44799), .Z(n48408) );
  XOR U47716 ( .A(n48409), .B(n48410), .Z(n44799) );
  ANDN U47717 ( .B(n48411), .A(n48412), .Z(n48409) );
  XNOR U47718 ( .A(n48413), .B(n48414), .Z(n46430) );
  ANDN U47719 ( .B(n48415), .A(n48416), .Z(n48413) );
  XOR U47720 ( .A(n48417), .B(n48418), .Z(n48407) );
  XOR U47721 ( .A(n44466), .B(n47404), .Z(n48418) );
  XNOR U47722 ( .A(n48419), .B(n48420), .Z(n47404) );
  NOR U47723 ( .A(n48421), .B(n48422), .Z(n48419) );
  XNOR U47724 ( .A(n48423), .B(n48424), .Z(n44466) );
  NOR U47725 ( .A(n48425), .B(n48426), .Z(n48423) );
  NOR U47726 ( .A(n41124), .B(n41125), .Z(n48404) );
  XOR U47727 ( .A(n48427), .B(n45519), .Z(n41125) );
  XNOR U47728 ( .A(n48088), .B(n44173), .Z(n41124) );
  XNOR U47729 ( .A(n48430), .B(n48431), .Z(n48088) );
  ANDN U47730 ( .B(n48432), .A(n48433), .Z(n48430) );
  XNOR U47731 ( .A(n48434), .B(n42274), .Z(n35523) );
  XOR U47732 ( .A(n48435), .B(n48436), .Z(n42274) );
  ANDN U47733 ( .B(n42275), .A(n43061), .Z(n48434) );
  XOR U47734 ( .A(n47797), .B(n45117), .Z(n43061) );
  IV U47735 ( .A(n42843), .Z(n45117) );
  XOR U47736 ( .A(n47144), .B(n48437), .Z(n42843) );
  XNOR U47737 ( .A(n48438), .B(n48439), .Z(n47144) );
  XOR U47738 ( .A(n47026), .B(n42653), .Z(n48439) );
  XOR U47739 ( .A(n48440), .B(n47122), .Z(n42653) );
  NOR U47740 ( .A(n47957), .B(n47121), .Z(n48440) );
  XOR U47741 ( .A(round_reg[1048]), .B(n48441), .Z(n47121) );
  IV U47742 ( .A(n47963), .Z(n47957) );
  XOR U47743 ( .A(round_reg[680]), .B(n48442), .Z(n47963) );
  XNOR U47744 ( .A(n48443), .B(n48444), .Z(n47026) );
  ANDN U47745 ( .B(n46962), .A(n47970), .Z(n48443) );
  XOR U47746 ( .A(n46600), .B(n48446), .Z(n48438) );
  XOR U47747 ( .A(n46715), .B(n47110), .Z(n48446) );
  XNOR U47748 ( .A(n4549), .B(n48448), .Z(n48447) );
  XOR U47749 ( .A(round_reg[1187]), .B(n48450), .Z(n47116) );
  XNOR U47750 ( .A(n48451), .B(n48342), .Z(n46715) );
  XOR U47751 ( .A(round_reg[1259]), .B(n48452), .Z(n47967) );
  XNOR U47752 ( .A(n48454), .B(n47125), .Z(n46600) );
  ANDN U47753 ( .B(n46968), .A(n47124), .Z(n48454) );
  XNOR U47754 ( .A(round_reg[1019]), .B(n48455), .Z(n47124) );
  XNOR U47755 ( .A(round_reg[908]), .B(n48456), .Z(n46968) );
  XNOR U47756 ( .A(n48457), .B(n48458), .Z(n47797) );
  NOR U47757 ( .A(n48459), .B(n48460), .Z(n48457) );
  XOR U47758 ( .A(n45781), .B(n47483), .Z(n42275) );
  XNOR U47759 ( .A(n48461), .B(n48462), .Z(n47483) );
  XNOR U47760 ( .A(n38521), .B(n48465), .Z(n48402) );
  XOR U47761 ( .A(n38539), .B(n40646), .Z(n48465) );
  XNOR U47762 ( .A(n48466), .B(n42267), .Z(n40646) );
  XOR U47763 ( .A(n46572), .B(n48467), .Z(n42267) );
  IV U47764 ( .A(n42860), .Z(n46572) );
  XOR U47765 ( .A(n48468), .B(n48469), .Z(n42860) );
  ANDN U47766 ( .B(n41136), .A(n42268), .Z(n48466) );
  XOR U47767 ( .A(n48225), .B(n44544), .Z(n42268) );
  IV U47768 ( .A(n47162), .Z(n44544) );
  XNOR U47769 ( .A(n48470), .B(n47516), .Z(n47162) );
  XNOR U47770 ( .A(n48471), .B(n48472), .Z(n47516) );
  XOR U47771 ( .A(n48473), .B(n47032), .Z(n48472) );
  XOR U47772 ( .A(n48474), .B(n48475), .Z(n47032) );
  NOR U47773 ( .A(n48476), .B(n48477), .Z(n48474) );
  XNOR U47774 ( .A(n48478), .B(n48479), .Z(n48471) );
  XOR U47775 ( .A(n45860), .B(n46737), .Z(n48479) );
  XNOR U47776 ( .A(n48480), .B(n48481), .Z(n46737) );
  ANDN U47777 ( .B(n48482), .A(n48483), .Z(n48480) );
  XNOR U47778 ( .A(n48484), .B(n48485), .Z(n45860) );
  ANDN U47779 ( .B(n48486), .A(n48487), .Z(n48484) );
  XOR U47780 ( .A(n48488), .B(n48489), .Z(n48225) );
  AND U47781 ( .A(n48490), .B(n48491), .Z(n48488) );
  XOR U47782 ( .A(n48492), .B(n43565), .Z(n41136) );
  XOR U47783 ( .A(n48493), .B(n48494), .Z(n43565) );
  XOR U47784 ( .A(n48495), .B(n42260), .Z(n38539) );
  XOR U47785 ( .A(n46041), .B(n44619), .Z(n42260) );
  XNOR U47786 ( .A(n48496), .B(n48497), .Z(n46041) );
  ANDN U47787 ( .B(n48498), .A(n48499), .Z(n48496) );
  ANDN U47788 ( .B(n42259), .A(n44148), .Z(n48495) );
  XNOR U47789 ( .A(n48500), .B(n42263), .Z(n38521) );
  XNOR U47790 ( .A(n48501), .B(n48502), .Z(n47331) );
  NOR U47791 ( .A(n47351), .B(n47352), .Z(n48501) );
  ANDN U47792 ( .B(n41130), .A(n41132), .Z(n48500) );
  XOR U47793 ( .A(n48503), .B(n47678), .Z(n41132) );
  XNOR U47794 ( .A(n48504), .B(n44528), .Z(n41130) );
  XOR U47795 ( .A(n48307), .B(n47683), .Z(n44528) );
  XNOR U47796 ( .A(n48505), .B(n48506), .Z(n47683) );
  XOR U47797 ( .A(n43705), .B(n46190), .Z(n48506) );
  XOR U47798 ( .A(n48507), .B(n46334), .Z(n46190) );
  XNOR U47799 ( .A(round_reg[407]), .B(n48508), .Z(n46334) );
  AND U47800 ( .A(n48509), .B(n46335), .Z(n48507) );
  XOR U47801 ( .A(n48510), .B(n46329), .Z(n43705) );
  ANDN U47802 ( .B(n48511), .A(n46328), .Z(n48510) );
  XOR U47803 ( .A(n44399), .B(n48512), .Z(n48505) );
  XOR U47804 ( .A(n43279), .B(n45825), .Z(n48512) );
  XNOR U47805 ( .A(n48513), .B(n46324), .Z(n45825) );
  XOR U47806 ( .A(round_reg[579]), .B(n48514), .Z(n46324) );
  XNOR U47807 ( .A(n48516), .B(n46338), .Z(n43279) );
  XNOR U47808 ( .A(round_reg[477]), .B(n48517), .Z(n46338) );
  ANDN U47809 ( .B(n46339), .A(n48518), .Z(n48516) );
  XNOR U47810 ( .A(n48519), .B(n47352), .Z(n44399) );
  XOR U47811 ( .A(round_reg[575]), .B(n48520), .Z(n47352) );
  XOR U47812 ( .A(n48522), .B(n48523), .Z(n48307) );
  XNOR U47813 ( .A(n45643), .B(n46257), .Z(n48523) );
  XOR U47814 ( .A(n48524), .B(n48525), .Z(n46257) );
  NOR U47815 ( .A(n48526), .B(n48527), .Z(n48524) );
  XNOR U47816 ( .A(n48528), .B(n48529), .Z(n45643) );
  XOR U47817 ( .A(n45942), .B(n48532), .Z(n48522) );
  XOR U47818 ( .A(n46318), .B(n42851), .Z(n48532) );
  XOR U47819 ( .A(n48533), .B(n48534), .Z(n42851) );
  XNOR U47820 ( .A(n48537), .B(n48538), .Z(n46318) );
  NOR U47821 ( .A(n48539), .B(n48540), .Z(n48537) );
  XNOR U47822 ( .A(n48541), .B(n48542), .Z(n45942) );
  XOR U47823 ( .A(n48545), .B(n42259), .Z(n41127) );
  XNOR U47824 ( .A(n48546), .B(n47809), .Z(n42259) );
  ANDN U47825 ( .B(n44148), .A(n45096), .Z(n48545) );
  IV U47826 ( .A(n44149), .Z(n45096) );
  XOR U47827 ( .A(n48547), .B(n44839), .Z(n44149) );
  IV U47828 ( .A(n48548), .Z(n44839) );
  XOR U47829 ( .A(n46384), .B(n46014), .Z(n44148) );
  XOR U47830 ( .A(n48549), .B(n47682), .Z(n46014) );
  XNOR U47831 ( .A(n48550), .B(n48551), .Z(n47682) );
  XNOR U47832 ( .A(n45280), .B(n47074), .Z(n48551) );
  XNOR U47833 ( .A(n48552), .B(n47089), .Z(n47074) );
  XOR U47834 ( .A(round_reg[1359]), .B(n48553), .Z(n47089) );
  AND U47835 ( .A(n46376), .B(n46375), .Z(n48552) );
  XOR U47836 ( .A(round_reg[983]), .B(n48554), .Z(n46375) );
  XNOR U47837 ( .A(n48555), .B(n47079), .Z(n45280) );
  XOR U47838 ( .A(round_reg[1579]), .B(n48452), .Z(n47079) );
  ANDN U47839 ( .B(n46379), .A(n46380), .Z(n48555) );
  XOR U47840 ( .A(round_reg[1215]), .B(n48520), .Z(n46379) );
  XOR U47841 ( .A(n45624), .B(n48556), .Z(n48550) );
  XNOR U47842 ( .A(n45770), .B(n41734), .Z(n48556) );
  XOR U47843 ( .A(n48557), .B(n47086), .Z(n41734) );
  XOR U47844 ( .A(round_reg[1453]), .B(n48558), .Z(n47086) );
  ANDN U47845 ( .B(n46386), .A(n46387), .Z(n48557) );
  XNOR U47846 ( .A(round_reg[1076]), .B(n48559), .Z(n46386) );
  XNOR U47847 ( .A(n48560), .B(n47092), .Z(n45770) );
  XOR U47848 ( .A(round_reg[1296]), .B(n48561), .Z(n47092) );
  ANDN U47849 ( .B(n47093), .A(n48562), .Z(n48560) );
  XNOR U47850 ( .A(n48563), .B(n47082), .Z(n45624) );
  XOR U47851 ( .A(round_reg[1514]), .B(n48564), .Z(n47082) );
  ANDN U47852 ( .B(n46686), .A(n48565), .Z(n48563) );
  XNOR U47853 ( .A(round_reg[1125]), .B(n48566), .Z(n46686) );
  XNOR U47854 ( .A(n48567), .B(n47093), .Z(n46384) );
  XOR U47855 ( .A(round_reg[1223]), .B(n48568), .Z(n47093) );
  XNOR U47856 ( .A(n47436), .B(n39475), .Z(n33761) );
  IV U47857 ( .A(n38277), .Z(n39475) );
  XOR U47858 ( .A(n41569), .B(n39985), .Z(n38277) );
  XNOR U47859 ( .A(n48569), .B(n48570), .Z(n39985) );
  XOR U47860 ( .A(n37967), .B(n38515), .Z(n48570) );
  XOR U47861 ( .A(n48571), .B(n48572), .Z(n38515) );
  AND U47862 ( .A(n43258), .B(n43257), .Z(n48571) );
  XOR U47863 ( .A(n48573), .B(n44841), .Z(n43258) );
  XOR U47864 ( .A(n48574), .B(n47356), .Z(n44841) );
  XNOR U47865 ( .A(n48575), .B(n48576), .Z(n47356) );
  XOR U47866 ( .A(n46081), .B(n46058), .Z(n48576) );
  XOR U47867 ( .A(n48577), .B(n48578), .Z(n46058) );
  ANDN U47868 ( .B(n48579), .A(n48580), .Z(n48577) );
  XNOR U47869 ( .A(n48581), .B(n48582), .Z(n46081) );
  ANDN U47870 ( .B(n48583), .A(n48584), .Z(n48581) );
  XNOR U47871 ( .A(n48309), .B(n48585), .Z(n48575) );
  XNOR U47872 ( .A(n45756), .B(n45215), .Z(n48585) );
  XOR U47873 ( .A(n48586), .B(n48587), .Z(n45215) );
  ANDN U47874 ( .B(n48588), .A(n48589), .Z(n48586) );
  XNOR U47875 ( .A(n48590), .B(n48591), .Z(n45756) );
  ANDN U47876 ( .B(n48592), .A(n48593), .Z(n48590) );
  XOR U47877 ( .A(n48594), .B(n48595), .Z(n48309) );
  ANDN U47878 ( .B(n48596), .A(n48597), .Z(n48594) );
  XNOR U47879 ( .A(n48598), .B(n41362), .Z(n37967) );
  ANDN U47880 ( .B(n41363), .A(n43266), .Z(n48598) );
  XOR U47881 ( .A(n48599), .B(n42160), .Z(n43266) );
  IV U47882 ( .A(n48600), .Z(n42160) );
  XOR U47883 ( .A(n43576), .B(n48601), .Z(n41363) );
  XOR U47884 ( .A(n48602), .B(n47029), .Z(n43576) );
  XNOR U47885 ( .A(n48603), .B(n48604), .Z(n47029) );
  XNOR U47886 ( .A(n47929), .B(n45718), .Z(n48604) );
  XOR U47887 ( .A(n48605), .B(n48606), .Z(n45718) );
  ANDN U47888 ( .B(n48607), .A(n47432), .Z(n48605) );
  XNOR U47889 ( .A(n48608), .B(n48609), .Z(n47929) );
  ANDN U47890 ( .B(n48610), .A(n48611), .Z(n48608) );
  XOR U47891 ( .A(n46296), .B(n48612), .Z(n48603) );
  XOR U47892 ( .A(n45655), .B(n48016), .Z(n48612) );
  XNOR U47893 ( .A(n48613), .B(n48614), .Z(n48016) );
  ANDN U47894 ( .B(n48615), .A(n47424), .Z(n48613) );
  XNOR U47895 ( .A(n48616), .B(n48617), .Z(n45655) );
  ANDN U47896 ( .B(n48618), .A(n47428), .Z(n48616) );
  XNOR U47897 ( .A(n48619), .B(n48620), .Z(n46296) );
  ANDN U47898 ( .B(n48621), .A(n47419), .Z(n48619) );
  XOR U47899 ( .A(n37057), .B(n48622), .Z(n48569) );
  XOR U47900 ( .A(n36938), .B(n40973), .Z(n48622) );
  XNOR U47901 ( .A(n48623), .B(n40980), .Z(n40973) );
  ANDN U47902 ( .B(n40981), .A(n44992), .Z(n48623) );
  XNOR U47903 ( .A(n42667), .B(n48624), .Z(n44992) );
  XNOR U47904 ( .A(n47843), .B(n47959), .Z(n42667) );
  XNOR U47905 ( .A(n48625), .B(n48626), .Z(n47959) );
  XNOR U47906 ( .A(n44930), .B(n43770), .Z(n48626) );
  XOR U47907 ( .A(n48627), .B(n48229), .Z(n43770) );
  ANDN U47908 ( .B(n48628), .A(n48629), .Z(n48627) );
  XOR U47909 ( .A(n48630), .B(n48242), .Z(n44930) );
  IV U47910 ( .A(n48631), .Z(n48242) );
  AND U47911 ( .A(n48632), .B(n48633), .Z(n48630) );
  XNOR U47912 ( .A(n44331), .B(n48634), .Z(n48625) );
  XOR U47913 ( .A(n45163), .B(n48635), .Z(n48634) );
  XOR U47914 ( .A(n48636), .B(n48238), .Z(n45163) );
  IV U47915 ( .A(n48637), .Z(n48238) );
  ANDN U47916 ( .B(n48638), .A(n48639), .Z(n48636) );
  XNOR U47917 ( .A(n48640), .B(n48233), .Z(n44331) );
  ANDN U47918 ( .B(n48641), .A(n48642), .Z(n48640) );
  XOR U47919 ( .A(n48643), .B(n48644), .Z(n47843) );
  XOR U47920 ( .A(n42222), .B(n48645), .Z(n48644) );
  XNOR U47921 ( .A(n48646), .B(n48647), .Z(n42222) );
  AND U47922 ( .A(n48481), .B(n48648), .Z(n48646) );
  XOR U47923 ( .A(n46394), .B(n48649), .Z(n48643) );
  XNOR U47924 ( .A(n46653), .B(n46885), .Z(n48649) );
  XNOR U47925 ( .A(n48650), .B(n48651), .Z(n46885) );
  AND U47926 ( .A(n48485), .B(n48652), .Z(n48650) );
  XNOR U47927 ( .A(n48653), .B(n48654), .Z(n46653) );
  ANDN U47928 ( .B(n48655), .A(n48656), .Z(n48653) );
  XNOR U47929 ( .A(n48657), .B(n48658), .Z(n46394) );
  AND U47930 ( .A(n48475), .B(n48659), .Z(n48657) );
  XNOR U47931 ( .A(n48273), .B(n43925), .Z(n40981) );
  XOR U47932 ( .A(n48660), .B(n48206), .Z(n48273) );
  ANDN U47933 ( .B(n48661), .A(n48662), .Z(n48660) );
  XNOR U47934 ( .A(n48663), .B(n40990), .Z(n36938) );
  ANDN U47935 ( .B(n43269), .A(n43268), .Z(n48663) );
  XOR U47936 ( .A(n48664), .B(n45011), .Z(n43268) );
  XOR U47937 ( .A(n46726), .B(n48665), .Z(n45011) );
  XNOR U47938 ( .A(n48666), .B(n48667), .Z(n46726) );
  XOR U47939 ( .A(n45518), .B(n46931), .Z(n48667) );
  XOR U47940 ( .A(n48668), .B(n48669), .Z(n46931) );
  ANDN U47941 ( .B(n48670), .A(n48671), .Z(n48668) );
  XNOR U47942 ( .A(n48672), .B(n48673), .Z(n45518) );
  ANDN U47943 ( .B(n48674), .A(n48675), .Z(n48672) );
  XOR U47944 ( .A(n47379), .B(n48676), .Z(n48666) );
  XOR U47945 ( .A(n48677), .B(n48427), .Z(n48676) );
  XNOR U47946 ( .A(n48678), .B(n48679), .Z(n48427) );
  ANDN U47947 ( .B(n48680), .A(n48681), .Z(n48678) );
  XNOR U47948 ( .A(n48682), .B(n48683), .Z(n47379) );
  ANDN U47949 ( .B(n48684), .A(n48685), .Z(n48682) );
  XOR U47950 ( .A(n48290), .B(n45497), .Z(n43269) );
  XNOR U47951 ( .A(n48686), .B(n48687), .Z(n48290) );
  ANDN U47952 ( .B(n48688), .A(n48689), .Z(n48686) );
  XNOR U47953 ( .A(n48690), .B(n40987), .Z(n37057) );
  ANDN U47954 ( .B(n43254), .A(n40986), .Z(n48690) );
  XNOR U47955 ( .A(n48478), .B(n47033), .Z(n40986) );
  IV U47956 ( .A(n45861), .Z(n47033) );
  XNOR U47957 ( .A(n48691), .B(n48655), .Z(n48478) );
  NOR U47958 ( .A(n48692), .B(n48693), .Z(n48691) );
  XOR U47959 ( .A(n48070), .B(n43341), .Z(n43254) );
  IV U47960 ( .A(n44710), .Z(n43341) );
  XOR U47961 ( .A(n47536), .B(n48694), .Z(n44710) );
  XOR U47962 ( .A(n48695), .B(n48696), .Z(n47536) );
  XNOR U47963 ( .A(n41875), .B(n45438), .Z(n48696) );
  XNOR U47964 ( .A(n48697), .B(n47199), .Z(n45438) );
  IV U47965 ( .A(n48698), .Z(n47199) );
  ANDN U47966 ( .B(n47200), .A(n48051), .Z(n48697) );
  XNOR U47967 ( .A(round_reg[1288]), .B(n48699), .Z(n47200) );
  XOR U47968 ( .A(n48700), .B(n47204), .Z(n41875) );
  AND U47969 ( .A(n48048), .B(n47205), .Z(n48700) );
  XNOR U47970 ( .A(round_reg[1571]), .B(n48701), .Z(n47205) );
  XNOR U47971 ( .A(n45850), .B(n48702), .Z(n48695) );
  XNOR U47972 ( .A(n45578), .B(n47173), .Z(n48702) );
  XNOR U47973 ( .A(n48703), .B(n48704), .Z(n47173) );
  ANDN U47974 ( .B(n48056), .A(n48054), .Z(n48703) );
  XNOR U47975 ( .A(n48705), .B(n47212), .Z(n45578) );
  ANDN U47976 ( .B(n47213), .A(n48044), .Z(n48705) );
  XNOR U47977 ( .A(round_reg[1351]), .B(n48706), .Z(n47213) );
  XNOR U47978 ( .A(n48707), .B(n47208), .Z(n45850) );
  AND U47979 ( .A(n48059), .B(n47209), .Z(n48707) );
  XNOR U47980 ( .A(round_reg[1506]), .B(n48708), .Z(n47209) );
  XNOR U47981 ( .A(n48709), .B(n48710), .Z(n48070) );
  ANDN U47982 ( .B(n48711), .A(n48712), .Z(n48709) );
  XOR U47983 ( .A(n48713), .B(n48714), .Z(n41569) );
  XOR U47984 ( .A(n39595), .B(n38443), .Z(n48714) );
  XOR U47985 ( .A(n48715), .B(n41394), .Z(n38443) );
  XOR U47986 ( .A(n48716), .B(n46032), .Z(n41394) );
  XOR U47987 ( .A(n46978), .B(n47579), .Z(n46032) );
  XNOR U47988 ( .A(n48717), .B(n48718), .Z(n47579) );
  XNOR U47989 ( .A(n46555), .B(n44903), .Z(n48718) );
  XOR U47990 ( .A(n48719), .B(n48720), .Z(n44903) );
  ANDN U47991 ( .B(n48721), .A(n48722), .Z(n48719) );
  XOR U47992 ( .A(n48723), .B(n48724), .Z(n46555) );
  ANDN U47993 ( .B(n48725), .A(n48726), .Z(n48723) );
  XNOR U47994 ( .A(n42547), .B(n48727), .Z(n48717) );
  XOR U47995 ( .A(n44685), .B(n47130), .Z(n48727) );
  XOR U47996 ( .A(n48728), .B(n48729), .Z(n47130) );
  ANDN U47997 ( .B(n48730), .A(n48731), .Z(n48728) );
  XOR U47998 ( .A(n48732), .B(n48733), .Z(n44685) );
  ANDN U47999 ( .B(n48734), .A(n48735), .Z(n48732) );
  XNOR U48000 ( .A(n48736), .B(n48737), .Z(n42547) );
  ANDN U48001 ( .B(n48738), .A(n48739), .Z(n48736) );
  XOR U48002 ( .A(n48740), .B(n48741), .Z(n46978) );
  XNOR U48003 ( .A(n46155), .B(n46504), .Z(n48741) );
  XNOR U48004 ( .A(n48742), .B(n48743), .Z(n46504) );
  ANDN U48005 ( .B(n48744), .A(n48745), .Z(n48742) );
  XOR U48006 ( .A(n48746), .B(n48747), .Z(n46155) );
  ANDN U48007 ( .B(n48748), .A(n48749), .Z(n48746) );
  XOR U48008 ( .A(n44761), .B(n48750), .Z(n48740) );
  XOR U48009 ( .A(n48751), .B(n45465), .Z(n48750) );
  XOR U48010 ( .A(n48752), .B(n48753), .Z(n45465) );
  NOR U48011 ( .A(n48754), .B(n48755), .Z(n48752) );
  XNOR U48012 ( .A(n48756), .B(n48757), .Z(n44761) );
  ANDN U48013 ( .B(n48758), .A(n48759), .Z(n48756) );
  NOR U48014 ( .A(n47440), .B(n43409), .Z(n48715) );
  XOR U48015 ( .A(n48760), .B(n44191), .Z(n43409) );
  XNOR U48016 ( .A(n48761), .B(n48762), .Z(n48311) );
  XNOR U48017 ( .A(n44938), .B(n48763), .Z(n48762) );
  XNOR U48018 ( .A(n48764), .B(n48765), .Z(n44938) );
  XOR U48019 ( .A(n43785), .B(n48766), .Z(n48761) );
  XOR U48020 ( .A(n45157), .B(n46288), .Z(n48766) );
  XNOR U48021 ( .A(n48767), .B(n48768), .Z(n46288) );
  ANDN U48022 ( .B(n48595), .A(n48596), .Z(n48767) );
  XNOR U48023 ( .A(n48769), .B(n48770), .Z(n45157) );
  ANDN U48024 ( .B(n48582), .A(n48583), .Z(n48769) );
  XNOR U48025 ( .A(n48771), .B(n48772), .Z(n43785) );
  XOR U48026 ( .A(n48774), .B(n42335), .Z(n47440) );
  IV U48027 ( .A(n45127), .Z(n42335) );
  XNOR U48028 ( .A(n48775), .B(n46678), .Z(n45127) );
  XOR U48029 ( .A(n48776), .B(n48777), .Z(n46678) );
  XNOR U48030 ( .A(n48778), .B(n45206), .Z(n48777) );
  XOR U48031 ( .A(n48779), .B(n48780), .Z(n45206) );
  ANDN U48032 ( .B(n48781), .A(n48782), .Z(n48779) );
  XOR U48033 ( .A(n43111), .B(n48783), .Z(n48776) );
  XOR U48034 ( .A(n42690), .B(n47463), .Z(n48783) );
  XOR U48035 ( .A(n48784), .B(n48785), .Z(n47463) );
  AND U48036 ( .A(n48786), .B(n48787), .Z(n48784) );
  XOR U48037 ( .A(n48788), .B(n48789), .Z(n42690) );
  ANDN U48038 ( .B(n48790), .A(n48791), .Z(n48788) );
  XNOR U48039 ( .A(n48792), .B(n48793), .Z(n43111) );
  ANDN U48040 ( .B(n48794), .A(n48795), .Z(n48792) );
  XNOR U48041 ( .A(n48796), .B(n41386), .Z(n39595) );
  XOR U48042 ( .A(n48797), .B(n43767), .Z(n41386) );
  XOR U48043 ( .A(n40001), .B(n48798), .Z(n48713) );
  XOR U48044 ( .A(n40049), .B(n40427), .Z(n48798) );
  XOR U48045 ( .A(n48799), .B(n43411), .Z(n40427) );
  XOR U48046 ( .A(n48800), .B(n44114), .Z(n43411) );
  ANDN U48047 ( .B(n43826), .A(n43398), .Z(n48799) );
  XNOR U48048 ( .A(n44693), .B(n48801), .Z(n43398) );
  XNOR U48049 ( .A(n48602), .B(n48802), .Z(n44693) );
  XOR U48050 ( .A(n48803), .B(n48804), .Z(n48602) );
  XNOR U48051 ( .A(n46925), .B(n45574), .Z(n48804) );
  XNOR U48052 ( .A(n48805), .B(n48033), .Z(n45574) );
  ANDN U48053 ( .B(n48032), .A(n46238), .Z(n48805) );
  XNOR U48054 ( .A(n48806), .B(n48022), .Z(n46925) );
  ANDN U48055 ( .B(n48021), .A(n46142), .Z(n48806) );
  XNOR U48056 ( .A(n45705), .B(n48807), .Z(n48803) );
  XOR U48057 ( .A(n47466), .B(n44532), .Z(n48807) );
  XNOR U48058 ( .A(n48808), .B(n48809), .Z(n44532) );
  ANDN U48059 ( .B(n48810), .A(n46146), .Z(n48808) );
  XNOR U48060 ( .A(n48811), .B(n48025), .Z(n47466) );
  ANDN U48061 ( .B(n48024), .A(n47153), .Z(n48811) );
  XNOR U48062 ( .A(n48812), .B(n48030), .Z(n45705) );
  ANDN U48063 ( .B(n48029), .A(n46136), .Z(n48812) );
  XOR U48064 ( .A(n48813), .B(n44513), .Z(n43826) );
  IV U48065 ( .A(n43600), .Z(n44513) );
  XOR U48066 ( .A(n48814), .B(n47056), .Z(n43600) );
  XOR U48067 ( .A(n48815), .B(n48816), .Z(n47056) );
  XNOR U48068 ( .A(n48817), .B(n43283), .Z(n48816) );
  XNOR U48069 ( .A(n48818), .B(n48819), .Z(n43283) );
  ANDN U48070 ( .B(n48820), .A(n48821), .Z(n48818) );
  XNOR U48071 ( .A(n44768), .B(n48822), .Z(n48815) );
  XOR U48072 ( .A(n46163), .B(n46541), .Z(n48822) );
  XNOR U48073 ( .A(n48823), .B(n48824), .Z(n46541) );
  ANDN U48074 ( .B(n48825), .A(n48826), .Z(n48823) );
  XNOR U48075 ( .A(n48827), .B(n48828), .Z(n46163) );
  AND U48076 ( .A(n48829), .B(n48830), .Z(n48827) );
  XNOR U48077 ( .A(n48831), .B(n48832), .Z(n44768) );
  ANDN U48078 ( .B(n48833), .A(n48834), .Z(n48831) );
  XNOR U48079 ( .A(n48835), .B(n41381), .Z(n40049) );
  XOR U48080 ( .A(n48296), .B(n45497), .Z(n41381) );
  XOR U48081 ( .A(n48836), .B(n47519), .Z(n45497) );
  XNOR U48082 ( .A(n48837), .B(n48838), .Z(n47519) );
  XNOR U48083 ( .A(n46597), .B(n46020), .Z(n48838) );
  XOR U48084 ( .A(n48839), .B(n48840), .Z(n46020) );
  ANDN U48085 ( .B(n48841), .A(n48842), .Z(n48839) );
  XOR U48086 ( .A(n48843), .B(n48844), .Z(n46597) );
  ANDN U48087 ( .B(n48845), .A(n48846), .Z(n48843) );
  XOR U48088 ( .A(n42847), .B(n48847), .Z(n48837) );
  XOR U48089 ( .A(n45682), .B(n47692), .Z(n48847) );
  XNOR U48090 ( .A(n48848), .B(n48849), .Z(n47692) );
  AND U48091 ( .A(n48850), .B(n48851), .Z(n48848) );
  XNOR U48092 ( .A(n48852), .B(n48853), .Z(n45682) );
  NOR U48093 ( .A(n48854), .B(n48855), .Z(n48852) );
  XOR U48094 ( .A(n48856), .B(n48857), .Z(n42847) );
  ANDN U48095 ( .B(n48858), .A(n48859), .Z(n48856) );
  XNOR U48096 ( .A(n48860), .B(n48861), .Z(n48296) );
  ANDN U48097 ( .B(n48862), .A(n48863), .Z(n48860) );
  ANDN U48098 ( .B(n43821), .A(n43402), .Z(n48835) );
  XNOR U48099 ( .A(n48864), .B(n44207), .Z(n43402) );
  XOR U48100 ( .A(n48865), .B(n44488), .Z(n43821) );
  XNOR U48101 ( .A(n48866), .B(n48867), .Z(n47248) );
  XNOR U48102 ( .A(n45449), .B(n42511), .Z(n48867) );
  XNOR U48103 ( .A(n48868), .B(n47627), .Z(n42511) );
  XOR U48104 ( .A(round_reg[717]), .B(n48869), .Z(n47627) );
  ANDN U48105 ( .B(n48870), .A(n48170), .Z(n48868) );
  XNOR U48106 ( .A(n48871), .B(n47613), .Z(n45449) );
  XNOR U48107 ( .A(round_reg[931]), .B(n48872), .Z(n47613) );
  XNOR U48108 ( .A(n45131), .B(n48874), .Z(n48866) );
  XOR U48109 ( .A(n45155), .B(n43677), .Z(n48874) );
  XNOR U48110 ( .A(n48875), .B(n47622), .Z(n43677) );
  XNOR U48111 ( .A(round_reg[860]), .B(n48876), .Z(n47622) );
  XNOR U48112 ( .A(n48878), .B(n47618), .Z(n45155) );
  XNOR U48113 ( .A(round_reg[703]), .B(n48879), .Z(n47618) );
  ANDN U48114 ( .B(n48880), .A(n48175), .Z(n48878) );
  XNOR U48115 ( .A(n48881), .B(n48182), .Z(n45131) );
  XNOR U48116 ( .A(n48884), .B(n41390), .Z(n40001) );
  XNOR U48117 ( .A(n48885), .B(n46198), .Z(n41390) );
  IV U48118 ( .A(n47529), .Z(n46198) );
  XNOR U48119 ( .A(n48886), .B(n46433), .Z(n47529) );
  XNOR U48120 ( .A(n48887), .B(n48888), .Z(n46433) );
  XOR U48121 ( .A(n48889), .B(n43098), .Z(n48888) );
  XOR U48122 ( .A(n48890), .B(n48891), .Z(n43098) );
  NOR U48123 ( .A(n48892), .B(n48893), .Z(n48890) );
  XOR U48124 ( .A(n45233), .B(n48894), .Z(n48887) );
  XOR U48125 ( .A(n42452), .B(n43720), .Z(n48894) );
  XNOR U48126 ( .A(n48895), .B(n48896), .Z(n43720) );
  XNOR U48127 ( .A(n48899), .B(n48900), .Z(n42452) );
  ANDN U48128 ( .B(n48901), .A(n48902), .Z(n48899) );
  XNOR U48129 ( .A(n48903), .B(n48904), .Z(n45233) );
  NOR U48130 ( .A(n48905), .B(n48906), .Z(n48903) );
  ANDN U48131 ( .B(n43834), .A(n43405), .Z(n48884) );
  XNOR U48132 ( .A(n48907), .B(n43965), .Z(n43405) );
  XNOR U48133 ( .A(n45786), .B(n46780), .Z(n43834) );
  XOR U48134 ( .A(n48908), .B(n48909), .Z(n46780) );
  ANDN U48135 ( .B(n48910), .A(n48332), .Z(n48908) );
  XOR U48136 ( .A(n48911), .B(n43817), .Z(n47436) );
  XOR U48137 ( .A(n48912), .B(n44571), .Z(n43817) );
  XNOR U48138 ( .A(n46872), .B(n48913), .Z(n44571) );
  XOR U48139 ( .A(n48914), .B(n48915), .Z(n46872) );
  XOR U48140 ( .A(n46440), .B(n46182), .Z(n48915) );
  XOR U48141 ( .A(n48916), .B(n48104), .Z(n46182) );
  AND U48142 ( .A(n48917), .B(n48105), .Z(n48916) );
  XNOR U48143 ( .A(n48918), .B(n48096), .Z(n46440) );
  XOR U48144 ( .A(n43523), .B(n48920), .Z(n48914) );
  XOR U48145 ( .A(n47575), .B(n45933), .Z(n48920) );
  XNOR U48146 ( .A(n48921), .B(n48091), .Z(n45933) );
  XNOR U48147 ( .A(n48923), .B(n48100), .Z(n47575) );
  AND U48148 ( .A(n48924), .B(n48101), .Z(n48923) );
  XNOR U48149 ( .A(n48925), .B(n48432), .Z(n43523) );
  ANDN U48150 ( .B(n43407), .A(n41384), .Z(n48911) );
  XOR U48151 ( .A(n48927), .B(n48928), .Z(n41384) );
  XOR U48152 ( .A(n48929), .B(n45339), .Z(n43407) );
  XNOR U48153 ( .A(n48930), .B(n48428), .Z(n45339) );
  XNOR U48154 ( .A(n48931), .B(n48932), .Z(n48428) );
  XNOR U48155 ( .A(n45840), .B(n46912), .Z(n48932) );
  XNOR U48156 ( .A(n48933), .B(n48934), .Z(n46912) );
  ANDN U48157 ( .B(n48095), .A(n48096), .Z(n48933) );
  XOR U48158 ( .A(round_reg[1585]), .B(n48935), .Z(n48096) );
  XOR U48159 ( .A(n48936), .B(n48937), .Z(n45840) );
  ANDN U48160 ( .B(n48431), .A(n48432), .Z(n48936) );
  XNOR U48161 ( .A(round_reg[1520]), .B(n48938), .Z(n48432) );
  XNOR U48162 ( .A(n44260), .B(n48939), .Z(n48931) );
  XOR U48163 ( .A(n43776), .B(n44231), .Z(n48939) );
  XOR U48164 ( .A(n48940), .B(n48941), .Z(n44231) );
  ANDN U48165 ( .B(n48099), .A(n48100), .Z(n48940) );
  XOR U48166 ( .A(round_reg[1459]), .B(n48942), .Z(n48100) );
  XOR U48167 ( .A(n48943), .B(n48944), .Z(n43776) );
  ANDN U48168 ( .B(n48090), .A(n48091), .Z(n48943) );
  XNOR U48169 ( .A(round_reg[1302]), .B(n48945), .Z(n48091) );
  XOR U48170 ( .A(n48946), .B(n48947), .Z(n44260) );
  ANDN U48171 ( .B(n48103), .A(n48104), .Z(n48946) );
  XOR U48172 ( .A(round_reg[1365]), .B(n48948), .Z(n48104) );
  XNOR U48173 ( .A(n48949), .B(n33765), .Z(n33700) );
  XOR U48174 ( .A(n38817), .B(n42651), .Z(n33765) );
  XNOR U48175 ( .A(n48950), .B(n40892), .Z(n42651) );
  AND U48176 ( .A(n41030), .B(n41642), .Z(n48950) );
  XOR U48177 ( .A(n48951), .B(n44608), .Z(n41030) );
  IV U48178 ( .A(n48123), .Z(n44608) );
  XNOR U48179 ( .A(n45062), .B(n41397), .Z(n38817) );
  XNOR U48180 ( .A(n48952), .B(n48953), .Z(n41397) );
  XOR U48181 ( .A(n36787), .B(n36951), .Z(n48953) );
  XOR U48182 ( .A(n48954), .B(n40891), .Z(n36951) );
  XOR U48183 ( .A(n43073), .B(n46473), .Z(n40891) );
  XNOR U48184 ( .A(n48955), .B(n48956), .Z(n46473) );
  ANDN U48185 ( .B(n46808), .A(n46809), .Z(n48955) );
  XNOR U48186 ( .A(round_reg[1358]), .B(n48957), .Z(n46809) );
  XNOR U48187 ( .A(n46947), .B(n48549), .Z(n43073) );
  XOR U48188 ( .A(n48958), .B(n48959), .Z(n48549) );
  XOR U48189 ( .A(n44985), .B(n48960), .Z(n48959) );
  XNOR U48190 ( .A(n48961), .B(n48369), .Z(n44985) );
  ANDN U48191 ( .B(n46475), .A(n46477), .Z(n48961) );
  XOR U48192 ( .A(round_reg[280]), .B(n48962), .Z(n46477) );
  XOR U48193 ( .A(n46311), .B(n48963), .Z(n48958) );
  XOR U48194 ( .A(n47810), .B(n45763), .Z(n48963) );
  XNOR U48195 ( .A(n48964), .B(n48357), .Z(n45763) );
  ANDN U48196 ( .B(n46480), .A(n46812), .Z(n48964) );
  IV U48197 ( .A(n46481), .Z(n46812) );
  XNOR U48198 ( .A(round_reg[28]), .B(n48965), .Z(n46481) );
  XNOR U48199 ( .A(n48966), .B(n48363), .Z(n47810) );
  ANDN U48200 ( .B(n46488), .A(n46490), .Z(n48966) );
  XOR U48201 ( .A(round_reg[114]), .B(n48967), .Z(n46490) );
  XNOR U48202 ( .A(n48968), .B(n48359), .Z(n46311) );
  ANDN U48203 ( .B(n48956), .A(n46808), .Z(n48968) );
  XOR U48204 ( .A(round_reg[173]), .B(n48558), .Z(n46808) );
  XOR U48205 ( .A(n48969), .B(n48970), .Z(n46947) );
  XOR U48206 ( .A(n43316), .B(n44821), .Z(n48970) );
  XOR U48207 ( .A(n48971), .B(n48972), .Z(n44821) );
  AND U48208 ( .A(n46608), .B(n46607), .Z(n48971) );
  XNOR U48209 ( .A(n48973), .B(n48974), .Z(n43316) );
  ANDN U48210 ( .B(n46611), .A(n46613), .Z(n48973) );
  XNOR U48211 ( .A(n42205), .B(n48975), .Z(n48969) );
  XOR U48212 ( .A(n47239), .B(n48976), .Z(n48975) );
  XNOR U48213 ( .A(n48977), .B(n48978), .Z(n47239) );
  ANDN U48214 ( .B(n46950), .A(n46952), .Z(n48977) );
  XOR U48215 ( .A(n48979), .B(n48980), .Z(n42205) );
  ANDN U48216 ( .B(n46621), .A(n46623), .Z(n48979) );
  ANDN U48217 ( .B(n40892), .A(n41642), .Z(n48954) );
  XOR U48218 ( .A(n48981), .B(n42868), .Z(n41642) );
  XOR U48219 ( .A(n48387), .B(n46185), .Z(n40892) );
  IV U48220 ( .A(n46501), .Z(n46185) );
  XNOR U48221 ( .A(n48982), .B(n47041), .Z(n48387) );
  ANDN U48222 ( .B(n48983), .A(n48984), .Z(n48982) );
  XOR U48223 ( .A(n48985), .B(n40882), .Z(n36787) );
  XOR U48224 ( .A(n48986), .B(n48548), .Z(n40882) );
  XOR U48225 ( .A(n48988), .B(n48989), .Z(n46684) );
  XNOR U48226 ( .A(n47023), .B(n46358), .Z(n48989) );
  XNOR U48227 ( .A(n48990), .B(n48991), .Z(n46358) );
  NOR U48228 ( .A(n48992), .B(n48993), .Z(n48990) );
  XNOR U48229 ( .A(n48994), .B(n48995), .Z(n47023) );
  ANDN U48230 ( .B(n48996), .A(n48997), .Z(n48994) );
  XNOR U48231 ( .A(n48998), .B(n48999), .Z(n48988) );
  XOR U48232 ( .A(n42497), .B(n46641), .Z(n48999) );
  XNOR U48233 ( .A(n49000), .B(n49001), .Z(n46641) );
  XNOR U48234 ( .A(n49004), .B(n49005), .Z(n42497) );
  NOR U48235 ( .A(n41651), .B(n40881), .Z(n48985) );
  XOR U48236 ( .A(n44688), .B(n49008), .Z(n40881) );
  IV U48237 ( .A(n48927), .Z(n44688) );
  XOR U48238 ( .A(n49009), .B(n46544), .Z(n48927) );
  XNOR U48239 ( .A(n49010), .B(n49011), .Z(n46544) );
  XNOR U48240 ( .A(n45480), .B(n45640), .Z(n49011) );
  XNOR U48241 ( .A(n49012), .B(n49013), .Z(n45640) );
  ANDN U48242 ( .B(n48209), .A(n49014), .Z(n49012) );
  XNOR U48243 ( .A(n49015), .B(n48280), .Z(n45480) );
  ANDN U48244 ( .B(n48281), .A(n49016), .Z(n49015) );
  XOR U48245 ( .A(n40844), .B(n49017), .Z(n49010) );
  XOR U48246 ( .A(n43582), .B(n46125), .Z(n49017) );
  XNOR U48247 ( .A(n49018), .B(n48276), .Z(n46125) );
  ANDN U48248 ( .B(n48213), .A(n48275), .Z(n49018) );
  XNOR U48249 ( .A(n49019), .B(n48284), .Z(n43582) );
  ANDN U48250 ( .B(n48200), .A(n48283), .Z(n49019) );
  XNOR U48251 ( .A(n49020), .B(n48661), .Z(n40844) );
  NOR U48252 ( .A(n49021), .B(n48204), .Z(n49020) );
  XOR U48253 ( .A(n49022), .B(n44026), .Z(n41651) );
  IV U48254 ( .A(n45308), .Z(n44026) );
  XOR U48255 ( .A(n35605), .B(n49023), .Z(n48952) );
  XOR U48256 ( .A(n35780), .B(n40859), .Z(n49023) );
  XNOR U48257 ( .A(n49024), .B(n40909), .Z(n40859) );
  XOR U48258 ( .A(n43587), .B(n49025), .Z(n40909) );
  ANDN U48259 ( .B(n40910), .A(n41647), .Z(n49024) );
  XOR U48260 ( .A(n49026), .B(n45753), .Z(n41647) );
  XOR U48261 ( .A(n46831), .B(n47844), .Z(n45753) );
  XNOR U48262 ( .A(n49027), .B(n49028), .Z(n47844) );
  XNOR U48263 ( .A(n49029), .B(n45349), .Z(n49028) );
  XOR U48264 ( .A(n49030), .B(n49031), .Z(n45349) );
  ANDN U48265 ( .B(n49032), .A(n49033), .Z(n49030) );
  XOR U48266 ( .A(n42856), .B(n49034), .Z(n49027) );
  XOR U48267 ( .A(n46232), .B(n49035), .Z(n49034) );
  XOR U48268 ( .A(n49036), .B(n49037), .Z(n46232) );
  NOR U48269 ( .A(n49038), .B(n47895), .Z(n49036) );
  XOR U48270 ( .A(n49039), .B(n49040), .Z(n42856) );
  NOR U48271 ( .A(n47901), .B(n49041), .Z(n49039) );
  IV U48272 ( .A(n49042), .Z(n47901) );
  XNOR U48273 ( .A(n49043), .B(n49044), .Z(n46831) );
  XNOR U48274 ( .A(n45232), .B(n49045), .Z(n49044) );
  XOR U48275 ( .A(n49046), .B(n49047), .Z(n45232) );
  AND U48276 ( .A(n49048), .B(n49049), .Z(n49046) );
  XNOR U48277 ( .A(n47325), .B(n49050), .Z(n49043) );
  XNOR U48278 ( .A(n45952), .B(n47034), .Z(n49050) );
  XNOR U48279 ( .A(n49051), .B(n49052), .Z(n47034) );
  ANDN U48280 ( .B(n49053), .A(n49054), .Z(n49051) );
  XNOR U48281 ( .A(n49055), .B(n49056), .Z(n45952) );
  NOR U48282 ( .A(n49057), .B(n49058), .Z(n49055) );
  XNOR U48283 ( .A(n49059), .B(n49060), .Z(n47325) );
  ANDN U48284 ( .B(n49061), .A(n49062), .Z(n49059) );
  XNOR U48285 ( .A(n48127), .B(n43552), .Z(n40910) );
  XNOR U48286 ( .A(n49063), .B(n49064), .Z(n43552) );
  XNOR U48287 ( .A(n49065), .B(n49066), .Z(n48127) );
  ANDN U48288 ( .B(n49067), .A(n49068), .Z(n49065) );
  XNOR U48289 ( .A(n49069), .B(n40885), .Z(n35780) );
  XNOR U48290 ( .A(n47874), .B(n41742), .Z(n40885) );
  XNOR U48291 ( .A(n46699), .B(n49070), .Z(n41742) );
  XNOR U48292 ( .A(n49071), .B(n49072), .Z(n46699) );
  XOR U48293 ( .A(n45809), .B(n43707), .Z(n49072) );
  XOR U48294 ( .A(n49073), .B(n47002), .Z(n43707) );
  XNOR U48295 ( .A(round_reg[69]), .B(n49074), .Z(n47002) );
  ANDN U48296 ( .B(n47003), .A(n47880), .Z(n49073) );
  XNOR U48297 ( .A(round_reg[1314]), .B(n49075), .Z(n47003) );
  XNOR U48298 ( .A(n49076), .B(n46855), .Z(n45809) );
  XOR U48299 ( .A(round_reg[299]), .B(n48452), .Z(n46855) );
  ANDN U48300 ( .B(n46856), .A(n47885), .Z(n49076) );
  XNOR U48301 ( .A(round_reg[1532]), .B(n49077), .Z(n46856) );
  XOR U48302 ( .A(n45094), .B(n49078), .Z(n49071) );
  XOR U48303 ( .A(n42525), .B(n45863), .Z(n49078) );
  XNOR U48304 ( .A(n49079), .B(n46869), .Z(n45863) );
  ANDN U48305 ( .B(n46870), .A(n47883), .Z(n49079) );
  XOR U48306 ( .A(round_reg[1471]), .B(n49081), .Z(n46870) );
  XNOR U48307 ( .A(n49082), .B(n46859), .Z(n42525) );
  XOR U48308 ( .A(round_reg[128]), .B(n49083), .Z(n46859) );
  ANDN U48309 ( .B(n46860), .A(n49084), .Z(n49082) );
  XNOR U48310 ( .A(n49085), .B(n46865), .Z(n45094) );
  XNOR U48311 ( .A(round_reg[47]), .B(n49086), .Z(n46865) );
  NOR U48312 ( .A(n47876), .B(n47877), .Z(n49085) );
  XOR U48313 ( .A(round_reg[1597]), .B(n49087), .Z(n47876) );
  XOR U48314 ( .A(n49088), .B(n46860), .Z(n47874) );
  XNOR U48315 ( .A(round_reg[1377]), .B(n49089), .Z(n46860) );
  ANDN U48316 ( .B(n49084), .A(n47014), .Z(n49088) );
  ANDN U48317 ( .B(n40886), .A(n41638), .Z(n49069) );
  XOR U48318 ( .A(n49090), .B(n43321), .Z(n41638) );
  IV U48319 ( .A(n48436), .Z(n43321) );
  XOR U48320 ( .A(n47468), .B(n49091), .Z(n48436) );
  XNOR U48321 ( .A(n49092), .B(n49093), .Z(n47468) );
  XNOR U48322 ( .A(n49094), .B(n45771), .Z(n49093) );
  XOR U48323 ( .A(n49095), .B(n49096), .Z(n45771) );
  ANDN U48324 ( .B(n49097), .A(n49098), .Z(n49095) );
  XNOR U48325 ( .A(n44184), .B(n49099), .Z(n49092) );
  XOR U48326 ( .A(n43078), .B(n46939), .Z(n49099) );
  XOR U48327 ( .A(n49100), .B(n49101), .Z(n46939) );
  XOR U48328 ( .A(n49104), .B(n49105), .Z(n43078) );
  ANDN U48329 ( .B(n49106), .A(n49107), .Z(n49104) );
  XOR U48330 ( .A(n49108), .B(n49109), .Z(n44184) );
  ANDN U48331 ( .B(n49110), .A(n49111), .Z(n49108) );
  XOR U48332 ( .A(n49112), .B(n45091), .Z(n40886) );
  XNOR U48333 ( .A(n49113), .B(n47259), .Z(n45091) );
  XOR U48334 ( .A(n49114), .B(n49115), .Z(n47259) );
  XNOR U48335 ( .A(n45329), .B(n45375), .Z(n49115) );
  XNOR U48336 ( .A(n49116), .B(n49117), .Z(n45375) );
  NOR U48337 ( .A(n47763), .B(n49118), .Z(n49116) );
  XNOR U48338 ( .A(n49119), .B(n49120), .Z(n45329) );
  NOR U48339 ( .A(n47768), .B(n49121), .Z(n49119) );
  XOR U48340 ( .A(n49122), .B(n49123), .Z(n49114) );
  XOR U48341 ( .A(n46169), .B(n44744), .Z(n49123) );
  XNOR U48342 ( .A(n49124), .B(n49125), .Z(n44744) );
  NOR U48343 ( .A(n47772), .B(n49126), .Z(n49124) );
  XNOR U48344 ( .A(n49127), .B(n49128), .Z(n46169) );
  AND U48345 ( .A(n47759), .B(n49129), .Z(n49127) );
  XOR U48346 ( .A(n49130), .B(n40896), .Z(n35605) );
  XNOR U48347 ( .A(n49131), .B(n45759), .Z(n40896) );
  NOR U48348 ( .A(n40895), .B(n41655), .Z(n49130) );
  XNOR U48349 ( .A(n47730), .B(n46702), .Z(n41655) );
  XNOR U48350 ( .A(n49132), .B(n49133), .Z(n47730) );
  AND U48351 ( .A(n49134), .B(n49135), .Z(n49132) );
  XOR U48352 ( .A(n46403), .B(n49136), .Z(n40895) );
  XNOR U48353 ( .A(n49137), .B(n49138), .Z(n48287) );
  XOR U48354 ( .A(n45412), .B(n46742), .Z(n49138) );
  XOR U48355 ( .A(n49139), .B(n48851), .Z(n46742) );
  ANDN U48356 ( .B(n49140), .A(n48850), .Z(n49139) );
  XNOR U48357 ( .A(n49141), .B(n48841), .Z(n45412) );
  ANDN U48358 ( .B(n49142), .A(n49143), .Z(n49141) );
  XOR U48359 ( .A(n47358), .B(n49144), .Z(n49137) );
  XOR U48360 ( .A(n47518), .B(n43718), .Z(n49144) );
  XOR U48361 ( .A(n49145), .B(n48859), .Z(n43718) );
  ANDN U48362 ( .B(n49146), .A(n48858), .Z(n49145) );
  XOR U48363 ( .A(n49147), .B(n48846), .Z(n47518) );
  ANDN U48364 ( .B(n49148), .A(n48845), .Z(n49147) );
  XOR U48365 ( .A(n49149), .B(n48855), .Z(n47358) );
  ANDN U48366 ( .B(n48854), .A(n49150), .Z(n49149) );
  XOR U48367 ( .A(n49151), .B(n49152), .Z(n46498) );
  XOR U48368 ( .A(n49153), .B(n49154), .Z(n49152) );
  XNOR U48369 ( .A(n47397), .B(n49155), .Z(n49151) );
  XNOR U48370 ( .A(n49156), .B(n49157), .Z(n49155) );
  XOR U48371 ( .A(n49158), .B(n49159), .Z(n47397) );
  ANDN U48372 ( .B(n49160), .A(n49161), .Z(n49158) );
  XOR U48373 ( .A(n49162), .B(n49163), .Z(n45062) );
  XOR U48374 ( .A(n37341), .B(n35154), .Z(n49163) );
  XOR U48375 ( .A(n49164), .B(n40875), .Z(n35154) );
  NOR U48376 ( .A(n40932), .B(n40876), .Z(n49164) );
  XOR U48377 ( .A(n49165), .B(n43323), .Z(n40876) );
  XOR U48378 ( .A(n46603), .B(n48166), .Z(n43323) );
  XNOR U48379 ( .A(n49166), .B(n49167), .Z(n48166) );
  XNOR U48380 ( .A(n46355), .B(n47606), .Z(n49167) );
  XNOR U48381 ( .A(n49168), .B(n49169), .Z(n47606) );
  ANDN U48382 ( .B(n47551), .A(n47552), .Z(n49168) );
  XOR U48383 ( .A(round_reg[1211]), .B(n49080), .Z(n47552) );
  XNOR U48384 ( .A(n49170), .B(n49171), .Z(n46355) );
  ANDN U48385 ( .B(n47556), .A(n47557), .Z(n49170) );
  XOR U48386 ( .A(round_reg[1219]), .B(n48514), .Z(n47557) );
  XOR U48387 ( .A(n44549), .B(n49172), .Z(n49166) );
  XOR U48388 ( .A(n45182), .B(n46787), .Z(n49172) );
  XNOR U48389 ( .A(n49173), .B(n49174), .Z(n46787) );
  ANDN U48390 ( .B(n47564), .A(n47566), .Z(n49173) );
  XNOR U48391 ( .A(round_reg[1121]), .B(n49175), .Z(n47566) );
  XNOR U48392 ( .A(n49176), .B(n49177), .Z(n45182) );
  ANDN U48393 ( .B(n47560), .A(n47561), .Z(n49176) );
  XOR U48394 ( .A(round_reg[1072]), .B(n49178), .Z(n47561) );
  XNOR U48395 ( .A(n49179), .B(n49180), .Z(n44549) );
  ANDN U48396 ( .B(n48184), .A(n47945), .Z(n49179) );
  XOR U48397 ( .A(round_reg[979]), .B(n49181), .Z(n47945) );
  XNOR U48398 ( .A(n49182), .B(n49183), .Z(n46603) );
  XOR U48399 ( .A(n46926), .B(n47462), .Z(n49183) );
  XOR U48400 ( .A(n49184), .B(n49185), .Z(n47462) );
  ANDN U48401 ( .B(n49186), .A(n49187), .Z(n49184) );
  XNOR U48402 ( .A(n49188), .B(n49189), .Z(n46926) );
  XOR U48403 ( .A(n45645), .B(n49192), .Z(n49182) );
  XOR U48404 ( .A(n49193), .B(n49194), .Z(n49192) );
  XNOR U48405 ( .A(n49195), .B(n49196), .Z(n45645) );
  XOR U48406 ( .A(n49199), .B(n44915), .Z(n40932) );
  IV U48407 ( .A(n45389), .Z(n44915) );
  XOR U48408 ( .A(n47997), .B(n47243), .Z(n45389) );
  XNOR U48409 ( .A(n49200), .B(n49201), .Z(n47243) );
  XOR U48410 ( .A(n46037), .B(n44825), .Z(n49201) );
  XOR U48411 ( .A(n49202), .B(n49203), .Z(n44825) );
  AND U48412 ( .A(n49204), .B(n49205), .Z(n49202) );
  XNOR U48413 ( .A(n49206), .B(n47019), .Z(n46037) );
  AND U48414 ( .A(n49207), .B(n47020), .Z(n49206) );
  XOR U48415 ( .A(n45652), .B(n49208), .Z(n49200) );
  XOR U48416 ( .A(n45596), .B(n44262), .Z(n49208) );
  XNOR U48417 ( .A(n49209), .B(n48498), .Z(n44262) );
  ANDN U48418 ( .B(n48499), .A(n49210), .Z(n49209) );
  XNOR U48419 ( .A(n49211), .B(n46051), .Z(n45596) );
  AND U48420 ( .A(n49212), .B(n46052), .Z(n49211) );
  XNOR U48421 ( .A(n49213), .B(n46047), .Z(n45652) );
  ANDN U48422 ( .B(n46048), .A(n49214), .Z(n49213) );
  XNOR U48423 ( .A(n49215), .B(n49216), .Z(n47997) );
  XOR U48424 ( .A(n43838), .B(n45936), .Z(n49216) );
  XOR U48425 ( .A(n49217), .B(n47297), .Z(n45936) );
  AND U48426 ( .A(n47377), .B(n47298), .Z(n49217) );
  XNOR U48427 ( .A(n49218), .B(n47290), .Z(n43838) );
  AND U48428 ( .A(n47374), .B(n47291), .Z(n49218) );
  XOR U48429 ( .A(n41656), .B(n49219), .Z(n49215) );
  XOR U48430 ( .A(n41729), .B(n44531), .Z(n49219) );
  XNOR U48431 ( .A(n49220), .B(n48082), .Z(n44531) );
  ANDN U48432 ( .B(n48083), .A(n47364), .Z(n49220) );
  XOR U48433 ( .A(n49221), .B(n49222), .Z(n41729) );
  ANDN U48434 ( .B(n49223), .A(n48345), .Z(n49221) );
  XNOR U48435 ( .A(n49224), .B(n47587), .Z(n41656) );
  ANDN U48436 ( .B(n47588), .A(n47368), .Z(n49224) );
  XNOR U48437 ( .A(n49225), .B(n40865), .Z(n37341) );
  NOR U48438 ( .A(n45075), .B(n43481), .Z(n49225) );
  XOR U48439 ( .A(n49226), .B(n42163), .Z(n43481) );
  XOR U48440 ( .A(n49227), .B(n43904), .Z(n45075) );
  XOR U48441 ( .A(n38736), .B(n49228), .Z(n49162) );
  XOR U48442 ( .A(n38877), .B(n39108), .Z(n49228) );
  XNOR U48443 ( .A(n49229), .B(n49230), .Z(n39108) );
  NOR U48444 ( .A(n41608), .B(n43488), .Z(n49229) );
  XNOR U48445 ( .A(n45151), .B(n47912), .Z(n41608) );
  XOR U48446 ( .A(n49231), .B(n49232), .Z(n47912) );
  AND U48447 ( .A(n47828), .B(n49233), .Z(n49231) );
  IV U48448 ( .A(n45992), .Z(n45151) );
  XNOR U48449 ( .A(n48406), .B(n48836), .Z(n45992) );
  XNOR U48450 ( .A(n49234), .B(n49235), .Z(n48836) );
  XNOR U48451 ( .A(n45730), .B(n48951), .Z(n49235) );
  XNOR U48452 ( .A(n49236), .B(n49237), .Z(n48951) );
  ANDN U48453 ( .B(n48687), .A(n48688), .Z(n49236) );
  XOR U48454 ( .A(n49238), .B(n49239), .Z(n45730) );
  NOR U48455 ( .A(n48294), .B(n48292), .Z(n49238) );
  XOR U48456 ( .A(n49240), .B(n49241), .Z(n49234) );
  XOR U48457 ( .A(n44607), .B(n48122), .Z(n49241) );
  XNOR U48458 ( .A(n49242), .B(n49243), .Z(n48122) );
  ANDN U48459 ( .B(n48304), .A(n48302), .Z(n49242) );
  XOR U48460 ( .A(n49244), .B(n49245), .Z(n44607) );
  XOR U48461 ( .A(n49246), .B(n49247), .Z(n48406) );
  XOR U48462 ( .A(n42449), .B(n44568), .Z(n49247) );
  XOR U48463 ( .A(n49248), .B(n47829), .Z(n44568) );
  ANDN U48464 ( .B(n49232), .A(n49233), .Z(n49248) );
  XNOR U48465 ( .A(n49249), .B(n47823), .Z(n42449) );
  NOR U48466 ( .A(n47920), .B(n47919), .Z(n49249) );
  XOR U48467 ( .A(n46577), .B(n49250), .Z(n49246) );
  XOR U48468 ( .A(n45744), .B(n45587), .Z(n49250) );
  XNOR U48469 ( .A(n49251), .B(n48164), .Z(n45587) );
  NOR U48470 ( .A(n47924), .B(n47922), .Z(n49251) );
  XNOR U48471 ( .A(n49252), .B(n47833), .Z(n45744) );
  ANDN U48472 ( .B(n47926), .A(n47927), .Z(n49252) );
  XNOR U48473 ( .A(n49253), .B(n49254), .Z(n46577) );
  ANDN U48474 ( .B(n47914), .A(n47916), .Z(n49253) );
  XNOR U48475 ( .A(n49255), .B(n40871), .Z(n38877) );
  NOR U48476 ( .A(n43493), .B(n40928), .Z(n49255) );
  XOR U48477 ( .A(n49240), .B(n48123), .Z(n40928) );
  XOR U48478 ( .A(n47693), .B(n46579), .Z(n48123) );
  XNOR U48479 ( .A(n49256), .B(n49257), .Z(n46579) );
  XOR U48480 ( .A(n49258), .B(n46075), .Z(n49257) );
  XNOR U48481 ( .A(n49259), .B(n49260), .Z(n46075) );
  AND U48482 ( .A(n48302), .B(n49243), .Z(n49259) );
  XOR U48483 ( .A(round_reg[924]), .B(n49261), .Z(n48302) );
  XOR U48484 ( .A(n42669), .B(n49262), .Z(n49256) );
  XNOR U48485 ( .A(n46511), .B(n47238), .Z(n49262) );
  XNOR U48486 ( .A(n49263), .B(n49264), .Z(n47238) );
  ANDN U48487 ( .B(n49237), .A(n48687), .Z(n49263) );
  XOR U48488 ( .A(round_reg[696]), .B(n49265), .Z(n48687) );
  XNOR U48489 ( .A(n49266), .B(n49267), .Z(n46511) );
  ANDN U48490 ( .B(n48298), .A(n49245), .Z(n49266) );
  XNOR U48491 ( .A(round_reg[853]), .B(n49268), .Z(n48298) );
  XNOR U48492 ( .A(n49269), .B(n49270), .Z(n42669) );
  ANDN U48493 ( .B(n48292), .A(n49239), .Z(n49269) );
  XOR U48494 ( .A(round_reg[710]), .B(n49271), .Z(n48292) );
  XOR U48495 ( .A(n49272), .B(n49273), .Z(n47693) );
  XNOR U48496 ( .A(n49274), .B(n49275), .Z(n49273) );
  XNOR U48497 ( .A(n45166), .B(n49276), .Z(n49272) );
  XOR U48498 ( .A(n45667), .B(n49277), .Z(n49276) );
  XOR U48499 ( .A(n49278), .B(n49279), .Z(n45667) );
  ANDN U48500 ( .B(n48846), .A(n48844), .Z(n49278) );
  XNOR U48501 ( .A(round_reg[102]), .B(n49280), .Z(n48846) );
  XNOR U48502 ( .A(n49281), .B(n49282), .Z(n45166) );
  XOR U48503 ( .A(round_reg[161]), .B(n49175), .Z(n48855) );
  XNOR U48504 ( .A(n49283), .B(n49284), .Z(n49240) );
  NOR U48505 ( .A(n48862), .B(n48861), .Z(n49283) );
  XOR U48506 ( .A(n49285), .B(n42524), .Z(n43493) );
  XNOR U48507 ( .A(n49286), .B(n41548), .Z(n38736) );
  XOR U48508 ( .A(n49287), .B(n43965), .Z(n40938) );
  XOR U48509 ( .A(n47360), .B(n47643), .Z(n43965) );
  XNOR U48510 ( .A(n49288), .B(n49289), .Z(n47643) );
  XNOR U48511 ( .A(n46003), .B(n42341), .Z(n49289) );
  XNOR U48512 ( .A(n49290), .B(n49291), .Z(n42341) );
  AND U48513 ( .A(n49292), .B(n49293), .Z(n49290) );
  XNOR U48514 ( .A(n49294), .B(n49295), .Z(n46003) );
  AND U48515 ( .A(n49296), .B(n49297), .Z(n49294) );
  XOR U48516 ( .A(n48106), .B(n49298), .Z(n49288) );
  XOR U48517 ( .A(n45246), .B(n47402), .Z(n49298) );
  XOR U48518 ( .A(n49299), .B(n49300), .Z(n47402) );
  XNOR U48519 ( .A(n49303), .B(n49304), .Z(n45246) );
  NOR U48520 ( .A(n49305), .B(n49306), .Z(n49303) );
  XNOR U48521 ( .A(n49307), .B(n49308), .Z(n48106) );
  NOR U48522 ( .A(n49309), .B(n49310), .Z(n49307) );
  XNOR U48523 ( .A(n49311), .B(n49312), .Z(n47360) );
  XNOR U48524 ( .A(n46357), .B(n47630), .Z(n49312) );
  XNOR U48525 ( .A(n49313), .B(n49204), .Z(n47630) );
  ANDN U48526 ( .B(n49314), .A(n49315), .Z(n49313) );
  XNOR U48527 ( .A(n49316), .B(n49212), .Z(n46357) );
  ANDN U48528 ( .B(n49317), .A(n46050), .Z(n49316) );
  XNOR U48529 ( .A(n49318), .B(n49319), .Z(n49311) );
  XNOR U48530 ( .A(n45370), .B(n45838), .Z(n49319) );
  XNOR U48531 ( .A(n49320), .B(n49210), .Z(n45838) );
  ANDN U48532 ( .B(n49321), .A(n48497), .Z(n49320) );
  XOR U48533 ( .A(n49322), .B(n49214), .Z(n45370) );
  IV U48534 ( .A(n49323), .Z(n49214) );
  NOR U48535 ( .A(n49324), .B(n46046), .Z(n49322) );
  XNOR U48536 ( .A(n49325), .B(n45734), .Z(n41549) );
  NOR U48537 ( .A(n33764), .B(n35918), .Z(n48949) );
  XOR U48538 ( .A(n37071), .B(n44363), .Z(n35918) );
  XOR U48539 ( .A(n49328), .B(n42918), .Z(n44363) );
  ANDN U48540 ( .B(n41328), .A(n45842), .Z(n49328) );
  IV U48541 ( .A(n41330), .Z(n45842) );
  XOR U48542 ( .A(n49329), .B(n44207), .Z(n41330) );
  XNOR U48543 ( .A(n49330), .B(n46694), .Z(n44207) );
  XOR U48544 ( .A(n49331), .B(n49332), .Z(n46694) );
  XOR U48545 ( .A(n42460), .B(n44028), .Z(n49332) );
  XOR U48546 ( .A(n49333), .B(n48143), .Z(n44028) );
  ANDN U48547 ( .B(n48144), .A(n49334), .Z(n49333) );
  XNOR U48548 ( .A(n49335), .B(n48131), .Z(n42460) );
  NOR U48549 ( .A(n48130), .B(n49336), .Z(n49335) );
  XOR U48550 ( .A(n47069), .B(n49337), .Z(n49331) );
  XOR U48551 ( .A(n45366), .B(n48124), .Z(n49337) );
  XNOR U48552 ( .A(n49338), .B(n48139), .Z(n48124) );
  ANDN U48553 ( .B(n48140), .A(n49339), .Z(n49338) );
  XNOR U48554 ( .A(n49340), .B(n48135), .Z(n45366) );
  ANDN U48555 ( .B(n48136), .A(n49341), .Z(n49340) );
  XNOR U48556 ( .A(n49342), .B(n49067), .Z(n47069) );
  AND U48557 ( .A(n49343), .B(n49068), .Z(n49342) );
  XOR U48558 ( .A(n49344), .B(n49345), .Z(n39841) );
  XNOR U48559 ( .A(n43497), .B(n42470), .Z(n49345) );
  XNOR U48560 ( .A(n49346), .B(n46230), .Z(n42470) );
  XOR U48561 ( .A(n49347), .B(n44864), .Z(n46230) );
  ANDN U48562 ( .B(n43988), .A(n43987), .Z(n49346) );
  XOR U48563 ( .A(n48153), .B(n47640), .Z(n43987) );
  XOR U48564 ( .A(n49348), .B(n49349), .Z(n48153) );
  ANDN U48565 ( .B(n49350), .A(n49351), .Z(n49348) );
  IV U48566 ( .A(n39504), .Z(n43988) );
  XNOR U48567 ( .A(n49354), .B(n47270), .Z(n47307) );
  ANDN U48568 ( .B(n48009), .A(n48008), .Z(n49354) );
  XNOR U48569 ( .A(n49355), .B(n43514), .Z(n43497) );
  XNOR U48570 ( .A(n43967), .B(n49356), .Z(n43514) );
  XNOR U48571 ( .A(n46319), .B(n46705), .Z(n43967) );
  XNOR U48572 ( .A(n49357), .B(n49358), .Z(n46705) );
  XOR U48573 ( .A(n47583), .B(n45591), .Z(n49358) );
  XOR U48574 ( .A(n49359), .B(n49360), .Z(n45591) );
  ANDN U48575 ( .B(n49361), .A(n49362), .Z(n49359) );
  XNOR U48576 ( .A(n49363), .B(n49364), .Z(n47583) );
  ANDN U48577 ( .B(n49365), .A(n49366), .Z(n49363) );
  XOR U48578 ( .A(n49367), .B(n49368), .Z(n49357) );
  XOR U48579 ( .A(n47455), .B(n49369), .Z(n49368) );
  XNOR U48580 ( .A(n49370), .B(n49371), .Z(n47455) );
  ANDN U48581 ( .B(n49372), .A(n49373), .Z(n49370) );
  XOR U48582 ( .A(n49374), .B(n49375), .Z(n46319) );
  XOR U48583 ( .A(n42418), .B(n42519), .Z(n49375) );
  XOR U48584 ( .A(n49376), .B(n49377), .Z(n42519) );
  ANDN U48585 ( .B(n48526), .A(n48525), .Z(n49376) );
  XNOR U48586 ( .A(n49378), .B(n49379), .Z(n42418) );
  ANDN U48587 ( .B(n48529), .A(n48531), .Z(n49378) );
  XOR U48588 ( .A(n46407), .B(n49380), .Z(n49374) );
  XOR U48589 ( .A(n44169), .B(n46025), .Z(n49380) );
  XNOR U48590 ( .A(n49381), .B(n49382), .Z(n46025) );
  ANDN U48591 ( .B(n48542), .A(n48544), .Z(n49381) );
  XNOR U48592 ( .A(n49383), .B(n49384), .Z(n44169) );
  AND U48593 ( .A(n48540), .B(n48538), .Z(n49383) );
  XNOR U48594 ( .A(n49385), .B(n49386), .Z(n46407) );
  NOR U48595 ( .A(n48536), .B(n48534), .Z(n49385) );
  AND U48596 ( .A(n39499), .B(n43513), .Z(n49355) );
  XOR U48597 ( .A(n43899), .B(n49387), .Z(n43513) );
  XNOR U48598 ( .A(n46989), .B(n44009), .Z(n39499) );
  XNOR U48599 ( .A(n49388), .B(n49389), .Z(n46989) );
  ANDN U48600 ( .B(n49390), .A(n48462), .Z(n49388) );
  XNOR U48601 ( .A(n40134), .B(n49391), .Z(n49344) );
  XOR U48602 ( .A(n41083), .B(n38960), .Z(n49391) );
  XNOR U48603 ( .A(n49392), .B(n43502), .Z(n38960) );
  IV U48604 ( .A(n46226), .Z(n43502) );
  XOR U48605 ( .A(n49393), .B(n46571), .Z(n46226) );
  ANDN U48606 ( .B(n43503), .A(n39512), .Z(n49392) );
  XOR U48607 ( .A(n49394), .B(n47991), .Z(n39512) );
  XOR U48608 ( .A(n48913), .B(n49395), .Z(n47991) );
  XNOR U48609 ( .A(n49396), .B(n49397), .Z(n48913) );
  XNOR U48610 ( .A(n49398), .B(n45674), .Z(n49397) );
  XOR U48611 ( .A(n49399), .B(n49400), .Z(n45674) );
  ANDN U48612 ( .B(n49401), .A(n49402), .Z(n49399) );
  XOR U48613 ( .A(n45639), .B(n49403), .Z(n49396) );
  XOR U48614 ( .A(n49404), .B(n43092), .Z(n49403) );
  XOR U48615 ( .A(n49405), .B(n49406), .Z(n43092) );
  ANDN U48616 ( .B(n49407), .A(n49408), .Z(n49405) );
  XOR U48617 ( .A(n49409), .B(n49410), .Z(n45639) );
  NOR U48618 ( .A(n49411), .B(n49412), .Z(n49409) );
  XOR U48619 ( .A(n45320), .B(n49413), .Z(n43503) );
  IV U48620 ( .A(n45630), .Z(n45320) );
  XNOR U48621 ( .A(n49414), .B(n43505), .Z(n41083) );
  XOR U48622 ( .A(n42504), .B(n49415), .Z(n43505) );
  AND U48623 ( .A(n43506), .B(n39508), .Z(n49414) );
  XNOR U48624 ( .A(n49416), .B(n45255), .Z(n39508) );
  XOR U48625 ( .A(n49417), .B(n45439), .Z(n43506) );
  IV U48626 ( .A(n45621), .Z(n45439) );
  XNOR U48627 ( .A(n49418), .B(n43511), .Z(n40134) );
  XNOR U48628 ( .A(n49419), .B(n44036), .Z(n43511) );
  AND U48629 ( .A(n40362), .B(n43510), .Z(n49418) );
  XOR U48630 ( .A(n49420), .B(n49156), .Z(n43510) );
  XOR U48631 ( .A(n49421), .B(n49422), .Z(n49156) );
  ANDN U48632 ( .B(n49423), .A(n49424), .Z(n49421) );
  XOR U48633 ( .A(n49274), .B(n45167), .Z(n40362) );
  XOR U48634 ( .A(n49425), .B(n49426), .Z(n49274) );
  ANDN U48635 ( .B(n48859), .A(n48857), .Z(n49425) );
  XOR U48636 ( .A(round_reg[268]), .B(n49427), .Z(n48859) );
  XOR U48637 ( .A(n49428), .B(n49429), .Z(n40086) );
  XNOR U48638 ( .A(n42904), .B(n36319), .Z(n49429) );
  XOR U48639 ( .A(n49430), .B(n42922), .Z(n36319) );
  XOR U48640 ( .A(n48381), .B(n45569), .Z(n42922) );
  XNOR U48641 ( .A(n49431), .B(n49432), .Z(n48381) );
  ANDN U48642 ( .B(n49433), .A(n47570), .Z(n49431) );
  ANDN U48643 ( .B(n43996), .A(n42921), .Z(n49430) );
  XOR U48644 ( .A(n45621), .B(n49434), .Z(n42921) );
  XNOR U48645 ( .A(n49435), .B(n41740), .Z(n43996) );
  IV U48646 ( .A(n46071), .Z(n41740) );
  XNOR U48647 ( .A(n49436), .B(n42925), .Z(n42904) );
  XOR U48648 ( .A(n49437), .B(n41649), .Z(n42925) );
  ANDN U48649 ( .B(n41332), .A(n42924), .Z(n49436) );
  XNOR U48650 ( .A(n49440), .B(n46571), .Z(n42924) );
  XOR U48651 ( .A(n48775), .B(n49441), .Z(n46571) );
  XOR U48652 ( .A(n49442), .B(n49443), .Z(n48775) );
  XOR U48653 ( .A(n46196), .B(n45394), .Z(n49443) );
  XNOR U48654 ( .A(n49444), .B(n49445), .Z(n45394) );
  ANDN U48655 ( .B(n49446), .A(n49447), .Z(n49444) );
  XOR U48656 ( .A(n49448), .B(n49449), .Z(n46196) );
  ANDN U48657 ( .B(n49450), .A(n49451), .Z(n49448) );
  XOR U48658 ( .A(n48195), .B(n49452), .Z(n49442) );
  XOR U48659 ( .A(n46285), .B(n47170), .Z(n49452) );
  XOR U48660 ( .A(n49453), .B(n49454), .Z(n47170) );
  ANDN U48661 ( .B(n49455), .A(n49456), .Z(n49453) );
  XNOR U48662 ( .A(n49457), .B(n49458), .Z(n46285) );
  ANDN U48663 ( .B(n49459), .A(n49460), .Z(n49457) );
  XOR U48664 ( .A(n49461), .B(n49462), .Z(n48195) );
  ANDN U48665 ( .B(n49463), .A(n49464), .Z(n49461) );
  XOR U48666 ( .A(n42855), .B(n49035), .Z(n41332) );
  XNOR U48667 ( .A(n49465), .B(n49466), .Z(n49035) );
  NOR U48668 ( .A(n49467), .B(n49468), .Z(n49465) );
  XOR U48669 ( .A(n41157), .B(n49469), .Z(n49428) );
  XNOR U48670 ( .A(n38424), .B(n38150), .Z(n49469) );
  XOR U48671 ( .A(n49470), .B(n42912), .Z(n38150) );
  IV U48672 ( .A(n45839), .Z(n42912) );
  XNOR U48673 ( .A(n49471), .B(n44114), .Z(n45839) );
  XOR U48674 ( .A(n49472), .B(n48190), .Z(n44114) );
  XNOR U48675 ( .A(n49473), .B(n49474), .Z(n48190) );
  XNOR U48676 ( .A(n49475), .B(n47473), .Z(n49474) );
  XNOR U48677 ( .A(n49476), .B(n49477), .Z(n47473) );
  ANDN U48678 ( .B(n49478), .A(n48724), .Z(n49476) );
  XOR U48679 ( .A(n46093), .B(n49479), .Z(n49473) );
  XOR U48680 ( .A(n45379), .B(n45248), .Z(n49479) );
  XOR U48681 ( .A(n49480), .B(n49481), .Z(n45248) );
  ANDN U48682 ( .B(n49482), .A(n48729), .Z(n49480) );
  XNOR U48683 ( .A(n49483), .B(n49484), .Z(n45379) );
  AND U48684 ( .A(n48737), .B(n49485), .Z(n49483) );
  XOR U48685 ( .A(n49486), .B(n49487), .Z(n46093) );
  ANDN U48686 ( .B(n49488), .A(n48720), .Z(n49486) );
  ANDN U48687 ( .B(n42913), .A(n41322), .Z(n49470) );
  XOR U48688 ( .A(n45858), .B(n49489), .Z(n41322) );
  IV U48689 ( .A(n46675), .Z(n45858) );
  XNOR U48690 ( .A(n47475), .B(n49009), .Z(n46675) );
  XNOR U48691 ( .A(n49490), .B(n49491), .Z(n49009) );
  XNOR U48692 ( .A(n48269), .B(n44855), .Z(n49491) );
  XNOR U48693 ( .A(n49492), .B(n49450), .Z(n44855) );
  ANDN U48694 ( .B(n49493), .A(n49494), .Z(n49492) );
  XNOR U48695 ( .A(n49495), .B(n49455), .Z(n48269) );
  ANDN U48696 ( .B(n49496), .A(n49497), .Z(n49495) );
  XNOR U48697 ( .A(n44920), .B(n49498), .Z(n49490) );
  XOR U48698 ( .A(n46790), .B(n46596), .Z(n49498) );
  XNOR U48699 ( .A(n49499), .B(n49463), .Z(n46596) );
  NOR U48700 ( .A(n49500), .B(n49501), .Z(n49499) );
  XNOR U48701 ( .A(n49502), .B(n49446), .Z(n46790) );
  ANDN U48702 ( .B(n49503), .A(n49504), .Z(n49502) );
  XNOR U48703 ( .A(n49505), .B(n49459), .Z(n44920) );
  ANDN U48704 ( .B(n49506), .A(n49507), .Z(n49505) );
  XOR U48705 ( .A(n49508), .B(n49509), .Z(n47475) );
  XNOR U48706 ( .A(n49419), .B(n44035), .Z(n49509) );
  XOR U48707 ( .A(n49510), .B(n48795), .Z(n44035) );
  ANDN U48708 ( .B(n49511), .A(n49512), .Z(n49510) );
  XNOR U48709 ( .A(n49513), .B(n48786), .Z(n49419) );
  AND U48710 ( .A(n49514), .B(n49515), .Z(n49513) );
  XOR U48711 ( .A(n44796), .B(n49516), .Z(n49508) );
  XNOR U48712 ( .A(n49517), .B(n46464), .Z(n49516) );
  XOR U48713 ( .A(n49518), .B(n48782), .Z(n46464) );
  ANDN U48714 ( .B(n49519), .A(n49520), .Z(n49518) );
  ANDN U48715 ( .B(n49522), .A(n49523), .Z(n49521) );
  XOR U48716 ( .A(n49524), .B(n42868), .Z(n42913) );
  IV U48717 ( .A(n49525), .Z(n42868) );
  XNOR U48718 ( .A(n49526), .B(n42917), .Z(n38424) );
  XNOR U48719 ( .A(n49420), .B(n49157), .Z(n42917) );
  XNOR U48720 ( .A(n49527), .B(n49528), .Z(n49157) );
  NOR U48721 ( .A(n49529), .B(n49530), .Z(n49527) );
  ANDN U48722 ( .B(n42918), .A(n41328), .Z(n49526) );
  XOR U48723 ( .A(n49369), .B(n47456), .Z(n41328) );
  IV U48724 ( .A(n45592), .Z(n47456) );
  XNOR U48725 ( .A(n49531), .B(n49532), .Z(n49369) );
  NOR U48726 ( .A(n49533), .B(n49534), .Z(n49531) );
  XNOR U48727 ( .A(n48473), .B(n45861), .Z(n42918) );
  XNOR U48728 ( .A(n49537), .B(n49538), .Z(n48473) );
  NOR U48729 ( .A(n49539), .B(n49540), .Z(n49537) );
  XNOR U48730 ( .A(n49541), .B(n42909), .Z(n41157) );
  XOR U48731 ( .A(n49542), .B(n42522), .Z(n42909) );
  IV U48732 ( .A(n45669), .Z(n42522) );
  XNOR U48733 ( .A(n49543), .B(n48469), .Z(n45669) );
  XNOR U48734 ( .A(n49544), .B(n49545), .Z(n48469) );
  XOR U48735 ( .A(n49546), .B(n44540), .Z(n49545) );
  XNOR U48736 ( .A(n49547), .B(n49548), .Z(n44540) );
  AND U48737 ( .A(n49133), .B(n49549), .Z(n49547) );
  XNOR U48738 ( .A(n46193), .B(n49550), .Z(n49544) );
  XOR U48739 ( .A(n49551), .B(n47072), .Z(n49550) );
  XNOR U48740 ( .A(n49552), .B(n49553), .Z(n47072) );
  ANDN U48741 ( .B(n49554), .A(n47726), .Z(n49552) );
  XNOR U48742 ( .A(n49555), .B(n49556), .Z(n46193) );
  ANDN U48743 ( .B(n49557), .A(n49558), .Z(n49555) );
  XOR U48744 ( .A(n46103), .B(n49559), .Z(n42910) );
  XNOR U48745 ( .A(n47688), .B(n45750), .Z(n46103) );
  XNOR U48746 ( .A(n49560), .B(n49561), .Z(n45750) );
  XOR U48747 ( .A(n46891), .B(n45224), .Z(n49561) );
  XOR U48748 ( .A(n49562), .B(n47102), .Z(n45224) );
  ANDN U48749 ( .B(n47103), .A(n49563), .Z(n49562) );
  XNOR U48750 ( .A(n49564), .B(n46908), .Z(n46891) );
  ANDN U48751 ( .B(n46909), .A(n48374), .Z(n49564) );
  XOR U48752 ( .A(n45811), .B(n49565), .Z(n49560) );
  XOR U48753 ( .A(n44181), .B(n44553), .Z(n49565) );
  XNOR U48754 ( .A(n49566), .B(n46904), .Z(n44553) );
  ANDN U48755 ( .B(n46905), .A(n48383), .Z(n49566) );
  XNOR U48756 ( .A(n49567), .B(n46898), .Z(n44181) );
  ANDN U48757 ( .B(n46899), .A(n48377), .Z(n49567) );
  XNOR U48758 ( .A(n49568), .B(n47571), .Z(n45811) );
  ANDN U48759 ( .B(n47572), .A(n49432), .Z(n49568) );
  XOR U48760 ( .A(n49569), .B(n49570), .Z(n47688) );
  XOR U48761 ( .A(n44973), .B(n45097), .Z(n49570) );
  XOR U48762 ( .A(n49571), .B(n47677), .Z(n45097) );
  NOR U48763 ( .A(n45869), .B(n47676), .Z(n49571) );
  XNOR U48764 ( .A(n49572), .B(n49573), .Z(n44973) );
  NOR U48765 ( .A(n45878), .B(n49574), .Z(n49572) );
  XOR U48766 ( .A(n46562), .B(n49575), .Z(n49569) );
  XOR U48767 ( .A(n42339), .B(n46626), .Z(n49575) );
  XNOR U48768 ( .A(n49576), .B(n47638), .Z(n46626) );
  NOR U48769 ( .A(n47637), .B(n49577), .Z(n49576) );
  XNOR U48770 ( .A(n49578), .B(n48186), .Z(n42339) );
  ANDN U48771 ( .B(n48187), .A(n45882), .Z(n49578) );
  XNOR U48772 ( .A(n49579), .B(n46760), .Z(n46562) );
  ANDN U48773 ( .B(n46761), .A(n45874), .Z(n49579) );
  XOR U48774 ( .A(n49580), .B(n48600), .Z(n41318) );
  XOR U48775 ( .A(n48493), .B(n49581), .Z(n48600) );
  XOR U48776 ( .A(n49582), .B(n49583), .Z(n48493) );
  XNOR U48777 ( .A(n49489), .B(n46676), .Z(n49583) );
  XOR U48778 ( .A(n49584), .B(n49512), .Z(n46676) );
  NOR U48779 ( .A(n49511), .B(n48793), .Z(n49584) );
  XNOR U48780 ( .A(n49585), .B(n49515), .Z(n49489) );
  ANDN U48781 ( .B(n48785), .A(n49514), .Z(n49585) );
  XOR U48782 ( .A(n46933), .B(n49586), .Z(n49582) );
  XOR U48783 ( .A(n46650), .B(n45859), .Z(n49586) );
  XNOR U48784 ( .A(n49587), .B(n49588), .Z(n45859) );
  ANDN U48785 ( .B(n49589), .A(n49590), .Z(n49587) );
  XOR U48786 ( .A(n49591), .B(n49520), .Z(n46650) );
  ANDN U48787 ( .B(n48780), .A(n49519), .Z(n49591) );
  XOR U48788 ( .A(n49592), .B(n49523), .Z(n46933) );
  ANDN U48789 ( .B(n48789), .A(n49522), .Z(n49592) );
  XOR U48790 ( .A(n38325), .B(n45040), .Z(n33764) );
  XNOR U48791 ( .A(n49593), .B(n44644), .Z(n45040) );
  ANDN U48792 ( .B(n41344), .A(n47601), .Z(n49593) );
  IV U48793 ( .A(n41346), .Z(n47601) );
  XNOR U48794 ( .A(n43722), .B(n48110), .Z(n41346) );
  XOR U48795 ( .A(n49594), .B(n49595), .Z(n48110) );
  XNOR U48796 ( .A(n39833), .B(n45906), .Z(n38325) );
  XNOR U48797 ( .A(n49596), .B(n49597), .Z(n45906) );
  XNOR U48798 ( .A(n40222), .B(n39288), .Z(n49597) );
  XOR U48799 ( .A(n49598), .B(n44645), .Z(n39288) );
  XNOR U48800 ( .A(n45786), .B(n46775), .Z(n44645) );
  XOR U48801 ( .A(n49599), .B(n49600), .Z(n46775) );
  ANDN U48802 ( .B(n49601), .A(n48336), .Z(n49599) );
  XOR U48803 ( .A(n49602), .B(n46450), .Z(n45786) );
  XNOR U48804 ( .A(n49603), .B(n49604), .Z(n46450) );
  XNOR U48805 ( .A(n46767), .B(n45424), .Z(n49604) );
  XNOR U48806 ( .A(n49605), .B(n49126), .Z(n45424) );
  ANDN U48807 ( .B(n47772), .A(n47773), .Z(n49605) );
  XOR U48808 ( .A(round_reg[94]), .B(n49606), .Z(n47772) );
  XNOR U48809 ( .A(n49607), .B(n49118), .Z(n46767) );
  ANDN U48810 ( .B(n47763), .A(n47765), .Z(n49607) );
  XNOR U48811 ( .A(round_reg[212]), .B(n49608), .Z(n47763) );
  XNOR U48812 ( .A(n44773), .B(n49609), .Z(n49603) );
  XNOR U48813 ( .A(n46353), .B(n47257), .Z(n49609) );
  XNOR U48814 ( .A(n49610), .B(n49129), .Z(n47257) );
  NOR U48815 ( .A(n47759), .B(n47761), .Z(n49610) );
  XOR U48816 ( .A(round_reg[8]), .B(n48699), .Z(n47759) );
  XNOR U48817 ( .A(n49611), .B(n49121), .Z(n46353) );
  XOR U48818 ( .A(round_reg[260]), .B(n49612), .Z(n47768) );
  XNOR U48819 ( .A(n49613), .B(n49614), .Z(n44773) );
  ANDN U48820 ( .B(n44644), .A(n41344), .Z(n49598) );
  XNOR U48821 ( .A(n49551), .B(n44541), .Z(n41344) );
  IV U48822 ( .A(n46194), .Z(n44541) );
  XNOR U48823 ( .A(n49615), .B(n49616), .Z(n49551) );
  NOR U48824 ( .A(n49617), .B(n47732), .Z(n49615) );
  XNOR U48825 ( .A(n44864), .B(n49618), .Z(n44644) );
  XNOR U48826 ( .A(n49619), .B(n46349), .Z(n44864) );
  XNOR U48827 ( .A(n49620), .B(n49621), .Z(n46349) );
  XNOR U48828 ( .A(n46936), .B(n43646), .Z(n49621) );
  XOR U48829 ( .A(n49622), .B(n46339), .Z(n43646) );
  XOR U48830 ( .A(round_reg[116]), .B(n49623), .Z(n46339) );
  ANDN U48831 ( .B(n48518), .A(n47337), .Z(n49622) );
  XOR U48832 ( .A(round_reg[282]), .B(n49625), .Z(n46328) );
  ANDN U48833 ( .B(n49626), .A(n48511), .Z(n49624) );
  IV U48834 ( .A(n49627), .Z(n48511) );
  XOR U48835 ( .A(n46538), .B(n49628), .Z(n49620) );
  XOR U48836 ( .A(n43101), .B(n47681), .Z(n49628) );
  XOR U48837 ( .A(n49629), .B(n46325), .Z(n47681) );
  XOR U48838 ( .A(round_reg[234]), .B(n48564), .Z(n46325) );
  NOR U48839 ( .A(n47339), .B(n48515), .Z(n49629) );
  XOR U48840 ( .A(n49630), .B(n47353), .Z(n43101) );
  XOR U48841 ( .A(round_reg[175]), .B(n49631), .Z(n47353) );
  ANDN U48842 ( .B(n48521), .A(n48502), .Z(n49630) );
  XNOR U48843 ( .A(n49632), .B(n46335), .Z(n46538) );
  XNOR U48844 ( .A(round_reg[30]), .B(n49633), .Z(n46335) );
  NOR U48845 ( .A(n48509), .B(n47333), .Z(n49632) );
  XOR U48846 ( .A(n49634), .B(n44655), .Z(n40222) );
  XOR U48847 ( .A(n49635), .B(n42662), .Z(n44655) );
  IV U48848 ( .A(n44186), .Z(n42662) );
  ANDN U48849 ( .B(n44654), .A(n41349), .Z(n49634) );
  XOR U48850 ( .A(n46166), .B(n49636), .Z(n41349) );
  XOR U48851 ( .A(n49637), .B(n49638), .Z(n46913) );
  XNOR U48852 ( .A(n42549), .B(n46001), .Z(n49638) );
  XOR U48853 ( .A(n49639), .B(n49640), .Z(n46001) );
  ANDN U48854 ( .B(n49641), .A(n49642), .Z(n49639) );
  XNOR U48855 ( .A(n49643), .B(n49402), .Z(n42549) );
  ANDN U48856 ( .B(n49644), .A(n49645), .Z(n49643) );
  XOR U48857 ( .A(n45895), .B(n49646), .Z(n49637) );
  XOR U48858 ( .A(n45981), .B(n46724), .Z(n49646) );
  XNOR U48859 ( .A(n49647), .B(n49408), .Z(n46724) );
  NOR U48860 ( .A(n49648), .B(n49649), .Z(n49647) );
  XNOR U48861 ( .A(n49650), .B(n49651), .Z(n45981) );
  ANDN U48862 ( .B(n49652), .A(n49653), .Z(n49650) );
  XNOR U48863 ( .A(n49654), .B(n49411), .Z(n45895) );
  NOR U48864 ( .A(n49655), .B(n49656), .Z(n49654) );
  XNOR U48865 ( .A(n49657), .B(n49658), .Z(n46706) );
  XOR U48866 ( .A(n46310), .B(n45010), .Z(n49658) );
  XOR U48867 ( .A(n49659), .B(n48670), .Z(n45010) );
  XNOR U48868 ( .A(n49661), .B(n48674), .Z(n46310) );
  XOR U48869 ( .A(n47811), .B(n49663), .Z(n49657) );
  XOR U48870 ( .A(n47169), .B(n48664), .Z(n49663) );
  XNOR U48871 ( .A(n49664), .B(n48680), .Z(n48664) );
  ANDN U48872 ( .B(n48681), .A(n49665), .Z(n49664) );
  XNOR U48873 ( .A(n49666), .B(n49667), .Z(n47169) );
  ANDN U48874 ( .B(n49668), .A(n49669), .Z(n49666) );
  XOR U48875 ( .A(n49670), .B(n48685), .Z(n47811) );
  NOR U48876 ( .A(n48684), .B(n49671), .Z(n49670) );
  IV U48877 ( .A(n49672), .Z(n48684) );
  XNOR U48878 ( .A(n48388), .B(n46501), .Z(n44654) );
  XOR U48879 ( .A(n49673), .B(n47699), .Z(n46501) );
  XNOR U48880 ( .A(n49674), .B(n49675), .Z(n47699) );
  XNOR U48881 ( .A(n44514), .B(n45888), .Z(n49675) );
  XOR U48882 ( .A(n49676), .B(n49677), .Z(n45888) );
  ANDN U48883 ( .B(n48826), .A(n49678), .Z(n49676) );
  XNOR U48884 ( .A(n49679), .B(n49680), .Z(n44514) );
  ANDN U48885 ( .B(n49681), .A(n49682), .Z(n49679) );
  XOR U48886 ( .A(n46750), .B(n49683), .Z(n49674) );
  XOR U48887 ( .A(n48813), .B(n43601), .Z(n49683) );
  XNOR U48888 ( .A(n49684), .B(n49685), .Z(n43601) );
  ANDN U48889 ( .B(n49686), .A(n48820), .Z(n49684) );
  XNOR U48890 ( .A(n49687), .B(n49688), .Z(n48813) );
  NOR U48891 ( .A(n48833), .B(n49689), .Z(n49687) );
  XNOR U48892 ( .A(n49690), .B(n48830), .Z(n46750) );
  NOR U48893 ( .A(n48829), .B(n49691), .Z(n49690) );
  XNOR U48894 ( .A(n49692), .B(n47045), .Z(n48388) );
  ANDN U48895 ( .B(n49693), .A(n49694), .Z(n49692) );
  XOR U48896 ( .A(n40197), .B(n49695), .Z(n49596) );
  XOR U48897 ( .A(n37886), .B(n38586), .Z(n49695) );
  XOR U48898 ( .A(n44659), .B(n47224), .Z(n44651) );
  XOR U48899 ( .A(n49697), .B(n49698), .Z(n47224) );
  ANDN U48900 ( .B(n49699), .A(n49700), .Z(n49697) );
  ANDN U48901 ( .B(n44652), .A(n41357), .Z(n49696) );
  XOR U48902 ( .A(n49701), .B(n45673), .Z(n41357) );
  XNOR U48903 ( .A(n49702), .B(n43327), .Z(n44652) );
  XOR U48904 ( .A(n49703), .B(n44648), .Z(n37886) );
  XOR U48905 ( .A(n49704), .B(n44741), .Z(n44648) );
  IV U48906 ( .A(n45123), .Z(n44741) );
  XOR U48907 ( .A(n49705), .B(n46920), .Z(n45123) );
  XNOR U48908 ( .A(n49706), .B(n49707), .Z(n46920) );
  XOR U48909 ( .A(n42671), .B(n46575), .Z(n49707) );
  XOR U48910 ( .A(n49708), .B(n47988), .Z(n46575) );
  XNOR U48911 ( .A(n49711), .B(n47982), .Z(n42671) );
  XOR U48912 ( .A(n46693), .B(n49714), .Z(n49706) );
  XOR U48913 ( .A(n43771), .B(n43339), .Z(n49714) );
  XNOR U48914 ( .A(n49715), .B(n47978), .Z(n43339) );
  NOR U48915 ( .A(n49716), .B(n49717), .Z(n49715) );
  XNOR U48916 ( .A(n49718), .B(n49719), .Z(n43771) );
  XNOR U48917 ( .A(n49722), .B(n49723), .Z(n46693) );
  ANDN U48918 ( .B(n44649), .A(n41340), .Z(n49703) );
  XOR U48919 ( .A(n49727), .B(n46414), .Z(n44649) );
  XOR U48920 ( .A(n48468), .B(n46873), .Z(n46414) );
  XNOR U48921 ( .A(n49728), .B(n49729), .Z(n46873) );
  XNOR U48922 ( .A(n48084), .B(n41593), .Z(n49729) );
  XOR U48923 ( .A(n49730), .B(n49731), .Z(n41593) );
  ANDN U48924 ( .B(n49732), .A(n49733), .Z(n49730) );
  XOR U48925 ( .A(n49734), .B(n49735), .Z(n48084) );
  ANDN U48926 ( .B(n49736), .A(n49737), .Z(n49734) );
  XNOR U48927 ( .A(n45711), .B(n49738), .Z(n49728) );
  XNOR U48928 ( .A(n44878), .B(n44322), .Z(n49738) );
  XNOR U48929 ( .A(n49739), .B(n49740), .Z(n44322) );
  ANDN U48930 ( .B(n49741), .A(n49742), .Z(n49739) );
  XNOR U48931 ( .A(n49743), .B(n49744), .Z(n44878) );
  NOR U48932 ( .A(n49745), .B(n49746), .Z(n49743) );
  XNOR U48933 ( .A(n49747), .B(n49748), .Z(n45711) );
  ANDN U48934 ( .B(n49749), .A(n49750), .Z(n49747) );
  XOR U48935 ( .A(n49751), .B(n49752), .Z(n48468) );
  XNOR U48936 ( .A(n46585), .B(n45219), .Z(n49752) );
  XNOR U48937 ( .A(n49753), .B(n49754), .Z(n45219) );
  NOR U48938 ( .A(n49755), .B(n49756), .Z(n49753) );
  XNOR U48939 ( .A(n49757), .B(n49758), .Z(n46585) );
  NOR U48940 ( .A(n49759), .B(n49760), .Z(n49757) );
  XNOR U48941 ( .A(n43328), .B(n49761), .Z(n49751) );
  XOR U48942 ( .A(n45178), .B(n49762), .Z(n49761) );
  XNOR U48943 ( .A(n49763), .B(n49764), .Z(n45178) );
  NOR U48944 ( .A(n49765), .B(n49766), .Z(n49763) );
  XNOR U48945 ( .A(n49767), .B(n49768), .Z(n43328) );
  NOR U48946 ( .A(n49769), .B(n49770), .Z(n49767) );
  XOR U48947 ( .A(n49771), .B(n44642), .Z(n40197) );
  XNOR U48948 ( .A(n49772), .B(n44410), .Z(n44642) );
  XOR U48949 ( .A(n49773), .B(n49774), .Z(n46850) );
  XNOR U48950 ( .A(n46515), .B(n45258), .Z(n49774) );
  XOR U48951 ( .A(n49775), .B(n47511), .Z(n45258) );
  ANDN U48952 ( .B(n47512), .A(n47859), .Z(n49775) );
  XNOR U48953 ( .A(n49776), .B(n47501), .Z(n46515) );
  ANDN U48954 ( .B(n47502), .A(n47856), .Z(n49776) );
  XNOR U48955 ( .A(n45421), .B(n49777), .Z(n49773) );
  XOR U48956 ( .A(n45309), .B(n44679), .Z(n49777) );
  XOR U48957 ( .A(n49778), .B(n47498), .Z(n44679) );
  NOR U48958 ( .A(n47867), .B(n47497), .Z(n49778) );
  XOR U48959 ( .A(n49779), .B(n47508), .Z(n45309) );
  NOR U48960 ( .A(n47870), .B(n47507), .Z(n49779) );
  XNOR U48961 ( .A(n49780), .B(n49781), .Z(n45421) );
  NOR U48962 ( .A(n47863), .B(n49782), .Z(n49780) );
  ANDN U48963 ( .B(n44641), .A(n41353), .Z(n49771) );
  XOR U48964 ( .A(n45778), .B(n47292), .Z(n41353) );
  XNOR U48965 ( .A(n49784), .B(n48347), .Z(n47292) );
  NOR U48966 ( .A(n49223), .B(n49222), .Z(n49784) );
  IV U48967 ( .A(n46421), .Z(n45778) );
  XOR U48968 ( .A(n49785), .B(n49353), .Z(n46421) );
  XOR U48969 ( .A(n49786), .B(n49787), .Z(n49353) );
  XOR U48970 ( .A(n44861), .B(n46391), .Z(n49787) );
  XOR U48971 ( .A(n49788), .B(n47365), .Z(n46391) );
  XOR U48972 ( .A(round_reg[536]), .B(n49789), .Z(n48082) );
  XOR U48973 ( .A(round_reg[898]), .B(n49790), .Z(n47366) );
  XNOR U48974 ( .A(n49791), .B(n47369), .Z(n44861) );
  ANDN U48975 ( .B(n47370), .A(n47587), .Z(n49791) );
  XOR U48976 ( .A(round_reg[432]), .B(n49178), .Z(n47587) );
  XOR U48977 ( .A(round_reg[794]), .B(n49792), .Z(n47370) );
  XOR U48978 ( .A(n47073), .B(n49793), .Z(n49786) );
  XOR U48979 ( .A(n46527), .B(n47359), .Z(n49793) );
  XNOR U48980 ( .A(n49794), .B(n47378), .Z(n47359) );
  XOR U48981 ( .A(round_reg[502]), .B(n49795), .Z(n47297) );
  XOR U48982 ( .A(round_reg[891]), .B(n49080), .Z(n47296) );
  XNOR U48983 ( .A(n49796), .B(n48346), .Z(n46527) );
  XOR U48984 ( .A(round_reg[670]), .B(n49797), .Z(n48347) );
  XNOR U48985 ( .A(round_reg[604]), .B(n49798), .Z(n49222) );
  XNOR U48986 ( .A(n49799), .B(n47375), .Z(n47073) );
  XNOR U48987 ( .A(round_reg[381]), .B(n49800), .Z(n47290) );
  XOR U48988 ( .A(round_reg[748]), .B(n49801), .Z(n47289) );
  XNOR U48989 ( .A(n47751), .B(n46054), .Z(n44641) );
  XNOR U48990 ( .A(n49802), .B(n49803), .Z(n47751) );
  ANDN U48991 ( .B(n49804), .A(n49805), .Z(n49802) );
  XOR U48992 ( .A(n49806), .B(n49807), .Z(n39833) );
  XNOR U48993 ( .A(n38632), .B(n40094), .Z(n49807) );
  XOR U48994 ( .A(n49808), .B(n40238), .Z(n40094) );
  XOR U48995 ( .A(n48778), .B(n42691), .Z(n40238) );
  XNOR U48996 ( .A(n49809), .B(n48196), .Z(n42691) );
  XOR U48997 ( .A(n49810), .B(n49811), .Z(n48196) );
  XNOR U48998 ( .A(n49812), .B(n46316), .Z(n49811) );
  XNOR U48999 ( .A(n49813), .B(n49500), .Z(n46316) );
  ANDN U49000 ( .B(n49464), .A(n49462), .Z(n49813) );
  XOR U49001 ( .A(n43915), .B(n49814), .Z(n49810) );
  XOR U49002 ( .A(n46033), .B(n47139), .Z(n49814) );
  XOR U49003 ( .A(n49815), .B(n49496), .Z(n47139) );
  ANDN U49004 ( .B(n49456), .A(n49454), .Z(n49815) );
  XOR U49005 ( .A(n49816), .B(n49506), .Z(n46033) );
  XOR U49006 ( .A(n49817), .B(n49493), .Z(n43915) );
  ANDN U49007 ( .B(n49451), .A(n49449), .Z(n49817) );
  XOR U49008 ( .A(n49818), .B(n49589), .Z(n48778) );
  ANDN U49009 ( .B(n49819), .A(n49820), .Z(n49818) );
  NOR U49010 ( .A(n40237), .B(n45332), .Z(n49808) );
  XOR U49011 ( .A(n49821), .B(n43767), .Z(n45332) );
  XNOR U49012 ( .A(n49822), .B(n42157), .Z(n40237) );
  XOR U49013 ( .A(n47459), .B(n49823), .Z(n42157) );
  XNOR U49014 ( .A(n49824), .B(n49825), .Z(n47459) );
  XNOR U49015 ( .A(n44683), .B(n47598), .Z(n49825) );
  XNOR U49016 ( .A(n49826), .B(n48181), .Z(n47598) );
  XOR U49017 ( .A(round_reg[401]), .B(n49827), .Z(n48181) );
  NOR U49018 ( .A(n49828), .B(n48882), .Z(n49826) );
  XOR U49019 ( .A(n49829), .B(n48170), .Z(n44683) );
  XOR U49020 ( .A(round_reg[350]), .B(n49633), .Z(n48170) );
  ANDN U49021 ( .B(n47625), .A(n48870), .Z(n49829) );
  XOR U49022 ( .A(n48865), .B(n49830), .Z(n49824) );
  XOR U49023 ( .A(n44487), .B(n47400), .Z(n49830) );
  XOR U49024 ( .A(n49831), .B(n48175), .Z(n47400) );
  XOR U49025 ( .A(round_reg[637]), .B(n49087), .Z(n48175) );
  XNOR U49026 ( .A(n49832), .B(n48172), .Z(n44487) );
  XOR U49027 ( .A(round_reg[471]), .B(n49833), .Z(n48172) );
  ANDN U49028 ( .B(n47621), .A(n48877), .Z(n49832) );
  IV U49029 ( .A(n49834), .Z(n48877) );
  XNOR U49030 ( .A(n49835), .B(n48178), .Z(n48865) );
  XOR U49031 ( .A(round_reg[569]), .B(n49836), .Z(n48178) );
  NOR U49032 ( .A(n47612), .B(n48873), .Z(n49835) );
  XOR U49033 ( .A(n49837), .B(n43291), .Z(n38632) );
  IV U49034 ( .A(n40229), .Z(n43291) );
  XOR U49035 ( .A(n49318), .B(n45371), .Z(n40229) );
  XNOR U49036 ( .A(n49838), .B(n49839), .Z(n48107) );
  XOR U49037 ( .A(n47679), .B(n49840), .Z(n49839) );
  XNOR U49038 ( .A(n49841), .B(n49842), .Z(n47679) );
  ANDN U49039 ( .B(n49295), .A(n49297), .Z(n49841) );
  XNOR U49040 ( .A(n49843), .B(n49844), .Z(n49838) );
  XOR U49041 ( .A(n48503), .B(n44505), .Z(n49844) );
  XOR U49042 ( .A(n49845), .B(n49846), .Z(n44505) );
  NOR U49043 ( .A(n49847), .B(n49293), .Z(n49845) );
  XNOR U49044 ( .A(n49848), .B(n49849), .Z(n48503) );
  ANDN U49045 ( .B(n49308), .A(n49850), .Z(n49848) );
  XNOR U49046 ( .A(n49851), .B(n49852), .Z(n48349) );
  XOR U49047 ( .A(n46300), .B(n44942), .Z(n49852) );
  XOR U49048 ( .A(n49853), .B(n49205), .Z(n44942) );
  NOR U49049 ( .A(n49204), .B(n49314), .Z(n49853) );
  XOR U49050 ( .A(round_reg[793]), .B(n49854), .Z(n49204) );
  XNOR U49051 ( .A(n49855), .B(n48499), .Z(n46300) );
  XOR U49052 ( .A(round_reg[1008]), .B(n49856), .Z(n48499) );
  ANDN U49053 ( .B(n49210), .A(n49321), .Z(n49855) );
  XOR U49054 ( .A(round_reg[897]), .B(n49857), .Z(n49210) );
  XOR U49055 ( .A(n46821), .B(n49858), .Z(n49851) );
  XOR U49056 ( .A(n43764), .B(n47242), .Z(n49858) );
  XNOR U49057 ( .A(n49859), .B(n46048), .Z(n47242) );
  XOR U49058 ( .A(round_reg[1248]), .B(n49860), .Z(n46048) );
  ANDN U49059 ( .B(n49324), .A(n49323), .Z(n49859) );
  XOR U49060 ( .A(round_reg[890]), .B(n49861), .Z(n49323) );
  XNOR U49061 ( .A(n49862), .B(n47020), .Z(n43764) );
  XOR U49062 ( .A(round_reg[1037]), .B(n49863), .Z(n47020) );
  NOR U49063 ( .A(n49864), .B(n49207), .Z(n49862) );
  XNOR U49064 ( .A(n49865), .B(n46052), .Z(n46821) );
  XOR U49065 ( .A(round_reg[1150]), .B(n49866), .Z(n46052) );
  NOR U49066 ( .A(n49212), .B(n49317), .Z(n49865) );
  XOR U49067 ( .A(round_reg[747]), .B(n49867), .Z(n49212) );
  XNOR U49068 ( .A(n49868), .B(n49207), .Z(n49318) );
  XOR U49069 ( .A(round_reg[669]), .B(n49869), .Z(n49207) );
  ANDN U49070 ( .B(n49864), .A(n47018), .Z(n49868) );
  NOR U49071 ( .A(n40228), .B(n42596), .Z(n49837) );
  XOR U49072 ( .A(n49870), .B(n43671), .Z(n42596) );
  XNOR U49073 ( .A(n49871), .B(n49872), .Z(n46583) );
  XNOR U49074 ( .A(n45132), .B(n44865), .Z(n49872) );
  XNOR U49075 ( .A(n49873), .B(n48535), .Z(n44865) );
  ANDN U49076 ( .B(n49874), .A(n49386), .Z(n49873) );
  XNOR U49077 ( .A(n49875), .B(n48527), .Z(n45132) );
  ANDN U49078 ( .B(n49876), .A(n49377), .Z(n49875) );
  XOR U49079 ( .A(n47472), .B(n49877), .Z(n49871) );
  XOR U49080 ( .A(n49347), .B(n49618), .Z(n49877) );
  XNOR U49081 ( .A(n49878), .B(n48543), .Z(n49618) );
  ANDN U49082 ( .B(n49879), .A(n49382), .Z(n49878) );
  XNOR U49083 ( .A(n49880), .B(n48530), .Z(n49347) );
  ANDN U49084 ( .B(n49881), .A(n49379), .Z(n49880) );
  XNOR U49085 ( .A(n49882), .B(n48539), .Z(n47472) );
  IV U49086 ( .A(n49883), .Z(n48539) );
  ANDN U49087 ( .B(n49884), .A(n49384), .Z(n49882) );
  XOR U49088 ( .A(n48248), .B(n43825), .Z(n40228) );
  IV U49089 ( .A(n44588), .Z(n43825) );
  XOR U49090 ( .A(n49886), .B(n49887), .Z(n48248) );
  AND U49091 ( .A(n49888), .B(n49889), .Z(n49886) );
  XOR U49092 ( .A(n39030), .B(n49890), .Z(n49806) );
  XOR U49093 ( .A(n36433), .B(n37671), .Z(n49890) );
  XNOR U49094 ( .A(n49891), .B(n40246), .Z(n37671) );
  XNOR U49095 ( .A(n46991), .B(n44009), .Z(n40246) );
  XNOR U49096 ( .A(n46698), .B(n49892), .Z(n44009) );
  XOR U49097 ( .A(n49893), .B(n49894), .Z(n46698) );
  XNOR U49098 ( .A(n45984), .B(n46849), .Z(n49894) );
  XOR U49099 ( .A(n49895), .B(n49782), .Z(n46849) );
  ANDN U49100 ( .B(n47863), .A(n47864), .Z(n49895) );
  XOR U49101 ( .A(round_reg[495]), .B(n49631), .Z(n47863) );
  XNOR U49102 ( .A(n49896), .B(n47512), .Z(n45984) );
  XNOR U49103 ( .A(round_reg[955]), .B(n49897), .Z(n47512) );
  ANDN U49104 ( .B(n47859), .A(n47860), .Z(n49896) );
  XOR U49105 ( .A(round_reg[529]), .B(n49898), .Z(n47859) );
  XNOR U49106 ( .A(n44507), .B(n49899), .Z(n49893) );
  XNOR U49107 ( .A(n43302), .B(n45719), .Z(n49899) );
  XNOR U49108 ( .A(n49900), .B(n47502), .Z(n45719) );
  XOR U49109 ( .A(round_reg[741]), .B(n49901), .Z(n47502) );
  ANDN U49110 ( .B(n47856), .A(n47857), .Z(n49900) );
  XNOR U49111 ( .A(round_reg[374]), .B(n49902), .Z(n47856) );
  XNOR U49112 ( .A(n49903), .B(n47497), .Z(n43302) );
  XOR U49113 ( .A(round_reg[787]), .B(n49904), .Z(n47497) );
  ANDN U49114 ( .B(n47867), .A(n47868), .Z(n49903) );
  XOR U49115 ( .A(round_reg[425]), .B(n49905), .Z(n47867) );
  XNOR U49116 ( .A(n49906), .B(n47507), .Z(n44507) );
  XNOR U49117 ( .A(round_reg[663]), .B(n48554), .Z(n47507) );
  ANDN U49118 ( .B(n47870), .A(n47871), .Z(n49906) );
  XNOR U49119 ( .A(round_reg[597]), .B(n49907), .Z(n47870) );
  XNOR U49120 ( .A(n49908), .B(n49909), .Z(n46991) );
  NOR U49121 ( .A(n49910), .B(n49911), .Z(n49908) );
  NOR U49122 ( .A(n40245), .B(n42604), .Z(n49891) );
  XOR U49123 ( .A(n45145), .B(n49912), .Z(n42604) );
  XOR U49124 ( .A(n45630), .B(n49913), .Z(n40245) );
  XNOR U49125 ( .A(n46038), .B(n49472), .Z(n45630) );
  XNOR U49126 ( .A(n49914), .B(n49915), .Z(n49472) );
  XOR U49127 ( .A(n49916), .B(n48318), .Z(n49915) );
  XOR U49128 ( .A(n49917), .B(n47658), .Z(n48318) );
  AND U49129 ( .A(n48114), .B(n49918), .Z(n49917) );
  XNOR U49130 ( .A(n47783), .B(n49919), .Z(n49914) );
  XOR U49131 ( .A(n47740), .B(n47406), .Z(n49919) );
  XNOR U49132 ( .A(n49920), .B(n47652), .Z(n47406) );
  ANDN U49133 ( .B(n49921), .A(n49595), .Z(n49920) );
  XNOR U49134 ( .A(n49922), .B(n47661), .Z(n47740) );
  ANDN U49135 ( .B(n49923), .A(n48116), .Z(n49922) );
  XNOR U49136 ( .A(n49924), .B(n47648), .Z(n47783) );
  AND U49137 ( .A(n49925), .B(n49926), .Z(n49924) );
  XOR U49138 ( .A(n49927), .B(n49928), .Z(n46038) );
  XNOR U49139 ( .A(n45520), .B(n46106), .Z(n49928) );
  XNOR U49140 ( .A(n49929), .B(n49302), .Z(n46106) );
  XNOR U49141 ( .A(n49932), .B(n49296), .Z(n45520) );
  XOR U49142 ( .A(n42152), .B(n49934), .Z(n49927) );
  XNOR U49143 ( .A(n44928), .B(n46410), .Z(n49934) );
  XNOR U49144 ( .A(n49935), .B(n49310), .Z(n46410) );
  AND U49145 ( .A(n49849), .B(n49936), .Z(n49935) );
  XNOR U49146 ( .A(n49937), .B(n49292), .Z(n44928) );
  ANDN U49147 ( .B(n49938), .A(n49846), .Z(n49937) );
  XNOR U49148 ( .A(n49939), .B(n49305), .Z(n42152) );
  ANDN U49149 ( .B(n49940), .A(n49941), .Z(n49939) );
  XOR U49150 ( .A(n49942), .B(n40242), .Z(n36433) );
  XOR U49151 ( .A(n48677), .B(n45519), .Z(n40242) );
  XNOR U49152 ( .A(n49943), .B(n49944), .Z(n49395) );
  XOR U49153 ( .A(n41739), .B(n45694), .Z(n49944) );
  XOR U49154 ( .A(n49945), .B(n49946), .Z(n45694) );
  AND U49155 ( .A(n48685), .B(n48683), .Z(n49945) );
  XOR U49156 ( .A(round_reg[1129]), .B(n49947), .Z(n48685) );
  XNOR U49157 ( .A(n49948), .B(n49949), .Z(n41739) );
  ANDN U49158 ( .B(n49950), .A(n49667), .Z(n49948) );
  XNOR U49159 ( .A(n49435), .B(n49951), .Z(n49943) );
  XNOR U49160 ( .A(n46070), .B(n49952), .Z(n49951) );
  XOR U49161 ( .A(n49953), .B(n49954), .Z(n46070) );
  ANDN U49162 ( .B(n48669), .A(n48670), .Z(n49953) );
  XOR U49163 ( .A(round_reg[987]), .B(n49955), .Z(n48670) );
  XOR U49164 ( .A(n49956), .B(n49957), .Z(n49435) );
  ANDN U49165 ( .B(n48673), .A(n48674), .Z(n49956) );
  XNOR U49166 ( .A(round_reg[1155]), .B(n49958), .Z(n48674) );
  XNOR U49167 ( .A(n49959), .B(n49960), .Z(n46584) );
  XNOR U49168 ( .A(n46419), .B(n45505), .Z(n49960) );
  XNOR U49169 ( .A(n49961), .B(n49962), .Z(n45505) );
  ANDN U49170 ( .B(n49963), .A(n49532), .Z(n49961) );
  XNOR U49171 ( .A(n49964), .B(n49965), .Z(n46419) );
  ANDN U49172 ( .B(n49966), .A(n49967), .Z(n49964) );
  XOR U49173 ( .A(n46718), .B(n49968), .Z(n49959) );
  XOR U49174 ( .A(n46264), .B(n49969), .Z(n49968) );
  XNOR U49175 ( .A(n49970), .B(n49971), .Z(n46264) );
  ANDN U49176 ( .B(n49972), .A(n49371), .Z(n49970) );
  XNOR U49177 ( .A(n49973), .B(n49974), .Z(n46718) );
  ANDN U49178 ( .B(n49975), .A(n49360), .Z(n49973) );
  XNOR U49179 ( .A(n49976), .B(n49950), .Z(n48677) );
  ANDN U49180 ( .B(n49667), .A(n49668), .Z(n49976) );
  XNOR U49181 ( .A(round_reg[1080]), .B(n49977), .Z(n49667) );
  ANDN U49182 ( .B(n40241), .A(n42608), .Z(n49942) );
  XNOR U49183 ( .A(n49978), .B(n49673), .Z(n45569) );
  XNOR U49184 ( .A(n49979), .B(n49980), .Z(n49673) );
  XOR U49185 ( .A(n47035), .B(n46060), .Z(n49980) );
  XOR U49186 ( .A(n49981), .B(n47054), .Z(n46060) );
  ANDN U49187 ( .B(n47055), .A(n48391), .Z(n49981) );
  XNOR U49188 ( .A(round_reg[44]), .B(n49982), .Z(n47055) );
  XNOR U49189 ( .A(n49983), .B(n47040), .Z(n47035) );
  ANDN U49190 ( .B(n47041), .A(n48983), .Z(n49983) );
  XNOR U49191 ( .A(round_reg[296]), .B(n49984), .Z(n47041) );
  XOR U49192 ( .A(n46368), .B(n49985), .Z(n49979) );
  XOR U49193 ( .A(n40848), .B(n43456), .Z(n49985) );
  XNOR U49194 ( .A(n49986), .B(n49987), .Z(n43456) );
  ANDN U49195 ( .B(n48394), .A(n48395), .Z(n49986) );
  XNOR U49196 ( .A(n49988), .B(n47044), .Z(n40848) );
  ANDN U49197 ( .B(n47045), .A(n49693), .Z(n49988) );
  XNOR U49198 ( .A(round_reg[66]), .B(n49989), .Z(n47045) );
  XNOR U49199 ( .A(n49990), .B(n47050), .Z(n46368) );
  ANDN U49200 ( .B(n47051), .A(n49991), .Z(n49990) );
  XOR U49201 ( .A(round_reg[189]), .B(n49992), .Z(n47051) );
  XNOR U49202 ( .A(n49993), .B(n49563), .Z(n48379) );
  ANDN U49203 ( .B(n49994), .A(n47101), .Z(n49993) );
  XOR U49204 ( .A(n49995), .B(n45673), .Z(n40241) );
  IV U49205 ( .A(n45415), .Z(n45673) );
  XNOR U49206 ( .A(n49998), .B(n43278), .Z(n39030) );
  IV U49207 ( .A(n40233), .Z(n43278) );
  XOR U49208 ( .A(n49999), .B(n44492), .Z(n40233) );
  IV U49209 ( .A(n41588), .Z(n44492) );
  XOR U49210 ( .A(n47721), .B(n50000), .Z(n41588) );
  XOR U49211 ( .A(n50001), .B(n50002), .Z(n47721) );
  XNOR U49212 ( .A(n44810), .B(n47096), .Z(n50002) );
  XNOR U49213 ( .A(n50003), .B(n49759), .Z(n47096) );
  XNOR U49214 ( .A(n50006), .B(n49770), .Z(n44810) );
  ANDN U49215 ( .B(n50007), .A(n50008), .Z(n50006) );
  XNOR U49216 ( .A(n45245), .B(n50009), .Z(n50001) );
  XOR U49217 ( .A(n46499), .B(n45286), .Z(n50009) );
  XOR U49218 ( .A(n50010), .B(n49766), .Z(n45286) );
  ANDN U49219 ( .B(n50011), .A(n50012), .Z(n50010) );
  XNOR U49220 ( .A(n50013), .B(n50014), .Z(n46499) );
  ANDN U49221 ( .B(n50015), .A(n50016), .Z(n50013) );
  XOR U49222 ( .A(n50017), .B(n49756), .Z(n45245) );
  NOR U49223 ( .A(n50018), .B(n50019), .Z(n50017) );
  ANDN U49224 ( .B(n42599), .A(n40232), .Z(n49998) );
  XOR U49225 ( .A(n49475), .B(n45249), .Z(n40232) );
  XOR U49226 ( .A(n45427), .B(n50020), .Z(n45249) );
  XOR U49227 ( .A(n50021), .B(n50022), .Z(n45427) );
  XNOR U49228 ( .A(n49701), .B(n49995), .Z(n50022) );
  XNOR U49229 ( .A(n50023), .B(n48754), .Z(n49995) );
  ANDN U49230 ( .B(n50024), .A(n50025), .Z(n50023) );
  XNOR U49231 ( .A(n50026), .B(n48759), .Z(n49701) );
  IV U49232 ( .A(n50027), .Z(n48759) );
  NOR U49233 ( .A(n50028), .B(n50029), .Z(n50026) );
  XOR U49234 ( .A(n45414), .B(n50030), .Z(n50021) );
  XOR U49235 ( .A(n45847), .B(n45672), .Z(n50030) );
  XNOR U49236 ( .A(n50031), .B(n48745), .Z(n45672) );
  ANDN U49237 ( .B(n50032), .A(n50033), .Z(n50031) );
  XNOR U49238 ( .A(n50034), .B(n50035), .Z(n45847) );
  XNOR U49239 ( .A(n50038), .B(n48749), .Z(n45414) );
  ANDN U49240 ( .B(n50039), .A(n50040), .Z(n50038) );
  XNOR U49241 ( .A(n50041), .B(n50042), .Z(n49475) );
  XOR U49242 ( .A(n31711), .B(n50043), .Z(n50042) );
  NANDN U49243 ( .A(n48733), .B(n50044), .Z(n50043) );
  ANDN U49244 ( .B(n4687), .A(rc_i[2]), .Z(n31711) );
  XOR U49245 ( .A(n47749), .B(n46054), .Z(n42599) );
  IV U49246 ( .A(n45236), .Z(n46054) );
  XOR U49247 ( .A(n46451), .B(n48017), .Z(n45236) );
  XNOR U49248 ( .A(n50045), .B(n50046), .Z(n48017) );
  XNOR U49249 ( .A(n45359), .B(n42320), .Z(n50046) );
  XOR U49250 ( .A(n50047), .B(n50048), .Z(n42320) );
  NOR U49251 ( .A(n48610), .B(n48609), .Z(n50047) );
  XOR U49252 ( .A(n50049), .B(n47421), .Z(n45359) );
  ANDN U49253 ( .B(n48620), .A(n48621), .Z(n50049) );
  XNOR U49254 ( .A(n46290), .B(n50050), .Z(n50045) );
  XNOR U49255 ( .A(n45160), .B(n44692), .Z(n50050) );
  XOR U49256 ( .A(n50051), .B(n47430), .Z(n44692) );
  ANDN U49257 ( .B(n48617), .A(n48618), .Z(n50051) );
  XNOR U49258 ( .A(n50052), .B(n47434), .Z(n45160) );
  ANDN U49259 ( .B(n48606), .A(n48607), .Z(n50052) );
  XOR U49260 ( .A(n50053), .B(n47426), .Z(n46290) );
  ANDN U49261 ( .B(n48614), .A(n48615), .Z(n50053) );
  XOR U49262 ( .A(n50054), .B(n50055), .Z(n46451) );
  XNOR U49263 ( .A(n50056), .B(n46124), .Z(n50055) );
  XOR U49264 ( .A(n50057), .B(n50058), .Z(n46124) );
  ANDN U49265 ( .B(n47753), .A(n47755), .Z(n50057) );
  XNOR U49266 ( .A(n48546), .B(n50059), .Z(n50054) );
  XNOR U49267 ( .A(n44198), .B(n47808), .Z(n50059) );
  XOR U49268 ( .A(n50060), .B(n50061), .Z(n47808) );
  ANDN U49269 ( .B(n50062), .A(n50063), .Z(n50060) );
  XNOR U49270 ( .A(n50064), .B(n50065), .Z(n44198) );
  ANDN U49271 ( .B(n49803), .A(n49804), .Z(n50064) );
  XOR U49272 ( .A(n50066), .B(n50067), .Z(n48546) );
  ANDN U49273 ( .B(n47746), .A(n47748), .Z(n50066) );
  XNOR U49274 ( .A(n50068), .B(n50062), .Z(n47749) );
  XOR U49275 ( .A(n50070), .B(n33752), .Z(n32979) );
  XOR U49276 ( .A(n39603), .B(n40977), .Z(n33752) );
  XNOR U49277 ( .A(n50071), .B(n44994), .Z(n40977) );
  ANDN U49278 ( .B(n48572), .A(n43257), .Z(n50071) );
  XOR U49279 ( .A(n43559), .B(n50072), .Z(n43257) );
  XNOR U49280 ( .A(n41995), .B(n41374), .Z(n39603) );
  XNOR U49281 ( .A(n50073), .B(n50074), .Z(n41374) );
  XNOR U49282 ( .A(n38864), .B(n39283), .Z(n50074) );
  XNOR U49283 ( .A(n50075), .B(n43270), .Z(n39283) );
  XOR U49284 ( .A(n45565), .B(n50076), .Z(n43270) );
  XNOR U49285 ( .A(n48189), .B(n49783), .Z(n45565) );
  XOR U49286 ( .A(n50077), .B(n50078), .Z(n49783) );
  XNOR U49287 ( .A(n47480), .B(n44881), .Z(n50078) );
  XNOR U49288 ( .A(n50079), .B(n47491), .Z(n44881) );
  IV U49289 ( .A(n50080), .Z(n47491) );
  ANDN U49290 ( .B(n47492), .A(n46993), .Z(n50079) );
  XOR U49291 ( .A(n50081), .B(n48464), .Z(n47480) );
  ANDN U49292 ( .B(n48463), .A(n49389), .Z(n50081) );
  XNOR U49293 ( .A(n46922), .B(n50082), .Z(n50077) );
  XNOR U49294 ( .A(n46887), .B(n46283), .Z(n50082) );
  XNOR U49295 ( .A(n50083), .B(n47486), .Z(n46283) );
  NOR U49296 ( .A(n46986), .B(n47485), .Z(n50083) );
  XOR U49297 ( .A(n50084), .B(n50085), .Z(n46887) );
  ANDN U49298 ( .B(n50086), .A(n49909), .Z(n50084) );
  XOR U49299 ( .A(n50087), .B(n50088), .Z(n46922) );
  ANDN U49300 ( .B(n50089), .A(n46982), .Z(n50087) );
  XOR U49301 ( .A(n50090), .B(n50091), .Z(n48189) );
  XOR U49302 ( .A(n45426), .B(n41885), .Z(n50091) );
  XNOR U49303 ( .A(n50092), .B(n50024), .Z(n41885) );
  ANDN U49304 ( .B(n50025), .A(n48753), .Z(n50092) );
  XOR U49305 ( .A(n50093), .B(n50037), .Z(n45426) );
  ANDN U49306 ( .B(n50036), .A(n50094), .Z(n50093) );
  XOR U49307 ( .A(n44863), .B(n50095), .Z(n50090) );
  XOR U49308 ( .A(n40852), .B(n43348), .Z(n50095) );
  XNOR U49309 ( .A(n50096), .B(n50097), .Z(n43348) );
  ANDN U49310 ( .B(n50029), .A(n48757), .Z(n50096) );
  XNOR U49311 ( .A(n50098), .B(n50032), .Z(n40852) );
  AND U49312 ( .A(n48743), .B(n50033), .Z(n50098) );
  XNOR U49313 ( .A(n50099), .B(n50039), .Z(n44863) );
  ANDN U49314 ( .B(n50040), .A(n48747), .Z(n50099) );
  ANDN U49315 ( .B(n40989), .A(n40990), .Z(n50075) );
  XNOR U49316 ( .A(n50100), .B(n43327), .Z(n40990) );
  XOR U49317 ( .A(n49812), .B(n43916), .Z(n40989) );
  XNOR U49318 ( .A(n50103), .B(n50104), .Z(n48494) );
  XNOR U49319 ( .A(n45115), .B(n49008), .Z(n50104) );
  XNOR U49320 ( .A(n50105), .B(n49501), .Z(n49008) );
  XOR U49321 ( .A(round_reg[310]), .B(n50106), .Z(n49500) );
  XOR U49322 ( .A(round_reg[1479]), .B(n50107), .Z(n49462) );
  XOR U49323 ( .A(n50108), .B(n50109), .Z(n45115) );
  ANDN U49324 ( .B(n49449), .A(n49493), .Z(n50108) );
  XOR U49325 ( .A(round_reg[58]), .B(n50110), .Z(n49493) );
  XOR U49326 ( .A(round_reg[1544]), .B(n50111), .Z(n49449) );
  XNOR U49327 ( .A(n48928), .B(n50112), .Z(n50103) );
  XOR U49328 ( .A(n45314), .B(n44689), .Z(n50112) );
  XOR U49329 ( .A(n50113), .B(n49503), .Z(n44689) );
  XOR U49330 ( .A(n50114), .B(n50115), .Z(n45314) );
  NOR U49331 ( .A(n49458), .B(n49506), .Z(n50114) );
  XOR U49332 ( .A(round_reg[198]), .B(n50116), .Z(n49506) );
  XOR U49333 ( .A(round_reg[1418]), .B(n50117), .Z(n49458) );
  XNOR U49334 ( .A(n50118), .B(n49497), .Z(n48928) );
  ANDN U49335 ( .B(n49454), .A(n49496), .Z(n50118) );
  XOR U49336 ( .A(round_reg[80]), .B(n50119), .Z(n49496) );
  XOR U49337 ( .A(round_reg[1325]), .B(n50120), .Z(n49454) );
  XOR U49338 ( .A(n50121), .B(n50122), .Z(n46595) );
  XNOR U49339 ( .A(n45843), .B(n45961), .Z(n50122) );
  XNOR U49340 ( .A(n50123), .B(n48275), .Z(n45961) );
  XOR U49341 ( .A(round_reg[1417]), .B(n50124), .Z(n48275) );
  NOR U49342 ( .A(n48214), .B(n48213), .Z(n50123) );
  XOR U49343 ( .A(round_reg[1040]), .B(n50119), .Z(n48213) );
  XOR U49344 ( .A(n50125), .B(n50126), .Z(n45843) );
  NOR U49345 ( .A(n48210), .B(n48209), .Z(n50125) );
  XOR U49346 ( .A(round_reg[1089]), .B(n50127), .Z(n48209) );
  XOR U49347 ( .A(n45442), .B(n50128), .Z(n50121) );
  XNOR U49348 ( .A(n46418), .B(n46542), .Z(n50128) );
  XNOR U49349 ( .A(n48283), .B(n50129), .Z(n46542) );
  XNOR U49350 ( .A(n4687), .B(n50130), .Z(n50129) );
  NANDN U49351 ( .A(n48200), .B(n48201), .Z(n50130) );
  XOR U49352 ( .A(round_reg[1179]), .B(n50131), .Z(n48200) );
  XOR U49353 ( .A(round_reg[1543]), .B(n50132), .Z(n48283) );
  XOR U49354 ( .A(n50133), .B(n48662), .Z(n46418) );
  IV U49355 ( .A(n49021), .Z(n48662) );
  XOR U49356 ( .A(round_reg[1324]), .B(n49982), .Z(n49021) );
  ANDN U49357 ( .B(n48204), .A(n50134), .Z(n50133) );
  XNOR U49358 ( .A(round_reg[1251]), .B(n48701), .Z(n48204) );
  XNOR U49359 ( .A(n50135), .B(n48281), .Z(n45442) );
  XNOR U49360 ( .A(round_reg[1387]), .B(n49867), .Z(n48281) );
  NOR U49361 ( .A(n48217), .B(n48218), .Z(n50135) );
  IV U49362 ( .A(n49016), .Z(n48217) );
  XOR U49363 ( .A(round_reg[1011]), .B(n50136), .Z(n49016) );
  XNOR U49364 ( .A(n50137), .B(n49504), .Z(n49812) );
  XNOR U49365 ( .A(round_reg[139]), .B(n50138), .Z(n49504) );
  ANDN U49366 ( .B(n49447), .A(n49445), .Z(n50137) );
  XOR U49367 ( .A(round_reg[1388]), .B(n50139), .Z(n49445) );
  IV U49368 ( .A(n50140), .Z(n49447) );
  XOR U49369 ( .A(n50141), .B(n43265), .Z(n38864) );
  XNOR U49370 ( .A(n43819), .B(n50142), .Z(n43265) );
  ANDN U49371 ( .B(n41361), .A(n41362), .Z(n50141) );
  XOR U49372 ( .A(n44504), .B(n49840), .Z(n41362) );
  XOR U49373 ( .A(n50145), .B(n49940), .Z(n49840) );
  AND U49374 ( .A(n49306), .B(n49304), .Z(n50145) );
  XNOR U49375 ( .A(n44743), .B(n49122), .Z(n41361) );
  XNOR U49376 ( .A(n50146), .B(n50147), .Z(n49122) );
  NOR U49377 ( .A(n47776), .B(n49614), .Z(n50146) );
  XOR U49378 ( .A(round_reg[153]), .B(n50148), .Z(n47776) );
  XNOR U49379 ( .A(n50149), .B(n50150), .Z(n48320) );
  XNOR U49380 ( .A(n50151), .B(n45084), .Z(n50150) );
  XNOR U49381 ( .A(n50152), .B(n47764), .Z(n45084) );
  AND U49382 ( .A(n49118), .B(n49117), .Z(n50152) );
  XOR U49383 ( .A(round_reg[621]), .B(n50153), .Z(n49118) );
  XOR U49384 ( .A(n47602), .B(n50154), .Z(n50149) );
  XOR U49385 ( .A(n47592), .B(n48343), .Z(n50154) );
  XNOR U49386 ( .A(n50155), .B(n47760), .Z(n48343) );
  ANDN U49387 ( .B(n49128), .A(n49129), .Z(n50155) );
  XOR U49388 ( .A(round_reg[385]), .B(n50156), .Z(n49129) );
  XOR U49389 ( .A(n50157), .B(n47774), .Z(n47592) );
  AND U49390 ( .A(n49126), .B(n49125), .Z(n50157) );
  XOR U49391 ( .A(round_reg[455]), .B(n50158), .Z(n49126) );
  XNOR U49392 ( .A(n50159), .B(n47778), .Z(n47602) );
  AND U49393 ( .A(n49614), .B(n50147), .Z(n50159) );
  XOR U49394 ( .A(round_reg[553]), .B(n48368), .Z(n49614) );
  XNOR U49395 ( .A(n50160), .B(n50161), .Z(n47414) );
  XNOR U49396 ( .A(n46874), .B(n45259), .Z(n50161) );
  XOR U49397 ( .A(n50162), .B(n49805), .Z(n45259) );
  ANDN U49398 ( .B(n50163), .A(n50065), .Z(n50162) );
  XNOR U49399 ( .A(n50164), .B(n48314), .Z(n46874) );
  XNOR U49400 ( .A(n46453), .B(n50167), .Z(n50160) );
  XOR U49401 ( .A(n45647), .B(n48263), .Z(n50167) );
  XNOR U49402 ( .A(n50168), .B(n50069), .Z(n48263) );
  ANDN U49403 ( .B(n50169), .A(n50061), .Z(n50168) );
  IV U49404 ( .A(n50170), .Z(n50061) );
  XNOR U49405 ( .A(n50171), .B(n47747), .Z(n45647) );
  ANDN U49406 ( .B(n50172), .A(n50067), .Z(n50171) );
  XNOR U49407 ( .A(n50173), .B(n47754), .Z(n46453) );
  ANDN U49408 ( .B(n50174), .A(n50058), .Z(n50173) );
  XOR U49409 ( .A(n39034), .B(n50175), .Z(n50073) );
  XOR U49410 ( .A(n40637), .B(n44988), .Z(n50175) );
  XNOR U49411 ( .A(n50176), .B(n43259), .Z(n44988) );
  XNOR U49412 ( .A(n49277), .B(n45167), .Z(n43259) );
  XOR U49413 ( .A(n50177), .B(n50178), .Z(n49277) );
  ANDN U49414 ( .B(n48849), .A(n48851), .Z(n50177) );
  XOR U49415 ( .A(round_reg[16]), .B(n48561), .Z(n48851) );
  ANDN U49416 ( .B(n44994), .A(n48572), .Z(n50176) );
  XOR U49417 ( .A(n43342), .B(n48147), .Z(n48572) );
  XOR U49418 ( .A(n50179), .B(n50180), .Z(n48147) );
  ANDN U49419 ( .B(n50181), .A(n50182), .Z(n50179) );
  IV U49420 ( .A(n47640), .Z(n43342) );
  XOR U49421 ( .A(n49064), .B(n50183), .Z(n47640) );
  XNOR U49422 ( .A(n50184), .B(n50185), .Z(n49064) );
  XOR U49423 ( .A(n45668), .B(n45407), .Z(n50185) );
  XOR U49424 ( .A(n50186), .B(n50187), .Z(n45407) );
  XNOR U49425 ( .A(n50188), .B(n50189), .Z(n45668) );
  NOR U49426 ( .A(n48156), .B(n48155), .Z(n50188) );
  XOR U49427 ( .A(n46791), .B(n50190), .Z(n50184) );
  XOR U49428 ( .A(n42521), .B(n49542), .Z(n50190) );
  XNOR U49429 ( .A(n50191), .B(n50192), .Z(n49542) );
  ANDN U49430 ( .B(n48149), .A(n48150), .Z(n50191) );
  XNOR U49431 ( .A(n50193), .B(n50194), .Z(n42521) );
  XNOR U49432 ( .A(n50195), .B(n50196), .Z(n46791) );
  ANDN U49433 ( .B(n50180), .A(n50181), .Z(n50195) );
  XOR U49434 ( .A(n48254), .B(n44588), .Z(n44994) );
  XOR U49435 ( .A(n50197), .B(n46428), .Z(n44588) );
  XNOR U49436 ( .A(n50198), .B(n50199), .Z(n46428) );
  XNOR U49437 ( .A(n45435), .B(n42215), .Z(n50199) );
  XNOR U49438 ( .A(n50200), .B(n50201), .Z(n42215) );
  ANDN U49439 ( .B(n48250), .A(n48251), .Z(n50200) );
  XNOR U49440 ( .A(n50202), .B(n50203), .Z(n45435) );
  XOR U49441 ( .A(n43652), .B(n50206), .Z(n50198) );
  XOR U49442 ( .A(n43928), .B(n43591), .Z(n50206) );
  XNOR U49443 ( .A(n50207), .B(n50208), .Z(n43591) );
  NOR U49444 ( .A(n48260), .B(n48262), .Z(n50207) );
  XNOR U49445 ( .A(n50209), .B(n50210), .Z(n43928) );
  XNOR U49446 ( .A(n50211), .B(n50212), .Z(n43652) );
  NOR U49447 ( .A(n50213), .B(n48258), .Z(n50211) );
  XOR U49448 ( .A(n50214), .B(n50205), .Z(n48254) );
  ANDN U49449 ( .B(n50204), .A(n50215), .Z(n50214) );
  XNOR U49450 ( .A(n50216), .B(n43255), .Z(n40637) );
  XNOR U49451 ( .A(n43865), .B(n50217), .Z(n43255) );
  XNOR U49452 ( .A(n46211), .B(n49996), .Z(n43865) );
  XNOR U49453 ( .A(n50218), .B(n50219), .Z(n49996) );
  XNOR U49454 ( .A(n45912), .B(n45129), .Z(n50219) );
  XNOR U49455 ( .A(n50220), .B(n48748), .Z(n45129) );
  ANDN U49456 ( .B(n48749), .A(n50039), .Z(n50220) );
  XNOR U49457 ( .A(round_reg[957]), .B(n49087), .Z(n50039) );
  XOR U49458 ( .A(round_reg[1004]), .B(n50221), .Z(n48749) );
  XNOR U49459 ( .A(n50222), .B(n50223), .Z(n45912) );
  ANDN U49460 ( .B(n50035), .A(n50037), .Z(n50222) );
  XOR U49461 ( .A(round_reg[743]), .B(n50224), .Z(n50037) );
  XOR U49462 ( .A(n45713), .B(n50225), .Z(n50218) );
  XOR U49463 ( .A(n44705), .B(n46977), .Z(n50225) );
  XNOR U49464 ( .A(n50226), .B(n48758), .Z(n46977) );
  ANDN U49465 ( .B(n50028), .A(n50027), .Z(n50226) );
  XNOR U49466 ( .A(round_reg[1033]), .B(n50227), .Z(n50027) );
  IV U49467 ( .A(n50097), .Z(n50028) );
  XOR U49468 ( .A(round_reg[665]), .B(n50228), .Z(n50097) );
  XNOR U49469 ( .A(n48755), .B(n50229), .Z(n44705) );
  XNOR U49470 ( .A(n11417), .B(n50230), .Z(n50229) );
  NANDN U49471 ( .A(n50024), .B(n48754), .Z(n50230) );
  XOR U49472 ( .A(round_reg[1172]), .B(n50231), .Z(n48754) );
  XOR U49473 ( .A(round_reg[789]), .B(n50232), .Z(n50024) );
  IV U49474 ( .A(rc_i[0]), .Z(n11417) );
  XNOR U49475 ( .A(n50233), .B(n48744), .Z(n45713) );
  ANDN U49476 ( .B(n48745), .A(n50032), .Z(n50233) );
  XOR U49477 ( .A(round_reg[886]), .B(n50234), .Z(n50032) );
  XOR U49478 ( .A(round_reg[1244]), .B(n49798), .Z(n48745) );
  XNOR U49479 ( .A(n50235), .B(n50236), .Z(n46211) );
  XOR U49480 ( .A(n48716), .B(n46741), .Z(n50236) );
  XOR U49481 ( .A(n50237), .B(n48738), .Z(n46741) );
  ANDN U49482 ( .B(n48739), .A(n49484), .Z(n50237) );
  XNOR U49483 ( .A(n50238), .B(n48734), .Z(n48716) );
  ANDN U49484 ( .B(n50041), .A(n50239), .Z(n50238) );
  XOR U49485 ( .A(n46289), .B(n50240), .Z(n50235) );
  XOR U49486 ( .A(n46031), .B(n46713), .Z(n50240) );
  XNOR U49487 ( .A(n50241), .B(n48725), .Z(n46713) );
  ANDN U49488 ( .B(n48726), .A(n49477), .Z(n50241) );
  XNOR U49489 ( .A(n50242), .B(n48730), .Z(n46031) );
  XNOR U49490 ( .A(n50243), .B(n48721), .Z(n46289) );
  ANDN U49491 ( .B(n49487), .A(n50244), .Z(n50243) );
  ANDN U49492 ( .B(n40985), .A(n40987), .Z(n50216) );
  XOR U49493 ( .A(n49094), .B(n46940), .Z(n40987) );
  XOR U49494 ( .A(n50246), .B(n50247), .Z(n47526) );
  XOR U49495 ( .A(n44751), .B(n47063), .Z(n50247) );
  XOR U49496 ( .A(n50248), .B(n50249), .Z(n47063) );
  XNOR U49497 ( .A(n50252), .B(n50253), .Z(n44751) );
  XOR U49498 ( .A(n46010), .B(n50256), .Z(n50246) );
  XOR U49499 ( .A(n50257), .B(n44522), .Z(n50256) );
  XNOR U49500 ( .A(n50258), .B(n50259), .Z(n44522) );
  NOR U49501 ( .A(n50260), .B(n50261), .Z(n50258) );
  XNOR U49502 ( .A(n50262), .B(n50263), .Z(n46010) );
  ANDN U49503 ( .B(n50264), .A(n50265), .Z(n50262) );
  XOR U49504 ( .A(n50266), .B(n50267), .Z(n49094) );
  ANDN U49505 ( .B(n50268), .A(n50269), .Z(n50266) );
  XOR U49506 ( .A(n50270), .B(n49525), .Z(n40985) );
  XOR U49507 ( .A(n46695), .B(n47253), .Z(n49525) );
  XNOR U49508 ( .A(n50271), .B(n50272), .Z(n47253) );
  XOR U49509 ( .A(n46930), .B(n45229), .Z(n50272) );
  XNOR U49510 ( .A(n50273), .B(n47719), .Z(n45229) );
  ANDN U49511 ( .B(n50274), .A(n50275), .Z(n50273) );
  XNOR U49512 ( .A(n50276), .B(n50277), .Z(n46930) );
  NOR U49513 ( .A(n50278), .B(n50279), .Z(n50276) );
  XNOR U49514 ( .A(n43775), .B(n50280), .Z(n50271) );
  XNOR U49515 ( .A(n45304), .B(n47971), .Z(n50280) );
  XOR U49516 ( .A(n50281), .B(n47709), .Z(n47971) );
  ANDN U49517 ( .B(n50282), .A(n50283), .Z(n50281) );
  XNOR U49518 ( .A(n50284), .B(n47715), .Z(n45304) );
  ANDN U49519 ( .B(n50285), .A(n50286), .Z(n50284) );
  XNOR U49520 ( .A(n50287), .B(n50288), .Z(n43775) );
  NOR U49521 ( .A(n50289), .B(n50290), .Z(n50287) );
  XNOR U49522 ( .A(n50291), .B(n50292), .Z(n46695) );
  XOR U49523 ( .A(n45340), .B(n46752), .Z(n50292) );
  XOR U49524 ( .A(n50293), .B(n47989), .Z(n46752) );
  ANDN U49525 ( .B(n47988), .A(n49710), .Z(n50293) );
  XOR U49526 ( .A(round_reg[656]), .B(n48561), .Z(n47988) );
  XOR U49527 ( .A(n50294), .B(n47981), .Z(n45340) );
  ANDN U49528 ( .B(n47982), .A(n49713), .Z(n50294) );
  XOR U49529 ( .A(round_reg[734]), .B(n49606), .Z(n47982) );
  XNOR U49530 ( .A(n42882), .B(n50295), .Z(n50291) );
  XOR U49531 ( .A(n45822), .B(n44407), .Z(n50295) );
  XNOR U49532 ( .A(n50296), .B(n50297), .Z(n44407) );
  ANDN U49533 ( .B(n47978), .A(n50298), .Z(n50296) );
  XOR U49534 ( .A(round_reg[948]), .B(n50299), .Z(n47978) );
  XOR U49535 ( .A(n50300), .B(n50301), .Z(n45822) );
  ANDN U49536 ( .B(n49719), .A(n49721), .Z(n50300) );
  XNOR U49537 ( .A(n50302), .B(n50303), .Z(n42882) );
  ANDN U49538 ( .B(n49723), .A(n49725), .Z(n50302) );
  IV U49539 ( .A(n50304), .Z(n49723) );
  XOR U49540 ( .A(n50305), .B(n43262), .Z(n39034) );
  XNOR U49541 ( .A(n48889), .B(n42453), .Z(n43262) );
  XNOR U49542 ( .A(n50306), .B(n48987), .Z(n42453) );
  XNOR U49543 ( .A(n50307), .B(n50308), .Z(n48987) );
  XOR U49544 ( .A(n46545), .B(n45801), .Z(n50308) );
  XNOR U49545 ( .A(n50309), .B(n49700), .Z(n45801) );
  AND U49546 ( .A(n50310), .B(n50311), .Z(n50309) );
  XNOR U49547 ( .A(n50312), .B(n47231), .Z(n46545) );
  NOR U49548 ( .A(n50313), .B(n50314), .Z(n50312) );
  XNOR U49549 ( .A(n50142), .B(n50315), .Z(n50307) );
  XOR U49550 ( .A(n46522), .B(n43820), .Z(n50315) );
  XOR U49551 ( .A(n50316), .B(n47222), .Z(n43820) );
  AND U49552 ( .A(n50317), .B(n50318), .Z(n50316) );
  XOR U49553 ( .A(n50319), .B(n47228), .Z(n46522) );
  XOR U49554 ( .A(n50322), .B(n50323), .Z(n50142) );
  ANDN U49555 ( .B(n50324), .A(n50325), .Z(n50322) );
  XOR U49556 ( .A(n50326), .B(n50327), .Z(n48889) );
  NOR U49557 ( .A(n50328), .B(n50329), .Z(n50326) );
  NOR U49558 ( .A(n40980), .B(n40979), .Z(n50305) );
  XOR U49559 ( .A(n50330), .B(n46443), .Z(n40979) );
  XOR U49560 ( .A(n50331), .B(n48429), .Z(n46443) );
  XOR U49561 ( .A(n50332), .B(n50333), .Z(n48429) );
  XNOR U49562 ( .A(n46299), .B(n46167), .Z(n50333) );
  XOR U49563 ( .A(n50334), .B(n49652), .Z(n46167) );
  ANDN U49564 ( .B(n50335), .A(n50336), .Z(n50334) );
  XNOR U49565 ( .A(n50337), .B(n49655), .Z(n46299) );
  AND U49566 ( .A(n49410), .B(n49656), .Z(n50337) );
  XNOR U49567 ( .A(n46590), .B(n50338), .Z(n50332) );
  XOR U49568 ( .A(n46254), .B(n49636), .Z(n50338) );
  XNOR U49569 ( .A(n50339), .B(n49645), .Z(n49636) );
  NOR U49570 ( .A(n50340), .B(n49644), .Z(n50339) );
  XNOR U49571 ( .A(n50341), .B(n49648), .Z(n46254) );
  AND U49572 ( .A(n49406), .B(n49649), .Z(n50341) );
  XNOR U49573 ( .A(n50342), .B(n49642), .Z(n46590) );
  ANDN U49574 ( .B(n50343), .A(n49641), .Z(n50342) );
  XOR U49575 ( .A(n45315), .B(n50344), .Z(n40980) );
  XOR U49576 ( .A(n50345), .B(n50346), .Z(n41995) );
  XNOR U49577 ( .A(n40375), .B(n37330), .Z(n50346) );
  XNOR U49578 ( .A(n50347), .B(n43250), .Z(n37330) );
  XOR U49579 ( .A(n49546), .B(n46194), .Z(n43250) );
  XNOR U49580 ( .A(n50348), .B(n50349), .Z(n46194) );
  XNOR U49581 ( .A(n50350), .B(n50351), .Z(n49546) );
  ANDN U49582 ( .B(n50352), .A(n47736), .Z(n50350) );
  ANDN U49583 ( .B(n42352), .A(n45003), .Z(n50347) );
  XOR U49584 ( .A(n50353), .B(n44119), .Z(n45003) );
  XNOR U49585 ( .A(n50354), .B(n47097), .Z(n44119) );
  XNOR U49586 ( .A(n50355), .B(n50356), .Z(n47097) );
  XNOR U49587 ( .A(n46255), .B(n44582), .Z(n50356) );
  XOR U49588 ( .A(n50357), .B(n49745), .Z(n44582) );
  AND U49589 ( .A(n50358), .B(n49746), .Z(n50357) );
  XNOR U49590 ( .A(n50359), .B(n49736), .Z(n46255) );
  AND U49591 ( .A(n50360), .B(n49737), .Z(n50359) );
  XOR U49592 ( .A(n44844), .B(n50361), .Z(n50355) );
  XOR U49593 ( .A(n45297), .B(n46871), .Z(n50361) );
  XNOR U49594 ( .A(n50362), .B(n49732), .Z(n46871) );
  ANDN U49595 ( .B(n49733), .A(n50363), .Z(n50362) );
  XNOR U49596 ( .A(n50364), .B(n49741), .Z(n45297) );
  AND U49597 ( .A(n50365), .B(n49742), .Z(n50364) );
  XNOR U49598 ( .A(n50366), .B(n49749), .Z(n44844) );
  ANDN U49599 ( .B(n49750), .A(n50367), .Z(n50366) );
  XOR U49600 ( .A(n44937), .B(n48763), .Z(n42352) );
  XOR U49601 ( .A(n50368), .B(n50369), .Z(n48763) );
  ANDN U49602 ( .B(n48578), .A(n48579), .Z(n50368) );
  IV U49603 ( .A(n43784), .Z(n44937) );
  XOR U49604 ( .A(n46683), .B(n47237), .Z(n43784) );
  XNOR U49605 ( .A(n50370), .B(n50371), .Z(n47237) );
  XNOR U49606 ( .A(n45921), .B(n46121), .Z(n50371) );
  XOR U49607 ( .A(n50372), .B(n50373), .Z(n46121) );
  ANDN U49608 ( .B(n50374), .A(n50375), .Z(n50372) );
  XNOR U49609 ( .A(n50376), .B(n50377), .Z(n45921) );
  ANDN U49610 ( .B(n50378), .A(n50379), .Z(n50376) );
  XNOR U49611 ( .A(n46026), .B(n50380), .Z(n50370) );
  XOR U49612 ( .A(n50381), .B(n47398), .Z(n50380) );
  XOR U49613 ( .A(n50382), .B(n50383), .Z(n47398) );
  ANDN U49614 ( .B(n50384), .A(n50385), .Z(n50382) );
  XOR U49615 ( .A(n50386), .B(n50387), .Z(n46026) );
  ANDN U49616 ( .B(n50388), .A(n50389), .Z(n50386) );
  XOR U49617 ( .A(n50390), .B(n50391), .Z(n46683) );
  XNOR U49618 ( .A(n43326), .B(n45954), .Z(n50391) );
  XNOR U49619 ( .A(n50392), .B(n50393), .Z(n45954) );
  ANDN U49620 ( .B(n48768), .A(n48595), .Z(n50392) );
  XOR U49621 ( .A(round_reg[814]), .B(n50394), .Z(n48595) );
  XNOR U49622 ( .A(n50395), .B(n50396), .Z(n43326) );
  ANDN U49623 ( .B(n48765), .A(n48587), .Z(n50395) );
  XOR U49624 ( .A(round_reg[918]), .B(n50397), .Z(n48587) );
  XNOR U49625 ( .A(n50100), .B(n50398), .Z(n50390) );
  XNOR U49626 ( .A(n45289), .B(n49702), .Z(n50398) );
  XOR U49627 ( .A(n50399), .B(n50400), .Z(n49702) );
  ANDN U49628 ( .B(n48772), .A(n48591), .Z(n50399) );
  XOR U49629 ( .A(round_reg[847]), .B(n50401), .Z(n48591) );
  XNOR U49630 ( .A(n50402), .B(n50403), .Z(n45289) );
  NOR U49631 ( .A(n48578), .B(n50369), .Z(n50402) );
  XNOR U49632 ( .A(round_reg[690]), .B(n50404), .Z(n48578) );
  XOR U49633 ( .A(n50405), .B(n50406), .Z(n50100) );
  ANDN U49634 ( .B(n48770), .A(n48582), .Z(n50405) );
  XOR U49635 ( .A(round_reg[704]), .B(n50407), .Z(n48582) );
  XOR U49636 ( .A(n50408), .B(n43239), .Z(n40375) );
  XOR U49637 ( .A(n49916), .B(n47407), .Z(n43239) );
  XNOR U49638 ( .A(n46411), .B(n50020), .Z(n47407) );
  XNOR U49639 ( .A(n50409), .B(n50410), .Z(n50020) );
  XOR U49640 ( .A(n43890), .B(n46225), .Z(n50410) );
  XNOR U49641 ( .A(n50411), .B(n48731), .Z(n46225) );
  XOR U49642 ( .A(round_reg[73]), .B(n50227), .Z(n48731) );
  NOR U49643 ( .A(n49481), .B(n49482), .Z(n50411) );
  XOR U49644 ( .A(round_reg[1318]), .B(n50412), .Z(n49481) );
  XNOR U49645 ( .A(n50413), .B(n50244), .Z(n43890) );
  IV U49646 ( .A(n48722), .Z(n50244) );
  XOR U49647 ( .A(round_reg[303]), .B(n50414), .Z(n48722) );
  NOR U49648 ( .A(n49487), .B(n49488), .Z(n50413) );
  XNOR U49649 ( .A(round_reg[1472]), .B(n50415), .Z(n49487) );
  XOR U49650 ( .A(n43866), .B(n50416), .Z(n50409) );
  XNOR U49651 ( .A(n45690), .B(n50217), .Z(n50416) );
  XNOR U49652 ( .A(n50417), .B(n50239), .Z(n50217) );
  IV U49653 ( .A(n48735), .Z(n50239) );
  XOR U49654 ( .A(round_reg[51]), .B(n50136), .Z(n48735) );
  NOR U49655 ( .A(n50044), .B(n50041), .Z(n50417) );
  XNOR U49656 ( .A(round_reg[1537]), .B(n49857), .Z(n50041) );
  XNOR U49657 ( .A(n50418), .B(n48726), .Z(n45690) );
  XNOR U49658 ( .A(round_reg[132]), .B(n50419), .Z(n48726) );
  ANDN U49659 ( .B(n49477), .A(n49478), .Z(n50418) );
  XOR U49660 ( .A(round_reg[1381]), .B(n49901), .Z(n49477) );
  XNOR U49661 ( .A(n50420), .B(n48739), .Z(n43866) );
  XOR U49662 ( .A(round_reg[255]), .B(n48520), .Z(n48739) );
  ANDN U49663 ( .B(n49484), .A(n49485), .Z(n50420) );
  XOR U49664 ( .A(round_reg[1411]), .B(n50421), .Z(n49484) );
  XOR U49665 ( .A(n50422), .B(n50423), .Z(n46411) );
  XNOR U49666 ( .A(n42332), .B(n45661), .Z(n50423) );
  XNOR U49667 ( .A(n50424), .B(n47666), .Z(n45661) );
  XOR U49668 ( .A(round_reg[745]), .B(n49905), .Z(n47666) );
  ANDN U49669 ( .B(n47665), .A(n50425), .Z(n50424) );
  XNOR U49670 ( .A(n50426), .B(n47657), .Z(n42332) );
  XNOR U49671 ( .A(round_reg[888]), .B(n50427), .Z(n47657) );
  ANDN U49672 ( .B(n47658), .A(n49918), .Z(n50426) );
  XOR U49673 ( .A(round_reg[499]), .B(n48942), .Z(n47658) );
  XNOR U49674 ( .A(n44162), .B(n50428), .Z(n50422) );
  XNOR U49675 ( .A(n44707), .B(n46209), .Z(n50428) );
  XNOR U49676 ( .A(n50429), .B(n47649), .Z(n46209) );
  NOR U49677 ( .A(n49926), .B(n47648), .Z(n50429) );
  XOR U49678 ( .A(round_reg[533]), .B(n50430), .Z(n47648) );
  XNOR U49679 ( .A(n50431), .B(n47653), .Z(n44707) );
  XOR U49680 ( .A(round_reg[791]), .B(n49833), .Z(n47653) );
  NOR U49681 ( .A(n49921), .B(n47652), .Z(n50431) );
  XNOR U49682 ( .A(round_reg[429]), .B(n50432), .Z(n47652) );
  XNOR U49683 ( .A(n50433), .B(n47662), .Z(n44162) );
  IV U49684 ( .A(n48117), .Z(n47662) );
  XOR U49685 ( .A(round_reg[667]), .B(n49955), .Z(n48117) );
  NOR U49686 ( .A(n49923), .B(n47661), .Z(n50433) );
  XNOR U49687 ( .A(round_reg[601]), .B(n50434), .Z(n47661) );
  XNOR U49688 ( .A(n50435), .B(n47665), .Z(n49916) );
  XNOR U49689 ( .A(round_reg[378]), .B(n50110), .Z(n47665) );
  ANDN U49690 ( .B(n50425), .A(n48119), .Z(n50435) );
  NOR U49691 ( .A(n45007), .B(n43006), .Z(n50408) );
  XOR U49692 ( .A(n49517), .B(n44797), .Z(n43006) );
  IV U49693 ( .A(n44036), .Z(n44797) );
  XNOR U49694 ( .A(n50436), .B(n48270), .Z(n44036) );
  XNOR U49695 ( .A(n50437), .B(n50438), .Z(n48270) );
  XOR U49696 ( .A(n49393), .B(n46570), .Z(n50438) );
  XNOR U49697 ( .A(n50439), .B(n50140), .Z(n46570) );
  XOR U49698 ( .A(round_reg[1012]), .B(n50440), .Z(n50140) );
  NOR U49699 ( .A(n49503), .B(n49446), .Z(n50439) );
  XNOR U49700 ( .A(round_reg[901]), .B(n50441), .Z(n49446) );
  XOR U49701 ( .A(round_reg[539]), .B(n50442), .Z(n49503) );
  XNOR U49702 ( .A(n50443), .B(n49451), .Z(n49393) );
  XNOR U49703 ( .A(round_reg[1180]), .B(n48876), .Z(n49451) );
  NOR U49704 ( .A(n50109), .B(n49450), .Z(n50443) );
  XOR U49705 ( .A(round_reg[797]), .B(n48517), .Z(n49450) );
  IV U49706 ( .A(n49494), .Z(n50109) );
  XOR U49707 ( .A(round_reg[435]), .B(n50444), .Z(n49494) );
  XNOR U49708 ( .A(n47022), .B(n50445), .Z(n50437) );
  XOR U49709 ( .A(n49440), .B(n43661), .Z(n50445) );
  XNOR U49710 ( .A(n50446), .B(n49456), .Z(n43661) );
  XNOR U49711 ( .A(round_reg[1252]), .B(n50447), .Z(n49456) );
  ANDN U49712 ( .B(n49497), .A(n49455), .Z(n50446) );
  XNOR U49713 ( .A(round_reg[894]), .B(n50448), .Z(n49455) );
  XOR U49714 ( .A(round_reg[505]), .B(n50449), .Z(n49497) );
  XNOR U49715 ( .A(n50450), .B(n49460), .Z(n49440) );
  XNOR U49716 ( .A(round_reg[1041]), .B(n49827), .Z(n49460) );
  IV U49717 ( .A(n50451), .Z(n49827) );
  NOR U49718 ( .A(n50115), .B(n49459), .Z(n50450) );
  XOR U49719 ( .A(round_reg[673]), .B(n50452), .Z(n49459) );
  IV U49720 ( .A(n49507), .Z(n50115) );
  XOR U49721 ( .A(round_reg[607]), .B(n50453), .Z(n49507) );
  XNOR U49722 ( .A(n50454), .B(n49464), .Z(n47022) );
  XNOR U49723 ( .A(round_reg[1090]), .B(n50455), .Z(n49464) );
  ANDN U49724 ( .B(n49501), .A(n49463), .Z(n50454) );
  XOR U49725 ( .A(round_reg[751]), .B(n50456), .Z(n49463) );
  XOR U49726 ( .A(round_reg[320]), .B(n50457), .Z(n49501) );
  XNOR U49727 ( .A(n50458), .B(n49820), .Z(n49517) );
  AND U49728 ( .A(n49590), .B(n49588), .Z(n50458) );
  XNOR U49729 ( .A(n48027), .B(n45635), .Z(n45007) );
  IV U49730 ( .A(n42659), .Z(n45635) );
  XNOR U49731 ( .A(n46292), .B(n50245), .Z(n42659) );
  XNOR U49732 ( .A(n50459), .B(n50460), .Z(n50245) );
  XNOR U49733 ( .A(n44498), .B(n45815), .Z(n50460) );
  XNOR U49734 ( .A(n50461), .B(n50462), .Z(n45815) );
  ANDN U49735 ( .B(n49096), .A(n49097), .Z(n50461) );
  XNOR U49736 ( .A(n50463), .B(n50464), .Z(n44498) );
  ANDN U49737 ( .B(n49105), .A(n49106), .Z(n50463) );
  XOR U49738 ( .A(n45354), .B(n50465), .Z(n50459) );
  XOR U49739 ( .A(n50466), .B(n44982), .Z(n50465) );
  XNOR U49740 ( .A(n50467), .B(n50468), .Z(n44982) );
  ANDN U49741 ( .B(n50267), .A(n50268), .Z(n50467) );
  XOR U49742 ( .A(n50469), .B(n50470), .Z(n45354) );
  XNOR U49743 ( .A(n50471), .B(n50472), .Z(n46292) );
  XOR U49744 ( .A(n45452), .B(n45740), .Z(n50472) );
  XOR U49745 ( .A(n50473), .B(n46148), .Z(n45740) );
  ANDN U49746 ( .B(n48809), .A(n46147), .Z(n50473) );
  XNOR U49747 ( .A(n50474), .B(n46137), .Z(n45452) );
  AND U49748 ( .A(n48030), .B(n46138), .Z(n50474) );
  XOR U49749 ( .A(round_reg[257]), .B(n49857), .Z(n46138) );
  XOR U49750 ( .A(round_reg[1490]), .B(n50475), .Z(n48030) );
  XOR U49751 ( .A(n45849), .B(n50476), .Z(n50471) );
  XOR U49752 ( .A(n45510), .B(n45892), .Z(n50476) );
  XNOR U49753 ( .A(n50477), .B(n47154), .Z(n45892) );
  XOR U49754 ( .A(round_reg[209]), .B(n49898), .Z(n47155) );
  XNOR U49755 ( .A(round_reg[1429]), .B(n50232), .Z(n48025) );
  XNOR U49756 ( .A(n50478), .B(n46143), .Z(n45510) );
  ANDN U49757 ( .B(n48022), .A(n46144), .Z(n50478) );
  XOR U49758 ( .A(round_reg[5]), .B(n50479), .Z(n46144) );
  XNOR U49759 ( .A(round_reg[1555]), .B(n50480), .Z(n48022) );
  XNOR U49760 ( .A(n50481), .B(n46239), .Z(n45849) );
  XOR U49761 ( .A(round_reg[150]), .B(n50482), .Z(n46240) );
  XOR U49762 ( .A(round_reg[1399]), .B(n50483), .Z(n48033) );
  XNOR U49763 ( .A(n50484), .B(n46147), .Z(n48027) );
  XOR U49764 ( .A(round_reg[91]), .B(n50485), .Z(n46147) );
  NOR U49765 ( .A(n48810), .B(n48809), .Z(n50484) );
  XOR U49766 ( .A(round_reg[1336]), .B(n50486), .Z(n48809) );
  XOR U49767 ( .A(n41715), .B(n50487), .Z(n50345) );
  XOR U49768 ( .A(n39133), .B(n38509), .Z(n50487) );
  XNOR U49769 ( .A(n50488), .B(n43248), .Z(n38509) );
  XNOR U49770 ( .A(n43091), .B(n49398), .Z(n43248) );
  XOR U49771 ( .A(n50489), .B(n50343), .Z(n49398) );
  ANDN U49772 ( .B(n49640), .A(n50490), .Z(n50489) );
  ANDN U49773 ( .B(n42348), .A(n45012), .Z(n50488) );
  XOR U49774 ( .A(n42540), .B(n47266), .Z(n45012) );
  ANDN U49775 ( .B(n50492), .A(n47310), .Z(n50491) );
  XNOR U49776 ( .A(n46594), .B(n48348), .Z(n42540) );
  XNOR U49777 ( .A(n50493), .B(n50494), .Z(n48348) );
  XOR U49778 ( .A(n46244), .B(n45388), .Z(n50494) );
  XOR U49779 ( .A(n50495), .B(n49223), .Z(n45388) );
  XNOR U49780 ( .A(round_reg[195]), .B(n49958), .Z(n49223) );
  ANDN U49781 ( .B(n48345), .A(n48346), .Z(n50495) );
  XNOR U49782 ( .A(round_reg[1038]), .B(n48957), .Z(n48346) );
  XNOR U49783 ( .A(round_reg[1415]), .B(n50158), .Z(n48345) );
  XNOR U49784 ( .A(n50496), .B(n48083), .Z(n46244) );
  XOR U49785 ( .A(round_reg[136]), .B(n50497), .Z(n48083) );
  XOR U49786 ( .A(round_reg[1009]), .B(n50498), .Z(n47365) );
  XOR U49787 ( .A(round_reg[1385]), .B(n49905), .Z(n47364) );
  XOR U49788 ( .A(n49199), .B(n50499), .Z(n50493) );
  XOR U49789 ( .A(n44914), .B(n46889), .Z(n50499) );
  XNOR U49790 ( .A(n50500), .B(n47298), .Z(n46889) );
  XNOR U49791 ( .A(round_reg[77]), .B(n48869), .Z(n47298) );
  NOR U49792 ( .A(n47377), .B(n47378), .Z(n50500) );
  XNOR U49793 ( .A(round_reg[1249]), .B(n50501), .Z(n47378) );
  XOR U49794 ( .A(round_reg[1322]), .B(n50502), .Z(n47377) );
  XNOR U49795 ( .A(n50503), .B(n47291), .Z(n44914) );
  XNOR U49796 ( .A(round_reg[307]), .B(n50504), .Z(n47291) );
  NOR U49797 ( .A(n47374), .B(n47375), .Z(n50503) );
  XOR U49798 ( .A(round_reg[1151]), .B(n49081), .Z(n47375) );
  XOR U49799 ( .A(round_reg[1476]), .B(n50505), .Z(n47374) );
  XNOR U49800 ( .A(n50506), .B(n47588), .Z(n49199) );
  XOR U49801 ( .A(round_reg[55]), .B(n50507), .Z(n47588) );
  ANDN U49802 ( .B(n47368), .A(n47369), .Z(n50506) );
  XNOR U49803 ( .A(round_reg[1177]), .B(n50508), .Z(n47369) );
  XNOR U49804 ( .A(round_reg[1541]), .B(n50509), .Z(n47368) );
  XOR U49805 ( .A(n50510), .B(n50511), .Z(n46594) );
  XNOR U49806 ( .A(n47172), .B(n44815), .Z(n50511) );
  XNOR U49807 ( .A(n50512), .B(n47305), .Z(n44815) );
  XOR U49808 ( .A(round_reg[795]), .B(n50513), .Z(n47305) );
  ANDN U49809 ( .B(n47278), .A(n48002), .Z(n50512) );
  IV U49810 ( .A(n47277), .Z(n48002) );
  XOR U49811 ( .A(round_reg[433]), .B(n50514), .Z(n47277) );
  XNOR U49812 ( .A(n50515), .B(n48009), .Z(n47172) );
  XNOR U49813 ( .A(round_reg[749]), .B(n50432), .Z(n48009) );
  NOR U49814 ( .A(n47269), .B(n47268), .Z(n50515) );
  XOR U49815 ( .A(round_reg[382]), .B(n50516), .Z(n47268) );
  XOR U49816 ( .A(n47996), .B(n50517), .Z(n50510) );
  XOR U49817 ( .A(n46111), .B(n47594), .Z(n50517) );
  XOR U49818 ( .A(n50518), .B(n47315), .Z(n47594) );
  XOR U49819 ( .A(round_reg[671]), .B(n50519), .Z(n47315) );
  ANDN U49820 ( .B(n47273), .A(n47274), .Z(n50518) );
  XOR U49821 ( .A(round_reg[605]), .B(n50520), .Z(n47273) );
  XOR U49822 ( .A(n50521), .B(n47312), .Z(n46111) );
  XOR U49823 ( .A(round_reg[892]), .B(n50522), .Z(n47312) );
  ANDN U49824 ( .B(n48005), .A(n50492), .Z(n50521) );
  XOR U49825 ( .A(round_reg[503]), .B(n50523), .Z(n48005) );
  XNOR U49826 ( .A(n50524), .B(n47303), .Z(n47996) );
  XOR U49827 ( .A(round_reg[899]), .B(n48514), .Z(n47303) );
  NOR U49828 ( .A(n47281), .B(n47283), .Z(n50524) );
  XOR U49829 ( .A(round_reg[537]), .B(n50508), .Z(n47281) );
  XOR U49830 ( .A(n50525), .B(n45759), .Z(n42348) );
  XOR U49831 ( .A(n47838), .B(n48243), .Z(n45759) );
  XOR U49832 ( .A(n50526), .B(n50527), .Z(n48243) );
  XNOR U49833 ( .A(n44925), .B(n43573), .Z(n50527) );
  XNOR U49834 ( .A(n50528), .B(n48692), .Z(n43573) );
  AND U49835 ( .A(n48654), .B(n48693), .Z(n50528) );
  XNOR U49836 ( .A(n50529), .B(n49540), .Z(n44925) );
  ANDN U49837 ( .B(n49539), .A(n50530), .Z(n50529) );
  XNOR U49838 ( .A(n45988), .B(n50531), .Z(n50526) );
  XOR U49839 ( .A(n47515), .B(n44229), .Z(n50531) );
  XNOR U49840 ( .A(n50532), .B(n48487), .Z(n44229) );
  NOR U49841 ( .A(n48486), .B(n48651), .Z(n50532) );
  XNOR U49842 ( .A(n50533), .B(n48483), .Z(n47515) );
  NOR U49843 ( .A(n48482), .B(n48647), .Z(n50533) );
  XOR U49844 ( .A(n50534), .B(n50535), .Z(n45988) );
  ANDN U49845 ( .B(n48477), .A(n48658), .Z(n50534) );
  XOR U49846 ( .A(n50536), .B(n50537), .Z(n47838) );
  XOR U49847 ( .A(n47886), .B(n46361), .Z(n50537) );
  XOR U49848 ( .A(n50538), .B(n50539), .Z(n46361) );
  ANDN U49849 ( .B(n49031), .A(n50540), .Z(n50538) );
  XNOR U49850 ( .A(n50541), .B(n47892), .Z(n47886) );
  NOR U49851 ( .A(n50542), .B(n49466), .Z(n50541) );
  XNOR U49852 ( .A(n47099), .B(n50543), .Z(n50536) );
  XOR U49853 ( .A(n47395), .B(n43679), .Z(n50543) );
  XNOR U49854 ( .A(n50544), .B(n47907), .Z(n43679) );
  ANDN U49855 ( .B(n50545), .A(n50546), .Z(n50544) );
  XNOR U49856 ( .A(n50547), .B(n47897), .Z(n47395) );
  ANDN U49857 ( .B(n49037), .A(n50548), .Z(n50547) );
  XNOR U49858 ( .A(n50549), .B(n47903), .Z(n47099) );
  ANDN U49859 ( .B(n49040), .A(n50550), .Z(n50549) );
  XNOR U49860 ( .A(n50551), .B(n43246), .Z(n39133) );
  XOR U49861 ( .A(n50552), .B(n43319), .Z(n43246) );
  XNOR U49862 ( .A(n50553), .B(n50554), .Z(n46532) );
  XNOR U49863 ( .A(n44556), .B(n41599), .Z(n50554) );
  XNOR U49864 ( .A(n50555), .B(n50556), .Z(n41599) );
  ANDN U49865 ( .B(n50557), .A(n47789), .Z(n50555) );
  XNOR U49866 ( .A(n50558), .B(n50559), .Z(n44556) );
  ANDN U49867 ( .B(n50560), .A(n47799), .Z(n50558) );
  XOR U49868 ( .A(n50561), .B(n50562), .Z(n50553) );
  XOR U49869 ( .A(n46915), .B(n44123), .Z(n50562) );
  XNOR U49870 ( .A(n50563), .B(n50564), .Z(n44123) );
  ANDN U49871 ( .B(n50565), .A(n47793), .Z(n50563) );
  XNOR U49872 ( .A(n50566), .B(n50567), .Z(n46915) );
  ANDN U49873 ( .B(n50568), .A(n47803), .Z(n50566) );
  ANDN U49874 ( .B(n45016), .A(n42359), .Z(n50551) );
  XOR U49875 ( .A(n47196), .B(n44673), .Z(n42359) );
  XNOR U49876 ( .A(n50571), .B(n50572), .Z(n48039) );
  XOR U49877 ( .A(n41730), .B(n46423), .Z(n50572) );
  XOR U49878 ( .A(n50573), .B(n50574), .Z(n46423) );
  ANDN U49879 ( .B(n47187), .A(n47188), .Z(n50573) );
  XNOR U49880 ( .A(n50575), .B(n50576), .Z(n41730) );
  ANDN U49881 ( .B(n47191), .A(n47192), .Z(n50575) );
  XNOR U49882 ( .A(n50577), .B(n50578), .Z(n50571) );
  XNOR U49883 ( .A(n45254), .B(n49416), .Z(n50578) );
  XNOR U49884 ( .A(n50579), .B(n50580), .Z(n49416) );
  ANDN U49885 ( .B(n47181), .A(n47182), .Z(n50579) );
  XNOR U49886 ( .A(n50581), .B(n50582), .Z(n45254) );
  AND U49887 ( .A(n48037), .B(n48035), .Z(n50581) );
  XNOR U49888 ( .A(n50583), .B(n50584), .Z(n47196) );
  AND U49889 ( .A(n48054), .B(n48704), .Z(n50583) );
  XOR U49890 ( .A(round_reg[1445]), .B(n48566), .Z(n48054) );
  XOR U49891 ( .A(n45348), .B(n49029), .Z(n45016) );
  XOR U49892 ( .A(n50585), .B(n50545), .Z(n49029) );
  NOR U49893 ( .A(n47905), .B(n50586), .Z(n50585) );
  IV U49894 ( .A(n50587), .Z(n47905) );
  IV U49895 ( .A(n42855), .Z(n45348) );
  XNOR U49896 ( .A(n50590), .B(n43242), .Z(n41715) );
  XOR U49897 ( .A(n50591), .B(n45082), .Z(n43242) );
  IV U49898 ( .A(n43287), .Z(n45082) );
  XOR U49899 ( .A(n49602), .B(n47355), .Z(n43287) );
  XNOR U49900 ( .A(n50592), .B(n50593), .Z(n47355) );
  XNOR U49901 ( .A(n50594), .B(n43544), .Z(n50593) );
  XNOR U49902 ( .A(n50595), .B(n50389), .Z(n43544) );
  AND U49903 ( .A(n50596), .B(n50597), .Z(n50595) );
  XOR U49904 ( .A(n45401), .B(n50598), .Z(n50592) );
  XOR U49905 ( .A(n44687), .B(n50599), .Z(n50598) );
  XNOR U49906 ( .A(n50600), .B(n50379), .Z(n44687) );
  XNOR U49907 ( .A(n50603), .B(n50385), .Z(n45401) );
  XOR U49908 ( .A(n50606), .B(n50607), .Z(n49602) );
  XOR U49909 ( .A(n49112), .B(n45956), .Z(n50607) );
  XOR U49910 ( .A(n50608), .B(n48326), .Z(n45956) );
  NOR U49911 ( .A(n46785), .B(n46784), .Z(n50608) );
  XNOR U49912 ( .A(n50609), .B(n48338), .Z(n49112) );
  NOR U49913 ( .A(n49600), .B(n49601), .Z(n50609) );
  XOR U49914 ( .A(n47667), .B(n50610), .Z(n50606) );
  XNOR U49915 ( .A(n46095), .B(n45090), .Z(n50610) );
  XOR U49916 ( .A(n50611), .B(n48330), .Z(n45090) );
  ANDN U49917 ( .B(n46777), .A(n46778), .Z(n50611) );
  XNOR U49918 ( .A(n50612), .B(n50613), .Z(n46095) );
  ANDN U49919 ( .B(n47531), .A(n47532), .Z(n50612) );
  XNOR U49920 ( .A(n50614), .B(n48334), .Z(n47667) );
  ANDN U49921 ( .B(n48909), .A(n48910), .Z(n50614) );
  ANDN U49922 ( .B(n45018), .A(n45457), .Z(n50590) );
  XNOR U49923 ( .A(n49275), .B(n45167), .Z(n45457) );
  XOR U49924 ( .A(n50615), .B(n46434), .Z(n45167) );
  XNOR U49925 ( .A(n50616), .B(n50617), .Z(n46434) );
  XOR U49926 ( .A(n46180), .B(n46459), .Z(n50617) );
  XNOR U49927 ( .A(n50618), .B(n49530), .Z(n46459) );
  NOR U49928 ( .A(n50619), .B(n50620), .Z(n50618) );
  XOR U49929 ( .A(n50621), .B(n50622), .Z(n46180) );
  ANDN U49930 ( .B(n50623), .A(n50624), .Z(n50621) );
  XNOR U49931 ( .A(n46172), .B(n50625), .Z(n50616) );
  XNOR U49932 ( .A(n50626), .B(n46765), .Z(n50625) );
  XOR U49933 ( .A(n50627), .B(n49160), .Z(n46765) );
  ANDN U49934 ( .B(n50628), .A(n50629), .Z(n50627) );
  XNOR U49935 ( .A(n50630), .B(n49423), .Z(n46172) );
  ANDN U49936 ( .B(n50631), .A(n50632), .Z(n50630) );
  XNOR U49937 ( .A(n50633), .B(n50634), .Z(n49275) );
  NOR U49938 ( .A(n48840), .B(n48841), .Z(n50633) );
  XOR U49939 ( .A(round_reg[220]), .B(n48876), .Z(n48841) );
  IV U49940 ( .A(n50635), .Z(n48876) );
  XNOR U49941 ( .A(n50636), .B(n50637), .Z(n49969) );
  ANDN U49942 ( .B(n50638), .A(n49364), .Z(n50636) );
  XNOR U49943 ( .A(n49619), .B(n50639), .Z(n45504) );
  XOR U49944 ( .A(n50640), .B(n50641), .Z(n49619) );
  XOR U49945 ( .A(n48504), .B(n44332), .Z(n50641) );
  XOR U49946 ( .A(n50642), .B(n48540), .Z(n44332) );
  XNOR U49947 ( .A(round_reg[646]), .B(n50643), .Z(n48540) );
  NOR U49948 ( .A(n49883), .B(n49884), .Z(n50642) );
  XNOR U49949 ( .A(round_reg[580]), .B(n49612), .Z(n49883) );
  XOR U49950 ( .A(n50644), .B(n48536), .Z(n48504) );
  XOR U49951 ( .A(round_reg[724]), .B(n50645), .Z(n48536) );
  ANDN U49952 ( .B(n48535), .A(n49874), .Z(n50644) );
  XNOR U49953 ( .A(round_reg[357]), .B(n50646), .Z(n48535) );
  XNOR U49954 ( .A(n46640), .B(n50647), .Z(n50640) );
  XOR U49955 ( .A(n44527), .B(n45284), .Z(n50647) );
  XOR U49956 ( .A(n50648), .B(n48531), .Z(n45284) );
  XOR U49957 ( .A(round_reg[770]), .B(n50455), .Z(n48531) );
  ANDN U49958 ( .B(n48530), .A(n49881), .Z(n50648) );
  XNOR U49959 ( .A(round_reg[408]), .B(n48441), .Z(n48530) );
  XOR U49960 ( .A(n50649), .B(n48544), .Z(n44527) );
  XOR U49961 ( .A(round_reg[867]), .B(n48450), .Z(n48544) );
  ANDN U49962 ( .B(n48543), .A(n49879), .Z(n50649) );
  XNOR U49963 ( .A(n50651), .B(n48526), .Z(n46640) );
  XNOR U49964 ( .A(round_reg[938]), .B(n48356), .Z(n48526) );
  ANDN U49965 ( .B(n48527), .A(n49876), .Z(n50651) );
  XOR U49966 ( .A(round_reg[512]), .B(n50415), .Z(n48527) );
  XNOR U49967 ( .A(n50652), .B(n33751), .Z(n35651) );
  XNOR U49968 ( .A(n35926), .B(n40862), .Z(n33751) );
  XNOR U49969 ( .A(n50653), .B(n41610), .Z(n40862) );
  AND U49970 ( .A(n43488), .B(n49230), .Z(n50653) );
  XNOR U49971 ( .A(n50654), .B(n45945), .Z(n43488) );
  XOR U49972 ( .A(n43685), .B(n40906), .Z(n35926) );
  XOR U49973 ( .A(n50655), .B(n50656), .Z(n40906) );
  XNOR U49974 ( .A(n34619), .B(n40923), .Z(n50656) );
  XNOR U49975 ( .A(n50657), .B(n43482), .Z(n40923) );
  XOR U49976 ( .A(n50658), .B(n44186), .Z(n43482) );
  XOR U49977 ( .A(n47932), .B(n48352), .Z(n44186) );
  XNOR U49978 ( .A(n50659), .B(n50660), .Z(n48352) );
  XNOR U49979 ( .A(n46159), .B(n50661), .Z(n50660) );
  XNOR U49980 ( .A(n50662), .B(n46622), .Z(n46159) );
  ANDN U49981 ( .B(n50663), .A(n48980), .Z(n50662) );
  XOR U49982 ( .A(n44473), .B(n50664), .Z(n50659) );
  XOR U49983 ( .A(n45506), .B(n46719), .Z(n50664) );
  XNOR U49984 ( .A(n50665), .B(n46951), .Z(n46719) );
  NOR U49985 ( .A(n48978), .B(n50666), .Z(n50665) );
  XNOR U49986 ( .A(n50667), .B(n46612), .Z(n45506) );
  NOR U49987 ( .A(n48974), .B(n50668), .Z(n50667) );
  XNOR U49988 ( .A(n50669), .B(n46609), .Z(n44473) );
  ANDN U49989 ( .B(n50670), .A(n48972), .Z(n50669) );
  XNOR U49990 ( .A(n50671), .B(n50672), .Z(n47932) );
  XOR U49991 ( .A(n47545), .B(n44511), .Z(n50672) );
  XOR U49992 ( .A(n50673), .B(n49197), .Z(n44511) );
  ANDN U49993 ( .B(n50674), .A(n50675), .Z(n50673) );
  XOR U49994 ( .A(n50676), .B(n50677), .Z(n47545) );
  XOR U49995 ( .A(n47065), .B(n50680), .Z(n50671) );
  XOR U49996 ( .A(n46404), .B(n46661), .Z(n50680) );
  XNOR U49997 ( .A(n50681), .B(n49187), .Z(n46661) );
  ANDN U49998 ( .B(n50682), .A(n50683), .Z(n50681) );
  XNOR U49999 ( .A(n50684), .B(n50685), .Z(n46404) );
  ANDN U50000 ( .B(n50686), .A(n50687), .Z(n50684) );
  XNOR U50001 ( .A(n50688), .B(n49190), .Z(n47065) );
  ANDN U50002 ( .B(n50689), .A(n50690), .Z(n50688) );
  ANDN U50003 ( .B(n40864), .A(n40865), .Z(n50657) );
  XOR U50004 ( .A(n45014), .B(n47983), .Z(n40865) );
  XNOR U50005 ( .A(n50691), .B(n50692), .Z(n47983) );
  ANDN U50006 ( .B(n50301), .A(n49719), .Z(n50691) );
  XOR U50007 ( .A(round_reg[877]), .B(n50693), .Z(n49719) );
  IV U50008 ( .A(n50694), .Z(n45014) );
  XNOR U50009 ( .A(n44767), .B(n48817), .Z(n40864) );
  XNOR U50010 ( .A(n50695), .B(n50696), .Z(n48817) );
  ANDN U50011 ( .B(n49682), .A(n50697), .Z(n50695) );
  IV U50012 ( .A(n43282), .Z(n44767) );
  XNOR U50013 ( .A(n50698), .B(n49705), .Z(n43282) );
  XNOR U50014 ( .A(n50699), .B(n50700), .Z(n49705) );
  XOR U50015 ( .A(n49524), .B(n50270), .Z(n50700) );
  XOR U50016 ( .A(n50701), .B(n50282), .Z(n50270) );
  ANDN U50017 ( .B(n50283), .A(n47707), .Z(n50701) );
  XOR U50018 ( .A(n50702), .B(n50289), .Z(n49524) );
  ANDN U50019 ( .B(n50290), .A(n47703), .Z(n50702) );
  XOR U50020 ( .A(n48981), .B(n50703), .Z(n50699) );
  XOR U50021 ( .A(n44551), .B(n42867), .Z(n50703) );
  XOR U50022 ( .A(n50704), .B(n50278), .Z(n42867) );
  ANDN U50023 ( .B(n50279), .A(n50705), .Z(n50704) );
  XNOR U50024 ( .A(n50706), .B(n50274), .Z(n44551) );
  ANDN U50025 ( .B(n50275), .A(n47717), .Z(n50706) );
  XNOR U50026 ( .A(n50707), .B(n50285), .Z(n48981) );
  ANDN U50027 ( .B(n50286), .A(n47713), .Z(n50707) );
  XOR U50028 ( .A(n50708), .B(n40933), .Z(n34619) );
  XOR U50029 ( .A(n43298), .B(n45867), .Z(n40933) );
  XNOR U50030 ( .A(n50709), .B(n49577), .Z(n45867) );
  NOR U50031 ( .A(n50710), .B(n47636), .Z(n50709) );
  XNOR U50032 ( .A(n49978), .B(n47004), .Z(n43298) );
  XNOR U50033 ( .A(n50711), .B(n50712), .Z(n47004) );
  XNOR U50034 ( .A(n48285), .B(n46104), .Z(n50712) );
  XOR U50035 ( .A(n50713), .B(n48187), .Z(n46104) );
  XNOR U50036 ( .A(round_reg[68]), .B(n50714), .Z(n48187) );
  XOR U50037 ( .A(round_reg[1313]), .B(n50715), .Z(n45882) );
  IV U50038 ( .A(n50716), .Z(n45883) );
  XNOR U50039 ( .A(n50717), .B(n47676), .Z(n48285) );
  XNOR U50040 ( .A(round_reg[46]), .B(n50718), .Z(n47676) );
  ANDN U50041 ( .B(n45869), .A(n45870), .Z(n50717) );
  XOR U50042 ( .A(round_reg[1596]), .B(n50719), .Z(n45869) );
  XNOR U50043 ( .A(n49559), .B(n50720), .Z(n50711) );
  XOR U50044 ( .A(n45140), .B(n42313), .Z(n50720) );
  XNOR U50045 ( .A(n50721), .B(n47637), .Z(n42313) );
  XNOR U50046 ( .A(round_reg[191]), .B(n49081), .Z(n47637) );
  ANDN U50047 ( .B(n49577), .A(n50722), .Z(n50721) );
  XOR U50048 ( .A(round_reg[1376]), .B(n50723), .Z(n49577) );
  XNOR U50049 ( .A(n50724), .B(n49574), .Z(n45140) );
  XOR U50050 ( .A(round_reg[1531]), .B(n49080), .Z(n45878) );
  IV U50051 ( .A(n50725), .Z(n45879) );
  XOR U50052 ( .A(n50726), .B(n46761), .Z(n49559) );
  XOR U50053 ( .A(round_reg[250]), .B(n50727), .Z(n46761) );
  ANDN U50054 ( .B(n45874), .A(n45876), .Z(n50726) );
  XNOR U50055 ( .A(round_reg[1470]), .B(n50728), .Z(n45874) );
  XOR U50056 ( .A(n50729), .B(n50730), .Z(n49978) );
  XOR U50057 ( .A(n43308), .B(n44480), .Z(n50730) );
  XOR U50058 ( .A(n50731), .B(n47103), .Z(n44480) );
  XNOR U50059 ( .A(round_reg[999]), .B(n50732), .Z(n47103) );
  ANDN U50060 ( .B(n49563), .A(n49994), .Z(n50731) );
  XNOR U50061 ( .A(round_reg[952]), .B(n50733), .Z(n49563) );
  XNOR U50062 ( .A(n50734), .B(n46905), .Z(n43308) );
  XOR U50063 ( .A(round_reg[1167]), .B(n50401), .Z(n46905) );
  ANDN U50064 ( .B(n48383), .A(n48384), .Z(n50734) );
  XNOR U50065 ( .A(round_reg[784]), .B(n50735), .Z(n48383) );
  XOR U50066 ( .A(n44948), .B(n50736), .Z(n50729) );
  XOR U50067 ( .A(n41744), .B(n45749), .Z(n50736) );
  XNOR U50068 ( .A(n50737), .B(n47572), .Z(n45749) );
  XOR U50069 ( .A(round_reg[1239]), .B(n50738), .Z(n47572) );
  ANDN U50070 ( .B(n49432), .A(n49433), .Z(n50737) );
  XOR U50071 ( .A(round_reg[881]), .B(n50739), .Z(n49432) );
  XNOR U50072 ( .A(n50740), .B(n46909), .Z(n41744) );
  XOR U50073 ( .A(round_reg[1028]), .B(n50741), .Z(n46909) );
  ANDN U50074 ( .B(n48374), .A(n48375), .Z(n50740) );
  XNOR U50075 ( .A(round_reg[660]), .B(n50742), .Z(n48374) );
  XNOR U50076 ( .A(n50743), .B(n46899), .Z(n44948) );
  XOR U50077 ( .A(round_reg[1141]), .B(n50744), .Z(n46899) );
  ANDN U50078 ( .B(n48377), .A(n48378), .Z(n50743) );
  XNOR U50079 ( .A(round_reg[738]), .B(n50745), .Z(n48377) );
  NOR U50080 ( .A(n40875), .B(n40874), .Z(n50708) );
  XNOR U50081 ( .A(n50151), .B(n47603), .Z(n40874) );
  IV U50082 ( .A(n45085), .Z(n47603) );
  XNOR U50083 ( .A(n50746), .B(n50747), .Z(n48265) );
  XNOR U50084 ( .A(n45296), .B(n47028), .Z(n50747) );
  XNOR U50085 ( .A(n50748), .B(n48315), .Z(n47028) );
  NOR U50086 ( .A(n50166), .B(n48314), .Z(n50748) );
  XOR U50087 ( .A(round_reg[620]), .B(n50749), .Z(n48314) );
  XNOR U50088 ( .A(n50750), .B(n47748), .Z(n45296) );
  XNOR U50089 ( .A(round_reg[764]), .B(n50751), .Z(n47748) );
  NOR U50090 ( .A(n47747), .B(n50172), .Z(n50750) );
  XOR U50091 ( .A(round_reg[333]), .B(n50752), .Z(n47747) );
  XOR U50092 ( .A(n46935), .B(n50753), .Z(n50746) );
  XOR U50093 ( .A(n45826), .B(n45005), .Z(n50753) );
  XNOR U50094 ( .A(n50754), .B(n50063), .Z(n45005) );
  XOR U50095 ( .A(round_reg[914]), .B(n50755), .Z(n50063) );
  NOR U50096 ( .A(n50069), .B(n50169), .Z(n50754) );
  XNOR U50097 ( .A(round_reg[552]), .B(n50756), .Z(n50069) );
  XNOR U50098 ( .A(n50757), .B(n49804), .Z(n45826) );
  XNOR U50099 ( .A(round_reg[843]), .B(n50758), .Z(n49804) );
  ANDN U50100 ( .B(n49805), .A(n50163), .Z(n50757) );
  XNOR U50101 ( .A(round_reg[454]), .B(n50759), .Z(n49805) );
  XNOR U50102 ( .A(n50760), .B(n47755), .Z(n46935) );
  XOR U50103 ( .A(round_reg[810]), .B(n50761), .Z(n47755) );
  NOR U50104 ( .A(n50174), .B(n47754), .Z(n50760) );
  XNOR U50105 ( .A(round_reg[384]), .B(n50407), .Z(n47754) );
  IV U50106 ( .A(n50762), .Z(n50174) );
  XOR U50107 ( .A(n50764), .B(n47770), .Z(n50151) );
  AND U50108 ( .A(n49121), .B(n49120), .Z(n50764) );
  XOR U50109 ( .A(round_reg[334]), .B(n50765), .Z(n49121) );
  XOR U50110 ( .A(n50257), .B(n44523), .Z(n40875) );
  XNOR U50111 ( .A(n50766), .B(n50767), .Z(n48437) );
  XOR U50112 ( .A(n46519), .B(n44746), .Z(n50767) );
  XOR U50113 ( .A(n50768), .B(n50769), .Z(n44746) );
  AND U50114 ( .A(n48460), .B(n48458), .Z(n50768) );
  XNOR U50115 ( .A(n50770), .B(n50568), .Z(n46519) );
  ANDN U50116 ( .B(n47803), .A(n50771), .Z(n50770) );
  XNOR U50117 ( .A(round_reg[206]), .B(n50772), .Z(n47803) );
  XOR U50118 ( .A(n46530), .B(n50773), .Z(n50766) );
  XOR U50119 ( .A(n45735), .B(n45402), .Z(n50773) );
  XNOR U50120 ( .A(n50774), .B(n50557), .Z(n45402) );
  AND U50121 ( .A(n47791), .B(n47789), .Z(n50774) );
  XOR U50122 ( .A(round_reg[2]), .B(n50775), .Z(n47789) );
  XNOR U50123 ( .A(n50776), .B(n50560), .Z(n45735) );
  XNOR U50124 ( .A(round_reg[318]), .B(n50777), .Z(n47799) );
  XNOR U50125 ( .A(n50778), .B(n50565), .Z(n46530) );
  AND U50126 ( .A(n47795), .B(n47793), .Z(n50778) );
  XNOR U50127 ( .A(round_reg[147]), .B(n49904), .Z(n47793) );
  XNOR U50128 ( .A(n50780), .B(n50781), .Z(n50257) );
  AND U50129 ( .A(n50782), .B(n50783), .Z(n50780) );
  XOR U50130 ( .A(n40902), .B(n50784), .Z(n50655) );
  XOR U50131 ( .A(n35591), .B(n39132), .Z(n50784) );
  XNOR U50132 ( .A(n50785), .B(n40929), .Z(n39132) );
  XOR U50133 ( .A(n50786), .B(n43713), .Z(n40929) );
  IV U50134 ( .A(n48401), .Z(n43713) );
  XOR U50135 ( .A(n50788), .B(n50789), .Z(n46100) );
  XOR U50136 ( .A(n45824), .B(n48573), .Z(n50789) );
  XOR U50137 ( .A(n50790), .B(n50791), .Z(n48573) );
  AND U50138 ( .A(n48995), .B(n50792), .Z(n50790) );
  XNOR U50139 ( .A(n50793), .B(n50794), .Z(n45824) );
  ANDN U50140 ( .B(n49001), .A(n50795), .Z(n50793) );
  XOR U50141 ( .A(n44840), .B(n50796), .Z(n50788) );
  XOR U50142 ( .A(n44885), .B(n45459), .Z(n50796) );
  XNOR U50143 ( .A(n50797), .B(n50798), .Z(n45459) );
  XNOR U50144 ( .A(n50801), .B(n50802), .Z(n44885) );
  ANDN U50145 ( .B(n48991), .A(n50803), .Z(n50801) );
  XNOR U50146 ( .A(n50804), .B(n50805), .Z(n44840) );
  AND U50147 ( .A(n49005), .B(n50806), .Z(n50804) );
  NOR U50148 ( .A(n40930), .B(n40871), .Z(n50785) );
  XOR U50149 ( .A(n45400), .B(n50599), .Z(n40871) );
  XNOR U50150 ( .A(n50807), .B(n50808), .Z(n50599) );
  IV U50151 ( .A(n43543), .Z(n45400) );
  XNOR U50152 ( .A(n48278), .B(n43925), .Z(n40930) );
  XNOR U50153 ( .A(n50811), .B(n50812), .Z(n49352) );
  XNOR U50154 ( .A(n45651), .B(n41640), .Z(n50812) );
  XOR U50155 ( .A(n50813), .B(n47278), .Z(n41640) );
  XOR U50156 ( .A(round_reg[56]), .B(n50486), .Z(n47278) );
  ANDN U50157 ( .B(n47279), .A(n47306), .Z(n50813) );
  XOR U50158 ( .A(round_reg[1178]), .B(n50814), .Z(n47306) );
  XNOR U50159 ( .A(round_reg[1542]), .B(n50815), .Z(n47279) );
  XNOR U50160 ( .A(n50816), .B(n47269), .Z(n45651) );
  XOR U50161 ( .A(round_reg[308]), .B(n50299), .Z(n47269) );
  AND U50162 ( .A(n48008), .B(n47270), .Z(n50816) );
  XNOR U50163 ( .A(round_reg[1477]), .B(n48453), .Z(n47270) );
  XNOR U50164 ( .A(round_reg[1088]), .B(n49083), .Z(n48008) );
  XOR U50165 ( .A(n46792), .B(n50817), .Z(n50811) );
  XOR U50166 ( .A(n45790), .B(n46277), .Z(n50817) );
  XNOR U50167 ( .A(n50818), .B(n47283), .Z(n46277) );
  XNOR U50168 ( .A(round_reg[137]), .B(n50124), .Z(n47283) );
  NOR U50169 ( .A(n47282), .B(n47302), .Z(n50818) );
  XNOR U50170 ( .A(round_reg[1010]), .B(n50404), .Z(n47302) );
  XOR U50171 ( .A(round_reg[1386]), .B(n50819), .Z(n47282) );
  XNOR U50172 ( .A(n50820), .B(n47274), .Z(n45790) );
  ANDN U50173 ( .B(n47275), .A(n47314), .Z(n50820) );
  XOR U50174 ( .A(round_reg[1039]), .B(n48553), .Z(n47314) );
  XOR U50175 ( .A(round_reg[1416]), .B(n50497), .Z(n47275) );
  XNOR U50176 ( .A(n50821), .B(n50492), .Z(n46792) );
  ANDN U50177 ( .B(n47310), .A(n47311), .Z(n50821) );
  XNOR U50178 ( .A(round_reg[1250]), .B(n50822), .Z(n47311) );
  XOR U50179 ( .A(round_reg[1323]), .B(n50823), .Z(n47310) );
  XOR U50180 ( .A(n50824), .B(n50825), .Z(n49441) );
  XNOR U50181 ( .A(n47262), .B(n44931), .Z(n50825) );
  XOR U50182 ( .A(n50826), .B(n48201), .Z(n44931) );
  XNOR U50183 ( .A(round_reg[796]), .B(n50827), .Z(n48201) );
  ANDN U50184 ( .B(n48202), .A(n48284), .Z(n50826) );
  XNOR U50185 ( .A(round_reg[57]), .B(n50828), .Z(n48284) );
  XNOR U50186 ( .A(round_reg[434]), .B(n50829), .Z(n48202) );
  XNOR U50187 ( .A(n50830), .B(n48210), .Z(n47262) );
  XNOR U50188 ( .A(round_reg[750]), .B(n50831), .Z(n48210) );
  ANDN U50189 ( .B(n48211), .A(n49013), .Z(n50830) );
  XOR U50190 ( .A(n44776), .B(n50832), .Z(n50824) );
  XOR U50191 ( .A(n46019), .B(n46094), .Z(n50832) );
  XNOR U50192 ( .A(n50833), .B(n48214), .Z(n46094) );
  XOR U50193 ( .A(round_reg[672]), .B(n50834), .Z(n48214) );
  XNOR U50194 ( .A(round_reg[197]), .B(n48453), .Z(n48276) );
  XOR U50195 ( .A(round_reg[606]), .B(n50835), .Z(n48215) );
  XNOR U50196 ( .A(n50836), .B(n50134), .Z(n46019) );
  IV U50197 ( .A(n48205), .Z(n50134) );
  XOR U50198 ( .A(round_reg[893]), .B(n50837), .Z(n48205) );
  ANDN U50199 ( .B(n48206), .A(n48661), .Z(n50836) );
  XOR U50200 ( .A(round_reg[79]), .B(n48553), .Z(n48661) );
  XOR U50201 ( .A(round_reg[504]), .B(n50838), .Z(n48206) );
  XNOR U50202 ( .A(n50839), .B(n48218), .Z(n44776) );
  XOR U50203 ( .A(round_reg[900]), .B(n49612), .Z(n48218) );
  ANDN U50204 ( .B(n48219), .A(n48280), .Z(n50839) );
  XOR U50205 ( .A(round_reg[138]), .B(n50117), .Z(n48280) );
  XOR U50206 ( .A(round_reg[538]), .B(n50814), .Z(n48219) );
  XNOR U50207 ( .A(n50840), .B(n48211), .Z(n48278) );
  XNOR U50208 ( .A(round_reg[383]), .B(n50841), .Z(n48211) );
  ANDN U50209 ( .B(n49013), .A(n50126), .Z(n50840) );
  IV U50210 ( .A(n49014), .Z(n50126) );
  XOR U50211 ( .A(round_reg[1478]), .B(n50116), .Z(n49014) );
  XNOR U50212 ( .A(round_reg[309]), .B(n50842), .Z(n49013) );
  XNOR U50213 ( .A(n50843), .B(n40939), .Z(n35591) );
  XOR U50214 ( .A(n46637), .B(n47898), .Z(n40939) );
  XOR U50215 ( .A(n50844), .B(n49032), .Z(n47898) );
  ANDN U50216 ( .B(n50539), .A(n50845), .Z(n50844) );
  IV U50217 ( .A(n44461), .Z(n46637) );
  XNOR U50218 ( .A(n50846), .B(n50847), .Z(n49536) );
  XNOR U50219 ( .A(n46088), .B(n49026), .Z(n50847) );
  XNOR U50220 ( .A(n50848), .B(n50586), .Z(n49026) );
  ANDN U50221 ( .B(n47907), .A(n50587), .Z(n50848) );
  XOR U50222 ( .A(round_reg[84]), .B(n50849), .Z(n50587) );
  XNOR U50223 ( .A(round_reg[1329]), .B(n50498), .Z(n47907) );
  XOR U50224 ( .A(n50850), .B(n50851), .Z(n46088) );
  AND U50225 ( .A(n47897), .B(n47895), .Z(n50850) );
  XOR U50226 ( .A(round_reg[202]), .B(n50852), .Z(n47895) );
  XOR U50227 ( .A(round_reg[1422]), .B(n50853), .Z(n47897) );
  XNOR U50228 ( .A(n46067), .B(n50854), .Z(n50846) );
  XOR U50229 ( .A(n45834), .B(n45752), .Z(n50854) );
  XNOR U50230 ( .A(n50855), .B(n49468), .Z(n45752) );
  ANDN U50231 ( .B(n49467), .A(n47892), .Z(n50855) );
  XOR U50232 ( .A(round_reg[1548]), .B(n48456), .Z(n47892) );
  IV U50233 ( .A(n49427), .Z(n48456) );
  IV U50234 ( .A(n47891), .Z(n49467) );
  XOR U50235 ( .A(round_reg[62]), .B(n50516), .Z(n47891) );
  XNOR U50236 ( .A(n50856), .B(n49041), .Z(n45834) );
  ANDN U50237 ( .B(n47903), .A(n49042), .Z(n50856) );
  XOR U50238 ( .A(round_reg[314]), .B(n50857), .Z(n49042) );
  XOR U50239 ( .A(round_reg[1483]), .B(n50758), .Z(n47903) );
  XNOR U50240 ( .A(n50858), .B(n49033), .Z(n46067) );
  NOR U50241 ( .A(n50539), .B(n49032), .Z(n50858) );
  XOR U50242 ( .A(round_reg[143]), .B(n50859), .Z(n49032) );
  XOR U50243 ( .A(round_reg[1392]), .B(n49178), .Z(n50539) );
  XNOR U50244 ( .A(n50860), .B(n50861), .Z(n48012) );
  XNOR U50245 ( .A(n45885), .B(n45501), .Z(n50861) );
  XOR U50246 ( .A(n50862), .B(n49049), .Z(n45501) );
  NOR U50247 ( .A(n50863), .B(n49048), .Z(n50862) );
  XNOR U50248 ( .A(n50864), .B(n50865), .Z(n45885) );
  NOR U50249 ( .A(n50866), .B(n50867), .Z(n50864) );
  XNOR U50250 ( .A(n46830), .B(n50868), .Z(n50860) );
  XOR U50251 ( .A(n43832), .B(n43655), .Z(n50868) );
  XNOR U50252 ( .A(n50869), .B(n49054), .Z(n43655) );
  ANDN U50253 ( .B(n50870), .A(n49053), .Z(n50869) );
  XNOR U50254 ( .A(n50871), .B(n49057), .Z(n43832) );
  AND U50255 ( .A(n50872), .B(n49058), .Z(n50871) );
  XNOR U50256 ( .A(n50873), .B(n49062), .Z(n46830) );
  ANDN U50257 ( .B(n50874), .A(n49061), .Z(n50873) );
  ANDN U50258 ( .B(n40940), .A(n41548), .Z(n50843) );
  XOR U50259 ( .A(n49762), .B(n43329), .Z(n41548) );
  XNOR U50260 ( .A(n50349), .B(n48085), .Z(n43329) );
  XNOR U50261 ( .A(n50875), .B(n50876), .Z(n48085) );
  XNOR U50262 ( .A(n45338), .B(n46351), .Z(n50876) );
  XNOR U50263 ( .A(n50877), .B(n50878), .Z(n46351) );
  NOR U50264 ( .A(n50879), .B(n49741), .Z(n50877) );
  XNOR U50265 ( .A(round_reg[240]), .B(n48938), .Z(n49741) );
  XNOR U50266 ( .A(n50880), .B(n50881), .Z(n45338) );
  ANDN U50267 ( .B(n49745), .A(n49744), .Z(n50880) );
  XOR U50268 ( .A(round_reg[122]), .B(n50882), .Z(n49745) );
  XNOR U50269 ( .A(n48929), .B(n50883), .Z(n50875) );
  XOR U50270 ( .A(n46307), .B(n46722), .Z(n50883) );
  XNOR U50271 ( .A(n50884), .B(n50885), .Z(n46722) );
  NOR U50272 ( .A(n49748), .B(n49749), .Z(n50884) );
  XOR U50273 ( .A(round_reg[181]), .B(n50744), .Z(n49749) );
  XNOR U50274 ( .A(n50886), .B(n50887), .Z(n46307) );
  ANDN U50275 ( .B(n49731), .A(n49732), .Z(n50886) );
  XNOR U50276 ( .A(round_reg[36]), .B(n50888), .Z(n49732) );
  XNOR U50277 ( .A(n50889), .B(n50890), .Z(n48929) );
  XOR U50278 ( .A(round_reg[288]), .B(n49860), .Z(n49736) );
  XOR U50279 ( .A(n50891), .B(n50892), .Z(n50349) );
  XOR U50280 ( .A(n43560), .B(n46007), .Z(n50892) );
  XNOR U50281 ( .A(n50893), .B(n50018), .Z(n46007) );
  XNOR U50282 ( .A(n50894), .B(n50005), .Z(n43560) );
  ANDN U50283 ( .B(n49760), .A(n50895), .Z(n50894) );
  XOR U50284 ( .A(n50072), .B(n50896), .Z(n50891) );
  XOR U50285 ( .A(n50897), .B(n44940), .Z(n50896) );
  XNOR U50286 ( .A(n50898), .B(n50012), .Z(n44940) );
  XNOR U50287 ( .A(n50899), .B(n50016), .Z(n50072) );
  NOR U50288 ( .A(n50900), .B(n50901), .Z(n50899) );
  XNOR U50289 ( .A(n50902), .B(n50901), .Z(n49762) );
  AND U50290 ( .A(n50014), .B(n50900), .Z(n50902) );
  XOR U50291 ( .A(n50903), .B(n43767), .Z(n40940) );
  XNOR U50292 ( .A(n50904), .B(n50905), .Z(n47694) );
  XOR U50293 ( .A(n45278), .B(n42876), .Z(n50905) );
  XOR U50294 ( .A(n50906), .B(n50628), .Z(n42876) );
  ANDN U50295 ( .B(n50629), .A(n49159), .Z(n50906) );
  XNOR U50296 ( .A(n50907), .B(n50623), .Z(n45278) );
  ANDN U50297 ( .B(n50624), .A(n50908), .Z(n50907) );
  XNOR U50298 ( .A(n46432), .B(n50909), .Z(n50904) );
  XOR U50299 ( .A(n45833), .B(n46097), .Z(n50909) );
  XOR U50300 ( .A(n50910), .B(n50911), .Z(n46097) );
  XNOR U50301 ( .A(n50914), .B(n50619), .Z(n45833) );
  XOR U50302 ( .A(n50915), .B(n50631), .Z(n46432) );
  AND U50303 ( .A(n49422), .B(n50632), .Z(n50915) );
  XNOR U50304 ( .A(n50916), .B(n50917), .Z(n46273) );
  XNOR U50305 ( .A(n46229), .B(n47528), .Z(n50917) );
  XNOR U50306 ( .A(n50918), .B(n48905), .Z(n47528) );
  AND U50307 ( .A(n50919), .B(n48906), .Z(n50918) );
  XOR U50308 ( .A(n50920), .B(n48898), .Z(n46229) );
  NOR U50309 ( .A(n48897), .B(n50921), .Z(n50920) );
  XNOR U50310 ( .A(n48885), .B(n50922), .Z(n50916) );
  XNOR U50311 ( .A(n46197), .B(n47390), .Z(n50922) );
  XNOR U50312 ( .A(n50923), .B(n48901), .Z(n47390) );
  ANDN U50313 ( .B(n48902), .A(n50924), .Z(n50923) );
  XNOR U50314 ( .A(n50925), .B(n48892), .Z(n46197) );
  ANDN U50315 ( .B(n48893), .A(n50926), .Z(n50925) );
  XNOR U50316 ( .A(n50927), .B(n50328), .Z(n48885) );
  AND U50317 ( .A(n50928), .B(n50329), .Z(n50927) );
  XNOR U50318 ( .A(n50929), .B(n41609), .Z(n40902) );
  XOR U50319 ( .A(n47724), .B(n44195), .Z(n41609) );
  IV U50320 ( .A(n46702), .Z(n44195) );
  XOR U50321 ( .A(n50183), .B(n47098), .Z(n46702) );
  XNOR U50322 ( .A(n50930), .B(n50931), .Z(n47098) );
  XOR U50323 ( .A(n47381), .B(n46413), .Z(n50931) );
  XNOR U50324 ( .A(n50932), .B(n49765), .Z(n46413) );
  XOR U50325 ( .A(round_reg[652]), .B(n50933), .Z(n49765) );
  ANDN U50326 ( .B(n49766), .A(n50011), .Z(n50932) );
  XOR U50327 ( .A(round_reg[586]), .B(n50934), .Z(n49766) );
  XNOR U50328 ( .A(n50935), .B(n50936), .Z(n47381) );
  ANDN U50329 ( .B(n49770), .A(n50007), .Z(n50935) );
  XOR U50330 ( .A(round_reg[363]), .B(n50823), .Z(n49770) );
  XNOR U50331 ( .A(n46446), .B(n50937), .Z(n50930) );
  XOR U50332 ( .A(n49727), .B(n47814), .Z(n50937) );
  XOR U50333 ( .A(n50938), .B(n49755), .Z(n47814) );
  XNOR U50334 ( .A(round_reg[944]), .B(n50939), .Z(n49755) );
  AND U50335 ( .A(n50019), .B(n49756), .Z(n50938) );
  XOR U50336 ( .A(round_reg[518]), .B(n50940), .Z(n49756) );
  XNOR U50337 ( .A(n50941), .B(n50900), .Z(n49727) );
  XOR U50338 ( .A(round_reg[873]), .B(n50942), .Z(n50900) );
  NOR U50339 ( .A(n50014), .B(n50015), .Z(n50941) );
  XOR U50340 ( .A(round_reg[484]), .B(n48449), .Z(n50014) );
  XNOR U50341 ( .A(n50943), .B(n49760), .Z(n46446) );
  XNOR U50342 ( .A(round_reg[776]), .B(n50497), .Z(n49760) );
  ANDN U50343 ( .B(n49759), .A(n50004), .Z(n50943) );
  XOR U50344 ( .A(round_reg[414]), .B(n49606), .Z(n49759) );
  XOR U50345 ( .A(n50944), .B(n50945), .Z(n50183) );
  XOR U50346 ( .A(n43779), .B(n46573), .Z(n50945) );
  XNOR U50347 ( .A(n50946), .B(n49554), .Z(n46573) );
  ANDN U50348 ( .B(n47726), .A(n47727), .Z(n50946) );
  XOR U50349 ( .A(round_reg[1160]), .B(n50947), .Z(n47726) );
  XNOR U50350 ( .A(n50948), .B(n49617), .Z(n43779) );
  ANDN U50351 ( .B(n47732), .A(n47734), .Z(n50948) );
  XNOR U50352 ( .A(round_reg[1085]), .B(n50949), .Z(n47732) );
  XOR U50353 ( .A(n47411), .B(n50950), .Z(n50944) );
  XOR U50354 ( .A(n42859), .B(n48467), .Z(n50950) );
  XNOR U50355 ( .A(n50951), .B(n49557), .Z(n48467) );
  ANDN U50356 ( .B(n49558), .A(n50952), .Z(n50951) );
  XNOR U50357 ( .A(n50953), .B(n50352), .Z(n42859) );
  XOR U50358 ( .A(round_reg[1134]), .B(n50394), .Z(n47736) );
  XNOR U50359 ( .A(n50954), .B(n49549), .Z(n47411) );
  NOR U50360 ( .A(n49135), .B(n49133), .Z(n50954) );
  XOR U50361 ( .A(round_reg[1232]), .B(n50955), .Z(n49133) );
  XOR U50362 ( .A(n50956), .B(n49558), .Z(n47724) );
  XNOR U50363 ( .A(round_reg[992]), .B(n50957), .Z(n49558) );
  AND U50364 ( .A(n50958), .B(n50952), .Z(n50956) );
  ANDN U50365 ( .B(n41610), .A(n49230), .Z(n50929) );
  XNOR U50366 ( .A(n50959), .B(n47632), .Z(n49230) );
  IV U50367 ( .A(n45814), .Z(n47632) );
  XOR U50368 ( .A(n50960), .B(n43472), .Z(n41610) );
  XNOR U50369 ( .A(n50348), .B(n50961), .Z(n43472) );
  XOR U50370 ( .A(n50962), .B(n50963), .Z(n50348) );
  XOR U50371 ( .A(n42165), .B(n47147), .Z(n50963) );
  XNOR U50372 ( .A(n50964), .B(n47728), .Z(n47147) );
  ANDN U50373 ( .B(n49553), .A(n49554), .Z(n50964) );
  XOR U50374 ( .A(round_reg[1588]), .B(n50299), .Z(n49554) );
  XOR U50375 ( .A(n50965), .B(n47737), .Z(n42165) );
  ANDN U50376 ( .B(n50351), .A(n50352), .Z(n50965) );
  XNOR U50377 ( .A(round_reg[1523]), .B(n50966), .Z(n50352) );
  XNOR U50378 ( .A(n45431), .B(n50967), .Z(n50962) );
  XOR U50379 ( .A(n46222), .B(n45393), .Z(n50967) );
  XNOR U50380 ( .A(n50968), .B(n47733), .Z(n45393) );
  ANDN U50381 ( .B(n49617), .A(n50969), .Z(n50968) );
  XNOR U50382 ( .A(round_reg[1462]), .B(n49795), .Z(n49617) );
  XNOR U50383 ( .A(n50970), .B(n49134), .Z(n46222) );
  NOR U50384 ( .A(n49548), .B(n49549), .Z(n50970) );
  XNOR U50385 ( .A(round_reg[1305]), .B(n50971), .Z(n49549) );
  XNOR U50386 ( .A(n50972), .B(n50958), .Z(n45431) );
  NOR U50387 ( .A(n49557), .B(n49556), .Z(n50972) );
  XNOR U50388 ( .A(round_reg[1368]), .B(n48441), .Z(n49557) );
  XOR U50389 ( .A(n50973), .B(n50974), .Z(n43685) );
  XNOR U50390 ( .A(n40508), .B(n38933), .Z(n50974) );
  XNOR U50391 ( .A(n50975), .B(n45225), .Z(n38933) );
  XOR U50392 ( .A(n41598), .B(n50561), .Z(n45225) );
  XNOR U50393 ( .A(n50976), .B(n50977), .Z(n50561) );
  ANDN U50394 ( .B(n50769), .A(n48458), .Z(n50976) );
  XNOR U50395 ( .A(round_reg[88]), .B(n48441), .Z(n48458) );
  IV U50396 ( .A(n50978), .Z(n48441) );
  IV U50397 ( .A(n44555), .Z(n41598) );
  XNOR U50398 ( .A(n46690), .B(n50979), .Z(n44555) );
  XOR U50399 ( .A(n50980), .B(n50981), .Z(n46690) );
  XNOR U50400 ( .A(n42500), .B(n44518), .Z(n50981) );
  XOR U50401 ( .A(n50982), .B(n47794), .Z(n44518) );
  ANDN U50402 ( .B(n50564), .A(n50565), .Z(n50982) );
  XOR U50403 ( .A(round_reg[547]), .B(n48450), .Z(n50565) );
  XOR U50404 ( .A(n50983), .B(n47790), .Z(n42500) );
  ANDN U50405 ( .B(n50556), .A(n50557), .Z(n50983) );
  XNOR U50406 ( .A(round_reg[443]), .B(n50984), .Z(n50557) );
  XNOR U50407 ( .A(n45947), .B(n50985), .Z(n50980) );
  XNOR U50408 ( .A(n46953), .B(n43347), .Z(n50985) );
  XNOR U50409 ( .A(n50986), .B(n48459), .Z(n43347) );
  ANDN U50410 ( .B(n50977), .A(n50769), .Z(n50986) );
  XNOR U50411 ( .A(round_reg[449]), .B(n50127), .Z(n50769) );
  XOR U50412 ( .A(n50987), .B(n47805), .Z(n46953) );
  ANDN U50413 ( .B(n50567), .A(n50568), .Z(n50987) );
  XNOR U50414 ( .A(round_reg[615]), .B(n50988), .Z(n50568) );
  XOR U50415 ( .A(n50989), .B(n47801), .Z(n45947) );
  ANDN U50416 ( .B(n50559), .A(n50560), .Z(n50989) );
  XNOR U50417 ( .A(round_reg[328]), .B(n48699), .Z(n50560) );
  ANDN U50418 ( .B(n43154), .A(n43155), .Z(n50975) );
  XOR U50419 ( .A(n46043), .B(n44619), .Z(n43155) );
  XOR U50420 ( .A(n49785), .B(n46412), .Z(n44619) );
  XNOR U50421 ( .A(n50990), .B(n50991), .Z(n46412) );
  XNOR U50422 ( .A(n47642), .B(n44460), .Z(n50991) );
  XNOR U50423 ( .A(n50992), .B(n49297), .Z(n44460) );
  XOR U50424 ( .A(round_reg[1383]), .B(n50224), .Z(n49297) );
  NOR U50425 ( .A(n49933), .B(n49296), .Z(n50992) );
  XOR U50426 ( .A(round_reg[1007]), .B(n49086), .Z(n49296) );
  XNOR U50427 ( .A(n49301), .B(n50993), .Z(n47642) );
  XNOR U50428 ( .A(n4687), .B(n50994), .Z(n50993) );
  OR U50429 ( .A(n49930), .B(n49302), .Z(n50994) );
  XOR U50430 ( .A(round_reg[1175]), .B(n50995), .Z(n49302) );
  IV U50431 ( .A(rc_i[1]), .Z(n4687) );
  XOR U50432 ( .A(n44916), .B(n50996), .Z(n50990) );
  XNOR U50433 ( .A(n44846), .B(n46149), .Z(n50996) );
  XNOR U50434 ( .A(n50997), .B(n49293), .Z(n46149) );
  XOR U50435 ( .A(round_reg[1413]), .B(n50998), .Z(n49293) );
  NOR U50436 ( .A(n49938), .B(n49292), .Z(n50997) );
  XOR U50437 ( .A(round_reg[1036]), .B(n50999), .Z(n49292) );
  XNOR U50438 ( .A(n51000), .B(n49306), .Z(n44846) );
  XOR U50439 ( .A(round_reg[1474]), .B(n51001), .Z(n49306) );
  XOR U50440 ( .A(round_reg[1149]), .B(n49992), .Z(n49305) );
  XNOR U50441 ( .A(n51002), .B(n49850), .Z(n44916) );
  IV U50442 ( .A(n49309), .Z(n49850) );
  XOR U50443 ( .A(round_reg[1320]), .B(n48442), .Z(n49309) );
  ANDN U50444 ( .B(n49310), .A(n49936), .Z(n51002) );
  XNOR U50445 ( .A(round_reg[1247]), .B(n50453), .Z(n49310) );
  XOR U50446 ( .A(n51003), .B(n51004), .Z(n49785) );
  XNOR U50447 ( .A(n43964), .B(n46258), .Z(n51004) );
  XOR U50448 ( .A(n51005), .B(n49324), .Z(n46258) );
  XNOR U50449 ( .A(round_reg[501]), .B(n50744), .Z(n49324) );
  ANDN U50450 ( .B(n46046), .A(n46047), .Z(n51005) );
  XOR U50451 ( .A(round_reg[1321]), .B(n51006), .Z(n46047) );
  XOR U50452 ( .A(round_reg[76]), .B(n51007), .Z(n46046) );
  XNOR U50453 ( .A(n51008), .B(n49864), .Z(n43964) );
  XOR U50454 ( .A(round_reg[603]), .B(n51009), .Z(n49864) );
  XNOR U50455 ( .A(round_reg[1414]), .B(n50759), .Z(n47019) );
  XOR U50456 ( .A(round_reg[194]), .B(n51010), .Z(n47018) );
  XOR U50457 ( .A(n49287), .B(n51011), .Z(n51003) );
  XOR U50458 ( .A(n44565), .B(n48907), .Z(n51011) );
  XNOR U50459 ( .A(n51012), .B(n49317), .Z(n48907) );
  XNOR U50460 ( .A(round_reg[380]), .B(n51013), .Z(n49317) );
  XNOR U50461 ( .A(round_reg[1475]), .B(n49958), .Z(n46051) );
  XOR U50462 ( .A(round_reg[306]), .B(n51014), .Z(n46050) );
  XNOR U50463 ( .A(n51015), .B(n49321), .Z(n44565) );
  XNOR U50464 ( .A(round_reg[535]), .B(n50995), .Z(n49321) );
  XNOR U50465 ( .A(round_reg[1384]), .B(n51016), .Z(n48498) );
  XOR U50466 ( .A(round_reg[135]), .B(n51017), .Z(n48497) );
  XNOR U50467 ( .A(n51018), .B(n49314), .Z(n49287) );
  XNOR U50468 ( .A(round_reg[431]), .B(n50456), .Z(n49314) );
  ANDN U50469 ( .B(n49315), .A(n49203), .Z(n51018) );
  XNOR U50470 ( .A(n51019), .B(n49315), .Z(n46043) );
  XOR U50471 ( .A(round_reg[54]), .B(n51020), .Z(n49315) );
  ANDN U50472 ( .B(n49203), .A(n49205), .Z(n51019) );
  XOR U50473 ( .A(round_reg[1176]), .B(n49789), .Z(n49205) );
  XOR U50474 ( .A(round_reg[1540]), .B(n49612), .Z(n49203) );
  XOR U50475 ( .A(n44520), .B(n51021), .Z(n43154) );
  XOR U50476 ( .A(n47321), .B(n51022), .Z(n44520) );
  XOR U50477 ( .A(n51023), .B(n51024), .Z(n47321) );
  XOR U50478 ( .A(n46999), .B(n45821), .Z(n51024) );
  XNOR U50479 ( .A(n51025), .B(n47562), .Z(n45821) );
  XOR U50480 ( .A(round_reg[640]), .B(n51026), .Z(n47562) );
  NOR U50481 ( .A(n49177), .B(n47936), .Z(n51025) );
  XNOR U50482 ( .A(n51027), .B(n47565), .Z(n46999) );
  XOR U50483 ( .A(round_reg[718]), .B(n48957), .Z(n47565) );
  ANDN U50484 ( .B(n47938), .A(n49174), .Z(n51027) );
  XOR U50485 ( .A(n44033), .B(n51028), .Z(n51023) );
  XOR U50486 ( .A(n46657), .B(n47457), .Z(n51028) );
  XNOR U50487 ( .A(n51029), .B(n47553), .Z(n47457) );
  XOR U50488 ( .A(round_reg[828]), .B(n51030), .Z(n47553) );
  ANDN U50489 ( .B(n47941), .A(n49169), .Z(n51029) );
  XNOR U50490 ( .A(n51031), .B(n47558), .Z(n46657) );
  ANDN U50491 ( .B(n47943), .A(n49171), .Z(n51031) );
  XNOR U50492 ( .A(n51033), .B(n47947), .Z(n44033) );
  XOR U50493 ( .A(round_reg[932]), .B(n50447), .Z(n47947) );
  ANDN U50494 ( .B(n47946), .A(n49180), .Z(n51033) );
  XOR U50495 ( .A(n51034), .B(n42086), .Z(n40508) );
  XNOR U50496 ( .A(n51035), .B(n46282), .Z(n42086) );
  IV U50497 ( .A(n46506), .Z(n46282) );
  ANDN U50498 ( .B(n43150), .A(n42085), .Z(n51034) );
  XNOR U50499 ( .A(n49420), .B(n49154), .Z(n42085) );
  XNOR U50500 ( .A(n51036), .B(n50908), .Z(n49154) );
  NOR U50501 ( .A(n50622), .B(n51037), .Z(n51036) );
  XOR U50502 ( .A(n48417), .B(n44800), .Z(n43150) );
  IV U50503 ( .A(n44467), .Z(n44800) );
  XNOR U50504 ( .A(n48038), .B(n46578), .Z(n44467) );
  XOR U50505 ( .A(n51038), .B(n51039), .Z(n46578) );
  XNOR U50506 ( .A(n46000), .B(n43666), .Z(n51039) );
  XNOR U50507 ( .A(n51040), .B(n47834), .Z(n43666) );
  ANDN U50508 ( .B(n47833), .A(n47926), .Z(n51040) );
  XOR U50509 ( .A(round_reg[1285]), .B(n51041), .Z(n47926) );
  XOR U50510 ( .A(round_reg[104]), .B(n51042), .Z(n47833) );
  XNOR U50511 ( .A(n51043), .B(n51044), .Z(n46000) );
  ANDN U50512 ( .B(n49254), .A(n47914), .Z(n51043) );
  XOR U50513 ( .A(round_reg[1348]), .B(n50741), .Z(n47914) );
  XOR U50514 ( .A(n43952), .B(n51045), .Z(n51038) );
  XNOR U50515 ( .A(n45093), .B(n47816), .Z(n51045) );
  XOR U50516 ( .A(n51046), .B(n48163), .Z(n47816) );
  AND U50517 ( .A(n47922), .B(n48164), .Z(n51046) );
  XNOR U50518 ( .A(round_reg[270]), .B(n51047), .Z(n48164) );
  XNOR U50519 ( .A(round_reg[1503]), .B(n51048), .Z(n47922) );
  XNOR U50520 ( .A(n51049), .B(n47824), .Z(n45093) );
  AND U50521 ( .A(n47919), .B(n47823), .Z(n51049) );
  XOR U50522 ( .A(round_reg[222]), .B(n51050), .Z(n47823) );
  XNOR U50523 ( .A(round_reg[1442]), .B(n51051), .Z(n47919) );
  XNOR U50524 ( .A(n51052), .B(n47830), .Z(n43952) );
  ANDN U50525 ( .B(n47829), .A(n49232), .Z(n51052) );
  XOR U50526 ( .A(round_reg[1568]), .B(n49860), .Z(n49232) );
  XNOR U50527 ( .A(round_reg[18]), .B(n51053), .Z(n47829) );
  XOR U50528 ( .A(n51054), .B(n51055), .Z(n48038) );
  XNOR U50529 ( .A(n44790), .B(n45445), .Z(n51055) );
  XOR U50530 ( .A(n51056), .B(n51057), .Z(n45445) );
  ANDN U50531 ( .B(n48410), .A(n48411), .Z(n51056) );
  XOR U50532 ( .A(n51058), .B(n51059), .Z(n44790) );
  AND U50533 ( .A(n48426), .B(n48424), .Z(n51058) );
  XNOR U50534 ( .A(n46827), .B(n51060), .Z(n51054) );
  XOR U50535 ( .A(n45142), .B(n43596), .Z(n51060) );
  XOR U50536 ( .A(n51061), .B(n51062), .Z(n43596) );
  ANDN U50537 ( .B(n51063), .A(n51064), .Z(n51061) );
  XOR U50538 ( .A(n51065), .B(n51066), .Z(n45142) );
  ANDN U50539 ( .B(n48420), .A(n51067), .Z(n51065) );
  XOR U50540 ( .A(n51068), .B(n51069), .Z(n46827) );
  ANDN U50541 ( .B(n48414), .A(n48415), .Z(n51068) );
  XNOR U50542 ( .A(n51070), .B(n51063), .Z(n48417) );
  ANDN U50543 ( .B(n51064), .A(n51071), .Z(n51070) );
  XOR U50544 ( .A(n40536), .B(n51072), .Z(n50973) );
  XOR U50545 ( .A(n42079), .B(n39237), .Z(n51072) );
  XNOR U50546 ( .A(n51073), .B(n42099), .Z(n39237) );
  XOR U50547 ( .A(n45145), .B(n51074), .Z(n42099) );
  AND U50548 ( .A(n43147), .B(n42100), .Z(n51073) );
  XOR U50549 ( .A(n51075), .B(n45397), .Z(n42100) );
  XOR U50550 ( .A(n46954), .B(n49091), .Z(n45397) );
  XNOR U50551 ( .A(n51076), .B(n51077), .Z(n49091) );
  XOR U50552 ( .A(n42405), .B(n47524), .Z(n51077) );
  XNOR U50553 ( .A(n51078), .B(n50783), .Z(n47524) );
  NOR U50554 ( .A(n50782), .B(n51079), .Z(n51078) );
  XOR U50555 ( .A(n51080), .B(n50251), .Z(n42405) );
  AND U50556 ( .A(n51081), .B(n50250), .Z(n51080) );
  XNOR U50557 ( .A(n45253), .B(n51082), .Z(n51076) );
  XOR U50558 ( .A(n46216), .B(n46204), .Z(n51082) );
  XNOR U50559 ( .A(n51083), .B(n50265), .Z(n46204) );
  NOR U50560 ( .A(n51084), .B(n50264), .Z(n51083) );
  XOR U50561 ( .A(n51085), .B(n50255), .Z(n46216) );
  NOR U50562 ( .A(n50254), .B(n51086), .Z(n51085) );
  XNOR U50563 ( .A(n51087), .B(n50260), .Z(n45253) );
  ANDN U50564 ( .B(n50261), .A(n51088), .Z(n51087) );
  XOR U50565 ( .A(n51089), .B(n51090), .Z(n46954) );
  XNOR U50566 ( .A(n46645), .B(n46923), .Z(n51090) );
  XOR U50567 ( .A(n51091), .B(n47800), .Z(n46923) );
  XNOR U50568 ( .A(round_reg[1487]), .B(n50401), .Z(n47800) );
  ANDN U50569 ( .B(n47801), .A(n50559), .Z(n51091) );
  XNOR U50570 ( .A(round_reg[759]), .B(n50483), .Z(n50559) );
  XOR U50571 ( .A(round_reg[1098]), .B(n50117), .Z(n47801) );
  XOR U50572 ( .A(n51092), .B(n47795), .Z(n46645) );
  XNOR U50573 ( .A(round_reg[1396]), .B(n49623), .Z(n47795) );
  ANDN U50574 ( .B(n47794), .A(n50564), .Z(n51092) );
  XOR U50575 ( .A(round_reg[909]), .B(n51093), .Z(n50564) );
  XOR U50576 ( .A(round_reg[1020]), .B(n51094), .Z(n47794) );
  XOR U50577 ( .A(n47159), .B(n51095), .Z(n51089) );
  XOR U50578 ( .A(n43597), .B(n47784), .Z(n51095) );
  XOR U50579 ( .A(n51096), .B(n48460), .Z(n47784) );
  XNOR U50580 ( .A(round_reg[1333]), .B(n51097), .Z(n48460) );
  ANDN U50581 ( .B(n48459), .A(n50977), .Z(n51096) );
  XNOR U50582 ( .A(round_reg[838]), .B(n50116), .Z(n50977) );
  XOR U50583 ( .A(round_reg[1260]), .B(n51098), .Z(n48459) );
  XNOR U50584 ( .A(n51099), .B(n50771), .Z(n43597) );
  IV U50585 ( .A(n47804), .Z(n50771) );
  XNOR U50586 ( .A(round_reg[1426]), .B(n51100), .Z(n47804) );
  ANDN U50587 ( .B(n47805), .A(n50567), .Z(n51099) );
  XOR U50588 ( .A(round_reg[681]), .B(n51006), .Z(n50567) );
  XOR U50589 ( .A(round_reg[1049]), .B(n51101), .Z(n47805) );
  XOR U50590 ( .A(n51102), .B(n47791), .Z(n47159) );
  XNOR U50591 ( .A(round_reg[1552]), .B(n51103), .Z(n47791) );
  ANDN U50592 ( .B(n47790), .A(n50556), .Z(n51102) );
  XNOR U50593 ( .A(round_reg[805]), .B(n48566), .Z(n50556) );
  XOR U50594 ( .A(round_reg[1188]), .B(n51104), .Z(n47790) );
  XOR U50595 ( .A(n42668), .B(n49258), .Z(n43147) );
  XNOR U50596 ( .A(n51105), .B(n51106), .Z(n49258) );
  XNOR U50597 ( .A(round_reg[820]), .B(n51107), .Z(n48861) );
  XNOR U50598 ( .A(n47817), .B(n50615), .Z(n42668) );
  XOR U50599 ( .A(n51108), .B(n51109), .Z(n50615) );
  XNOR U50600 ( .A(n43903), .B(n49227), .Z(n51109) );
  XNOR U50601 ( .A(n51110), .B(n49142), .Z(n49227) );
  ANDN U50602 ( .B(n48840), .A(n50634), .Z(n51110) );
  IV U50603 ( .A(n51111), .Z(n50634) );
  XOR U50604 ( .A(round_reg[629]), .B(n50842), .Z(n48840) );
  XNOR U50605 ( .A(n51112), .B(n49146), .Z(n43903) );
  ANDN U50606 ( .B(n48857), .A(n51113), .Z(n51112) );
  XOR U50607 ( .A(round_reg[342]), .B(n48945), .Z(n48857) );
  XOR U50608 ( .A(n45852), .B(n51114), .Z(n51108) );
  XOR U50609 ( .A(n51115), .B(n48220), .Z(n51114) );
  XNOR U50610 ( .A(n51116), .B(n49148), .Z(n48220) );
  ANDN U50611 ( .B(n48844), .A(n51117), .Z(n51116) );
  XOR U50612 ( .A(round_reg[463]), .B(n50859), .Z(n48844) );
  XNOR U50613 ( .A(n51118), .B(n49150), .Z(n45852) );
  NOR U50614 ( .A(n48853), .B(n49282), .Z(n51118) );
  XOR U50615 ( .A(round_reg[561]), .B(n50739), .Z(n48853) );
  XNOR U50616 ( .A(n51119), .B(n51120), .Z(n47817) );
  XNOR U50617 ( .A(n45662), .B(n47779), .Z(n51120) );
  XNOR U50618 ( .A(n51121), .B(n48863), .Z(n47779) );
  IV U50619 ( .A(n51122), .Z(n48863) );
  ANDN U50620 ( .B(n51106), .A(n49284), .Z(n51121) );
  XNOR U50621 ( .A(round_reg[1203]), .B(n50966), .Z(n49284) );
  XNOR U50622 ( .A(n51123), .B(n48689), .Z(n45662) );
  ANDN U50623 ( .B(n49264), .A(n49237), .Z(n51123) );
  XOR U50624 ( .A(round_reg[1064]), .B(n51042), .Z(n49237) );
  XOR U50625 ( .A(n44858), .B(n51124), .Z(n51119) );
  XOR U50626 ( .A(n51125), .B(n46589), .Z(n51124) );
  XNOR U50627 ( .A(n51126), .B(n48303), .Z(n46589) );
  NOR U50628 ( .A(n49260), .B(n49243), .Z(n51126) );
  XNOR U50629 ( .A(round_reg[971]), .B(n51127), .Z(n49243) );
  IV U50630 ( .A(n51128), .Z(n49260) );
  XOR U50631 ( .A(n51129), .B(n48293), .Z(n44858) );
  AND U50632 ( .A(n49239), .B(n49270), .Z(n51129) );
  XOR U50633 ( .A(round_reg[1113]), .B(n49854), .Z(n49239) );
  XNOR U50634 ( .A(n51130), .B(n42089), .Z(n42079) );
  XOR U50635 ( .A(n48323), .B(n44201), .Z(n42089) );
  XOR U50636 ( .A(n51131), .B(n50763), .Z(n44201) );
  XNOR U50637 ( .A(n51132), .B(n51133), .Z(n50763) );
  XNOR U50638 ( .A(n47741), .B(n46034), .Z(n51133) );
  XNOR U50639 ( .A(n51134), .B(n47761), .Z(n46034) );
  XOR U50640 ( .A(round_reg[1558]), .B(n50397), .Z(n47761) );
  NOR U50641 ( .A(n47760), .B(n49128), .Z(n51134) );
  XOR U50642 ( .A(round_reg[811]), .B(n51135), .Z(n49128) );
  XNOR U50643 ( .A(round_reg[1194]), .B(n48564), .Z(n47760) );
  XNOR U50644 ( .A(n51136), .B(n47777), .Z(n47741) );
  XOR U50645 ( .A(round_reg[1402]), .B(n51137), .Z(n47777) );
  ANDN U50646 ( .B(n47778), .A(n50147), .Z(n51136) );
  XOR U50647 ( .A(round_reg[915]), .B(n50480), .Z(n50147) );
  XOR U50648 ( .A(round_reg[962]), .B(n50775), .Z(n47778) );
  XOR U50649 ( .A(n45746), .B(n51138), .Z(n51132) );
  XOR U50650 ( .A(n46246), .B(n43084), .Z(n51138) );
  XNOR U50651 ( .A(n51139), .B(n47773), .Z(n43084) );
  XOR U50652 ( .A(round_reg[1339]), .B(n48455), .Z(n47773) );
  XNOR U50653 ( .A(round_reg[844]), .B(n51140), .Z(n49125) );
  XOR U50654 ( .A(round_reg[1266]), .B(n51014), .Z(n47774) );
  IV U50655 ( .A(n51141), .Z(n51014) );
  XNOR U50656 ( .A(n51142), .B(n47769), .Z(n46246) );
  XNOR U50657 ( .A(round_reg[1493]), .B(n50430), .Z(n47769) );
  XNOR U50658 ( .A(round_reg[765]), .B(n50949), .Z(n49120) );
  XOR U50659 ( .A(round_reg[1104]), .B(n51143), .Z(n47770) );
  XNOR U50660 ( .A(n51144), .B(n47765), .Z(n45746) );
  XNOR U50661 ( .A(round_reg[1432]), .B(n51145), .Z(n47765) );
  NOR U50662 ( .A(n47764), .B(n49117), .Z(n51144) );
  XNOR U50663 ( .A(round_reg[687]), .B(n49086), .Z(n49117) );
  IV U50664 ( .A(n51146), .Z(n49086) );
  XOR U50665 ( .A(round_reg[1055]), .B(n51147), .Z(n47764) );
  XNOR U50666 ( .A(n51148), .B(n47533), .Z(n48323) );
  ANDN U50667 ( .B(n51149), .A(n50613), .Z(n51148) );
  ANDN U50668 ( .B(n42090), .A(n43159), .Z(n51130) );
  XOR U50669 ( .A(n51115), .B(n45853), .Z(n43159) );
  IV U50670 ( .A(n43904), .Z(n45853) );
  XOR U50671 ( .A(n51150), .B(n51151), .Z(n43904) );
  XNOR U50672 ( .A(n51152), .B(n49140), .Z(n51115) );
  XOR U50673 ( .A(round_reg[393]), .B(n50227), .Z(n48849) );
  XOR U50674 ( .A(n48645), .B(n46886), .Z(n42090) );
  XOR U50675 ( .A(n51153), .B(n50589), .Z(n46886) );
  XOR U50676 ( .A(n51154), .B(n51155), .Z(n50589) );
  XNOR U50677 ( .A(n45703), .B(n44758), .Z(n51155) );
  XNOR U50678 ( .A(n51156), .B(n50548), .Z(n44758) );
  IV U50679 ( .A(n47896), .Z(n50548) );
  XOR U50680 ( .A(round_reg[1045]), .B(n48948), .Z(n47896) );
  ANDN U50681 ( .B(n49038), .A(n49037), .Z(n51156) );
  XOR U50682 ( .A(round_reg[677]), .B(n50646), .Z(n49037) );
  IV U50683 ( .A(n50851), .Z(n49038) );
  XOR U50684 ( .A(round_reg[611]), .B(n48872), .Z(n50851) );
  XOR U50685 ( .A(n51157), .B(n47902), .Z(n45703) );
  IV U50686 ( .A(n50550), .Z(n47902) );
  XOR U50687 ( .A(round_reg[1094]), .B(n50759), .Z(n50550) );
  ANDN U50688 ( .B(n49041), .A(n49040), .Z(n51157) );
  XOR U50689 ( .A(round_reg[755]), .B(n50444), .Z(n49040) );
  XNOR U50690 ( .A(round_reg[324]), .B(n51158), .Z(n49041) );
  XNOR U50691 ( .A(n46734), .B(n51159), .Z(n51154) );
  XNOR U50692 ( .A(n47837), .B(n46890), .Z(n51159) );
  XOR U50693 ( .A(n51160), .B(n47893), .Z(n46890) );
  IV U50694 ( .A(n50542), .Z(n47893) );
  XOR U50695 ( .A(round_reg[1184]), .B(n51161), .Z(n50542) );
  AND U50696 ( .A(n49468), .B(n49466), .Z(n51160) );
  XNOR U50697 ( .A(round_reg[801]), .B(n49175), .Z(n49466) );
  XOR U50698 ( .A(round_reg[439]), .B(n50483), .Z(n49468) );
  XNOR U50699 ( .A(n51162), .B(n47906), .Z(n47837) );
  IV U50700 ( .A(n50546), .Z(n47906) );
  XOR U50701 ( .A(round_reg[1256]), .B(n49984), .Z(n50546) );
  ANDN U50702 ( .B(n50586), .A(n50545), .Z(n51162) );
  XNOR U50703 ( .A(round_reg[834]), .B(n51010), .Z(n50545) );
  XNOR U50704 ( .A(round_reg[509]), .B(n49992), .Z(n50586) );
  XOR U50705 ( .A(n51163), .B(n50845), .Z(n46734) );
  IV U50706 ( .A(n50540), .Z(n50845) );
  XOR U50707 ( .A(round_reg[1016]), .B(n50486), .Z(n50540) );
  ANDN U50708 ( .B(n49033), .A(n49031), .Z(n51163) );
  XOR U50709 ( .A(round_reg[905]), .B(n51164), .Z(n49031) );
  XNOR U50710 ( .A(round_reg[543]), .B(n51048), .Z(n49033) );
  XOR U50711 ( .A(n51165), .B(n50530), .Z(n48645) );
  ANDN U50712 ( .B(n49538), .A(n51166), .Z(n51165) );
  XNOR U50713 ( .A(n51167), .B(n42096), .Z(n40536) );
  XOR U50714 ( .A(n51168), .B(n43540), .Z(n42096) );
  IV U50715 ( .A(n47388), .Z(n43540) );
  XNOR U50716 ( .A(n51169), .B(n51170), .Z(n46914) );
  XNOR U50717 ( .A(n50344), .B(n42457), .Z(n51170) );
  XOR U50718 ( .A(n51171), .B(n48924), .Z(n42457) );
  ANDN U50719 ( .B(n48941), .A(n48099), .Z(n51171) );
  XOR U50720 ( .A(round_reg[239]), .B(n51172), .Z(n48099) );
  XOR U50721 ( .A(n51173), .B(n48926), .Z(n50344) );
  XNOR U50722 ( .A(n45512), .B(n51174), .Z(n51169) );
  XOR U50723 ( .A(n51175), .B(n45316), .Z(n51174) );
  XNOR U50724 ( .A(n51176), .B(n48922), .Z(n45316) );
  ANDN U50725 ( .B(n48944), .A(n48090), .Z(n51176) );
  XOR U50726 ( .A(round_reg[121]), .B(n51177), .Z(n48090) );
  XNOR U50727 ( .A(n51178), .B(n48919), .Z(n45512) );
  NOR U50728 ( .A(n48934), .B(n48095), .Z(n51178) );
  XOR U50729 ( .A(round_reg[35]), .B(n51179), .Z(n48095) );
  XOR U50730 ( .A(n51180), .B(n51181), .Z(n50000) );
  XOR U50731 ( .A(n46105), .B(n44118), .Z(n51181) );
  XOR U50732 ( .A(n51182), .B(n49750), .Z(n44118) );
  XNOR U50733 ( .A(round_reg[1366]), .B(n51183), .Z(n49750) );
  ANDN U50734 ( .B(n50367), .A(n50885), .Z(n51182) );
  XNOR U50735 ( .A(n51184), .B(n49742), .Z(n46105) );
  XNOR U50736 ( .A(round_reg[1460]), .B(n51185), .Z(n49742) );
  NOR U50737 ( .A(n50878), .B(n50365), .Z(n51184) );
  XOR U50738 ( .A(n50353), .B(n51186), .Z(n51180) );
  XOR U50739 ( .A(n46669), .B(n47261), .Z(n51186) );
  XNOR U50740 ( .A(n51187), .B(n49733), .Z(n47261) );
  XNOR U50741 ( .A(round_reg[1586]), .B(n51141), .Z(n49733) );
  ANDN U50742 ( .B(n50363), .A(n50887), .Z(n51187) );
  XNOR U50743 ( .A(n51188), .B(n49737), .Z(n46669) );
  XOR U50744 ( .A(round_reg[1521]), .B(n50739), .Z(n49737) );
  ANDN U50745 ( .B(n50890), .A(n50360), .Z(n51188) );
  XNOR U50746 ( .A(n51189), .B(n49746), .Z(n50353) );
  XOR U50747 ( .A(round_reg[1303]), .B(n48554), .Z(n49746) );
  NOR U50748 ( .A(n50881), .B(n50358), .Z(n51189) );
  ANDN U50749 ( .B(n42095), .A(n43701), .Z(n51167) );
  XOR U50750 ( .A(n47678), .B(n49843), .Z(n43701) );
  XNOR U50751 ( .A(n51190), .B(n49931), .Z(n49843) );
  ANDN U50752 ( .B(n49301), .A(n49300), .Z(n51190) );
  XNOR U50753 ( .A(round_reg[1539]), .B(n48514), .Z(n49301) );
  IV U50754 ( .A(n44504), .Z(n47678) );
  XOR U50755 ( .A(n51191), .B(n47244), .Z(n44504) );
  XNOR U50756 ( .A(n51192), .B(n51193), .Z(n47244) );
  XOR U50757 ( .A(n45631), .B(n49913), .Z(n51193) );
  XNOR U50758 ( .A(n51194), .B(n49930), .Z(n49913) );
  XNOR U50759 ( .A(round_reg[792]), .B(n51145), .Z(n49930) );
  ANDN U50760 ( .B(n49300), .A(n49931), .Z(n51194) );
  XOR U50761 ( .A(round_reg[430]), .B(n50831), .Z(n49931) );
  XOR U50762 ( .A(round_reg[53]), .B(n51195), .Z(n49300) );
  XNOR U50763 ( .A(n51196), .B(n49941), .Z(n45631) );
  XOR U50764 ( .A(round_reg[746]), .B(n50819), .Z(n49941) );
  NOR U50765 ( .A(n49304), .B(n49940), .Z(n51196) );
  XNOR U50766 ( .A(round_reg[379]), .B(n48455), .Z(n49940) );
  XOR U50767 ( .A(round_reg[305]), .B(n48935), .Z(n49304) );
  XOR U50768 ( .A(n47024), .B(n51197), .Z(n51192) );
  XOR U50769 ( .A(n45319), .B(n49413), .Z(n51197) );
  XNOR U50770 ( .A(n51198), .B(n49933), .Z(n49413) );
  XOR U50771 ( .A(round_reg[896]), .B(n51199), .Z(n49933) );
  NOR U50772 ( .A(n49295), .B(n49842), .Z(n51198) );
  XNOR U50773 ( .A(round_reg[534]), .B(n51200), .Z(n49842) );
  XOR U50774 ( .A(round_reg[134]), .B(n51201), .Z(n49295) );
  XNOR U50775 ( .A(n51202), .B(n49938), .Z(n45319) );
  XOR U50776 ( .A(round_reg[668]), .B(n48965), .Z(n49938) );
  ANDN U50777 ( .B(n49846), .A(n49291), .Z(n51202) );
  IV U50778 ( .A(n49847), .Z(n49291) );
  XOR U50779 ( .A(round_reg[193]), .B(n51203), .Z(n49847) );
  XNOR U50780 ( .A(round_reg[602]), .B(n49625), .Z(n49846) );
  XNOR U50781 ( .A(n51204), .B(n49936), .Z(n47024) );
  XOR U50782 ( .A(round_reg[889]), .B(n49836), .Z(n49936) );
  NOR U50783 ( .A(n49308), .B(n49849), .Z(n51204) );
  XOR U50784 ( .A(round_reg[500]), .B(n51185), .Z(n49849) );
  XNOR U50785 ( .A(round_reg[75]), .B(n51205), .Z(n49308) );
  XNOR U50786 ( .A(n51206), .B(n42163), .Z(n42095) );
  XNOR U50787 ( .A(n46672), .B(n47537), .Z(n42163) );
  XNOR U50788 ( .A(n51207), .B(n51208), .Z(n47537) );
  XNOR U50789 ( .A(n46797), .B(n44908), .Z(n51208) );
  XOR U50790 ( .A(n51209), .B(n47182), .Z(n44908) );
  XOR U50791 ( .A(round_reg[1116]), .B(n50827), .Z(n47182) );
  ANDN U50792 ( .B(n47183), .A(n51210), .Z(n51209) );
  XOR U50793 ( .A(n51211), .B(n47178), .Z(n46797) );
  ANDN U50794 ( .B(n47179), .A(n51212), .Z(n51211) );
  XNOR U50795 ( .A(n40857), .B(n51213), .Z(n51207) );
  XNOR U50796 ( .A(n45810), .B(n43931), .Z(n51213) );
  XNOR U50797 ( .A(n51214), .B(n47192), .Z(n43931) );
  XOR U50798 ( .A(round_reg[1206]), .B(n50234), .Z(n47192) );
  ANDN U50799 ( .B(n47193), .A(n51215), .Z(n51214) );
  XOR U50800 ( .A(n51216), .B(n47188), .Z(n45810) );
  XOR U50801 ( .A(round_reg[1067]), .B(n51217), .Z(n47188) );
  ANDN U50802 ( .B(n47189), .A(n51218), .Z(n51216) );
  XNOR U50803 ( .A(n51219), .B(n48037), .Z(n40857) );
  XOR U50804 ( .A(round_reg[1278]), .B(n50777), .Z(n48037) );
  NOR U50805 ( .A(n51220), .B(n48036), .Z(n51219) );
  XNOR U50806 ( .A(n51221), .B(n51222), .Z(n46672) );
  XNOR U50807 ( .A(n48405), .B(n45965), .Z(n51222) );
  XNOR U50808 ( .A(n51223), .B(n48421), .Z(n45965) );
  IV U50809 ( .A(n51067), .Z(n48421) );
  XOR U50810 ( .A(round_reg[632]), .B(n51224), .Z(n51067) );
  ANDN U50811 ( .B(n48422), .A(n51225), .Z(n51223) );
  XNOR U50812 ( .A(n51226), .B(n48426), .Z(n48405) );
  XNOR U50813 ( .A(round_reg[564]), .B(n51227), .Z(n48426) );
  ANDN U50814 ( .B(n48425), .A(n51228), .Z(n51226) );
  XNOR U50815 ( .A(n41750), .B(n51229), .Z(n51221) );
  XNOR U50816 ( .A(n46660), .B(n44580), .Z(n51229) );
  XNOR U50817 ( .A(n51230), .B(n48411), .Z(n44580) );
  XNOR U50818 ( .A(round_reg[345]), .B(n50971), .Z(n48411) );
  ANDN U50819 ( .B(n48412), .A(n51231), .Z(n51230) );
  XOR U50820 ( .A(n51232), .B(n48415), .Z(n46660) );
  XOR U50821 ( .A(round_reg[466]), .B(n51100), .Z(n48415) );
  ANDN U50822 ( .B(n48416), .A(n51233), .Z(n51232) );
  XOR U50823 ( .A(n51234), .B(n51064), .Z(n41750) );
  XOR U50824 ( .A(round_reg[396]), .B(n51007), .Z(n51064) );
  ANDN U50825 ( .B(n51071), .A(n51235), .Z(n51234) );
  NOR U50826 ( .A(n38841), .B(n35232), .Z(n50652) );
  XOR U50827 ( .A(n45572), .B(n39278), .Z(n35232) );
  XOR U50828 ( .A(n39417), .B(n42225), .Z(n39278) );
  XNOR U50829 ( .A(n51236), .B(n51237), .Z(n42225) );
  XNOR U50830 ( .A(n37920), .B(n39422), .Z(n51237) );
  XOR U50831 ( .A(n51238), .B(n41052), .Z(n39422) );
  XNOR U50832 ( .A(n51239), .B(n46506), .Z(n41052) );
  XOR U50833 ( .A(n50961), .B(n46921), .Z(n46506) );
  XNOR U50834 ( .A(n51240), .B(n51241), .Z(n46921) );
  XOR U50835 ( .A(n46083), .B(n44206), .Z(n51241) );
  XNOR U50836 ( .A(n51242), .B(n48140), .Z(n44206) );
  XOR U50837 ( .A(round_reg[126]), .B(n51243), .Z(n48140) );
  ANDN U50838 ( .B(n49339), .A(n51244), .Z(n51242) );
  XNOR U50839 ( .A(n51245), .B(n48130), .Z(n46083) );
  XOR U50840 ( .A(round_reg[244]), .B(n51246), .Z(n48130) );
  ANDN U50841 ( .B(n49336), .A(n51247), .Z(n51245) );
  XNOR U50842 ( .A(n42515), .B(n51248), .Z(n51240) );
  XOR U50843 ( .A(n49329), .B(n48864), .Z(n51248) );
  XOR U50844 ( .A(n51249), .B(n49068), .Z(n48864) );
  XOR U50845 ( .A(round_reg[292]), .B(n50447), .Z(n49068) );
  IV U50846 ( .A(n51250), .Z(n50447) );
  ANDN U50847 ( .B(n51251), .A(n49343), .Z(n51249) );
  XOR U50848 ( .A(n51252), .B(n48144), .Z(n49329) );
  XOR U50849 ( .A(round_reg[185]), .B(n51253), .Z(n48144) );
  AND U50850 ( .A(n51254), .B(n49334), .Z(n51252) );
  XOR U50851 ( .A(n51255), .B(n48136), .Z(n42515) );
  XNOR U50852 ( .A(round_reg[40]), .B(n48442), .Z(n48136) );
  ANDN U50853 ( .B(n49341), .A(n51256), .Z(n51255) );
  XNOR U50854 ( .A(n51257), .B(n51258), .Z(n50961) );
  XNOR U50855 ( .A(n51259), .B(n49025), .Z(n51258) );
  XNOR U50856 ( .A(n51260), .B(n51261), .Z(n49025) );
  ANDN U50857 ( .B(n51262), .A(n50187), .Z(n51260) );
  XOR U50858 ( .A(n43588), .B(n51263), .Z(n51257) );
  XNOR U50859 ( .A(n51264), .B(n44670), .Z(n51263) );
  XNOR U50860 ( .A(n51265), .B(n50182), .Z(n44670) );
  ANDN U50861 ( .B(n51266), .A(n50196), .Z(n51265) );
  XNOR U50862 ( .A(n51267), .B(n48151), .Z(n43588) );
  ANDN U50863 ( .B(n51268), .A(n50192), .Z(n51267) );
  ANDN U50864 ( .B(n41051), .A(n45196), .Z(n51238) );
  IV U50865 ( .A(n42008), .Z(n45196) );
  XOR U50866 ( .A(n51269), .B(n45973), .Z(n42008) );
  IV U50867 ( .A(n42504), .Z(n45973) );
  XOR U50868 ( .A(n47887), .B(n47476), .Z(n42504) );
  XOR U50869 ( .A(n51270), .B(n51271), .Z(n47476) );
  XOR U50870 ( .A(n49726), .B(n51074), .Z(n51271) );
  XNOR U50871 ( .A(n51272), .B(n51273), .Z(n51074) );
  ANDN U50872 ( .B(n51274), .A(n51275), .Z(n51272) );
  XNOR U50873 ( .A(n51276), .B(n47953), .Z(n49726) );
  XOR U50874 ( .A(n49912), .B(n51279), .Z(n51270) );
  XOR U50875 ( .A(n45144), .B(n51280), .Z(n51279) );
  XOR U50876 ( .A(n51281), .B(n46837), .Z(n45144) );
  ANDN U50877 ( .B(n51282), .A(n51283), .Z(n51281) );
  XNOR U50878 ( .A(n51284), .B(n51285), .Z(n49912) );
  ANDN U50879 ( .B(n51286), .A(n51287), .Z(n51284) );
  XOR U50880 ( .A(n51288), .B(n51289), .Z(n47887) );
  XNOR U50881 ( .A(n44979), .B(n46879), .Z(n51289) );
  XNOR U50882 ( .A(n51290), .B(n49058), .Z(n46879) );
  XNOR U50883 ( .A(round_reg[1044]), .B(n50849), .Z(n49058) );
  ANDN U50884 ( .B(n51291), .A(n50872), .Z(n51290) );
  XOR U50885 ( .A(n51292), .B(n49061), .Z(n44979) );
  XOR U50886 ( .A(round_reg[1093]), .B(n51293), .Z(n49061) );
  NOR U50887 ( .A(n51294), .B(n50874), .Z(n51292) );
  XOR U50888 ( .A(n48010), .B(n51295), .Z(n51288) );
  XNOR U50889 ( .A(n45582), .B(n46729), .Z(n51295) );
  XOR U50890 ( .A(n51296), .B(n49053), .Z(n46729) );
  XOR U50891 ( .A(round_reg[1255]), .B(n50988), .Z(n49053) );
  ANDN U50892 ( .B(n51297), .A(n50870), .Z(n51296) );
  XNOR U50893 ( .A(n51298), .B(n49048), .Z(n45582) );
  XNOR U50894 ( .A(round_reg[1015]), .B(n50507), .Z(n49048) );
  ANDN U50895 ( .B(n51299), .A(n51300), .Z(n51298) );
  XOR U50896 ( .A(n51301), .B(n50867), .Z(n48010) );
  ANDN U50897 ( .B(n50866), .A(n51302), .Z(n51301) );
  XOR U50898 ( .A(n46164), .B(n46841), .Z(n41051) );
  XNOR U50899 ( .A(n51303), .B(n51304), .Z(n46841) );
  ANDN U50900 ( .B(n51305), .A(n51285), .Z(n51303) );
  XOR U50901 ( .A(n51306), .B(n41056), .Z(n37920) );
  XOR U50902 ( .A(n44203), .B(n47710), .Z(n41056) );
  XNOR U50903 ( .A(n51307), .B(n50705), .Z(n47710) );
  AND U50904 ( .A(n50277), .B(n51308), .Z(n51307) );
  IV U50905 ( .A(n44869), .Z(n44203) );
  XOR U50906 ( .A(n48814), .B(n48193), .Z(n44869) );
  XNOR U50907 ( .A(n51309), .B(n51310), .Z(n48193) );
  XNOR U50908 ( .A(n46344), .B(n45641), .Z(n51310) );
  XNOR U50909 ( .A(n51311), .B(n50298), .Z(n45641) );
  IV U50910 ( .A(n49716), .Z(n50298) );
  XNOR U50911 ( .A(round_reg[522]), .B(n50852), .Z(n49716) );
  ANDN U50912 ( .B(n49717), .A(n47976), .Z(n51311) );
  XNOR U50913 ( .A(n51312), .B(n49710), .Z(n46344) );
  XOR U50914 ( .A(round_reg[590]), .B(n51313), .Z(n49710) );
  NOR U50915 ( .A(n49709), .B(n47987), .Z(n51312) );
  IV U50916 ( .A(n51314), .Z(n49709) );
  XOR U50917 ( .A(n42209), .B(n51315), .Z(n51309) );
  XOR U50918 ( .A(n46919), .B(n44603), .Z(n51315) );
  XNOR U50919 ( .A(n51316), .B(n49721), .Z(n44603) );
  XOR U50920 ( .A(round_reg[488]), .B(n51317), .Z(n49721) );
  ANDN U50921 ( .B(n49720), .A(n50692), .Z(n51316) );
  XNOR U50922 ( .A(n51318), .B(n49725), .Z(n46919) );
  NOR U50923 ( .A(n49724), .B(n51319), .Z(n51318) );
  IV U50924 ( .A(n51320), .Z(n49724) );
  XNOR U50925 ( .A(n51321), .B(n49713), .Z(n42209) );
  XOR U50926 ( .A(round_reg[367]), .B(n51146), .Z(n49713) );
  ANDN U50927 ( .B(n49712), .A(n47980), .Z(n51321) );
  XOR U50928 ( .A(n51322), .B(n51323), .Z(n48814) );
  XNOR U50929 ( .A(n49704), .B(n47673), .Z(n51323) );
  XNOR U50930 ( .A(n51324), .B(n50290), .Z(n47673) );
  XOR U50931 ( .A(round_reg[1025]), .B(n50156), .Z(n50290) );
  ANDN U50932 ( .B(n47703), .A(n47704), .Z(n51324) );
  XOR U50933 ( .A(round_reg[657]), .B(n51325), .Z(n47703) );
  XNOR U50934 ( .A(n51326), .B(n50275), .Z(n49704) );
  XOR U50935 ( .A(round_reg[1138]), .B(n51327), .Z(n50275) );
  ANDN U50936 ( .B(n47717), .A(n47718), .Z(n51326) );
  XNOR U50937 ( .A(round_reg[735]), .B(n51147), .Z(n47717) );
  XOR U50938 ( .A(n45122), .B(n51328), .Z(n51322) );
  XOR U50939 ( .A(n44740), .B(n46746), .Z(n51328) );
  XNOR U50940 ( .A(n51329), .B(n50279), .Z(n46746) );
  ANDN U50941 ( .B(n50705), .A(n51308), .Z(n51329) );
  XOR U50942 ( .A(round_reg[781]), .B(n51330), .Z(n50705) );
  XNOR U50943 ( .A(n51331), .B(n50286), .Z(n44740) );
  XOR U50944 ( .A(round_reg[1236]), .B(n51332), .Z(n50286) );
  ANDN U50945 ( .B(n47713), .A(n47714), .Z(n51331) );
  XOR U50946 ( .A(round_reg[878]), .B(n51333), .Z(n47713) );
  XNOR U50947 ( .A(n51334), .B(n50283), .Z(n45122) );
  XOR U50948 ( .A(round_reg[996]), .B(n51335), .Z(n50283) );
  ANDN U50949 ( .B(n47707), .A(n47708), .Z(n51334) );
  XOR U50950 ( .A(round_reg[949]), .B(n51336), .Z(n47707) );
  ANDN U50951 ( .B(n41055), .A(n42228), .Z(n51306) );
  XOR U50952 ( .A(n47118), .B(n43815), .Z(n42228) );
  XOR U50953 ( .A(n48470), .B(n50979), .Z(n43815) );
  XNOR U50954 ( .A(n51337), .B(n51338), .Z(n50979) );
  XNOR U50955 ( .A(n46534), .B(n45830), .Z(n51338) );
  XNOR U50956 ( .A(n51339), .B(n46973), .Z(n45830) );
  XNOR U50957 ( .A(round_reg[448]), .B(n49083), .Z(n46973) );
  ANDN U50958 ( .B(n46974), .A(n48342), .Z(n51339) );
  XOR U50959 ( .A(round_reg[1332]), .B(n50440), .Z(n48342) );
  XNOR U50960 ( .A(round_reg[87]), .B(n48508), .Z(n46974) );
  XNOR U50961 ( .A(n51340), .B(n47958), .Z(n46534) );
  XNOR U50962 ( .A(round_reg[614]), .B(n51341), .Z(n47958) );
  ANDN U50963 ( .B(n47120), .A(n47122), .Z(n51340) );
  XOR U50964 ( .A(round_reg[1425]), .B(n51342), .Z(n47122) );
  XOR U50965 ( .A(round_reg[205]), .B(n51343), .Z(n47120) );
  XNOR U50966 ( .A(n44857), .B(n51344), .Z(n51337) );
  XOR U50967 ( .A(n43894), .B(n45276), .Z(n51344) );
  XOR U50968 ( .A(n51345), .B(n46960), .Z(n45276) );
  XOR U50969 ( .A(round_reg[442]), .B(n51137), .Z(n46960) );
  ANDN U50970 ( .B(n46959), .A(n47115), .Z(n51345) );
  XOR U50971 ( .A(round_reg[1551]), .B(n51346), .Z(n47115) );
  XOR U50972 ( .A(round_reg[1]), .B(n51347), .Z(n46959) );
  XOR U50973 ( .A(n51348), .B(n46964), .Z(n43894) );
  XOR U50974 ( .A(round_reg[327]), .B(n51349), .Z(n46964) );
  ANDN U50975 ( .B(n46963), .A(n48444), .Z(n51348) );
  IV U50976 ( .A(n51350), .Z(n48444) );
  XOR U50977 ( .A(n51351), .B(n46970), .Z(n44857) );
  XOR U50978 ( .A(round_reg[546]), .B(n51352), .Z(n46970) );
  ANDN U50979 ( .B(n46969), .A(n47125), .Z(n51351) );
  XNOR U50980 ( .A(round_reg[1395]), .B(n50444), .Z(n47125) );
  XOR U50981 ( .A(round_reg[146]), .B(n51100), .Z(n46969) );
  XOR U50982 ( .A(n51353), .B(n51354), .Z(n48470) );
  XOR U50983 ( .A(n42523), .B(n49285), .Z(n51354) );
  XOR U50984 ( .A(n51355), .B(n48629), .Z(n49285) );
  AND U50985 ( .A(n48228), .B(n48227), .Z(n51355) );
  XNOR U50986 ( .A(n51356), .B(n51357), .Z(n42523) );
  XOR U50987 ( .A(n41584), .B(n51358), .Z(n51353) );
  XOR U50988 ( .A(n47322), .B(n51359), .Z(n51358) );
  XOR U50989 ( .A(n51360), .B(n48632), .Z(n47322) );
  XOR U50990 ( .A(n51361), .B(n48641), .Z(n41584) );
  NOR U50991 ( .A(n48234), .B(n48232), .Z(n51361) );
  XNOR U50992 ( .A(n51362), .B(n46963), .Z(n47118) );
  XNOR U50993 ( .A(round_reg[317]), .B(n49087), .Z(n46963) );
  IV U50994 ( .A(n51363), .Z(n49087) );
  ANDN U50995 ( .B(n47970), .A(n51350), .Z(n51362) );
  XOR U50996 ( .A(round_reg[1486]), .B(n50772), .Z(n51350) );
  XNOR U50997 ( .A(round_reg[1097]), .B(n51364), .Z(n47970) );
  XOR U50998 ( .A(n45781), .B(n47489), .Z(n41055) );
  XNOR U50999 ( .A(n51365), .B(n46983), .Z(n47489) );
  XOR U51000 ( .A(n36304), .B(n51366), .Z(n51236) );
  XNOR U51001 ( .A(n41039), .B(n38890), .Z(n51366) );
  XNOR U51002 ( .A(n51367), .B(n46664), .Z(n38890) );
  XNOR U51003 ( .A(n51368), .B(n51259), .Z(n46664) );
  XOR U51004 ( .A(n51369), .B(n48161), .Z(n51259) );
  ANDN U51005 ( .B(n51370), .A(n50194), .Z(n51369) );
  AND U51006 ( .A(n41948), .B(n41950), .Z(n51367) );
  XNOR U51007 ( .A(n50626), .B(n46181), .Z(n41950) );
  XNOR U51008 ( .A(n51150), .B(n50306), .Z(n46181) );
  XNOR U51009 ( .A(n51371), .B(n51372), .Z(n50306) );
  XNOR U51010 ( .A(n46297), .B(n44338), .Z(n51372) );
  XNOR U51011 ( .A(n51373), .B(n51374), .Z(n44338) );
  ANDN U51012 ( .B(n48900), .A(n48901), .Z(n51373) );
  XOR U51013 ( .A(round_reg[1061]), .B(n49901), .Z(n48901) );
  XOR U51014 ( .A(n51375), .B(n51376), .Z(n46297) );
  AND U51015 ( .A(n48892), .B(n48891), .Z(n51375) );
  XOR U51016 ( .A(round_reg[968]), .B(n48699), .Z(n48892) );
  IV U51017 ( .A(n51377), .Z(n48699) );
  XNOR U51018 ( .A(n45916), .B(n51378), .Z(n51371) );
  XNOR U51019 ( .A(n51379), .B(n45816), .Z(n51378) );
  XNOR U51020 ( .A(n51380), .B(n51381), .Z(n45816) );
  ANDN U51021 ( .B(n48896), .A(n48898), .Z(n51380) );
  XOR U51022 ( .A(round_reg[1272]), .B(n51224), .Z(n48898) );
  XOR U51023 ( .A(n51382), .B(n51383), .Z(n45916) );
  XNOR U51024 ( .A(round_reg[1110]), .B(n50482), .Z(n48905) );
  XOR U51025 ( .A(n51384), .B(n51385), .Z(n51150) );
  XOR U51026 ( .A(n46496), .B(n46276), .Z(n51385) );
  XNOR U51027 ( .A(n51386), .B(n51037), .Z(n46276) );
  ANDN U51028 ( .B(n50622), .A(n50623), .Z(n51386) );
  XOR U51029 ( .A(round_reg[219]), .B(n50442), .Z(n50623) );
  XOR U51030 ( .A(round_reg[628]), .B(n50299), .Z(n50622) );
  NOR U51031 ( .A(n50911), .B(n51389), .Z(n51387) );
  XNOR U51032 ( .A(n44401), .B(n51390), .Z(n51384) );
  XOR U51033 ( .A(n44013), .B(n45462), .Z(n51390) );
  XNOR U51034 ( .A(n51391), .B(n51392), .Z(n45462) );
  NOR U51035 ( .A(n50628), .B(n49160), .Z(n51391) );
  XNOR U51036 ( .A(round_reg[392]), .B(n51393), .Z(n49160) );
  XOR U51037 ( .A(round_reg[15]), .B(n48362), .Z(n50628) );
  AND U51038 ( .A(n50619), .B(n49530), .Z(n51394) );
  XOR U51039 ( .A(round_reg[462]), .B(n51395), .Z(n49530) );
  XNOR U51040 ( .A(round_reg[101]), .B(n49901), .Z(n50619) );
  XNOR U51041 ( .A(n51396), .B(n49424), .Z(n44401) );
  NOR U51042 ( .A(n49423), .B(n50631), .Z(n51396) );
  XOR U51043 ( .A(round_reg[160]), .B(n51397), .Z(n50631) );
  XOR U51044 ( .A(round_reg[560]), .B(n48938), .Z(n49423) );
  XNOR U51045 ( .A(n51398), .B(n51389), .Z(n50626) );
  ANDN U51046 ( .B(n50911), .A(n50912), .Z(n51398) );
  XOR U51047 ( .A(round_reg[267]), .B(n51399), .Z(n50911) );
  XNOR U51048 ( .A(n49404), .B(n43091), .Z(n41948) );
  XOR U51049 ( .A(n51400), .B(n47576), .Z(n43091) );
  XOR U51050 ( .A(n51401), .B(n51402), .Z(n47576) );
  XOR U51051 ( .A(n46442), .B(n50330), .Z(n51402) );
  XNOR U51052 ( .A(n51403), .B(n50336), .Z(n50330) );
  IV U51053 ( .A(n49653), .Z(n50336) );
  XOR U51054 ( .A(round_reg[988]), .B(n48965), .Z(n49653) );
  ANDN U51055 ( .B(n51404), .A(n50335), .Z(n51403) );
  XNOR U51056 ( .A(n51405), .B(n49656), .Z(n46442) );
  XNOR U51057 ( .A(round_reg[1156]), .B(n50505), .Z(n49656) );
  ANDN U51058 ( .B(n49412), .A(n49410), .Z(n51405) );
  XOR U51059 ( .A(round_reg[773]), .B(n51293), .Z(n49410) );
  XOR U51060 ( .A(n47441), .B(n51406), .Z(n51401) );
  XOR U51061 ( .A(n44590), .B(n43467), .Z(n51406) );
  XOR U51062 ( .A(n51407), .B(n49644), .Z(n43467) );
  XNOR U51063 ( .A(round_reg[1081]), .B(n51177), .Z(n49644) );
  ANDN U51064 ( .B(n50340), .A(n49401), .Z(n51407) );
  IV U51065 ( .A(n49400), .Z(n50340) );
  XOR U51066 ( .A(round_reg[649]), .B(n51408), .Z(n49400) );
  XOR U51067 ( .A(n51409), .B(n49641), .Z(n44590) );
  XNOR U51068 ( .A(round_reg[1130]), .B(n50761), .Z(n49641) );
  ANDN U51069 ( .B(n50490), .A(n50343), .Z(n51409) );
  XOR U51070 ( .A(round_reg[727]), .B(n48508), .Z(n50343) );
  XNOR U51071 ( .A(n51410), .B(n49649), .Z(n47441) );
  XNOR U51072 ( .A(round_reg[1228]), .B(n49427), .Z(n49649) );
  NOR U51073 ( .A(n49406), .B(n49407), .Z(n51410) );
  XOR U51074 ( .A(round_reg[870]), .B(n51411), .Z(n49406) );
  XOR U51075 ( .A(n51412), .B(n50335), .Z(n49404) );
  XOR U51076 ( .A(round_reg[941]), .B(n50153), .Z(n50335) );
  NOR U51077 ( .A(n49651), .B(n51404), .Z(n51412) );
  XOR U51078 ( .A(n51413), .B(n41059), .Z(n41039) );
  XNOR U51079 ( .A(n48998), .B(n42498), .Z(n41059) );
  XOR U51080 ( .A(n50143), .B(n50101), .Z(n42498) );
  XNOR U51081 ( .A(n51414), .B(n51415), .Z(n50101) );
  XOR U51082 ( .A(n51416), .B(n46644), .Z(n51415) );
  XOR U51083 ( .A(n51417), .B(n48597), .Z(n46644) );
  NOR U51084 ( .A(n50393), .B(n48768), .Z(n51417) );
  XOR U51085 ( .A(round_reg[1197]), .B(n50693), .Z(n48768) );
  XOR U51086 ( .A(n44025), .B(n51418), .Z(n51414) );
  XOR U51087 ( .A(n49022), .B(n45307), .Z(n51418) );
  XNOR U51088 ( .A(n51419), .B(n48584), .Z(n45307) );
  NOR U51089 ( .A(n51420), .B(n48770), .Z(n51419) );
  XNOR U51090 ( .A(round_reg[1107]), .B(n49904), .Z(n48770) );
  XNOR U51091 ( .A(n51421), .B(n48593), .Z(n49022) );
  ANDN U51092 ( .B(n50400), .A(n48772), .Z(n51421) );
  XOR U51093 ( .A(round_reg[1269]), .B(n51336), .Z(n48772) );
  XNOR U51094 ( .A(n51422), .B(n48589), .Z(n44025) );
  NOR U51095 ( .A(n48765), .B(n50396), .Z(n51422) );
  XOR U51096 ( .A(round_reg[965]), .B(n51041), .Z(n48765) );
  XOR U51097 ( .A(n51423), .B(n51424), .Z(n50143) );
  XOR U51098 ( .A(n43712), .B(n48400), .Z(n51424) );
  XOR U51099 ( .A(n51425), .B(n50792), .Z(n48400) );
  NOR U51100 ( .A(n51426), .B(n48995), .Z(n51425) );
  XNOR U51101 ( .A(round_reg[625]), .B(n48935), .Z(n48995) );
  XOR U51102 ( .A(n51427), .B(n50795), .Z(n43712) );
  NOR U51103 ( .A(n49003), .B(n49001), .Z(n51427) );
  XNOR U51104 ( .A(round_reg[338]), .B(n51428), .Z(n49001) );
  XOR U51105 ( .A(n50786), .B(n51429), .Z(n51423) );
  XOR U51106 ( .A(n45731), .B(n45086), .Z(n51429) );
  XNOR U51107 ( .A(n51430), .B(n50800), .Z(n45086) );
  ANDN U51108 ( .B(n51431), .A(n50799), .Z(n51430) );
  XNOR U51109 ( .A(n51432), .B(n51433), .Z(n45731) );
  ANDN U51110 ( .B(n48993), .A(n48991), .Z(n51432) );
  XNOR U51111 ( .A(round_reg[459]), .B(n51434), .Z(n48991) );
  XNOR U51112 ( .A(n51435), .B(n50806), .Z(n50786) );
  NOR U51113 ( .A(n49007), .B(n49005), .Z(n51435) );
  XNOR U51114 ( .A(round_reg[557]), .B(n50693), .Z(n49005) );
  XNOR U51115 ( .A(n51436), .B(n50799), .Z(n48998) );
  XNOR U51116 ( .A(round_reg[389]), .B(n51437), .Z(n50799) );
  ANDN U51117 ( .B(n51438), .A(n51431), .Z(n51436) );
  ANDN U51118 ( .B(n41060), .A(n41957), .Z(n51413) );
  XOR U51119 ( .A(n50897), .B(n43559), .Z(n41957) );
  XOR U51120 ( .A(n48930), .B(n47149), .Z(n43559) );
  XNOR U51121 ( .A(n51439), .B(n51440), .Z(n47149) );
  XNOR U51122 ( .A(n46548), .B(n49999), .Z(n51440) );
  XOR U51123 ( .A(n51441), .B(n50011), .Z(n49999) );
  XOR U51124 ( .A(round_reg[241]), .B(n50739), .Z(n50011) );
  AND U51125 ( .A(n49764), .B(n50012), .Z(n51441) );
  XOR U51126 ( .A(round_reg[1461]), .B(n50744), .Z(n50012) );
  XOR U51127 ( .A(round_reg[1084]), .B(n50751), .Z(n49764) );
  XNOR U51128 ( .A(n51442), .B(n50019), .Z(n46548) );
  XNOR U51129 ( .A(round_reg[182]), .B(n49795), .Z(n50019) );
  ANDN U51130 ( .B(n50018), .A(n49754), .Z(n51442) );
  XOR U51131 ( .A(round_reg[991]), .B(n50519), .Z(n49754) );
  XNOR U51132 ( .A(round_reg[1367]), .B(n48508), .Z(n50018) );
  IV U51133 ( .A(n51443), .Z(n48508) );
  XOR U51134 ( .A(n45932), .B(n51444), .Z(n51439) );
  XOR U51135 ( .A(n41587), .B(n44491), .Z(n51444) );
  XNOR U51136 ( .A(n51445), .B(n50015), .Z(n44491) );
  XNOR U51137 ( .A(round_reg[123]), .B(n50984), .Z(n50015) );
  AND U51138 ( .A(n50901), .B(n50016), .Z(n51445) );
  XOR U51139 ( .A(round_reg[1304]), .B(n51446), .Z(n50016) );
  XNOR U51140 ( .A(round_reg[1231]), .B(n51346), .Z(n50901) );
  XNOR U51141 ( .A(n51447), .B(n50004), .Z(n41587) );
  XNOR U51142 ( .A(round_reg[37]), .B(n50646), .Z(n50004) );
  ANDN U51143 ( .B(n50895), .A(n50005), .Z(n51447) );
  XOR U51144 ( .A(round_reg[1587]), .B(n50504), .Z(n50005) );
  IV U51145 ( .A(n49758), .Z(n50895) );
  XOR U51146 ( .A(round_reg[1159]), .B(n51448), .Z(n49758) );
  XNOR U51147 ( .A(n51449), .B(n50007), .Z(n45932) );
  XNOR U51148 ( .A(round_reg[289]), .B(n50501), .Z(n50007) );
  AND U51149 ( .A(n49768), .B(n50008), .Z(n51449) );
  XOR U51150 ( .A(n51450), .B(n51451), .Z(n48930) );
  XOR U51151 ( .A(n43539), .B(n47387), .Z(n51451) );
  XOR U51152 ( .A(n51452), .B(n50367), .Z(n47387) );
  XNOR U51153 ( .A(round_reg[990]), .B(n49633), .Z(n50367) );
  AND U51154 ( .A(n49748), .B(n50885), .Z(n51452) );
  XOR U51155 ( .A(round_reg[943]), .B(n50414), .Z(n50885) );
  XOR U51156 ( .A(round_reg[517]), .B(n48453), .Z(n49748) );
  XNOR U51157 ( .A(n51453), .B(n50363), .Z(n43539) );
  XNOR U51158 ( .A(round_reg[1158]), .B(n50116), .Z(n50363) );
  IV U51159 ( .A(n50940), .Z(n50116) );
  XOR U51160 ( .A(n51454), .B(n51455), .Z(n50940) );
  ANDN U51161 ( .B(n50887), .A(n49731), .Z(n51453) );
  XOR U51162 ( .A(round_reg[413]), .B(n51456), .Z(n49731) );
  XOR U51163 ( .A(round_reg[775]), .B(n51017), .Z(n50887) );
  IV U51164 ( .A(n50158), .Z(n51017) );
  XOR U51165 ( .A(n44529), .B(n51457), .Z(n51450) );
  XOR U51166 ( .A(n46564), .B(n51168), .Z(n51457) );
  XOR U51167 ( .A(n51458), .B(n50358), .Z(n51168) );
  XOR U51168 ( .A(round_reg[1230]), .B(n51047), .Z(n50358) );
  XOR U51169 ( .A(round_reg[872]), .B(n50756), .Z(n50881) );
  XNOR U51170 ( .A(round_reg[483]), .B(n51459), .Z(n49744) );
  XOR U51171 ( .A(n51460), .B(n50365), .Z(n46564) );
  XOR U51172 ( .A(round_reg[1083]), .B(n50984), .Z(n50365) );
  XOR U51173 ( .A(round_reg[651]), .B(n51461), .Z(n50878) );
  IV U51174 ( .A(n49740), .Z(n50879) );
  XOR U51175 ( .A(round_reg[585]), .B(n51462), .Z(n49740) );
  XOR U51176 ( .A(n51463), .B(n50360), .Z(n44529) );
  XNOR U51177 ( .A(round_reg[1132]), .B(n48365), .Z(n50360) );
  NOR U51178 ( .A(n49735), .B(n50890), .Z(n51463) );
  XNOR U51179 ( .A(round_reg[729]), .B(n51101), .Z(n50890) );
  XOR U51180 ( .A(round_reg[362]), .B(n51464), .Z(n49735) );
  XNOR U51181 ( .A(n51465), .B(n50008), .Z(n50897) );
  XOR U51182 ( .A(round_reg[1522]), .B(n51466), .Z(n50008) );
  NOR U51183 ( .A(n50936), .B(n49768), .Z(n51465) );
  XOR U51184 ( .A(round_reg[1133]), .B(n51467), .Z(n49768) );
  IV U51185 ( .A(n49769), .Z(n50936) );
  XNOR U51186 ( .A(round_reg[730]), .B(n51468), .Z(n49769) );
  XNOR U51187 ( .A(n50577), .B(n45255), .Z(n41060) );
  IV U51188 ( .A(n41731), .Z(n45255) );
  XOR U51189 ( .A(n46829), .B(n49327), .Z(n41731) );
  XNOR U51190 ( .A(n51469), .B(n51470), .Z(n49327) );
  XOR U51191 ( .A(n41882), .B(n46253), .Z(n51470) );
  XOR U51192 ( .A(n51471), .B(n51212), .Z(n46253) );
  NOR U51193 ( .A(n47177), .B(n51472), .Z(n51471) );
  XNOR U51194 ( .A(n51473), .B(n51215), .Z(n41882) );
  XNOR U51195 ( .A(round_reg[1570]), .B(n50822), .Z(n47191) );
  XOR U51196 ( .A(n44560), .B(n51474), .Z(n51469) );
  XOR U51197 ( .A(n46280), .B(n51475), .Z(n51474) );
  XNOR U51198 ( .A(n51476), .B(n51218), .Z(n46280) );
  ANDN U51199 ( .B(n50574), .A(n47187), .Z(n51476) );
  XNOR U51200 ( .A(round_reg[1444]), .B(n48449), .Z(n47187) );
  XNOR U51201 ( .A(n51477), .B(n51210), .Z(n44560) );
  ANDN U51202 ( .B(n50580), .A(n47181), .Z(n51477) );
  XOR U51203 ( .A(round_reg[1505]), .B(n51478), .Z(n47181) );
  XNOR U51204 ( .A(n51479), .B(n51480), .Z(n46829) );
  XOR U51205 ( .A(n45819), .B(n43541), .Z(n51480) );
  XOR U51206 ( .A(n51481), .B(n51225), .Z(n43541) );
  ANDN U51207 ( .B(n51066), .A(n48420), .Z(n51481) );
  XNOR U51208 ( .A(round_reg[698]), .B(n50110), .Z(n48420) );
  XNOR U51209 ( .A(n51482), .B(n51231), .Z(n45819) );
  ANDN U51210 ( .B(n51057), .A(n48410), .Z(n51482) );
  XNOR U51211 ( .A(round_reg[712]), .B(n51483), .Z(n48410) );
  XOR U51212 ( .A(n41648), .B(n51484), .Z(n51479) );
  XOR U51213 ( .A(n49437), .B(n44947), .Z(n51484) );
  XNOR U51214 ( .A(n51485), .B(n51228), .Z(n44947) );
  ANDN U51215 ( .B(n51059), .A(n48424), .Z(n51485) );
  XNOR U51216 ( .A(round_reg[926]), .B(n51486), .Z(n48424) );
  XNOR U51217 ( .A(n51487), .B(n51233), .Z(n49437) );
  ANDN U51218 ( .B(n51069), .A(n48414), .Z(n51487) );
  XNOR U51219 ( .A(round_reg[855]), .B(n50995), .Z(n48414) );
  XNOR U51220 ( .A(n51488), .B(n51235), .Z(n41648) );
  NOR U51221 ( .A(n51489), .B(n51063), .Z(n51488) );
  XOR U51222 ( .A(round_reg[822]), .B(n49795), .Z(n51063) );
  XNOR U51223 ( .A(n51490), .B(n51472), .Z(n50577) );
  ANDN U51224 ( .B(n47177), .A(n47178), .Z(n51490) );
  XOR U51225 ( .A(round_reg[974]), .B(n51491), .Z(n47178) );
  XNOR U51226 ( .A(round_reg[1350]), .B(n49271), .Z(n47177) );
  XNOR U51227 ( .A(n51492), .B(n41046), .Z(n36304) );
  XNOR U51228 ( .A(n44659), .B(n47218), .Z(n41046) );
  XNOR U51229 ( .A(n51493), .B(n51494), .Z(n47218) );
  ANDN U51230 ( .B(n51495), .A(n50323), .Z(n51493) );
  IV U51231 ( .A(n51496), .Z(n50323) );
  XOR U51232 ( .A(n48574), .B(n46272), .Z(n44659) );
  XNOR U51233 ( .A(n51497), .B(n51498), .Z(n46272) );
  XNOR U51234 ( .A(n45372), .B(n46424), .Z(n51498) );
  XOR U51235 ( .A(n51499), .B(n50320), .Z(n46424) );
  NOR U51236 ( .A(n47227), .B(n47226), .Z(n51499) );
  XNOR U51237 ( .A(n51500), .B(n50317), .Z(n45372) );
  ANDN U51238 ( .B(n47220), .A(n47221), .Z(n51500) );
  XNOR U51239 ( .A(n45357), .B(n51501), .Z(n51497) );
  XOR U51240 ( .A(n43534), .B(n51502), .Z(n51501) );
  XNOR U51241 ( .A(n51503), .B(n50310), .Z(n43534) );
  ANDN U51242 ( .B(n49698), .A(n49699), .Z(n51503) );
  XOR U51243 ( .A(n51504), .B(n50313), .Z(n45357) );
  ANDN U51244 ( .B(n47230), .A(n47232), .Z(n51504) );
  XOR U51245 ( .A(n51505), .B(n51506), .Z(n48574) );
  XNOR U51246 ( .A(n46265), .B(n44190), .Z(n51506) );
  XNOR U51247 ( .A(n51507), .B(n49006), .Z(n44190) );
  ANDN U51248 ( .B(n50805), .A(n50806), .Z(n51507) );
  XOR U51249 ( .A(round_reg[919]), .B(n50738), .Z(n50806) );
  XNOR U51250 ( .A(n51508), .B(n51438), .Z(n46265) );
  ANDN U51251 ( .B(n50798), .A(n50800), .Z(n51508) );
  XOR U51252 ( .A(round_reg[815]), .B(n49631), .Z(n50800) );
  XNOR U51253 ( .A(n47585), .B(n51509), .Z(n51505) );
  XOR U51254 ( .A(n45410), .B(n48760), .Z(n51509) );
  XOR U51255 ( .A(n51510), .B(n51511), .Z(n48760) );
  AND U51256 ( .A(n50795), .B(n50794), .Z(n51510) );
  XOR U51257 ( .A(round_reg[705]), .B(n51512), .Z(n50795) );
  XOR U51258 ( .A(n51513), .B(n51514), .Z(n45410) );
  ANDN U51259 ( .B(n50791), .A(n50792), .Z(n51513) );
  XOR U51260 ( .A(round_reg[691]), .B(n50136), .Z(n50792) );
  XOR U51261 ( .A(n51515), .B(n48992), .Z(n47585) );
  ANDN U51262 ( .B(n50802), .A(n51433), .Z(n51515) );
  IV U51263 ( .A(n50803), .Z(n51433) );
  XOR U51264 ( .A(round_reg[848]), .B(n51516), .Z(n50803) );
  ANDN U51265 ( .B(n41047), .A(n41954), .Z(n51492) );
  XOR U51266 ( .A(n47335), .B(n42395), .Z(n41954) );
  XOR U51267 ( .A(n46550), .B(n49885), .Z(n42395) );
  XNOR U51268 ( .A(n51517), .B(n51518), .Z(n49885) );
  XNOR U51269 ( .A(n45413), .B(n42308), .Z(n51518) );
  XOR U51270 ( .A(n51519), .B(n48521), .Z(n42308) );
  XNOR U51271 ( .A(round_reg[1360]), .B(n50119), .Z(n48521) );
  AND U51272 ( .A(n47351), .B(n48502), .Z(n51519) );
  XOR U51273 ( .A(round_reg[984]), .B(n51446), .Z(n48502) );
  XOR U51274 ( .A(round_reg[937]), .B(n51520), .Z(n47351) );
  XNOR U51275 ( .A(n51521), .B(n48509), .Z(n45413) );
  XOR U51276 ( .A(round_reg[1580]), .B(n50749), .Z(n48509) );
  ANDN U51277 ( .B(n47333), .A(n46333), .Z(n51521) );
  XOR U51278 ( .A(round_reg[1152]), .B(n50415), .Z(n47333) );
  XNOR U51279 ( .A(n46347), .B(n51522), .Z(n51517) );
  XOR U51280 ( .A(n42544), .B(n46113), .Z(n51522) );
  XNOR U51281 ( .A(n51523), .B(n48518), .Z(n46113) );
  XOR U51282 ( .A(round_reg[1297]), .B(n51325), .Z(n48518) );
  AND U51283 ( .A(n46337), .B(n47337), .Z(n51523) );
  XNOR U51284 ( .A(round_reg[1224]), .B(n50111), .Z(n47337) );
  XOR U51285 ( .A(round_reg[866]), .B(n48708), .Z(n46337) );
  XOR U51286 ( .A(n51524), .B(n48515), .Z(n42544) );
  XOR U51287 ( .A(round_reg[1454]), .B(n51525), .Z(n48515) );
  ANDN U51288 ( .B(n47339), .A(n46323), .Z(n51524) );
  XOR U51289 ( .A(round_reg[645]), .B(n51041), .Z(n46323) );
  IV U51290 ( .A(n50479), .Z(n51041) );
  XOR U51291 ( .A(round_reg[1077]), .B(n51526), .Z(n47339) );
  XOR U51292 ( .A(n51527), .B(n49627), .Z(n46347) );
  XOR U51293 ( .A(round_reg[1515]), .B(n51528), .Z(n49627) );
  NOR U51294 ( .A(n46327), .B(n49626), .Z(n51527) );
  XOR U51295 ( .A(n51529), .B(n51530), .Z(n46550) );
  XNOR U51296 ( .A(n46370), .B(n45701), .Z(n51530) );
  XNOR U51297 ( .A(n51531), .B(n46687), .Z(n45701) );
  IV U51298 ( .A(n48565), .Z(n46687) );
  XOR U51299 ( .A(round_reg[722]), .B(n51532), .Z(n48565) );
  ANDN U51300 ( .B(n46688), .A(n47081), .Z(n51531) );
  XOR U51301 ( .A(round_reg[281]), .B(n50434), .Z(n47081) );
  XNOR U51302 ( .A(round_reg[355]), .B(n51533), .Z(n46688) );
  XNOR U51303 ( .A(n51534), .B(n46376), .Z(n46370) );
  XOR U51304 ( .A(round_reg[936]), .B(n49984), .Z(n46376) );
  IV U51305 ( .A(n51535), .Z(n49984) );
  ANDN U51306 ( .B(n46377), .A(n47088), .Z(n51534) );
  XOR U51307 ( .A(round_reg[174]), .B(n50394), .Z(n47088) );
  XOR U51308 ( .A(round_reg[574]), .B(n50448), .Z(n46377) );
  XNOR U51309 ( .A(n44592), .B(n51536), .Z(n51529) );
  XNOR U51310 ( .A(n44217), .B(n45754), .Z(n51536) );
  XNOR U51311 ( .A(n51537), .B(n46387), .Z(n45754) );
  XNOR U51312 ( .A(round_reg[644]), .B(n51538), .Z(n46387) );
  ANDN U51313 ( .B(n46388), .A(n47085), .Z(n51537) );
  XOR U51314 ( .A(round_reg[233]), .B(n50942), .Z(n47085) );
  XNOR U51315 ( .A(round_reg[578]), .B(n51539), .Z(n46388) );
  XOR U51316 ( .A(n51540), .B(n46380), .Z(n44217) );
  XOR U51317 ( .A(round_reg[768]), .B(n49083), .Z(n46380) );
  ANDN U51318 ( .B(n46381), .A(n47343), .Z(n51540) );
  XOR U51319 ( .A(round_reg[29]), .B(n51541), .Z(n47343) );
  XOR U51320 ( .A(round_reg[406]), .B(n51542), .Z(n46381) );
  XOR U51321 ( .A(n51543), .B(n48562), .Z(n44592) );
  XOR U51322 ( .A(round_reg[865]), .B(n51478), .Z(n48562) );
  NOR U51323 ( .A(n47091), .B(n47349), .Z(n51543) );
  XOR U51324 ( .A(round_reg[476]), .B(n51544), .Z(n47349) );
  XOR U51325 ( .A(round_reg[115]), .B(n51545), .Z(n47091) );
  XOR U51326 ( .A(n51546), .B(n49626), .Z(n47335) );
  XNOR U51327 ( .A(round_reg[1126]), .B(n51547), .Z(n49626) );
  XOR U51328 ( .A(round_reg[723]), .B(n51548), .Z(n46327) );
  XOR U51329 ( .A(round_reg[356]), .B(n50888), .Z(n46329) );
  XNOR U51330 ( .A(n44497), .B(n50466), .Z(n41047) );
  XNOR U51331 ( .A(n51549), .B(n51550), .Z(n50466) );
  ANDN U51332 ( .B(n49109), .A(n49110), .Z(n51549) );
  IV U51333 ( .A(n45353), .Z(n44497) );
  XOR U51334 ( .A(n45893), .B(n50779), .Z(n45353) );
  XNOR U51335 ( .A(n51551), .B(n51552), .Z(n50779) );
  XOR U51336 ( .A(n50552), .B(n45384), .Z(n51552) );
  XOR U51337 ( .A(n51553), .B(n51554), .Z(n45384) );
  ANDN U51338 ( .B(n50253), .A(n50255), .Z(n51553) );
  XOR U51339 ( .A(round_reg[616]), .B(n51535), .Z(n50255) );
  XNOR U51340 ( .A(n51555), .B(n51556), .Z(n50552) );
  AND U51341 ( .A(n50260), .B(n50259), .Z(n51555) );
  XNOR U51342 ( .A(round_reg[329]), .B(n51557), .Z(n50260) );
  XOR U51343 ( .A(n45347), .B(n51558), .Z(n51551) );
  XOR U51344 ( .A(n44179), .B(n43318), .Z(n51558) );
  XNOR U51345 ( .A(n51559), .B(n51560), .Z(n43318) );
  AND U51346 ( .A(n50265), .B(n50263), .Z(n51559) );
  XOR U51347 ( .A(round_reg[548]), .B(n51561), .Z(n50265) );
  XNOR U51348 ( .A(n51562), .B(n51563), .Z(n44179) );
  XNOR U51349 ( .A(round_reg[450]), .B(n51564), .Z(n50783) );
  XNOR U51350 ( .A(n51565), .B(n51566), .Z(n45347) );
  ANDN U51351 ( .B(n50249), .A(n50251), .Z(n51565) );
  XOR U51352 ( .A(round_reg[444]), .B(n51567), .Z(n50251) );
  XOR U51353 ( .A(n51568), .B(n51569), .Z(n45893) );
  XOR U51354 ( .A(n50654), .B(n42821), .Z(n51569) );
  XOR U51355 ( .A(n51570), .B(n51571), .Z(n42821) );
  NOR U51356 ( .A(n49101), .B(n50470), .Z(n51570) );
  XOR U51357 ( .A(round_reg[1190]), .B(n51572), .Z(n49101) );
  XNOR U51358 ( .A(n51573), .B(n51574), .Z(n50654) );
  ANDN U51359 ( .B(n50462), .A(n49096), .Z(n51573) );
  XNOR U51360 ( .A(round_reg[1051]), .B(n50485), .Z(n49096) );
  XOR U51361 ( .A(n51575), .B(n51576), .Z(n51568) );
  XNOR U51362 ( .A(n45944), .B(n47806), .Z(n51576) );
  XNOR U51363 ( .A(n51577), .B(n51578), .Z(n47806) );
  ANDN U51364 ( .B(n50468), .A(n50267), .Z(n51577) );
  XOR U51365 ( .A(round_reg[1100]), .B(n51579), .Z(n50267) );
  XOR U51366 ( .A(n51580), .B(n51581), .Z(n45944) );
  ANDN U51367 ( .B(n50464), .A(n49105), .Z(n51580) );
  XOR U51368 ( .A(round_reg[1262]), .B(n51582), .Z(n49105) );
  XOR U51369 ( .A(n51583), .B(n51584), .Z(n39417) );
  XNOR U51370 ( .A(n39554), .B(n40047), .Z(n51584) );
  XOR U51371 ( .A(n51585), .B(n41785), .Z(n40047) );
  XOR U51372 ( .A(n51359), .B(n42524), .Z(n41785) );
  XOR U51373 ( .A(n46536), .B(n49535), .Z(n42524) );
  XNOR U51374 ( .A(n51586), .B(n51587), .Z(n49535) );
  XNOR U51375 ( .A(n46008), .B(n43862), .Z(n51587) );
  XOR U51376 ( .A(n51588), .B(n51166), .Z(n43862) );
  ANDN U51377 ( .B(n49540), .A(n49538), .Z(n51588) );
  XNOR U51378 ( .A(round_reg[678]), .B(n51589), .Z(n49538) );
  XOR U51379 ( .A(round_reg[612]), .B(n51250), .Z(n49540) );
  XNOR U51380 ( .A(n51590), .B(n48648), .Z(n46008) );
  ANDN U51381 ( .B(n48483), .A(n48481), .Z(n51590) );
  XOR U51382 ( .A(round_reg[756]), .B(n48559), .Z(n48481) );
  XOR U51383 ( .A(round_reg[325]), .B(n50479), .Z(n48483) );
  XNOR U51384 ( .A(n51591), .B(n51592), .Z(n50479) );
  XOR U51385 ( .A(n47842), .B(n51593), .Z(n51586) );
  XOR U51386 ( .A(n44595), .B(n44780), .Z(n51593) );
  XNOR U51387 ( .A(n51594), .B(n48652), .Z(n44780) );
  ANDN U51388 ( .B(n48487), .A(n48485), .Z(n51594) );
  XOR U51389 ( .A(round_reg[802]), .B(n51595), .Z(n48485) );
  XOR U51390 ( .A(round_reg[440]), .B(n49977), .Z(n48487) );
  XOR U51391 ( .A(n51596), .B(n48656), .Z(n44595) );
  XNOR U51392 ( .A(round_reg[835]), .B(n51597), .Z(n48655) );
  XOR U51393 ( .A(round_reg[510]), .B(n50728), .Z(n48692) );
  XNOR U51394 ( .A(n51598), .B(n48659), .Z(n47842) );
  NOR U51395 ( .A(n50535), .B(n48475), .Z(n51598) );
  XOR U51396 ( .A(round_reg[906]), .B(n51599), .Z(n48475) );
  IV U51397 ( .A(n48476), .Z(n50535) );
  XOR U51398 ( .A(round_reg[544]), .B(n51161), .Z(n48476) );
  XOR U51399 ( .A(n51600), .B(n51601), .Z(n46536) );
  XNOR U51400 ( .A(n48624), .B(n44233), .Z(n51601) );
  XOR U51401 ( .A(n51602), .B(n48642), .Z(n44233) );
  ANDN U51402 ( .B(n48232), .A(n48641), .Z(n51602) );
  XOR U51403 ( .A(round_reg[1550]), .B(n51047), .Z(n48641) );
  XNOR U51404 ( .A(round_reg[1186]), .B(n51352), .Z(n48232) );
  XNOR U51405 ( .A(n51603), .B(n48628), .Z(n48624) );
  ANDN U51406 ( .B(n48629), .A(n48227), .Z(n51603) );
  XOR U51407 ( .A(round_reg[1047]), .B(n51443), .Z(n48227) );
  XOR U51408 ( .A(n51604), .B(n51605), .Z(n51443) );
  XNOR U51409 ( .A(round_reg[1424]), .B(n50735), .Z(n48629) );
  XOR U51410 ( .A(n46696), .B(n51606), .Z(n51600) );
  XOR U51411 ( .A(n42666), .B(n46036), .Z(n51606) );
  XNOR U51412 ( .A(n51607), .B(n48638), .Z(n46036) );
  ANDN U51413 ( .B(n48639), .A(n48236), .Z(n51607) );
  XNOR U51414 ( .A(n51608), .B(n48633), .Z(n42666) );
  NOR U51415 ( .A(n48240), .B(n48632), .Z(n51608) );
  XOR U51416 ( .A(round_reg[1394]), .B(n50829), .Z(n48632) );
  XOR U51417 ( .A(round_reg[1018]), .B(n51609), .Z(n48240) );
  XNOR U51418 ( .A(n51610), .B(n51611), .Z(n46696) );
  ANDN U51419 ( .B(n51357), .A(n48489), .Z(n51610) );
  XOR U51420 ( .A(round_reg[1096]), .B(n50497), .Z(n48489) );
  XNOR U51421 ( .A(n51612), .B(n48639), .Z(n51359) );
  XOR U51422 ( .A(round_reg[1331]), .B(n50136), .Z(n48639) );
  ANDN U51423 ( .B(n48236), .A(n48237), .Z(n51612) );
  XOR U51424 ( .A(round_reg[1258]), .B(n48356), .Z(n48236) );
  AND U51425 ( .A(n42844), .B(n40120), .Z(n51585) );
  XOR U51426 ( .A(n51613), .B(n44681), .Z(n40120) );
  IV U51427 ( .A(n45828), .Z(n44681) );
  XNOR U51428 ( .A(n51614), .B(n51615), .Z(n47972) );
  XOR U51429 ( .A(n46429), .B(n45513), .Z(n51615) );
  XOR U51430 ( .A(n51616), .B(n47708), .Z(n45513) );
  XNOR U51431 ( .A(round_reg[523]), .B(n50758), .Z(n47708) );
  ANDN U51432 ( .B(n47709), .A(n50282), .Z(n51616) );
  XOR U51433 ( .A(round_reg[1372]), .B(n51617), .Z(n50282) );
  XNOR U51434 ( .A(round_reg[187]), .B(n51618), .Z(n47709) );
  XNOR U51435 ( .A(n51619), .B(n47704), .Z(n46429) );
  XOR U51436 ( .A(round_reg[591]), .B(n51346), .Z(n47704) );
  ANDN U51437 ( .B(n50289), .A(n50288), .Z(n51619) );
  IV U51438 ( .A(n47705), .Z(n50288) );
  XOR U51439 ( .A(round_reg[246]), .B(n50234), .Z(n47705) );
  XOR U51440 ( .A(round_reg[1466]), .B(n51620), .Z(n50289) );
  XOR U51441 ( .A(n42502), .B(n51621), .Z(n51614) );
  XOR U51442 ( .A(n46153), .B(n46882), .Z(n51621) );
  XNOR U51443 ( .A(n51622), .B(n47714), .Z(n46882) );
  XNOR U51444 ( .A(round_reg[489]), .B(n49947), .Z(n47714) );
  ANDN U51445 ( .B(n47715), .A(n50285), .Z(n51622) );
  XNOR U51446 ( .A(round_reg[1309]), .B(n49869), .Z(n50285) );
  XOR U51447 ( .A(round_reg[64]), .B(n50407), .Z(n47715) );
  XNOR U51448 ( .A(n51623), .B(n51308), .Z(n46153) );
  XOR U51449 ( .A(round_reg[419]), .B(n51624), .Z(n51308) );
  ANDN U51450 ( .B(n50278), .A(n50277), .Z(n51623) );
  XOR U51451 ( .A(round_reg[42]), .B(n50502), .Z(n50277) );
  XOR U51452 ( .A(round_reg[1592]), .B(n50733), .Z(n50278) );
  XNOR U51453 ( .A(n51625), .B(n47718), .Z(n42502) );
  XOR U51454 ( .A(round_reg[368]), .B(n49856), .Z(n47718) );
  ANDN U51455 ( .B(n47719), .A(n50274), .Z(n51625) );
  XNOR U51456 ( .A(round_reg[1527]), .B(n51626), .Z(n50274) );
  XOR U51457 ( .A(round_reg[294]), .B(n51341), .Z(n47719) );
  XNOR U51458 ( .A(n51627), .B(n51628), .Z(n47995) );
  XNOR U51459 ( .A(n45928), .B(n44499), .Z(n51628) );
  XOR U51460 ( .A(n51629), .B(n48826), .Z(n44499) );
  XOR U51461 ( .A(round_reg[1026]), .B(n51630), .Z(n48826) );
  AND U51462 ( .A(n51631), .B(n49678), .Z(n51629) );
  XNOR U51463 ( .A(round_reg[1139]), .B(n48942), .Z(n49682) );
  ANDN U51464 ( .B(n51633), .A(n49681), .Z(n51632) );
  XNOR U51465 ( .A(n47449), .B(n51634), .Z(n51627) );
  XOR U51466 ( .A(n47538), .B(n47698), .Z(n51634) );
  XNOR U51467 ( .A(n51635), .B(n48829), .Z(n47698) );
  XNOR U51468 ( .A(round_reg[1165]), .B(n51343), .Z(n48829) );
  AND U51469 ( .A(n51636), .B(n49691), .Z(n51635) );
  XNOR U51470 ( .A(n51637), .B(n48820), .Z(n47538) );
  XOR U51471 ( .A(round_reg[1237]), .B(n49907), .Z(n48820) );
  NOR U51472 ( .A(n51638), .B(n49686), .Z(n51637) );
  XNOR U51473 ( .A(n51639), .B(n48833), .Z(n47449) );
  XNOR U51474 ( .A(round_reg[997]), .B(n51640), .Z(n48833) );
  AND U51475 ( .A(n51641), .B(n49689), .Z(n51639) );
  XNOR U51476 ( .A(n51368), .B(n51264), .Z(n42844) );
  XOR U51477 ( .A(n51642), .B(n48157), .Z(n51264) );
  ANDN U51478 ( .B(n51643), .A(n50189), .Z(n51642) );
  IV U51479 ( .A(n43587), .Z(n51368) );
  XNOR U51480 ( .A(n49330), .B(n47148), .Z(n43587) );
  XNOR U51481 ( .A(n51644), .B(n51645), .Z(n47148) );
  XOR U51482 ( .A(n45220), .B(n47245), .Z(n51645) );
  XOR U51483 ( .A(n51646), .B(n47734), .Z(n47245) );
  XNOR U51484 ( .A(round_reg[653]), .B(n50752), .Z(n47734) );
  ANDN U51485 ( .B(n50969), .A(n47733), .Z(n51646) );
  XOR U51486 ( .A(round_reg[587]), .B(n51647), .Z(n47733) );
  IV U51487 ( .A(n49616), .Z(n50969) );
  XOR U51488 ( .A(round_reg[242]), .B(n51466), .Z(n49616) );
  XNOR U51489 ( .A(n51648), .B(n47738), .Z(n45220) );
  XNOR U51490 ( .A(round_reg[731]), .B(n50485), .Z(n47738) );
  NOR U51491 ( .A(n47737), .B(n50351), .Z(n51648) );
  XOR U51492 ( .A(round_reg[364]), .B(n49982), .Z(n47737) );
  XOR U51493 ( .A(n47720), .B(n51649), .Z(n51644) );
  XOR U51494 ( .A(n47544), .B(n47324), .Z(n51649) );
  XNOR U51495 ( .A(n51650), .B(n47727), .Z(n47324) );
  XNOR U51496 ( .A(round_reg[777]), .B(n50124), .Z(n47727) );
  NOR U51497 ( .A(n47728), .B(n49553), .Z(n51650) );
  XNOR U51498 ( .A(round_reg[38]), .B(n50412), .Z(n49553) );
  XOR U51499 ( .A(round_reg[415]), .B(n51147), .Z(n47728) );
  XNOR U51500 ( .A(n51651), .B(n49135), .Z(n47544) );
  XOR U51501 ( .A(round_reg[874]), .B(n48564), .Z(n49135) );
  ANDN U51502 ( .B(n49548), .A(n49134), .Z(n51651) );
  XOR U51503 ( .A(round_reg[485]), .B(n48566), .Z(n49134) );
  XOR U51504 ( .A(round_reg[124]), .B(n50751), .Z(n49548) );
  IV U51505 ( .A(n51567), .Z(n50751) );
  XNOR U51506 ( .A(n51652), .B(n50952), .Z(n47720) );
  XOR U51507 ( .A(round_reg[945]), .B(n48935), .Z(n50952) );
  ANDN U51508 ( .B(n49556), .A(n50958), .Z(n51652) );
  XOR U51509 ( .A(round_reg[519]), .B(n50107), .Z(n50958) );
  XNOR U51510 ( .A(round_reg[183]), .B(n50523), .Z(n49556) );
  XOR U51511 ( .A(n51653), .B(n51654), .Z(n49330) );
  XOR U51512 ( .A(n46674), .B(n46249), .Z(n51654) );
  XOR U51513 ( .A(n51655), .B(n49350), .Z(n46249) );
  XNOR U51514 ( .A(round_reg[1369]), .B(n51656), .Z(n49350) );
  NOR U51515 ( .A(n51261), .B(n51262), .Z(n51655) );
  IV U51516 ( .A(n49351), .Z(n51261) );
  XOR U51517 ( .A(round_reg[993]), .B(n50715), .Z(n49351) );
  XNOR U51518 ( .A(n51657), .B(n48160), .Z(n46674) );
  XNOR U51519 ( .A(round_reg[1589]), .B(n50842), .Z(n48160) );
  IV U51520 ( .A(n51336), .Z(n50842) );
  XOR U51521 ( .A(n51658), .B(n51659), .Z(n51336) );
  XOR U51522 ( .A(round_reg[1161]), .B(n51660), .Z(n48161) );
  XOR U51523 ( .A(n46730), .B(n51661), .Z(n51653) );
  XOR U51524 ( .A(n46553), .B(n45202), .Z(n51661) );
  XNOR U51525 ( .A(n51662), .B(n48150), .Z(n45202) );
  XOR U51526 ( .A(round_reg[1306]), .B(n51663), .Z(n48150) );
  ANDN U51527 ( .B(n48151), .A(n51268), .Z(n51662) );
  XNOR U51528 ( .A(round_reg[1233]), .B(n51664), .Z(n48151) );
  XNOR U51529 ( .A(n51665), .B(n48156), .Z(n46553) );
  XOR U51530 ( .A(round_reg[1463]), .B(n50523), .Z(n48156) );
  XOR U51531 ( .A(round_reg[1086]), .B(n51243), .Z(n48157) );
  XNOR U51532 ( .A(n51666), .B(n50181), .Z(n46730) );
  XNOR U51533 ( .A(round_reg[1524]), .B(n51246), .Z(n50181) );
  ANDN U51534 ( .B(n50182), .A(n51266), .Z(n51666) );
  XOR U51535 ( .A(round_reg[1135]), .B(n49631), .Z(n50182) );
  XOR U51536 ( .A(n51667), .B(n41792), .Z(n39554) );
  XOR U51537 ( .A(n51475), .B(n41883), .Z(n41792) );
  XNOR U51538 ( .A(n51668), .B(n51669), .Z(n47454) );
  XOR U51539 ( .A(n42162), .B(n51206), .Z(n51669) );
  XOR U51540 ( .A(n51670), .B(n47189), .Z(n51206) );
  XOR U51541 ( .A(round_reg[699]), .B(n48455), .Z(n47189) );
  ANDN U51542 ( .B(n51218), .A(n50574), .Z(n51670) );
  XOR U51543 ( .A(round_reg[224]), .B(n51671), .Z(n50574) );
  XNOR U51544 ( .A(round_reg[633]), .B(n51672), .Z(n51218) );
  XNOR U51545 ( .A(n51673), .B(n47183), .Z(n42162) );
  XOR U51546 ( .A(round_reg[713]), .B(n50227), .Z(n47183) );
  XNOR U51547 ( .A(round_reg[272]), .B(n50955), .Z(n50580) );
  XOR U51548 ( .A(round_reg[346]), .B(n51663), .Z(n51210) );
  XOR U51549 ( .A(n44265), .B(n51674), .Z(n51668) );
  XOR U51550 ( .A(n47250), .B(n49226), .Z(n51674) );
  XNOR U51551 ( .A(n51675), .B(n47193), .Z(n49226) );
  XOR U51552 ( .A(round_reg[823]), .B(n50523), .Z(n47193) );
  ANDN U51553 ( .B(n51215), .A(n50576), .Z(n51675) );
  XOR U51554 ( .A(round_reg[20]), .B(n51676), .Z(n50576) );
  XNOR U51555 ( .A(round_reg[397]), .B(n48869), .Z(n51215) );
  XOR U51556 ( .A(n51677), .B(n48036), .Z(n47250) );
  XNOR U51557 ( .A(round_reg[856]), .B(n49789), .Z(n48036) );
  AND U51558 ( .A(n50582), .B(n51220), .Z(n51677) );
  XNOR U51559 ( .A(n51678), .B(n47179), .Z(n44265) );
  XNOR U51560 ( .A(round_reg[927]), .B(n50453), .Z(n47179) );
  AND U51561 ( .A(n51472), .B(n51212), .Z(n51678) );
  XOR U51562 ( .A(round_reg[565]), .B(n51679), .Z(n51212) );
  XOR U51563 ( .A(n51682), .B(n51683), .Z(n49438) );
  XNOR U51564 ( .A(n46359), .B(n43312), .Z(n51683) );
  XNOR U51565 ( .A(n51684), .B(n51071), .Z(n43312) );
  XNOR U51566 ( .A(round_reg[19]), .B(n51685), .Z(n51071) );
  ANDN U51567 ( .B(n51235), .A(n51062), .Z(n51684) );
  IV U51568 ( .A(n51489), .Z(n51062) );
  XNOR U51569 ( .A(round_reg[1205]), .B(n51679), .Z(n51489) );
  XNOR U51570 ( .A(round_reg[1569]), .B(n50501), .Z(n51235) );
  XNOR U51571 ( .A(n51686), .B(n48422), .Z(n46359) );
  XNOR U51572 ( .A(round_reg[223]), .B(n51687), .Z(n48422) );
  ANDN U51573 ( .B(n51225), .A(n51066), .Z(n51686) );
  XOR U51574 ( .A(round_reg[1066]), .B(n51688), .Z(n51066) );
  XOR U51575 ( .A(round_reg[1443]), .B(n51459), .Z(n51225) );
  XOR U51576 ( .A(n46670), .B(n51689), .Z(n51682) );
  XNOR U51577 ( .A(n46509), .B(n45736), .Z(n51689) );
  XOR U51578 ( .A(n51690), .B(n48416), .Z(n45736) );
  XOR U51579 ( .A(round_reg[105]), .B(n49905), .Z(n48416) );
  ANDN U51580 ( .B(n51233), .A(n51069), .Z(n51690) );
  XOR U51581 ( .A(round_reg[1277]), .B(n51363), .Z(n51069) );
  XOR U51582 ( .A(n51691), .B(n51692), .Z(n51363) );
  XOR U51583 ( .A(round_reg[1286]), .B(n50643), .Z(n51233) );
  XNOR U51584 ( .A(n51693), .B(n48412), .Z(n46509) );
  XOR U51585 ( .A(round_reg[271]), .B(n51346), .Z(n48412) );
  ANDN U51586 ( .B(n51231), .A(n51057), .Z(n51693) );
  XOR U51587 ( .A(round_reg[1115]), .B(n51694), .Z(n51057) );
  XNOR U51588 ( .A(round_reg[1504]), .B(n51161), .Z(n51231) );
  XNOR U51589 ( .A(n51695), .B(n48425), .Z(n46670) );
  XNOR U51590 ( .A(round_reg[164]), .B(n48449), .Z(n48425) );
  ANDN U51591 ( .B(n51228), .A(n51059), .Z(n51695) );
  XOR U51592 ( .A(round_reg[973]), .B(n51696), .Z(n51059) );
  XNOR U51593 ( .A(round_reg[1349]), .B(n49074), .Z(n51228) );
  XNOR U51594 ( .A(n51697), .B(n51220), .Z(n51475) );
  XNOR U51595 ( .A(round_reg[467]), .B(n49904), .Z(n51220) );
  IV U51596 ( .A(n51698), .Z(n49904) );
  NOR U51597 ( .A(n48035), .B(n50582), .Z(n51697) );
  XNOR U51598 ( .A(round_reg[106]), .B(n51688), .Z(n50582) );
  XNOR U51599 ( .A(round_reg[1287]), .B(n51699), .Z(n48035) );
  AND U51600 ( .A(n42857), .B(n41941), .Z(n51667) );
  XOR U51601 ( .A(n47985), .B(n50694), .Z(n41941) );
  XOR U51602 ( .A(n49063), .B(n46884), .Z(n50694) );
  XOR U51603 ( .A(n51700), .B(n51701), .Z(n46884) );
  XNOR U51604 ( .A(n45362), .B(n43087), .Z(n51701) );
  XOR U51605 ( .A(n51702), .B(n49720), .Z(n43087) );
  XOR U51606 ( .A(round_reg[127]), .B(n51703), .Z(n49720) );
  ANDN U51607 ( .B(n50692), .A(n50301), .Z(n51702) );
  XOR U51608 ( .A(round_reg[1235]), .B(n50480), .Z(n50301) );
  XOR U51609 ( .A(round_reg[1308]), .B(n48965), .Z(n50692) );
  XOR U51610 ( .A(n51704), .B(n51320), .Z(n45362) );
  XOR U51611 ( .A(round_reg[41]), .B(n51006), .Z(n51320) );
  XNOR U51612 ( .A(n44934), .B(n51705), .Z(n51700) );
  XOR U51613 ( .A(n48192), .B(n43849), .Z(n51705) );
  XNOR U51614 ( .A(n51706), .B(n49712), .Z(n43849) );
  XNOR U51615 ( .A(round_reg[293]), .B(n51707), .Z(n49712) );
  ANDN U51616 ( .B(n47980), .A(n47981), .Z(n51706) );
  XOR U51617 ( .A(round_reg[1137]), .B(n51708), .Z(n47981) );
  XOR U51618 ( .A(round_reg[1526]), .B(n50234), .Z(n47980) );
  XNOR U51619 ( .A(n51709), .B(n49717), .Z(n48192) );
  XNOR U51620 ( .A(round_reg[186]), .B(n51620), .Z(n49717) );
  ANDN U51621 ( .B(n47976), .A(n47977), .Z(n51709) );
  IV U51622 ( .A(n50297), .Z(n47977) );
  XOR U51623 ( .A(round_reg[995]), .B(n51533), .Z(n50297) );
  XNOR U51624 ( .A(round_reg[1371]), .B(n50485), .Z(n47976) );
  IV U51625 ( .A(n51710), .Z(n50485) );
  XOR U51626 ( .A(n51711), .B(n51314), .Z(n44934) );
  XOR U51627 ( .A(round_reg[245]), .B(n51679), .Z(n51314) );
  AND U51628 ( .A(n47989), .B(n47987), .Z(n51711) );
  XNOR U51629 ( .A(round_reg[1465]), .B(n50449), .Z(n47987) );
  XNOR U51630 ( .A(round_reg[1024]), .B(n50407), .Z(n47989) );
  XOR U51631 ( .A(n51712), .B(n51713), .Z(n49063) );
  XNOR U51632 ( .A(n45313), .B(n45558), .Z(n51713) );
  XNOR U51633 ( .A(n51714), .B(n51715), .Z(n45558) );
  NOR U51634 ( .A(n48131), .B(n48129), .Z(n51714) );
  XOR U51635 ( .A(round_reg[589]), .B(n51093), .Z(n48131) );
  XNOR U51636 ( .A(n51716), .B(n51251), .Z(n45313) );
  NOR U51637 ( .A(n51717), .B(n49067), .Z(n51716) );
  XOR U51638 ( .A(round_reg[366]), .B(n50718), .Z(n49067) );
  XNOR U51639 ( .A(n51718), .B(n51719), .Z(n51712) );
  XNOR U51640 ( .A(n45153), .B(n42674), .Z(n51719) );
  XNOR U51641 ( .A(n51720), .B(n51254), .Z(n42674) );
  NOR U51642 ( .A(n48142), .B(n48143), .Z(n51720) );
  XNOR U51643 ( .A(round_reg[521]), .B(n51721), .Z(n48143) );
  XNOR U51644 ( .A(n51722), .B(n51244), .Z(n45153) );
  ANDN U51645 ( .B(n48138), .A(n48139), .Z(n51722) );
  XOR U51646 ( .A(round_reg[487]), .B(n51723), .Z(n48139) );
  XNOR U51647 ( .A(n51724), .B(n51319), .Z(n47985) );
  XNOR U51648 ( .A(round_reg[1591]), .B(n51725), .Z(n51319) );
  ANDN U51649 ( .B(n50304), .A(n50303), .Z(n51724) );
  XOR U51650 ( .A(round_reg[1163]), .B(n50758), .Z(n50303) );
  IV U51651 ( .A(n51726), .Z(n50758) );
  XOR U51652 ( .A(round_reg[780]), .B(n51727), .Z(n50304) );
  XNOR U51653 ( .A(n48976), .B(n42206), .Z(n42857) );
  XNOR U51654 ( .A(n47320), .B(n51728), .Z(n42206) );
  XOR U51655 ( .A(n51729), .B(n51730), .Z(n47320) );
  XNOR U51656 ( .A(n45742), .B(n47931), .Z(n51730) );
  XNOR U51657 ( .A(n51731), .B(n50675), .Z(n47931) );
  NOR U51658 ( .A(n49196), .B(n50674), .Z(n51731) );
  XOR U51659 ( .A(n51732), .B(n50679), .Z(n45742) );
  ANDN U51660 ( .B(n50678), .A(n51733), .Z(n51732) );
  XNOR U51661 ( .A(n45420), .B(n51734), .Z(n51729) );
  XNOR U51662 ( .A(n47697), .B(n42324), .Z(n51734) );
  XNOR U51663 ( .A(n51735), .B(n50686), .Z(n42324) );
  ANDN U51664 ( .B(n50687), .A(n51736), .Z(n51735) );
  XOR U51665 ( .A(n51737), .B(n50682), .Z(n47697) );
  ANDN U51666 ( .B(n50683), .A(n49185), .Z(n51737) );
  XOR U51667 ( .A(n51738), .B(n50689), .Z(n45420) );
  ANDN U51668 ( .B(n50690), .A(n49189), .Z(n51738) );
  XNOR U51669 ( .A(n51739), .B(n51740), .Z(n48976) );
  ANDN U51670 ( .B(n46617), .A(n46618), .Z(n51739) );
  XOR U51671 ( .A(n35368), .B(n51741), .Z(n51583) );
  XOR U51672 ( .A(n38976), .B(n40327), .Z(n51741) );
  XOR U51673 ( .A(n51742), .B(n41796), .Z(n40327) );
  XOR U51674 ( .A(n46164), .B(n46839), .Z(n41796) );
  XNOR U51675 ( .A(n51743), .B(n51744), .Z(n46839) );
  ANDN U51676 ( .B(n51745), .A(n51273), .Z(n51743) );
  XOR U51677 ( .A(n49809), .B(n51746), .Z(n46164) );
  XOR U51678 ( .A(n51747), .B(n51748), .Z(n49809) );
  XNOR U51679 ( .A(n43564), .B(n46529), .Z(n51748) );
  XNOR U51680 ( .A(n51749), .B(n49514), .Z(n46529) );
  XOR U51681 ( .A(round_reg[798]), .B(n50650), .Z(n49514) );
  NOR U51682 ( .A(n48787), .B(n48785), .Z(n51749) );
  XOR U51683 ( .A(round_reg[436]), .B(n48559), .Z(n48785) );
  IV U51684 ( .A(n49623), .Z(n48559) );
  XOR U51685 ( .A(n51750), .B(n51751), .Z(n49623) );
  XNOR U51686 ( .A(n51752), .B(n49522), .Z(n43564) );
  XNOR U51687 ( .A(round_reg[752]), .B(n49178), .Z(n49522) );
  ANDN U51688 ( .B(n48791), .A(n48789), .Z(n51752) );
  XNOR U51689 ( .A(round_reg[321]), .B(n51347), .Z(n48789) );
  XNOR U51690 ( .A(n47068), .B(n51753), .Z(n51747) );
  XOR U51691 ( .A(n48492), .B(n43783), .Z(n51753) );
  XNOR U51692 ( .A(n51754), .B(n49590), .Z(n43783) );
  XOR U51693 ( .A(round_reg[674]), .B(n49075), .Z(n49590) );
  NOR U51694 ( .A(n49819), .B(n49589), .Z(n51754) );
  XNOR U51695 ( .A(round_reg[608]), .B(n49860), .Z(n49589) );
  XNOR U51696 ( .A(n51755), .B(n49519), .Z(n48492) );
  XNOR U51697 ( .A(round_reg[895]), .B(n48520), .Z(n49519) );
  NOR U51698 ( .A(n48781), .B(n48780), .Z(n51755) );
  XOR U51699 ( .A(round_reg[506]), .B(n51620), .Z(n48780) );
  XNOR U51700 ( .A(n51756), .B(n49511), .Z(n47068) );
  XOR U51701 ( .A(round_reg[902]), .B(n50815), .Z(n49511) );
  ANDN U51702 ( .B(n48793), .A(n48794), .Z(n51756) );
  XNOR U51703 ( .A(round_reg[540]), .B(n50635), .Z(n48793) );
  AND U51704 ( .A(n39573), .B(n42861), .Z(n51742) );
  XNOR U51705 ( .A(n44663), .B(n47047), .Z(n42861) );
  XOR U51706 ( .A(n51757), .B(n51758), .Z(n47047) );
  ANDN U51707 ( .B(n49987), .A(n48394), .Z(n51757) );
  XNOR U51708 ( .A(round_reg[248]), .B(n50427), .Z(n48394) );
  XOR U51709 ( .A(n50698), .B(n46892), .Z(n44663) );
  XOR U51710 ( .A(n51759), .B(n51760), .Z(n46892) );
  XOR U51711 ( .A(n44559), .B(n51761), .Z(n51760) );
  XNOR U51712 ( .A(n51762), .B(n48392), .Z(n44559) );
  NOR U51713 ( .A(n47054), .B(n47053), .Z(n51762) );
  XOR U51714 ( .A(round_reg[421]), .B(n49901), .Z(n47054) );
  XOR U51715 ( .A(n46085), .B(n51765), .Z(n51759) );
  XOR U51716 ( .A(n43957), .B(n51766), .Z(n51765) );
  XNOR U51717 ( .A(n51767), .B(n48396), .Z(n43957) );
  NOR U51718 ( .A(n49987), .B(n51758), .Z(n51767) );
  XNOR U51719 ( .A(round_reg[593]), .B(n51664), .Z(n49987) );
  XNOR U51720 ( .A(n51768), .B(n48984), .Z(n46085) );
  NOR U51721 ( .A(n47039), .B(n47040), .Z(n51768) );
  XNOR U51722 ( .A(round_reg[370]), .B(n50404), .Z(n47040) );
  IV U51723 ( .A(n51769), .Z(n47039) );
  XOR U51724 ( .A(n51770), .B(n51771), .Z(n50698) );
  XNOR U51725 ( .A(n46976), .B(n46119), .Z(n51771) );
  XOR U51726 ( .A(n51772), .B(n51636), .Z(n46119) );
  NOR U51727 ( .A(n48828), .B(n48830), .Z(n51772) );
  XOR U51728 ( .A(round_reg[1593]), .B(n51773), .Z(n48830) );
  XOR U51729 ( .A(n51774), .B(n51633), .Z(n46976) );
  NOR U51730 ( .A(n49680), .B(n50696), .Z(n51774) );
  IV U51731 ( .A(n50697), .Z(n49680) );
  XOR U51732 ( .A(round_reg[1528]), .B(n50427), .Z(n50697) );
  XOR U51733 ( .A(n46308), .B(n51775), .Z(n51770) );
  XOR U51734 ( .A(n46801), .B(n47251), .Z(n51775) );
  XOR U51735 ( .A(n51776), .B(n51631), .Z(n47251) );
  NOR U51736 ( .A(n48825), .B(n48824), .Z(n51776) );
  IV U51737 ( .A(n49677), .Z(n48825) );
  XOR U51738 ( .A(round_reg[1467]), .B(n51618), .Z(n49677) );
  XNOR U51739 ( .A(n51777), .B(n51638), .Z(n46801) );
  NOR U51740 ( .A(n49685), .B(n48819), .Z(n51777) );
  IV U51741 ( .A(n48821), .Z(n49685) );
  XOR U51742 ( .A(round_reg[1310]), .B(n49633), .Z(n48821) );
  IV U51743 ( .A(n49797), .Z(n49633) );
  XOR U51744 ( .A(n51778), .B(n51779), .Z(n49797) );
  XOR U51745 ( .A(n51780), .B(n51641), .Z(n46308) );
  NOR U51746 ( .A(n49688), .B(n48832), .Z(n51780) );
  IV U51747 ( .A(n48834), .Z(n49688) );
  XOR U51748 ( .A(round_reg[1373]), .B(n51781), .Z(n48834) );
  XNOR U51749 ( .A(n51502), .B(n45358), .Z(n39573) );
  XOR U51750 ( .A(n48886), .B(n48773), .Z(n45358) );
  XOR U51751 ( .A(n51782), .B(n51783), .Z(n48773) );
  XNOR U51752 ( .A(n45741), .B(n46682), .Z(n51783) );
  XOR U51753 ( .A(n51784), .B(n51431), .Z(n46682) );
  XOR U51754 ( .A(round_reg[12]), .B(n50933), .Z(n51431) );
  NOR U51755 ( .A(n51438), .B(n50798), .Z(n51784) );
  XOR U51756 ( .A(round_reg[1198]), .B(n51333), .Z(n50798) );
  XOR U51757 ( .A(round_reg[1562]), .B(n49625), .Z(n51438) );
  XNOR U51758 ( .A(n51785), .B(n51426), .Z(n45741) );
  IV U51759 ( .A(n48997), .Z(n51426) );
  XNOR U51760 ( .A(round_reg[216]), .B(n49789), .Z(n48997) );
  NOR U51761 ( .A(n48996), .B(n50791), .Z(n51785) );
  XOR U51762 ( .A(round_reg[1059]), .B(n51624), .Z(n50791) );
  IV U51763 ( .A(n51514), .Z(n48996) );
  XOR U51764 ( .A(round_reg[1436]), .B(n50827), .Z(n51514) );
  XOR U51765 ( .A(n45623), .B(n51786), .Z(n51782) );
  XOR U51766 ( .A(n43593), .B(n45334), .Z(n51786) );
  XNOR U51767 ( .A(n51787), .B(n49003), .Z(n45334) );
  XOR U51768 ( .A(round_reg[264]), .B(n51788), .Z(n49003) );
  NOR U51769 ( .A(n49002), .B(n50794), .Z(n51787) );
  XOR U51770 ( .A(round_reg[1108]), .B(n51789), .Z(n50794) );
  IV U51771 ( .A(n51511), .Z(n49002) );
  XOR U51772 ( .A(round_reg[1497]), .B(n51790), .Z(n51511) );
  XOR U51773 ( .A(n51791), .B(n48993), .Z(n43593) );
  XOR U51774 ( .A(round_reg[98]), .B(n50745), .Z(n48993) );
  XOR U51775 ( .A(round_reg[1270]), .B(n50106), .Z(n50802) );
  XOR U51776 ( .A(round_reg[1343]), .B(n48879), .Z(n48992) );
  XNOR U51777 ( .A(n51792), .B(n49007), .Z(n45623) );
  NOR U51778 ( .A(n49006), .B(n50805), .Z(n51792) );
  XOR U51779 ( .A(round_reg[966]), .B(n50643), .Z(n50805) );
  XOR U51780 ( .A(round_reg[1406]), .B(n51793), .Z(n49006) );
  XOR U51781 ( .A(n51794), .B(n51795), .Z(n48886) );
  XOR U51782 ( .A(n44838), .B(n48547), .Z(n51795) );
  XOR U51783 ( .A(n51796), .B(n50318), .Z(n48547) );
  NOR U51784 ( .A(n50317), .B(n47220), .Z(n51796) );
  XNOR U51785 ( .A(round_reg[217]), .B(n50508), .Z(n47220) );
  XOR U51786 ( .A(round_reg[626]), .B(n51141), .Z(n50317) );
  XNOR U51787 ( .A(n51797), .B(n50311), .Z(n44838) );
  NOR U51788 ( .A(n49698), .B(n50310), .Z(n51797) );
  XOR U51789 ( .A(round_reg[339]), .B(n51685), .Z(n50310) );
  IV U51790 ( .A(n49181), .Z(n51685) );
  XOR U51791 ( .A(round_reg[265]), .B(n51462), .Z(n49698) );
  XOR U51792 ( .A(n48986), .B(n51798), .Z(n51794) );
  XOR U51793 ( .A(n45264), .B(n45958), .Z(n51798) );
  NOR U51794 ( .A(n51800), .B(n50324), .Z(n51799) );
  IV U51795 ( .A(n51494), .Z(n51800) );
  XNOR U51796 ( .A(n51801), .B(n50321), .Z(n45264) );
  AND U51797 ( .A(n47226), .B(n50320), .Z(n51801) );
  XOR U51798 ( .A(round_reg[460]), .B(n51579), .Z(n50320) );
  XNOR U51799 ( .A(round_reg[99]), .B(n51624), .Z(n47226) );
  XOR U51800 ( .A(n51802), .B(n50314), .Z(n48986) );
  XNOR U51801 ( .A(round_reg[158]), .B(n50650), .Z(n47230) );
  XOR U51802 ( .A(round_reg[558]), .B(n51333), .Z(n50313) );
  XNOR U51803 ( .A(n51803), .B(n50324), .Z(n51502) );
  XOR U51804 ( .A(round_reg[390]), .B(n49271), .Z(n50324) );
  NOR U51805 ( .A(n51494), .B(n51495), .Z(n51803) );
  XOR U51806 ( .A(round_reg[13]), .B(n50752), .Z(n51494) );
  XOR U51807 ( .A(n51804), .B(n41794), .Z(n38976) );
  XOR U51808 ( .A(n49194), .B(n45646), .Z(n41794) );
  XNOR U51809 ( .A(n51805), .B(n51736), .Z(n49194) );
  AND U51810 ( .A(n42853), .B(n41615), .Z(n51804) );
  XNOR U51811 ( .A(n51379), .B(n45915), .Z(n41615) );
  IV U51812 ( .A(n44337), .Z(n45915) );
  XOR U51813 ( .A(n46497), .B(n50144), .Z(n44337) );
  XNOR U51814 ( .A(n51807), .B(n51808), .Z(n50144) );
  XOR U51815 ( .A(n44669), .B(n46098), .Z(n51808) );
  XOR U51816 ( .A(n51809), .B(n47227), .Z(n46098) );
  XNOR U51817 ( .A(round_reg[1280]), .B(n50457), .Z(n47227) );
  ANDN U51818 ( .B(n47228), .A(n50321), .Z(n51809) );
  XOR U51819 ( .A(round_reg[849]), .B(n49898), .Z(n50321) );
  XOR U51820 ( .A(round_reg[1271]), .B(n51810), .Z(n47228) );
  XNOR U51821 ( .A(n51811), .B(n47232), .Z(n44669) );
  XOR U51822 ( .A(round_reg[1407]), .B(n51703), .Z(n47232) );
  ANDN U51823 ( .B(n50314), .A(n47231), .Z(n51811) );
  XOR U51824 ( .A(round_reg[967]), .B(n51699), .Z(n47231) );
  XOR U51825 ( .A(round_reg[920]), .B(n51812), .Z(n50314) );
  XOR U51826 ( .A(n45468), .B(n51813), .Z(n51807) );
  XOR U51827 ( .A(n45658), .B(n43845), .Z(n51813) );
  XNOR U51828 ( .A(n51814), .B(n49699), .Z(n43845) );
  XOR U51829 ( .A(round_reg[1498]), .B(n50814), .Z(n49699) );
  ANDN U51830 ( .B(n49700), .A(n50311), .Z(n51814) );
  XNOR U51831 ( .A(round_reg[706]), .B(n49989), .Z(n50311) );
  XOR U51832 ( .A(round_reg[1109]), .B(n50232), .Z(n49700) );
  XNOR U51833 ( .A(n51815), .B(n47221), .Z(n45658) );
  XNOR U51834 ( .A(round_reg[1437]), .B(n48517), .Z(n47221) );
  ANDN U51835 ( .B(n47222), .A(n50318), .Z(n51815) );
  XOR U51836 ( .A(round_reg[692]), .B(n50440), .Z(n50318) );
  XOR U51837 ( .A(round_reg[1060]), .B(n51816), .Z(n47222) );
  XNOR U51838 ( .A(n51817), .B(n51495), .Z(n45468) );
  XOR U51839 ( .A(round_reg[1563]), .B(n51009), .Z(n51495) );
  ANDN U51840 ( .B(n50325), .A(n51496), .Z(n51817) );
  XNOR U51841 ( .A(round_reg[1199]), .B(n51172), .Z(n51496) );
  XOR U51842 ( .A(round_reg[816]), .B(n51818), .Z(n50325) );
  XOR U51843 ( .A(n51819), .B(n51820), .Z(n46497) );
  XOR U51844 ( .A(n45779), .B(n47214), .Z(n51820) );
  XOR U51845 ( .A(n51821), .B(n50921), .Z(n47214) );
  ANDN U51846 ( .B(n51381), .A(n48896), .Z(n51821) );
  XOR U51847 ( .A(round_reg[1281]), .B(n51347), .Z(n48896) );
  XNOR U51848 ( .A(n51822), .B(n50924), .Z(n45779) );
  NOR U51849 ( .A(n51374), .B(n48900), .Z(n51822) );
  XNOR U51850 ( .A(round_reg[1438]), .B(n50650), .Z(n48900) );
  IV U51851 ( .A(n51823), .Z(n51374) );
  XOR U51852 ( .A(n46937), .B(n51824), .Z(n51819) );
  XOR U51853 ( .A(n46703), .B(n45553), .Z(n51824) );
  XOR U51854 ( .A(n51825), .B(n50928), .Z(n45553) );
  ANDN U51855 ( .B(n50327), .A(n51826), .Z(n51825) );
  XOR U51856 ( .A(n51827), .B(n50919), .Z(n46703) );
  ANDN U51857 ( .B(n51383), .A(n48904), .Z(n51827) );
  XNOR U51858 ( .A(round_reg[1499]), .B(n50131), .Z(n48904) );
  XNOR U51859 ( .A(n51828), .B(n50926), .Z(n46937) );
  ANDN U51860 ( .B(n51376), .A(n48891), .Z(n51828) );
  XOR U51861 ( .A(round_reg[1344]), .B(n50407), .Z(n48891) );
  XNOR U51862 ( .A(n51829), .B(n51830), .Z(n50407) );
  XNOR U51863 ( .A(n51831), .B(n51826), .Z(n51379) );
  ANDN U51864 ( .B(n50328), .A(n50327), .Z(n51831) );
  XOR U51865 ( .A(round_reg[1564]), .B(n49261), .Z(n50327) );
  XOR U51866 ( .A(round_reg[1200]), .B(n48938), .Z(n50328) );
  XOR U51867 ( .A(n45781), .B(n47488), .Z(n42853) );
  XNOR U51868 ( .A(n51832), .B(n49911), .Z(n47488) );
  IV U51869 ( .A(n45481), .Z(n45781) );
  XOR U51870 ( .A(n51833), .B(n49997), .Z(n45481) );
  XOR U51871 ( .A(n51834), .B(n51835), .Z(n49997) );
  XOR U51872 ( .A(n45261), .B(n43961), .Z(n51835) );
  XNOR U51873 ( .A(n51836), .B(n49910), .Z(n43961) );
  ANDN U51874 ( .B(n49911), .A(n50085), .Z(n51836) );
  XOR U51875 ( .A(round_reg[253]), .B(n51837), .Z(n50085) );
  XOR U51876 ( .A(round_reg[598]), .B(n50397), .Z(n49911) );
  XNOR U51877 ( .A(n51838), .B(n49390), .Z(n45261) );
  ANDN U51878 ( .B(n48462), .A(n48464), .Z(n51838) );
  XOR U51879 ( .A(round_reg[301]), .B(n51839), .Z(n48464) );
  XOR U51880 ( .A(round_reg[375]), .B(n50507), .Z(n48462) );
  XNOR U51881 ( .A(n44941), .B(n51840), .Z(n51834) );
  XNOR U51882 ( .A(n46822), .B(n41746), .Z(n51840) );
  XNOR U51883 ( .A(n51841), .B(n51842), .Z(n41746) );
  NOR U51884 ( .A(n46987), .B(n47486), .Z(n51841) );
  XOR U51885 ( .A(round_reg[49]), .B(n50498), .Z(n47486) );
  XOR U51886 ( .A(round_reg[426]), .B(n50819), .Z(n46987) );
  IV U51887 ( .A(n51688), .Z(n50819) );
  XOR U51888 ( .A(n51843), .B(n51844), .Z(n51688) );
  XOR U51889 ( .A(n51845), .B(n51846), .Z(n46822) );
  ANDN U51890 ( .B(n46995), .A(n50080), .Z(n51845) );
  XOR U51891 ( .A(round_reg[71]), .B(n51847), .Z(n50080) );
  XNOR U51892 ( .A(round_reg[496]), .B(n51818), .Z(n46995) );
  XOR U51893 ( .A(n51848), .B(n46984), .Z(n44941) );
  ANDN U51894 ( .B(n46983), .A(n50088), .Z(n51848) );
  XOR U51895 ( .A(round_reg[130]), .B(n50455), .Z(n50088) );
  IV U51896 ( .A(n51564), .Z(n50455) );
  XNOR U51897 ( .A(round_reg[530]), .B(n50475), .Z(n46983) );
  XNOR U51898 ( .A(n51849), .B(n41787), .Z(n35368) );
  XOR U51899 ( .A(n49952), .B(n46071), .Z(n41787) );
  XOR U51900 ( .A(n51400), .B(n50639), .Z(n46071) );
  XNOR U51901 ( .A(n51850), .B(n51851), .Z(n50639) );
  XNOR U51902 ( .A(n45627), .B(n45361), .Z(n51851) );
  XNOR U51903 ( .A(n51852), .B(n49373), .Z(n45361) );
  XNOR U51904 ( .A(n51853), .B(n49534), .Z(n45627) );
  ANDN U51905 ( .B(n49962), .A(n49963), .Z(n51853) );
  XOR U51906 ( .A(n47241), .B(n51854), .Z(n51850) );
  XOR U51907 ( .A(n45302), .B(n48306), .Z(n51854) );
  XNOR U51908 ( .A(n51855), .B(n49366), .Z(n48306) );
  ANDN U51909 ( .B(n50637), .A(n50638), .Z(n51855) );
  XNOR U51910 ( .A(n51856), .B(n51857), .Z(n45302) );
  XNOR U51911 ( .A(n51858), .B(n49362), .Z(n47241) );
  XOR U51912 ( .A(n51859), .B(n51860), .Z(n51400) );
  XOR U51913 ( .A(n46503), .B(n45901), .Z(n51860) );
  XOR U51914 ( .A(n51861), .B(n49662), .Z(n45901) );
  ANDN U51915 ( .B(n49957), .A(n48673), .Z(n51861) );
  XOR U51916 ( .A(round_reg[1583]), .B(n50414), .Z(n48673) );
  XNOR U51917 ( .A(n51862), .B(n49671), .Z(n46503) );
  ANDN U51918 ( .B(n49946), .A(n48683), .Z(n51862) );
  XOR U51919 ( .A(round_reg[1518]), .B(n51333), .Z(n48683) );
  XOR U51920 ( .A(n51863), .B(n51864), .Z(n51859) );
  XOR U51921 ( .A(n46082), .B(n51865), .Z(n51864) );
  XNOR U51922 ( .A(n51866), .B(n49665), .Z(n46082) );
  ANDN U51923 ( .B(n51867), .A(n48679), .Z(n51866) );
  XNOR U51924 ( .A(n51868), .B(n51867), .Z(n49952) );
  ANDN U51925 ( .B(n48679), .A(n48680), .Z(n51868) );
  XNOR U51926 ( .A(round_reg[1227]), .B(n51647), .Z(n48680) );
  XNOR U51927 ( .A(round_reg[1300]), .B(n50742), .Z(n48679) );
  AND U51928 ( .A(n39566), .B(n42848), .Z(n51849) );
  XNOR U51929 ( .A(n51869), .B(n42848), .Z(n45572) );
  XNOR U51930 ( .A(n47447), .B(n51870), .Z(n42848) );
  IV U51931 ( .A(n43899), .Z(n47447) );
  XOR U51932 ( .A(n47107), .B(n48883), .Z(n43899) );
  XNOR U51933 ( .A(n51871), .B(n51872), .Z(n48883) );
  XOR U51934 ( .A(n45657), .B(n44699), .Z(n51872) );
  XOR U51935 ( .A(n51873), .B(n49889), .Z(n44699) );
  XOR U51936 ( .A(round_reg[23]), .B(n48554), .Z(n49889) );
  ANDN U51937 ( .B(n51874), .A(n49888), .Z(n51873) );
  XNOR U51938 ( .A(n51875), .B(n48258), .Z(n45657) );
  XOR U51939 ( .A(round_reg[109]), .B(n50432), .Z(n48258) );
  NOR U51940 ( .A(n48257), .B(n51876), .Z(n51875) );
  XOR U51941 ( .A(n47836), .B(n51877), .Z(n51871) );
  XOR U51942 ( .A(n43561), .B(n48244), .Z(n51877) );
  XNOR U51943 ( .A(n51878), .B(n48251), .Z(n48244) );
  XOR U51944 ( .A(round_reg[275]), .B(n50480), .Z(n48251) );
  AND U51945 ( .A(n51879), .B(n48252), .Z(n51878) );
  XNOR U51946 ( .A(n51880), .B(n48262), .Z(n43561) );
  XOR U51947 ( .A(round_reg[227]), .B(n48450), .Z(n48262) );
  NOR U51948 ( .A(n48261), .B(n51881), .Z(n51880) );
  XNOR U51949 ( .A(n51882), .B(n50204), .Z(n47836) );
  XNOR U51950 ( .A(round_reg[168]), .B(n51883), .Z(n50204) );
  ANDN U51951 ( .B(n50215), .A(n51884), .Z(n51882) );
  XOR U51952 ( .A(n51885), .B(n51886), .Z(n47107) );
  XOR U51953 ( .A(n45637), .B(n51887), .Z(n51886) );
  XNOR U51954 ( .A(n51888), .B(n51889), .Z(n45637) );
  ANDN U51955 ( .B(n51890), .A(n48067), .Z(n51888) );
  XOR U51956 ( .A(n42300), .B(n51891), .Z(n51885) );
  XOR U51957 ( .A(n42317), .B(n47470), .Z(n51891) );
  XNOR U51958 ( .A(n51892), .B(n51893), .Z(n47470) );
  NOR U51959 ( .A(n48063), .B(n51894), .Z(n51892) );
  XNOR U51960 ( .A(n51895), .B(n51896), .Z(n42317) );
  ANDN U51961 ( .B(n51897), .A(n48077), .Z(n51895) );
  XNOR U51962 ( .A(n51898), .B(n51899), .Z(n42300) );
  ANDN U51963 ( .B(n51900), .A(n48073), .Z(n51898) );
  NOR U51964 ( .A(n39567), .B(n39566), .Z(n51869) );
  XNOR U51965 ( .A(n45154), .B(n51718), .Z(n39566) );
  XOR U51966 ( .A(n51901), .B(n51256), .Z(n51718) );
  NOR U51967 ( .A(n51902), .B(n48135), .Z(n51901) );
  XNOR U51968 ( .A(round_reg[417]), .B(n49089), .Z(n48135) );
  XOR U51969 ( .A(n49543), .B(n48194), .Z(n45154) );
  XOR U51970 ( .A(n51903), .B(n51904), .Z(n48194) );
  XOR U51971 ( .A(n46505), .B(n51239), .Z(n51904) );
  XOR U51972 ( .A(n51905), .B(n49341), .Z(n51239) );
  XOR U51973 ( .A(round_reg[1590]), .B(n50106), .Z(n49341) );
  ANDN U51974 ( .B(n51256), .A(n48134), .Z(n51905) );
  IV U51975 ( .A(n51902), .Z(n48134) );
  XOR U51976 ( .A(round_reg[779]), .B(n50138), .Z(n51902) );
  XOR U51977 ( .A(round_reg[1162]), .B(n50852), .Z(n51256) );
  XNOR U51978 ( .A(n51906), .B(n49336), .Z(n46505) );
  XNOR U51979 ( .A(round_reg[1464]), .B(n51907), .Z(n49336) );
  ANDN U51980 ( .B(n48129), .A(n51715), .Z(n51906) );
  IV U51981 ( .A(n51247), .Z(n51715) );
  XOR U51982 ( .A(round_reg[1087]), .B(n51703), .Z(n51247) );
  XNOR U51983 ( .A(round_reg[655]), .B(n48362), .Z(n48129) );
  XOR U51984 ( .A(n46281), .B(n51908), .Z(n51903) );
  XOR U51985 ( .A(n51035), .B(n47840), .Z(n51908) );
  XOR U51986 ( .A(n51909), .B(n49343), .Z(n47840) );
  XNOR U51987 ( .A(round_reg[1525]), .B(n51679), .Z(n49343) );
  NOR U51988 ( .A(n49066), .B(n51251), .Z(n51909) );
  IV U51989 ( .A(n51717), .Z(n49066) );
  XOR U51990 ( .A(round_reg[733]), .B(n51781), .Z(n51717) );
  XNOR U51991 ( .A(n51910), .B(n49339), .Z(n51035) );
  XOR U51992 ( .A(round_reg[1307]), .B(n49955), .Z(n49339) );
  ANDN U51993 ( .B(n51244), .A(n48138), .Z(n51910) );
  XOR U51994 ( .A(round_reg[876]), .B(n51911), .Z(n48138) );
  XOR U51995 ( .A(round_reg[1234]), .B(n50755), .Z(n51244) );
  XNOR U51996 ( .A(n51912), .B(n49334), .Z(n46281) );
  XOR U51997 ( .A(round_reg[1370]), .B(n51468), .Z(n49334) );
  ANDN U51998 ( .B(n48142), .A(n51254), .Z(n51912) );
  XOR U51999 ( .A(round_reg[994]), .B(n49075), .Z(n51254) );
  XOR U52000 ( .A(round_reg[947]), .B(n50504), .Z(n48142) );
  XOR U52001 ( .A(n51913), .B(n51914), .Z(n49543) );
  XOR U52002 ( .A(n46087), .B(n50960), .Z(n51914) );
  XOR U52003 ( .A(n51915), .B(n51266), .Z(n50960) );
  XOR U52004 ( .A(round_reg[732]), .B(n51617), .Z(n51266) );
  ANDN U52005 ( .B(n50196), .A(n50180), .Z(n51915) );
  XOR U52006 ( .A(round_reg[291]), .B(n48872), .Z(n50180) );
  IV U52007 ( .A(n48701), .Z(n48872) );
  XNOR U52008 ( .A(round_reg[365]), .B(n50120), .Z(n50196) );
  XNOR U52009 ( .A(n51918), .B(n51268), .Z(n46087) );
  XOR U52010 ( .A(round_reg[875]), .B(n51528), .Z(n51268) );
  ANDN U52011 ( .B(n50192), .A(n48149), .Z(n51918) );
  XOR U52012 ( .A(round_reg[486]), .B(n51547), .Z(n50192) );
  XOR U52013 ( .A(n43554), .B(n51919), .Z(n51913) );
  XOR U52014 ( .A(n44561), .B(n43471), .Z(n51919) );
  XNOR U52015 ( .A(n51920), .B(n51643), .Z(n43471) );
  XNOR U52016 ( .A(round_reg[654]), .B(n50765), .Z(n51643) );
  AND U52017 ( .A(n48155), .B(n50189), .Z(n51920) );
  XNOR U52018 ( .A(round_reg[588]), .B(n49427), .Z(n50189) );
  XOR U52019 ( .A(round_reg[243]), .B(n50966), .Z(n48155) );
  XNOR U52020 ( .A(n51923), .B(n51262), .Z(n44561) );
  XNOR U52021 ( .A(round_reg[946]), .B(n51141), .Z(n51262) );
  ANDN U52022 ( .B(n50187), .A(n49349), .Z(n51923) );
  XOR U52023 ( .A(round_reg[184]), .B(n50838), .Z(n49349) );
  IV U52024 ( .A(n51907), .Z(n50838) );
  XOR U52025 ( .A(round_reg[520]), .B(n50947), .Z(n50187) );
  XNOR U52026 ( .A(n51926), .B(n51370), .Z(n43554) );
  XOR U52027 ( .A(round_reg[778]), .B(n50117), .Z(n51370) );
  ANDN U52028 ( .B(n50194), .A(n48159), .Z(n51926) );
  XOR U52029 ( .A(round_reg[39]), .B(n51927), .Z(n48159) );
  XNOR U52030 ( .A(round_reg[416]), .B(n51928), .Z(n50194) );
  XNOR U52031 ( .A(n51175), .B(n45315), .Z(n39567) );
  XNOR U52032 ( .A(n46725), .B(n50354), .Z(n45315) );
  XOR U52033 ( .A(n51929), .B(n51930), .Z(n50354) );
  XOR U52034 ( .A(n43556), .B(n48912), .Z(n51930) );
  XOR U52035 ( .A(n51931), .B(n48105), .Z(n48912) );
  XNOR U52036 ( .A(round_reg[989]), .B(n49869), .Z(n48105) );
  NOR U52037 ( .A(n48947), .B(n48917), .Z(n51931) );
  IV U52038 ( .A(n51932), .Z(n48947) );
  XNOR U52039 ( .A(n51933), .B(n48101), .Z(n43556) );
  XNOR U52040 ( .A(round_reg[1082]), .B(n50882), .Z(n48101) );
  NOR U52041 ( .A(n48941), .B(n48924), .Z(n51933) );
  XOR U52042 ( .A(round_reg[650]), .B(n51934), .Z(n48924) );
  XOR U52043 ( .A(round_reg[584]), .B(n51788), .Z(n48941) );
  XOR U52044 ( .A(n45211), .B(n51935), .Z(n51929) );
  XOR U52045 ( .A(n44570), .B(n47328), .Z(n51935) );
  XNOR U52046 ( .A(n51936), .B(n48097), .Z(n47328) );
  XNOR U52047 ( .A(round_reg[1157]), .B(n48453), .Z(n48097) );
  XOR U52048 ( .A(n51937), .B(n51938), .Z(n48453) );
  ANDN U52049 ( .B(n48934), .A(n48919), .Z(n51936) );
  XOR U52050 ( .A(round_reg[774]), .B(n50759), .Z(n48919) );
  IV U52051 ( .A(n51201), .Z(n50759) );
  XOR U52052 ( .A(n51592), .B(n51939), .Z(n51201) );
  XOR U52053 ( .A(n51940), .B(n51941), .Z(n51592) );
  XNOR U52054 ( .A(round_reg[1349]), .B(round_reg[1029]), .Z(n51941) );
  XOR U52055 ( .A(round_reg[389]), .B(n51942), .Z(n51940) );
  XOR U52056 ( .A(round_reg[709]), .B(round_reg[69]), .Z(n51942) );
  XNOR U52057 ( .A(round_reg[412]), .B(n51617), .Z(n48934) );
  XNOR U52058 ( .A(n51943), .B(n48433), .Z(n44570) );
  XOR U52059 ( .A(round_reg[1131]), .B(n51135), .Z(n48433) );
  NOR U52060 ( .A(n48937), .B(n48926), .Z(n51943) );
  XNOR U52061 ( .A(round_reg[728]), .B(n50978), .Z(n48926) );
  XNOR U52062 ( .A(n51944), .B(n51945), .Z(n50978) );
  XOR U52063 ( .A(round_reg[361]), .B(n51006), .Z(n48937) );
  XNOR U52064 ( .A(n51946), .B(n48092), .Z(n45211) );
  XOR U52065 ( .A(round_reg[1229]), .B(n51093), .Z(n48092) );
  NOR U52066 ( .A(n48922), .B(n48944), .Z(n51946) );
  XOR U52067 ( .A(round_reg[482]), .B(n51051), .Z(n48944) );
  XOR U52068 ( .A(round_reg[871]), .B(n51947), .Z(n48922) );
  XOR U52069 ( .A(n51948), .B(n51949), .Z(n46725) );
  XOR U52070 ( .A(n49394), .B(n47990), .Z(n51949) );
  XOR U52071 ( .A(n51950), .B(n49412), .Z(n47990) );
  XNOR U52072 ( .A(round_reg[411]), .B(n51710), .Z(n49412) );
  XOR U52073 ( .A(round_reg[1584]), .B(n51953), .Z(n49655) );
  XOR U52074 ( .A(round_reg[34]), .B(n51954), .Z(n49411) );
  XNOR U52075 ( .A(n51955), .B(n50490), .Z(n49394) );
  XOR U52076 ( .A(round_reg[360]), .B(n48442), .Z(n50490) );
  ANDN U52077 ( .B(n49642), .A(n49640), .Z(n51955) );
  XOR U52078 ( .A(round_reg[286]), .B(n51486), .Z(n49640) );
  XNOR U52079 ( .A(round_reg[1519]), .B(n51172), .Z(n49642) );
  XOR U52080 ( .A(n44471), .B(n51956), .Z(n51948) );
  XNOR U52081 ( .A(n43715), .B(n45757), .Z(n51956) );
  XOR U52082 ( .A(n51957), .B(n49401), .Z(n45757) );
  XOR U52083 ( .A(round_reg[583]), .B(n48568), .Z(n49401) );
  IV U52084 ( .A(n50132), .Z(n48568) );
  XOR U52085 ( .A(round_reg[238]), .B(n51333), .Z(n49402) );
  XOR U52086 ( .A(n51958), .B(n51959), .Z(n51333) );
  XNOR U52087 ( .A(round_reg[1458]), .B(n51327), .Z(n49645) );
  XNOR U52088 ( .A(n51960), .B(n49407), .Z(n43715) );
  AND U52089 ( .A(n49648), .B(n49408), .Z(n51960) );
  XNOR U52090 ( .A(round_reg[120]), .B(n49977), .Z(n49408) );
  XOR U52091 ( .A(round_reg[1301]), .B(n51961), .Z(n49648) );
  XOR U52092 ( .A(n51962), .B(n51404), .Z(n44471) );
  XOR U52093 ( .A(round_reg[515]), .B(n49958), .Z(n51404) );
  IV U52094 ( .A(n51597), .Z(n49958) );
  XNOR U52095 ( .A(n51963), .B(n51964), .Z(n51597) );
  ANDN U52096 ( .B(n49651), .A(n49652), .Z(n51962) );
  XOR U52097 ( .A(round_reg[1364]), .B(n50645), .Z(n49652) );
  IV U52098 ( .A(n50849), .Z(n50645) );
  XOR U52099 ( .A(round_reg[179]), .B(n48942), .Z(n49651) );
  XNOR U52100 ( .A(n51965), .B(n48917), .Z(n51175) );
  XNOR U52101 ( .A(round_reg[942]), .B(n51582), .Z(n48917) );
  NOR U52102 ( .A(n51932), .B(n48103), .Z(n51965) );
  XOR U52103 ( .A(round_reg[180]), .B(n51107), .Z(n48103) );
  IV U52104 ( .A(n51185), .Z(n51107) );
  XOR U52105 ( .A(round_reg[516]), .B(n50505), .Z(n51932) );
  XOR U52106 ( .A(n41411), .B(n39099), .Z(n38841) );
  IV U52107 ( .A(n38826), .Z(n39099) );
  XOR U52108 ( .A(n39700), .B(n42122), .Z(n38826) );
  XOR U52109 ( .A(n51966), .B(n51967), .Z(n42122) );
  XNOR U52110 ( .A(n45019), .B(n38355), .Z(n51967) );
  XNOR U52111 ( .A(n51968), .B(n45024), .Z(n38355) );
  XOR U52112 ( .A(n43543), .B(n50594), .Z(n45024) );
  XNOR U52113 ( .A(n51969), .B(n50375), .Z(n50594) );
  ANDN U52114 ( .B(n51970), .A(n51971), .Z(n51969) );
  XNOR U52115 ( .A(n49113), .B(n48310), .Z(n43543) );
  XNOR U52116 ( .A(n51972), .B(n51973), .Z(n48310) );
  XOR U52117 ( .A(n47133), .B(n45663), .Z(n51973) );
  XOR U52118 ( .A(n51974), .B(n51975), .Z(n45663) );
  ANDN U52119 ( .B(n50808), .A(n50810), .Z(n51974) );
  XNOR U52120 ( .A(n51976), .B(n50374), .Z(n47133) );
  AND U52121 ( .A(n51971), .B(n50375), .Z(n51976) );
  XOR U52122 ( .A(round_reg[214]), .B(n51200), .Z(n50375) );
  XOR U52123 ( .A(n47064), .B(n51977), .Z(n51972) );
  XOR U52124 ( .A(n47235), .B(n46576), .Z(n51977) );
  XNOR U52125 ( .A(n51978), .B(n50388), .Z(n46576) );
  ANDN U52126 ( .B(n50389), .A(n50597), .Z(n51978) );
  XNOR U52127 ( .A(round_reg[10]), .B(n51934), .Z(n50389) );
  XNOR U52128 ( .A(n51979), .B(n50378), .Z(n47235) );
  ANDN U52129 ( .B(n50379), .A(n50602), .Z(n51979) );
  XNOR U52130 ( .A(round_reg[262]), .B(n50815), .Z(n50379) );
  XNOR U52131 ( .A(n51980), .B(n50384), .Z(n47064) );
  ANDN U52132 ( .B(n50385), .A(n50605), .Z(n51980) );
  XNOR U52133 ( .A(round_reg[155]), .B(n50513), .Z(n50385) );
  XOR U52134 ( .A(n51981), .B(n51982), .Z(n49113) );
  XNOR U52135 ( .A(n48319), .B(n44569), .Z(n51982) );
  XNOR U52136 ( .A(n51983), .B(n48333), .Z(n44569) );
  ANDN U52137 ( .B(n48334), .A(n48909), .Z(n51983) );
  XNOR U52138 ( .A(round_reg[916]), .B(n51984), .Z(n48909) );
  XNOR U52139 ( .A(n51986), .B(n48329), .Z(n48319) );
  XOR U52140 ( .A(round_reg[812]), .B(n48365), .Z(n46777) );
  XOR U52141 ( .A(round_reg[1195]), .B(n51528), .Z(n48330) );
  XOR U52142 ( .A(n45941), .B(n51987), .Z(n51981) );
  XOR U52143 ( .A(n45311), .B(n44224), .Z(n51987) );
  XNOR U52144 ( .A(n51988), .B(n48325), .Z(n44224) );
  AND U52145 ( .A(n46784), .B(n48326), .Z(n51988) );
  XOR U52146 ( .A(round_reg[1056]), .B(n50723), .Z(n48326) );
  IV U52147 ( .A(n51928), .Z(n50723) );
  XNOR U52148 ( .A(round_reg[688]), .B(n49856), .Z(n46784) );
  XNOR U52149 ( .A(n51989), .B(n51149), .Z(n45311) );
  ANDN U52150 ( .B(n50613), .A(n47531), .Z(n51989) );
  XOR U52151 ( .A(round_reg[845]), .B(n51343), .Z(n47531) );
  XOR U52152 ( .A(round_reg[1267]), .B(n51990), .Z(n50613) );
  XNOR U52153 ( .A(n51991), .B(n48337), .Z(n45941) );
  AND U52154 ( .A(n49600), .B(n48338), .Z(n51991) );
  XOR U52155 ( .A(round_reg[1105]), .B(n51342), .Z(n48338) );
  XOR U52156 ( .A(round_reg[766]), .B(n51793), .Z(n49600) );
  AND U52157 ( .A(n44714), .B(n44722), .Z(n51968) );
  XOR U52158 ( .A(n40840), .B(n47610), .Z(n44722) );
  XNOR U52159 ( .A(n51992), .B(n49828), .Z(n47610) );
  AND U52160 ( .A(n48182), .B(n48180), .Z(n51992) );
  XOR U52161 ( .A(round_reg[827]), .B(n51618), .Z(n48182) );
  IV U52162 ( .A(n45723), .Z(n40840) );
  XNOR U52163 ( .A(n51993), .B(n51994), .Z(n51022) );
  XOR U52164 ( .A(n45488), .B(n49822), .Z(n51994) );
  XNOR U52165 ( .A(n51995), .B(n48882), .Z(n49822) );
  XNOR U52166 ( .A(round_reg[24]), .B(n51446), .Z(n48882) );
  ANDN U52167 ( .B(n49828), .A(n48180), .Z(n51995) );
  XNOR U52168 ( .A(round_reg[1210]), .B(n49861), .Z(n48180) );
  XOR U52169 ( .A(round_reg[1574]), .B(n51341), .Z(n49828) );
  XNOR U52170 ( .A(n51996), .B(n49834), .Z(n45488) );
  XOR U52171 ( .A(round_reg[110]), .B(n51997), .Z(n49834) );
  ANDN U52172 ( .B(n47623), .A(n47621), .Z(n51996) );
  XOR U52173 ( .A(round_reg[1291]), .B(n51127), .Z(n47621) );
  XOR U52174 ( .A(round_reg[1218]), .B(n51539), .Z(n47623) );
  XNOR U52175 ( .A(n47695), .B(n51998), .Z(n51993) );
  XOR U52176 ( .A(n46569), .B(n42156), .Z(n51998) );
  XNOR U52177 ( .A(n51999), .B(n48870), .Z(n42156) );
  XOR U52178 ( .A(round_reg[276]), .B(n51984), .Z(n48870) );
  NOR U52179 ( .A(n47625), .B(n47626), .Z(n51999) );
  XNOR U52180 ( .A(round_reg[1120]), .B(n52000), .Z(n47626) );
  XOR U52181 ( .A(round_reg[1509]), .B(n52001), .Z(n47625) );
  XNOR U52182 ( .A(n52002), .B(n48880), .Z(n46569) );
  XOR U52183 ( .A(round_reg[228]), .B(n51561), .Z(n48880) );
  ANDN U52184 ( .B(n47619), .A(n47617), .Z(n52002) );
  XOR U52185 ( .A(round_reg[1448]), .B(n51883), .Z(n47617) );
  XOR U52186 ( .A(round_reg[1071]), .B(n50456), .Z(n47619) );
  XNOR U52187 ( .A(n52003), .B(n48873), .Z(n47695) );
  XOR U52188 ( .A(round_reg[169]), .B(n49947), .Z(n48873) );
  ANDN U52189 ( .B(n47612), .A(n48177), .Z(n52003) );
  IV U52190 ( .A(n47614), .Z(n48177) );
  XOR U52191 ( .A(round_reg[978]), .B(n51053), .Z(n47614) );
  XOR U52192 ( .A(round_reg[1354]), .B(n52004), .Z(n47612) );
  XOR U52193 ( .A(n52005), .B(n52006), .Z(n45437) );
  XOR U52194 ( .A(n46341), .B(n52007), .Z(n52006) );
  XNOR U52195 ( .A(n52008), .B(n51879), .Z(n46341) );
  ANDN U52196 ( .B(n50201), .A(n48250), .Z(n52008) );
  XOR U52197 ( .A(round_reg[349]), .B(n51541), .Z(n48250) );
  IV U52198 ( .A(n49869), .Z(n51541) );
  XOR U52199 ( .A(n52009), .B(n52010), .Z(n49869) );
  XOR U52200 ( .A(n42512), .B(n52011), .Z(n52005) );
  XNOR U52201 ( .A(n47027), .B(n52012), .Z(n52011) );
  XNOR U52202 ( .A(n52013), .B(n51876), .Z(n47027) );
  ANDN U52203 ( .B(n50212), .A(n48256), .Z(n52013) );
  IV U52204 ( .A(n50213), .Z(n48256) );
  XNOR U52205 ( .A(round_reg[470]), .B(n50482), .Z(n50213) );
  XNOR U52206 ( .A(n52014), .B(n51884), .Z(n42512) );
  ANDN U52207 ( .B(n50203), .A(n50205), .Z(n52014) );
  XOR U52208 ( .A(round_reg[568]), .B(n52015), .Z(n50205) );
  XNOR U52209 ( .A(n51761), .B(n46086), .Z(n44714) );
  IV U52210 ( .A(n43958), .Z(n46086) );
  XOR U52211 ( .A(n52016), .B(n48399), .Z(n51761) );
  ANDN U52212 ( .B(n47049), .A(n47050), .Z(n52016) );
  XOR U52213 ( .A(round_reg[525]), .B(n51343), .Z(n47050) );
  XNOR U52214 ( .A(n52017), .B(n45031), .Z(n45019) );
  XOR U52215 ( .A(n49367), .B(n45592), .Z(n45031) );
  XOR U52216 ( .A(n46408), .B(n48665), .Z(n45592) );
  XNOR U52217 ( .A(n52018), .B(n52019), .Z(n48665) );
  XNOR U52218 ( .A(n46582), .B(n45275), .Z(n52019) );
  XNOR U52219 ( .A(n52020), .B(n49966), .Z(n45275) );
  XNOR U52220 ( .A(round_reg[647]), .B(n51699), .Z(n49966) );
  ANDN U52221 ( .B(n49967), .A(n52021), .Z(n52020) );
  XNOR U52222 ( .A(n52022), .B(n49972), .Z(n46582) );
  XOR U52223 ( .A(round_reg[939]), .B(n48452), .Z(n49972) );
  ANDN U52224 ( .B(n49371), .A(n49372), .Z(n52022) );
  XNOR U52225 ( .A(round_reg[513]), .B(n51203), .Z(n49371) );
  XOR U52226 ( .A(n45408), .B(n52023), .Z(n52018) );
  XNOR U52227 ( .A(n46259), .B(n43331), .Z(n52023) );
  XOR U52228 ( .A(n52024), .B(n50638), .Z(n43331) );
  XOR U52229 ( .A(round_reg[868]), .B(n51104), .Z(n50638) );
  ANDN U52230 ( .B(n49364), .A(n49365), .Z(n52024) );
  XNOR U52231 ( .A(round_reg[479]), .B(n52025), .Z(n49364) );
  XNOR U52232 ( .A(n52026), .B(n49975), .Z(n46259) );
  XOR U52233 ( .A(round_reg[725]), .B(n48948), .Z(n49975) );
  ANDN U52234 ( .B(n49360), .A(n49361), .Z(n52026) );
  XNOR U52235 ( .A(round_reg[358]), .B(n50412), .Z(n49360) );
  XNOR U52236 ( .A(n52027), .B(n49963), .Z(n45408) );
  XNOR U52237 ( .A(round_reg[771]), .B(n52028), .Z(n49963) );
  AND U52238 ( .A(n49533), .B(n49532), .Z(n52027) );
  XNOR U52239 ( .A(round_reg[409]), .B(n51656), .Z(n49532) );
  XNOR U52240 ( .A(n52029), .B(n52030), .Z(n46408) );
  XOR U52241 ( .A(n46170), .B(n43670), .Z(n52030) );
  XOR U52242 ( .A(n52031), .B(n49879), .Z(n43670) );
  XNOR U52243 ( .A(round_reg[117]), .B(n52032), .Z(n49879) );
  ANDN U52244 ( .B(n49382), .A(n48542), .Z(n52031) );
  XNOR U52245 ( .A(round_reg[1225]), .B(n51164), .Z(n48542) );
  XOR U52246 ( .A(round_reg[1298]), .B(n51428), .Z(n49382) );
  XNOR U52247 ( .A(n52033), .B(n49874), .Z(n46170) );
  XOR U52248 ( .A(round_reg[283]), .B(n51009), .Z(n49874) );
  AND U52249 ( .A(n48534), .B(n49386), .Z(n52033) );
  XOR U52250 ( .A(round_reg[1516]), .B(n51911), .Z(n49386) );
  XOR U52251 ( .A(round_reg[1127]), .B(n52034), .Z(n48534) );
  XOR U52252 ( .A(n46492), .B(n52035), .Z(n52029) );
  XOR U52253 ( .A(n49870), .B(n44489), .Z(n52035) );
  XNOR U52254 ( .A(n52036), .B(n49884), .Z(n44489) );
  XOR U52255 ( .A(round_reg[235]), .B(n51528), .Z(n49884) );
  ANDN U52256 ( .B(n49384), .A(n48538), .Z(n52036) );
  XNOR U52257 ( .A(round_reg[1078]), .B(n48445), .Z(n48538) );
  XOR U52258 ( .A(round_reg[1455]), .B(n49631), .Z(n49384) );
  XOR U52259 ( .A(n52037), .B(n52038), .Z(n49631) );
  XNOR U52260 ( .A(n52039), .B(n49876), .Z(n49870) );
  XNOR U52261 ( .A(round_reg[176]), .B(n51818), .Z(n49876) );
  AND U52262 ( .A(n48525), .B(n49377), .Z(n52039) );
  XNOR U52263 ( .A(round_reg[1361]), .B(n50451), .Z(n49377) );
  XOR U52264 ( .A(round_reg[985]), .B(n50971), .Z(n48525) );
  IV U52265 ( .A(n50228), .Z(n50971) );
  XNOR U52266 ( .A(n52040), .B(n49881), .Z(n46492) );
  XNOR U52267 ( .A(round_reg[31]), .B(n52041), .Z(n49881) );
  ANDN U52268 ( .B(n49379), .A(n48529), .Z(n52040) );
  XNOR U52269 ( .A(round_reg[1153]), .B(n51203), .Z(n48529) );
  XNOR U52270 ( .A(round_reg[1581]), .B(n50153), .Z(n49379) );
  XNOR U52271 ( .A(n52042), .B(n49967), .Z(n49367) );
  XNOR U52272 ( .A(round_reg[581]), .B(n50509), .Z(n49967) );
  IV U52273 ( .A(n50441), .Z(n50509) );
  ANDN U52274 ( .B(n52021), .A(n51857), .Z(n52042) );
  ANDN U52275 ( .B(n44447), .A(n45032), .Z(n52017) );
  XOR U52276 ( .A(n45231), .B(n49045), .Z(n45032) );
  XOR U52277 ( .A(n52043), .B(n52044), .Z(n49045) );
  ANDN U52278 ( .B(n50867), .A(n50865), .Z(n52043) );
  XOR U52279 ( .A(round_reg[1183]), .B(n51687), .Z(n50867) );
  IV U52280 ( .A(n45953), .Z(n45231) );
  XNOR U52281 ( .A(n52045), .B(n52046), .Z(n50588) );
  XNOR U52282 ( .A(n47567), .B(n50959), .Z(n52046) );
  AND U52283 ( .A(n49054), .B(n49052), .Z(n52047) );
  XNOR U52284 ( .A(round_reg[1328]), .B(n49856), .Z(n49054) );
  ANDN U52285 ( .B(n49057), .A(n49056), .Z(n52048) );
  XNOR U52286 ( .A(round_reg[1421]), .B(n51330), .Z(n49057) );
  XOR U52287 ( .A(n47631), .B(n52049), .Z(n52045) );
  XOR U52288 ( .A(n45813), .B(n52050), .Z(n52049) );
  XNOR U52289 ( .A(n52051), .B(n51294), .Z(n45813) );
  ANDN U52290 ( .B(n49062), .A(n49060), .Z(n52051) );
  XNOR U52291 ( .A(round_reg[1482]), .B(n50852), .Z(n49062) );
  XOR U52292 ( .A(n52052), .B(n51299), .Z(n47631) );
  NOR U52293 ( .A(n49049), .B(n49047), .Z(n52052) );
  XOR U52294 ( .A(round_reg[1391]), .B(n52053), .Z(n49049) );
  XNOR U52295 ( .A(n52054), .B(n52055), .Z(n51746) );
  XNOR U52296 ( .A(n49580), .B(n45636), .Z(n52055) );
  XOR U52297 ( .A(n52056), .B(n51287), .Z(n45636) );
  ANDN U52298 ( .B(n51304), .A(n51305), .Z(n52056) );
  XOR U52299 ( .A(n52057), .B(n52058), .Z(n49580) );
  ANDN U52300 ( .B(n46845), .A(n46843), .Z(n52057) );
  XNOR U52301 ( .A(n42159), .B(n52059), .Z(n52054) );
  XOR U52302 ( .A(n48599), .B(n46636), .Z(n52059) );
  XNOR U52303 ( .A(n52060), .B(n51274), .Z(n46636) );
  XNOR U52304 ( .A(n52061), .B(n51277), .Z(n48599) );
  ANDN U52305 ( .B(n47954), .A(n47952), .Z(n52061) );
  XNOR U52306 ( .A(n52062), .B(n51282), .Z(n42159) );
  ANDN U52307 ( .B(n46838), .A(n46836), .Z(n52062) );
  IV U52308 ( .A(n52063), .Z(n46838) );
  XNOR U52309 ( .A(n43722), .B(n48111), .Z(n44447) );
  XNOR U52310 ( .A(n52064), .B(n49925), .Z(n48111) );
  XOR U52311 ( .A(round_reg[959]), .B(n52065), .Z(n47649) );
  XOR U52312 ( .A(n47131), .B(n51191), .Z(n43722) );
  XOR U52313 ( .A(n52066), .B(n52067), .Z(n51191) );
  XOR U52314 ( .A(n44113), .B(n49471), .Z(n52067) );
  XOR U52315 ( .A(n52068), .B(n49918), .Z(n49471) );
  XOR U52316 ( .A(round_reg[74]), .B(n52004), .Z(n49918) );
  NOR U52317 ( .A(n48114), .B(n47656), .Z(n52068) );
  XNOR U52318 ( .A(round_reg[1246]), .B(n51486), .Z(n47656) );
  XOR U52319 ( .A(round_reg[1319]), .B(n50732), .Z(n48114) );
  XNOR U52320 ( .A(n52069), .B(n49926), .Z(n44113) );
  XNOR U52321 ( .A(round_reg[133]), .B(n51293), .Z(n49926) );
  NOR U52322 ( .A(n49925), .B(n47647), .Z(n52069) );
  XOR U52323 ( .A(round_reg[1006]), .B(n50718), .Z(n47647) );
  XNOR U52324 ( .A(round_reg[1382]), .B(n49280), .Z(n49925) );
  XOR U52325 ( .A(n47158), .B(n52070), .Z(n52066) );
  XOR U52326 ( .A(n48800), .B(n45712), .Z(n52070) );
  XNOR U52327 ( .A(n52071), .B(n50425), .Z(n45712) );
  XNOR U52328 ( .A(round_reg[304]), .B(n51953), .Z(n50425) );
  ANDN U52329 ( .B(n48119), .A(n47664), .Z(n52071) );
  XNOR U52330 ( .A(round_reg[1148]), .B(n52072), .Z(n47664) );
  XOR U52331 ( .A(round_reg[1473]), .B(n52073), .Z(n48119) );
  XNOR U52332 ( .A(n52074), .B(n49921), .Z(n48800) );
  XOR U52333 ( .A(round_reg[52]), .B(n50440), .Z(n49921) );
  ANDN U52334 ( .B(n49595), .A(n47651), .Z(n52074) );
  XOR U52335 ( .A(round_reg[1174]), .B(n51200), .Z(n47651) );
  XOR U52336 ( .A(round_reg[1538]), .B(n49790), .Z(n49595) );
  IV U52337 ( .A(n51539), .Z(n49790) );
  XNOR U52338 ( .A(n52075), .B(n49923), .Z(n47158) );
  XOR U52339 ( .A(round_reg[192]), .B(n50415), .Z(n49923) );
  ANDN U52340 ( .B(n48116), .A(n47660), .Z(n52075) );
  XNOR U52341 ( .A(round_reg[1035]), .B(n51205), .Z(n47660) );
  XOR U52342 ( .A(round_reg[1412]), .B(n52076), .Z(n48116) );
  XOR U52343 ( .A(n52077), .B(n52078), .Z(n47131) );
  XNOR U52344 ( .A(n47589), .B(n47634), .Z(n52078) );
  XNOR U52345 ( .A(n52079), .B(n50044), .Z(n47634) );
  XOR U52346 ( .A(round_reg[1173]), .B(n49268), .Z(n50044) );
  ANDN U52347 ( .B(n48733), .A(n48734), .Z(n52079) );
  XNOR U52348 ( .A(round_reg[428]), .B(n50139), .Z(n48734) );
  XOR U52349 ( .A(round_reg[790]), .B(n50482), .Z(n48733) );
  XNOR U52350 ( .A(n52080), .B(n49485), .Z(n47589) );
  XOR U52351 ( .A(round_reg[1034]), .B(n52004), .Z(n49485) );
  NOR U52352 ( .A(n48737), .B(n48738), .Z(n52080) );
  XNOR U52353 ( .A(round_reg[600]), .B(n51812), .Z(n48738) );
  XOR U52354 ( .A(round_reg[666]), .B(n52081), .Z(n48737) );
  XOR U52355 ( .A(n44038), .B(n52082), .Z(n52077) );
  XOR U52356 ( .A(n45494), .B(n48188), .Z(n52082) );
  XNOR U52357 ( .A(n52083), .B(n49488), .Z(n48188) );
  XOR U52358 ( .A(round_reg[1147]), .B(n52084), .Z(n49488) );
  ANDN U52359 ( .B(n48720), .A(n48721), .Z(n52083) );
  XNOR U52360 ( .A(round_reg[377]), .B(n50828), .Z(n48721) );
  XOR U52361 ( .A(round_reg[744]), .B(n51042), .Z(n48720) );
  XNOR U52362 ( .A(n52085), .B(n49482), .Z(n45494) );
  XOR U52363 ( .A(round_reg[1245]), .B(n50520), .Z(n49482) );
  ANDN U52364 ( .B(n48729), .A(n48730), .Z(n52085) );
  XNOR U52365 ( .A(round_reg[498]), .B(n52086), .Z(n48730) );
  XOR U52366 ( .A(round_reg[887]), .B(n52087), .Z(n48729) );
  XNOR U52367 ( .A(n52088), .B(n49478), .Z(n44038) );
  XOR U52368 ( .A(round_reg[1005]), .B(n52089), .Z(n49478) );
  ANDN U52369 ( .B(n48724), .A(n48725), .Z(n52088) );
  XNOR U52370 ( .A(round_reg[532]), .B(n49608), .Z(n48725) );
  XOR U52371 ( .A(round_reg[958]), .B(n52090), .Z(n48724) );
  XNOR U52372 ( .A(n39173), .B(n52091), .Z(n51966) );
  XOR U52373 ( .A(n38484), .B(n35578), .Z(n52091) );
  XNOR U52374 ( .A(n52092), .B(n45026), .Z(n35578) );
  XOR U52375 ( .A(n47417), .B(n46158), .Z(n45026) );
  IV U52376 ( .A(n43337), .Z(n46158) );
  XOR U52377 ( .A(n48264), .B(n47151), .Z(n43337) );
  XNOR U52378 ( .A(n52093), .B(n52094), .Z(n47151) );
  XNOR U52379 ( .A(n48801), .B(n46115), .Z(n52094) );
  XNOR U52380 ( .A(n52095), .B(n48024), .Z(n46115) );
  XOR U52381 ( .A(round_reg[1052]), .B(n51617), .Z(n48024) );
  ANDN U52382 ( .B(n47153), .A(n47154), .Z(n52095) );
  XOR U52383 ( .A(round_reg[618]), .B(n48356), .Z(n47154) );
  XNOR U52384 ( .A(round_reg[684]), .B(n49982), .Z(n47153) );
  IV U52385 ( .A(n50221), .Z(n49982) );
  XOR U52386 ( .A(n52096), .B(n52097), .Z(n50221) );
  XNOR U52387 ( .A(n52098), .B(n48029), .Z(n48801) );
  XOR U52388 ( .A(round_reg[1101]), .B(n51330), .Z(n48029) );
  XNOR U52389 ( .A(round_reg[331]), .B(n51127), .Z(n46137) );
  XOR U52390 ( .A(round_reg[762]), .B(n51137), .Z(n46136) );
  IV U52391 ( .A(n50882), .Z(n51137) );
  XOR U52392 ( .A(n52099), .B(n52100), .Z(n50882) );
  XOR U52393 ( .A(n46174), .B(n52101), .Z(n52093) );
  XOR U52394 ( .A(n45321), .B(n44694), .Z(n52101) );
  XNOR U52395 ( .A(n52102), .B(n48032), .Z(n44694) );
  XNOR U52396 ( .A(round_reg[1023]), .B(n50841), .Z(n48032) );
  ANDN U52397 ( .B(n46238), .A(n46239), .Z(n52102) );
  XNOR U52398 ( .A(round_reg[550]), .B(n51411), .Z(n46239) );
  XNOR U52399 ( .A(round_reg[912]), .B(n50955), .Z(n46238) );
  XNOR U52400 ( .A(n52103), .B(n48810), .Z(n45321) );
  XOR U52401 ( .A(round_reg[1263]), .B(n50414), .Z(n48810) );
  ANDN U52402 ( .B(n46146), .A(n46148), .Z(n52103) );
  XNOR U52403 ( .A(round_reg[452]), .B(n50419), .Z(n46148) );
  XNOR U52404 ( .A(round_reg[841]), .B(n51721), .Z(n46146) );
  XNOR U52405 ( .A(n52104), .B(n48021), .Z(n46174) );
  XNOR U52406 ( .A(round_reg[1191]), .B(n51947), .Z(n48021) );
  ANDN U52407 ( .B(n46142), .A(n46143), .Z(n52104) );
  XNOR U52408 ( .A(round_reg[446]), .B(n51793), .Z(n46143) );
  IV U52409 ( .A(n51243), .Z(n51793) );
  XNOR U52410 ( .A(n52106), .B(n52107), .Z(n51692) );
  XNOR U52411 ( .A(round_reg[1341]), .B(round_reg[1021]), .Z(n52107) );
  XOR U52412 ( .A(round_reg[381]), .B(n52108), .Z(n52106) );
  XOR U52413 ( .A(round_reg[701]), .B(round_reg[61]), .Z(n52108) );
  XNOR U52414 ( .A(round_reg[808]), .B(n51883), .Z(n46142) );
  XOR U52415 ( .A(n52109), .B(n52110), .Z(n48264) );
  XNOR U52416 ( .A(n44255), .B(n45502), .Z(n52110) );
  XNOR U52417 ( .A(n52111), .B(n48621), .Z(n45502) );
  XOR U52418 ( .A(round_reg[6]), .B(n50643), .Z(n48621) );
  ANDN U52419 ( .B(n47419), .A(n47420), .Z(n52111) );
  XOR U52420 ( .A(round_reg[1556]), .B(n51332), .Z(n47419) );
  XNOR U52421 ( .A(n52112), .B(n48615), .Z(n44255) );
  XNOR U52422 ( .A(round_reg[151]), .B(n52113), .Z(n48615) );
  ANDN U52423 ( .B(n47424), .A(n47425), .Z(n52112) );
  XOR U52424 ( .A(n44566), .B(n52114), .Z(n52109) );
  XOR U52425 ( .A(n43575), .B(n48601), .Z(n52114) );
  XNOR U52426 ( .A(n52115), .B(n48607), .Z(n48601) );
  XOR U52427 ( .A(round_reg[92]), .B(n51617), .Z(n48607) );
  XOR U52428 ( .A(n52116), .B(n52117), .Z(n51617) );
  ANDN U52429 ( .B(n47432), .A(n47433), .Z(n52115) );
  XNOR U52430 ( .A(n52118), .B(n48610), .Z(n43575) );
  XNOR U52431 ( .A(round_reg[210]), .B(n50475), .Z(n48610) );
  ANDN U52432 ( .B(n48611), .A(n52119), .Z(n52118) );
  XNOR U52433 ( .A(n52120), .B(n48618), .Z(n44566) );
  XNOR U52434 ( .A(round_reg[258]), .B(n51539), .Z(n48618) );
  ANDN U52435 ( .B(n47428), .A(n47429), .Z(n52120) );
  XOR U52436 ( .A(round_reg[1491]), .B(n52123), .Z(n47428) );
  XNOR U52437 ( .A(n52124), .B(n48611), .Z(n47417) );
  XOR U52438 ( .A(round_reg[1430]), .B(n50482), .Z(n48611) );
  XNOR U52439 ( .A(n52125), .B(n52126), .Z(n50482) );
  ANDN U52440 ( .B(n52119), .A(n50048), .Z(n52124) );
  ANDN U52441 ( .B(n44725), .A(n44451), .Z(n52092) );
  XOR U52442 ( .A(n47825), .B(n43829), .Z(n44451) );
  XOR U52443 ( .A(n52127), .B(n49439), .Z(n43829) );
  XNOR U52444 ( .A(n52128), .B(n52129), .Z(n49439) );
  XNOR U52445 ( .A(n41653), .B(n45265), .Z(n52129) );
  XNOR U52446 ( .A(n52130), .B(n47924), .Z(n45265) );
  XOR U52447 ( .A(round_reg[1114]), .B(n49792), .Z(n47924) );
  NOR U52448 ( .A(n47923), .B(n48163), .Z(n52130) );
  XOR U52449 ( .A(round_reg[344]), .B(n51446), .Z(n48163) );
  XOR U52450 ( .A(round_reg[711]), .B(n48706), .Z(n47923) );
  XNOR U52451 ( .A(n52131), .B(n49233), .Z(n41653) );
  XOR U52452 ( .A(round_reg[1204]), .B(n51227), .Z(n49233) );
  NOR U52453 ( .A(n47830), .B(n47828), .Z(n52131) );
  XNOR U52454 ( .A(round_reg[821]), .B(n50744), .Z(n47828) );
  XNOR U52455 ( .A(round_reg[395]), .B(n51205), .Z(n47830) );
  XNOR U52456 ( .A(n47908), .B(n52134), .Z(n52128) );
  XNOR U52457 ( .A(n43604), .B(n46911), .Z(n52134) );
  XOR U52458 ( .A(n52135), .B(n47927), .Z(n46911) );
  XOR U52459 ( .A(round_reg[1276]), .B(n50719), .Z(n47927) );
  ANDN U52460 ( .B(n47832), .A(n47834), .Z(n52135) );
  XOR U52461 ( .A(round_reg[465]), .B(n51342), .Z(n47834) );
  XOR U52462 ( .A(round_reg[854]), .B(n51200), .Z(n47832) );
  XNOR U52463 ( .A(n52136), .B(n47920), .Z(n43604) );
  XOR U52464 ( .A(round_reg[1065]), .B(n49905), .Z(n47920) );
  XNOR U52465 ( .A(n52137), .B(n52138), .Z(n49905) );
  NOR U52466 ( .A(n47824), .B(n47822), .Z(n52136) );
  XOR U52467 ( .A(round_reg[697]), .B(n50828), .Z(n47822) );
  XOR U52468 ( .A(round_reg[631]), .B(n51810), .Z(n47824) );
  XOR U52469 ( .A(n52139), .B(n47916), .Z(n47908) );
  XNOR U52470 ( .A(round_reg[972]), .B(n50933), .Z(n47916) );
  NOR U52471 ( .A(n51044), .B(n47915), .Z(n52139) );
  XOR U52472 ( .A(n52140), .B(n47915), .Z(n47825) );
  XNOR U52473 ( .A(round_reg[925]), .B(n50520), .Z(n47915) );
  XOR U52474 ( .A(round_reg[163]), .B(n51459), .Z(n49254) );
  XNOR U52475 ( .A(round_reg[563]), .B(n50966), .Z(n51044) );
  XNOR U52476 ( .A(n52012), .B(n42513), .Z(n44725) );
  XNOR U52477 ( .A(n52141), .B(n51874), .Z(n52012) );
  ANDN U52478 ( .B(n50210), .A(n49887), .Z(n52141) );
  XOR U52479 ( .A(round_reg[400]), .B(n52142), .Z(n49887) );
  XNOR U52480 ( .A(n52143), .B(n47513), .Z(n38484) );
  XOR U52481 ( .A(n51887), .B(n42301), .Z(n47513) );
  XNOR U52482 ( .A(n52144), .B(n52145), .Z(n50570) );
  XOR U52483 ( .A(n46800), .B(n49325), .Z(n52145) );
  XNOR U52484 ( .A(n52146), .B(n48055), .Z(n49325) );
  XOR U52485 ( .A(round_reg[225]), .B(n51478), .Z(n48704) );
  XOR U52486 ( .A(n52147), .B(n48058), .Z(n46800) );
  XNOR U52487 ( .A(round_reg[273]), .B(n52148), .Z(n47208) );
  XOR U52488 ( .A(n41643), .B(n52149), .Z(n52144) );
  XOR U52489 ( .A(n45733), .B(n46462), .Z(n52149) );
  XNOR U52490 ( .A(n52150), .B(n48052), .Z(n46462) );
  ANDN U52491 ( .B(n47198), .A(n48698), .Z(n52150) );
  XOR U52492 ( .A(round_reg[107]), .B(n51217), .Z(n48698) );
  IV U52493 ( .A(n49867), .Z(n51217) );
  XNOR U52494 ( .A(n52151), .B(n48045), .Z(n45733) );
  XNOR U52495 ( .A(round_reg[166]), .B(n51547), .Z(n47212) );
  XOR U52496 ( .A(n52152), .B(n48047), .Z(n41643) );
  ANDN U52497 ( .B(n47203), .A(n47204), .Z(n52152) );
  XOR U52498 ( .A(round_reg[21]), .B(n52153), .Z(n47204) );
  XNOR U52499 ( .A(n52154), .B(n52155), .Z(n48245) );
  XOR U52500 ( .A(n45120), .B(n46201), .Z(n52155) );
  XOR U52501 ( .A(n52156), .B(n48075), .Z(n46201) );
  ANDN U52502 ( .B(n51899), .A(n51900), .Z(n52156) );
  XNOR U52503 ( .A(n52157), .B(n48065), .Z(n45120) );
  AND U52504 ( .A(n51894), .B(n51893), .Z(n52157) );
  XNOR U52505 ( .A(n52158), .B(n52159), .Z(n52154) );
  XOR U52506 ( .A(n46708), .B(n46876), .Z(n52159) );
  XOR U52507 ( .A(n52160), .B(n48079), .Z(n46876) );
  ANDN U52508 ( .B(n51896), .A(n51897), .Z(n52160) );
  XOR U52509 ( .A(n52161), .B(n48712), .Z(n46708) );
  ANDN U52510 ( .B(n52162), .A(n52163), .Z(n52161) );
  XOR U52511 ( .A(n52164), .B(n52162), .Z(n51887) );
  ANDN U52512 ( .B(n52163), .A(n48710), .Z(n52164) );
  ANDN U52513 ( .B(n44727), .A(n44437), .Z(n52143) );
  IV U52514 ( .A(n44728), .Z(n44437) );
  XOR U52515 ( .A(n51863), .B(n45902), .Z(n44728) );
  XNOR U52516 ( .A(n52165), .B(n49660), .Z(n51863) );
  ANDN U52517 ( .B(n49954), .A(n48669), .Z(n52165) );
  XNOR U52518 ( .A(round_reg[1363]), .B(n52166), .Z(n48669) );
  XOR U52519 ( .A(n49193), .B(n45646), .Z(n44727) );
  XOR U52520 ( .A(n46948), .B(n47607), .Z(n45646) );
  XNOR U52521 ( .A(n52167), .B(n52168), .Z(n47607) );
  XOR U52522 ( .A(n45301), .B(n47593), .Z(n52168) );
  XNOR U52523 ( .A(n52169), .B(n47941), .Z(n47593) );
  XOR U52524 ( .A(round_reg[402]), .B(n51532), .Z(n47941) );
  ANDN U52525 ( .B(n49169), .A(n47551), .Z(n52169) );
  XOR U52526 ( .A(round_reg[1575]), .B(n52170), .Z(n47551) );
  XOR U52527 ( .A(round_reg[25]), .B(n50228), .Z(n49169) );
  XOR U52528 ( .A(n52171), .B(n52172), .Z(n50228) );
  XOR U52529 ( .A(n52173), .B(n47938), .Z(n45301) );
  XNOR U52530 ( .A(round_reg[351]), .B(n52041), .Z(n47938) );
  ANDN U52531 ( .B(n49174), .A(n47564), .Z(n52173) );
  XOR U52532 ( .A(round_reg[1510]), .B(n51572), .Z(n47564) );
  IV U52533 ( .A(n51411), .Z(n51572) );
  XNOR U52534 ( .A(round_reg[277]), .B(n49907), .Z(n49174) );
  XOR U52535 ( .A(n51021), .B(n52174), .Z(n52167) );
  XOR U52536 ( .A(n47391), .B(n44521), .Z(n52174) );
  XNOR U52537 ( .A(n52175), .B(n47943), .Z(n44521) );
  XNOR U52538 ( .A(round_reg[472]), .B(n51145), .Z(n47943) );
  ANDN U52539 ( .B(n49171), .A(n47556), .Z(n52175) );
  XOR U52540 ( .A(round_reg[1292]), .B(n52176), .Z(n47556) );
  XNOR U52541 ( .A(round_reg[111]), .B(n50456), .Z(n49171) );
  IV U52542 ( .A(n52053), .Z(n50456) );
  XOR U52543 ( .A(n52177), .B(n52178), .Z(n52053) );
  XNOR U52544 ( .A(n52179), .B(n47946), .Z(n47391) );
  XNOR U52545 ( .A(round_reg[570]), .B(n49861), .Z(n47946) );
  ANDN U52546 ( .B(n49180), .A(n48184), .Z(n52179) );
  XNOR U52547 ( .A(round_reg[1355]), .B(n51205), .Z(n48184) );
  XOR U52548 ( .A(round_reg[170]), .B(n50761), .Z(n49180) );
  XOR U52549 ( .A(n52180), .B(n47936), .Z(n51021) );
  XOR U52550 ( .A(round_reg[638]), .B(n50777), .Z(n47936) );
  ANDN U52551 ( .B(n49177), .A(n47560), .Z(n52180) );
  XOR U52552 ( .A(round_reg[1449]), .B(n52181), .Z(n47560) );
  XNOR U52553 ( .A(round_reg[229]), .B(n52001), .Z(n49177) );
  XOR U52554 ( .A(n52182), .B(n52183), .Z(n46948) );
  XNOR U52555 ( .A(n47319), .B(n44329), .Z(n52183) );
  XNOR U52556 ( .A(n52184), .B(n50683), .Z(n44329) );
  XOR U52557 ( .A(round_reg[1073]), .B(n50514), .Z(n50683) );
  ANDN U52558 ( .B(n49185), .A(n49186), .Z(n52184) );
  XOR U52559 ( .A(round_reg[641]), .B(n51347), .Z(n49185) );
  XNOR U52560 ( .A(n52185), .B(n50690), .Z(n47319) );
  XNOR U52561 ( .A(round_reg[1122]), .B(n51595), .Z(n50690) );
  ANDN U52562 ( .B(n49189), .A(n49191), .Z(n52185) );
  XOR U52563 ( .A(round_reg[719]), .B(n48553), .Z(n49189) );
  XOR U52564 ( .A(n46160), .B(n52186), .Z(n52182) );
  XOR U52565 ( .A(n46118), .B(n44226), .Z(n52186) );
  XNOR U52566 ( .A(n52187), .B(n50678), .Z(n44226) );
  XNOR U52567 ( .A(round_reg[1212]), .B(n49077), .Z(n50678) );
  ANDN U52568 ( .B(n51733), .A(n52188), .Z(n52187) );
  XNOR U52569 ( .A(n52189), .B(n50687), .Z(n46118) );
  XOR U52570 ( .A(round_reg[1220]), .B(n49612), .Z(n50687) );
  XNOR U52571 ( .A(n52190), .B(n52191), .Z(n49612) );
  ANDN U52572 ( .B(n51736), .A(n51806), .Z(n52189) );
  XOR U52573 ( .A(round_reg[862]), .B(n51050), .Z(n51736) );
  XOR U52574 ( .A(n52192), .B(n50674), .Z(n46160) );
  XOR U52575 ( .A(round_reg[980]), .B(n50742), .Z(n50674) );
  ANDN U52576 ( .B(n49196), .A(n49198), .Z(n52192) );
  XNOR U52577 ( .A(round_reg[933]), .B(n51707), .Z(n49196) );
  XNOR U52578 ( .A(n52193), .B(n51733), .Z(n49193) );
  XOR U52579 ( .A(round_reg[829]), .B(n49992), .Z(n51733) );
  AND U52580 ( .A(n50677), .B(n52188), .Z(n52193) );
  XNOR U52581 ( .A(n52194), .B(n46558), .Z(n39173) );
  XOR U52582 ( .A(n44472), .B(n50661), .Z(n46558) );
  XNOR U52583 ( .A(n52195), .B(n46619), .Z(n50661) );
  ANDN U52584 ( .B(n52196), .A(n51740), .Z(n52195) );
  XNOR U52585 ( .A(n47546), .B(n46804), .Z(n44472) );
  XNOR U52586 ( .A(n52197), .B(n52198), .Z(n46804) );
  XNOR U52587 ( .A(n46057), .B(n45283), .Z(n52198) );
  XOR U52588 ( .A(n52199), .B(n46618), .Z(n45283) );
  XOR U52589 ( .A(round_reg[1074]), .B(n48967), .Z(n46618) );
  IV U52590 ( .A(n50829), .Z(n48967) );
  ANDN U52591 ( .B(n46619), .A(n52196), .Z(n52199) );
  XOR U52592 ( .A(round_reg[642]), .B(n50775), .Z(n46619) );
  XOR U52593 ( .A(n52200), .B(n46952), .Z(n46057) );
  XOR U52594 ( .A(round_reg[1221]), .B(n50441), .Z(n46952) );
  AND U52595 ( .A(n50666), .B(n46951), .Z(n52200) );
  XNOR U52596 ( .A(round_reg[863]), .B(n51687), .Z(n46951) );
  IV U52597 ( .A(n51048), .Z(n51687) );
  XOR U52598 ( .A(n52201), .B(n52202), .Z(n51048) );
  XNOR U52599 ( .A(n46602), .B(n52203), .Z(n52197) );
  XOR U52600 ( .A(n45679), .B(n44317), .Z(n52203) );
  XNOR U52601 ( .A(n52204), .B(n46608), .Z(n44317) );
  XOR U52602 ( .A(round_reg[1213]), .B(n50837), .Z(n46608) );
  ANDN U52603 ( .B(n46609), .A(n50670), .Z(n52204) );
  XOR U52604 ( .A(round_reg[830]), .B(n49866), .Z(n46609) );
  IV U52605 ( .A(n50728), .Z(n49866) );
  XOR U52606 ( .A(n52205), .B(n46613), .Z(n45679) );
  XOR U52607 ( .A(round_reg[981]), .B(n52153), .Z(n46613) );
  AND U52608 ( .A(n50668), .B(n46612), .Z(n52205) );
  XOR U52609 ( .A(round_reg[934]), .B(n51341), .Z(n46612) );
  XOR U52610 ( .A(n52206), .B(n46623), .Z(n46602) );
  XOR U52611 ( .A(round_reg[1123]), .B(n51459), .Z(n46623) );
  ANDN U52612 ( .B(n46622), .A(n50663), .Z(n52206) );
  XNOR U52613 ( .A(round_reg[720]), .B(n50119), .Z(n46622) );
  IV U52614 ( .A(n52142), .Z(n50119) );
  XOR U52615 ( .A(n52207), .B(n52208), .Z(n52142) );
  XOR U52616 ( .A(n52209), .B(n52210), .Z(n47546) );
  XNOR U52617 ( .A(n45336), .B(n44827), .Z(n52210) );
  XOR U52618 ( .A(n52211), .B(n52188), .Z(n44827) );
  XOR U52619 ( .A(round_reg[403]), .B(n51548), .Z(n52188) );
  NOR U52620 ( .A(n50679), .B(n50677), .Z(n52211) );
  XOR U52621 ( .A(round_reg[26]), .B(n52081), .Z(n50677) );
  XOR U52622 ( .A(round_reg[1576]), .B(n51535), .Z(n50679) );
  XOR U52623 ( .A(n52137), .B(n52212), .Z(n51535) );
  XOR U52624 ( .A(n52213), .B(n52214), .Z(n52137) );
  XNOR U52625 ( .A(round_reg[1320]), .B(round_reg[1000]), .Z(n52214) );
  XOR U52626 ( .A(round_reg[360]), .B(n52215), .Z(n52213) );
  XOR U52627 ( .A(round_reg[680]), .B(round_reg[40]), .Z(n52215) );
  XOR U52628 ( .A(n52216), .B(n49191), .Z(n45336) );
  XOR U52629 ( .A(round_reg[352]), .B(n50834), .Z(n49191) );
  ANDN U52630 ( .B(n49190), .A(n50689), .Z(n52216) );
  XOR U52631 ( .A(round_reg[278]), .B(n50397), .Z(n49190) );
  XOR U52632 ( .A(n49165), .B(n52217), .Z(n52209) );
  XNOR U52633 ( .A(n43322), .B(n45227), .Z(n52217) );
  XOR U52634 ( .A(n52218), .B(n49198), .Z(n45227) );
  XOR U52635 ( .A(round_reg[571]), .B(n49080), .Z(n49198) );
  XNOR U52636 ( .A(n52219), .B(n52220), .Z(n52099) );
  XNOR U52637 ( .A(round_reg[1466]), .B(round_reg[1146]), .Z(n52220) );
  XOR U52638 ( .A(round_reg[186]), .B(n52221), .Z(n52219) );
  XOR U52639 ( .A(round_reg[826]), .B(round_reg[506]), .Z(n52221) );
  AND U52640 ( .A(n50675), .B(n49197), .Z(n52218) );
  XOR U52641 ( .A(round_reg[171]), .B(n51135), .Z(n49197) );
  XOR U52642 ( .A(round_reg[1356]), .B(n50999), .Z(n50675) );
  XNOR U52643 ( .A(n52223), .B(n51806), .Z(n43322) );
  XOR U52644 ( .A(round_reg[473]), .B(n50148), .Z(n51806) );
  ANDN U52645 ( .B(n50685), .A(n50686), .Z(n52223) );
  XNOR U52646 ( .A(round_reg[1293]), .B(n50752), .Z(n50686) );
  IV U52647 ( .A(n51696), .Z(n50752) );
  XOR U52648 ( .A(round_reg[112]), .B(n49178), .Z(n50685) );
  XNOR U52649 ( .A(n52226), .B(n52227), .Z(n49178) );
  XNOR U52650 ( .A(n52228), .B(n49186), .Z(n49165) );
  XNOR U52651 ( .A(round_reg[639]), .B(n52065), .Z(n49186) );
  ANDN U52652 ( .B(n49187), .A(n50682), .Z(n52228) );
  XOR U52653 ( .A(round_reg[1450]), .B(n50761), .Z(n50682) );
  XNOR U52654 ( .A(round_reg[230]), .B(n51411), .Z(n49187) );
  XNOR U52655 ( .A(n51763), .B(n52229), .Z(n51411) );
  XOR U52656 ( .A(n52230), .B(n52231), .Z(n51763) );
  XNOR U52657 ( .A(round_reg[1445]), .B(round_reg[1125]), .Z(n52231) );
  XOR U52658 ( .A(round_reg[165]), .B(n52232), .Z(n52230) );
  XOR U52659 ( .A(round_reg[805]), .B(round_reg[485]), .Z(n52232) );
  ANDN U52660 ( .B(n44720), .A(n44441), .Z(n52194) );
  XOR U52661 ( .A(n51575), .B(n45945), .Z(n44441) );
  IV U52662 ( .A(n42822), .Z(n45945) );
  XOR U52663 ( .A(n47150), .B(n50569), .Z(n42822) );
  XOR U52664 ( .A(n52233), .B(n52234), .Z(n50569) );
  XNOR U52665 ( .A(n46689), .B(n46154), .Z(n52234) );
  XNOR U52666 ( .A(n52235), .B(n51088), .Z(n46154) );
  ANDN U52667 ( .B(n51556), .A(n50259), .Z(n52235) );
  XNOR U52668 ( .A(round_reg[760]), .B(n49977), .Z(n50259) );
  XNOR U52669 ( .A(n52236), .B(n52237), .Z(n49977) );
  XNOR U52670 ( .A(n52238), .B(n51084), .Z(n46689) );
  ANDN U52671 ( .B(n51560), .A(n50263), .Z(n52238) );
  XNOR U52672 ( .A(round_reg[910]), .B(n51047), .Z(n50263) );
  IV U52673 ( .A(n51313), .Z(n51047) );
  XNOR U52674 ( .A(n52239), .B(n52240), .Z(n51313) );
  XNOR U52675 ( .A(n42509), .B(n52241), .Z(n52233) );
  XOR U52676 ( .A(n45147), .B(n44577), .Z(n52241) );
  XNOR U52677 ( .A(n52242), .B(n51079), .Z(n44577) );
  ANDN U52678 ( .B(n51563), .A(n50781), .Z(n52242) );
  XOR U52679 ( .A(round_reg[839]), .B(n51448), .Z(n50781) );
  XNOR U52680 ( .A(n52243), .B(n51086), .Z(n45147) );
  ANDN U52681 ( .B(n51554), .A(n50253), .Z(n52243) );
  XNOR U52682 ( .A(round_reg[682]), .B(n50502), .Z(n50253) );
  IV U52683 ( .A(n51464), .Z(n50502) );
  XNOR U52684 ( .A(n52244), .B(n51081), .Z(n42509) );
  ANDN U52685 ( .B(n51566), .A(n50249), .Z(n52244) );
  XOR U52686 ( .A(round_reg[806]), .B(n51547), .Z(n50249) );
  XOR U52687 ( .A(n52245), .B(n52246), .Z(n47150) );
  XNOR U52688 ( .A(n49434), .B(n52247), .Z(n52246) );
  XNOR U52689 ( .A(n52248), .B(n49098), .Z(n49434) );
  ANDN U52690 ( .B(n51574), .A(n50462), .Z(n52248) );
  XOR U52691 ( .A(round_reg[1428]), .B(n51789), .Z(n50462) );
  XNOR U52692 ( .A(n45622), .B(n52249), .Z(n52245) );
  XOR U52693 ( .A(n49417), .B(n45440), .Z(n52249) );
  XNOR U52694 ( .A(n52250), .B(n50269), .Z(n45440) );
  ANDN U52695 ( .B(n51578), .A(n50468), .Z(n52250) );
  XOR U52696 ( .A(round_reg[1489]), .B(n49898), .Z(n50468) );
  XNOR U52697 ( .A(n52251), .B(n49111), .Z(n49417) );
  ANDN U52698 ( .B(n52252), .A(n51550), .Z(n52251) );
  XNOR U52699 ( .A(n52253), .B(n49103), .Z(n45622) );
  AND U52700 ( .A(n50470), .B(n51571), .Z(n52253) );
  XNOR U52701 ( .A(round_reg[1554]), .B(n50755), .Z(n50470) );
  XNOR U52702 ( .A(n52254), .B(n52252), .Z(n51575) );
  ANDN U52703 ( .B(n51550), .A(n49109), .Z(n52254) );
  XOR U52704 ( .A(round_reg[1022]), .B(n52255), .Z(n49109) );
  XNOR U52705 ( .A(round_reg[1398]), .B(n48445), .Z(n51550) );
  XOR U52706 ( .A(n45145), .B(n51280), .Z(n44720) );
  XOR U52707 ( .A(n52256), .B(n46844), .Z(n51280) );
  ANDN U52708 ( .B(n52257), .A(n52258), .Z(n52256) );
  XNOR U52709 ( .A(n50436), .B(n48011), .Z(n45145) );
  XOR U52710 ( .A(n52259), .B(n52260), .Z(n48011) );
  XNOR U52711 ( .A(n46677), .B(n46203), .Z(n52260) );
  XOR U52712 ( .A(n52261), .B(n46845), .Z(n46203) );
  XOR U52713 ( .A(round_reg[799]), .B(n52025), .Z(n46845) );
  ANDN U52714 ( .B(n52258), .A(n46844), .Z(n52261) );
  XOR U52715 ( .A(round_reg[437]), .B(n52032), .Z(n46844) );
  XNOR U52716 ( .A(n52262), .B(n52063), .Z(n46677) );
  XOR U52717 ( .A(round_reg[753]), .B(n50514), .Z(n52063) );
  ANDN U52718 ( .B(n51283), .A(n46837), .Z(n52262) );
  XNOR U52719 ( .A(round_reg[322]), .B(n50775), .Z(n46837) );
  XOR U52720 ( .A(n42305), .B(n52263), .Z(n52259) );
  XOR U52721 ( .A(n46250), .B(n46547), .Z(n52263) );
  XOR U52722 ( .A(n52264), .B(n47954), .Z(n46547) );
  XOR U52723 ( .A(round_reg[675]), .B(n51533), .Z(n47954) );
  NOR U52724 ( .A(n51278), .B(n47953), .Z(n52264) );
  XNOR U52725 ( .A(round_reg[609]), .B(n52265), .Z(n47953) );
  XNOR U52726 ( .A(n52266), .B(n51745), .Z(n46250) );
  XOR U52727 ( .A(round_reg[832]), .B(n50415), .Z(n51745) );
  XOR U52728 ( .A(n52267), .B(n52268), .Z(n50415) );
  ANDN U52729 ( .B(n51273), .A(n52269), .Z(n52266) );
  XNOR U52730 ( .A(round_reg[507]), .B(n51618), .Z(n51273) );
  IV U52731 ( .A(n52084), .Z(n51618) );
  XOR U52732 ( .A(n52270), .B(n52271), .Z(n52084) );
  XNOR U52733 ( .A(n52272), .B(n51305), .Z(n42305) );
  XNOR U52734 ( .A(round_reg[903]), .B(n50132), .Z(n51305) );
  ANDN U52735 ( .B(n51285), .A(n51286), .Z(n52272) );
  XNOR U52736 ( .A(round_reg[541]), .B(n51032), .Z(n51285) );
  XOR U52737 ( .A(n52273), .B(n52274), .Z(n50436) );
  XNOR U52738 ( .A(n48339), .B(n46417), .Z(n52274) );
  XOR U52739 ( .A(n52275), .B(n48791), .Z(n46417) );
  XOR U52740 ( .A(round_reg[311]), .B(n51725), .Z(n48791) );
  IV U52741 ( .A(n51810), .Z(n51725) );
  ANDN U52742 ( .B(n49523), .A(n48790), .Z(n52275) );
  XNOR U52743 ( .A(round_reg[1480]), .B(n50947), .Z(n48790) );
  XOR U52744 ( .A(round_reg[1091]), .B(n52028), .Z(n49523) );
  XNOR U52745 ( .A(n52276), .B(n49819), .Z(n48339) );
  XNOR U52746 ( .A(round_reg[199]), .B(n50107), .Z(n49819) );
  IV U52747 ( .A(n51448), .Z(n50107) );
  ANDN U52748 ( .B(n49820), .A(n49588), .Z(n52276) );
  XOR U52749 ( .A(round_reg[1042]), .B(n51532), .Z(n49588) );
  XNOR U52750 ( .A(round_reg[1419]), .B(n50138), .Z(n49820) );
  XOR U52751 ( .A(n45126), .B(n52279), .Z(n52273) );
  XOR U52752 ( .A(n48774), .B(n42334), .Z(n52279) );
  XNOR U52753 ( .A(n52280), .B(n48781), .Z(n42334) );
  XNOR U52754 ( .A(round_reg[81]), .B(n50451), .Z(n48781) );
  XOR U52755 ( .A(round_reg[1326]), .B(n50718), .Z(n48782) );
  XOR U52756 ( .A(round_reg[1253]), .B(n51707), .Z(n49520) );
  XNOR U52757 ( .A(n52281), .B(n48794), .Z(n48774) );
  XNOR U52758 ( .A(round_reg[140]), .B(n51727), .Z(n48794) );
  AND U52759 ( .A(n49512), .B(n48795), .Z(n52281) );
  XOR U52760 ( .A(round_reg[1389]), .B(n50432), .Z(n48795) );
  XOR U52761 ( .A(round_reg[1013]), .B(n51195), .Z(n49512) );
  XNOR U52762 ( .A(n52282), .B(n48787), .Z(n45126) );
  XOR U52763 ( .A(round_reg[59]), .B(n48455), .Z(n48787) );
  XNOR U52764 ( .A(n52283), .B(n52284), .Z(n48455) );
  NOR U52765 ( .A(n49515), .B(n48786), .Z(n52282) );
  XOR U52766 ( .A(round_reg[1545]), .B(n51164), .Z(n48786) );
  IV U52767 ( .A(n51462), .Z(n51164) );
  XNOR U52768 ( .A(round_reg[1181]), .B(n51032), .Z(n49515) );
  XOR U52769 ( .A(n52287), .B(n52288), .Z(n39700) );
  XOR U52770 ( .A(n37074), .B(n38173), .Z(n52288) );
  XOR U52771 ( .A(n52289), .B(n44094), .Z(n38173) );
  XNOR U52772 ( .A(n48751), .B(n45466), .Z(n44094) );
  IV U52773 ( .A(n44762), .Z(n45466) );
  XOR U52774 ( .A(n49892), .B(n47132), .Z(n44762) );
  XOR U52775 ( .A(n52290), .B(n52291), .Z(n47132) );
  XNOR U52776 ( .A(n46242), .B(n46123), .Z(n52291) );
  XNOR U52777 ( .A(n52292), .B(n50033), .Z(n46123) );
  XOR U52778 ( .A(round_reg[497]), .B(n51708), .Z(n50033) );
  NOR U52779 ( .A(n48743), .B(n48744), .Z(n52292) );
  XNOR U52780 ( .A(round_reg[1317]), .B(n50646), .Z(n48744) );
  IV U52781 ( .A(n51640), .Z(n50646) );
  XOR U52782 ( .A(n52293), .B(n52294), .Z(n51640) );
  XOR U52783 ( .A(round_reg[72]), .B(n51483), .Z(n48743) );
  IV U52784 ( .A(n51393), .Z(n51483) );
  XNOR U52785 ( .A(n52295), .B(n50036), .Z(n46242) );
  XNOR U52786 ( .A(round_reg[376]), .B(n50486), .Z(n50036) );
  IV U52787 ( .A(n49265), .Z(n50486) );
  XOR U52788 ( .A(n52296), .B(n52297), .Z(n49265) );
  XOR U52789 ( .A(n50076), .B(n52298), .Z(n52290) );
  XOR U52790 ( .A(n45580), .B(n45566), .Z(n52298) );
  XNOR U52791 ( .A(n52299), .B(n50029), .Z(n45566) );
  XOR U52792 ( .A(round_reg[599]), .B(n50738), .Z(n50029) );
  ANDN U52793 ( .B(n48757), .A(n48758), .Z(n52299) );
  XNOR U52794 ( .A(round_reg[1410]), .B(n51564), .Z(n48758) );
  XOR U52795 ( .A(round_reg[254]), .B(n50448), .Z(n48757) );
  XNOR U52796 ( .A(n52302), .B(n50040), .Z(n45580) );
  XNOR U52797 ( .A(round_reg[531]), .B(n52303), .Z(n50040) );
  ANDN U52798 ( .B(n48747), .A(n48748), .Z(n52302) );
  XNOR U52799 ( .A(round_reg[1380]), .B(n52304), .Z(n48748) );
  XOR U52800 ( .A(round_reg[131]), .B(n50421), .Z(n48747) );
  XNOR U52801 ( .A(n52305), .B(n50025), .Z(n50076) );
  XNOR U52802 ( .A(round_reg[427]), .B(n49867), .Z(n50025) );
  XOR U52803 ( .A(n52306), .B(n52307), .Z(n49867) );
  XNOR U52804 ( .A(round_reg[1536]), .B(n51199), .Z(n48755) );
  XOR U52805 ( .A(n52308), .B(n52309), .Z(n49892) );
  XOR U52806 ( .A(n44695), .B(n44409), .Z(n52309) );
  XOR U52807 ( .A(n52310), .B(n50089), .Z(n44409) );
  XOR U52808 ( .A(round_reg[1379]), .B(n51624), .Z(n50089) );
  ANDN U52809 ( .B(n46982), .A(n46984), .Z(n52310) );
  XOR U52810 ( .A(round_reg[956]), .B(n50719), .Z(n46984) );
  XOR U52811 ( .A(round_reg[1003]), .B(n50823), .Z(n46982) );
  XNOR U52812 ( .A(n47485), .B(n52311), .Z(n44695) );
  XNOR U52813 ( .A(n4549), .B(n52312), .Z(n52311) );
  NANDN U52814 ( .A(n51842), .B(n46986), .Z(n52312) );
  XOR U52815 ( .A(round_reg[1171]), .B(n52123), .Z(n46986) );
  IV U52816 ( .A(n46988), .Z(n51842) );
  XNOR U52817 ( .A(round_reg[788]), .B(n51789), .Z(n46988) );
  IV U52818 ( .A(rc_i[2]), .Z(n4549) );
  XNOR U52819 ( .A(round_reg[1599]), .B(n52313), .Z(n47485) );
  XOR U52820 ( .A(n49772), .B(n52314), .Z(n52308) );
  XOR U52821 ( .A(n42336), .B(n45761), .Z(n52314) );
  XNOR U52822 ( .A(n52315), .B(n47492), .Z(n45761) );
  XOR U52823 ( .A(round_reg[1316]), .B(n51335), .Z(n47492) );
  ANDN U52824 ( .B(n46993), .A(n51846), .Z(n52315) );
  IV U52825 ( .A(n46994), .Z(n51846) );
  XNOR U52826 ( .A(round_reg[885]), .B(n51679), .Z(n46994) );
  XOR U52827 ( .A(n51750), .B(n52316), .Z(n51679) );
  XOR U52828 ( .A(n52317), .B(n52318), .Z(n51750) );
  XNOR U52829 ( .A(round_reg[1460]), .B(round_reg[1140]), .Z(n52318) );
  XOR U52830 ( .A(round_reg[180]), .B(n52319), .Z(n52317) );
  XOR U52831 ( .A(round_reg[820]), .B(round_reg[500]), .Z(n52319) );
  XOR U52832 ( .A(round_reg[1243]), .B(n51009), .Z(n46993) );
  XNOR U52833 ( .A(n52320), .B(n50086), .Z(n42336) );
  XNOR U52834 ( .A(round_reg[1409]), .B(n50127), .Z(n50086) );
  XNOR U52835 ( .A(round_reg[664]), .B(n51446), .Z(n49910) );
  XOR U52836 ( .A(n52321), .B(n52322), .Z(n51446) );
  XOR U52837 ( .A(round_reg[1032]), .B(n51393), .Z(n49909) );
  XNOR U52838 ( .A(n52323), .B(n48463), .Z(n49772) );
  XOR U52839 ( .A(round_reg[1534]), .B(n50448), .Z(n48463) );
  XOR U52840 ( .A(round_reg[742]), .B(n49280), .Z(n49390) );
  XOR U52841 ( .A(round_reg[1145]), .B(n51253), .Z(n49389) );
  XOR U52842 ( .A(n52324), .B(n50094), .Z(n48751) );
  XOR U52843 ( .A(round_reg[302]), .B(n51582), .Z(n50094) );
  ANDN U52844 ( .B(n50223), .A(n50035), .Z(n52324) );
  XOR U52845 ( .A(round_reg[1535]), .B(n48520), .Z(n50223) );
  XOR U52846 ( .A(n52325), .B(n52105), .Z(n48520) );
  XNOR U52847 ( .A(n52326), .B(n52327), .Z(n52105) );
  XNOR U52848 ( .A(round_reg[1470]), .B(round_reg[1150]), .Z(n52327) );
  XOR U52849 ( .A(round_reg[190]), .B(n52328), .Z(n52326) );
  XOR U52850 ( .A(round_reg[830]), .B(round_reg[510]), .Z(n52328) );
  ANDN U52851 ( .B(n41415), .A(n41417), .Z(n52289) );
  XOR U52852 ( .A(n52007), .B(n42513), .Z(n41417) );
  XNOR U52853 ( .A(n52329), .B(n52330), .Z(n49823) );
  XOR U52854 ( .A(n46788), .B(n47448), .Z(n52330) );
  XOR U52855 ( .A(n52331), .B(n49888), .Z(n47448) );
  XOR U52856 ( .A(round_reg[1573]), .B(n51707), .Z(n49888) );
  IV U52857 ( .A(n52332), .Z(n51707) );
  NOR U52858 ( .A(n50210), .B(n51874), .Z(n52331) );
  XNOR U52859 ( .A(round_reg[1209]), .B(n49836), .Z(n51874) );
  XNOR U52860 ( .A(round_reg[826]), .B(n51620), .Z(n50210) );
  XNOR U52861 ( .A(n52333), .B(n52334), .Z(n51620) );
  XNOR U52862 ( .A(n52335), .B(n48257), .Z(n46788) );
  XOR U52863 ( .A(round_reg[1290]), .B(n51934), .Z(n48257) );
  IV U52864 ( .A(n52336), .Z(n51934) );
  ANDN U52865 ( .B(n51876), .A(n50212), .Z(n52335) );
  XNOR U52866 ( .A(round_reg[859]), .B(n50131), .Z(n50212) );
  IV U52867 ( .A(n50442), .Z(n50131) );
  XOR U52868 ( .A(n52337), .B(n52338), .Z(n50442) );
  XOR U52869 ( .A(round_reg[1217]), .B(n49857), .Z(n51876) );
  XOR U52870 ( .A(n43900), .B(n52339), .Z(n52329) );
  XOR U52871 ( .A(n51870), .B(n49387), .Z(n52339) );
  XNOR U52872 ( .A(n52340), .B(n50215), .Z(n49387) );
  XOR U52873 ( .A(round_reg[1353]), .B(n50227), .Z(n50215) );
  XNOR U52874 ( .A(round_reg[930]), .B(n50822), .Z(n50203) );
  XOR U52875 ( .A(round_reg[977]), .B(n51325), .Z(n51884) );
  XOR U52876 ( .A(n52343), .B(n48261), .Z(n51870) );
  XOR U52877 ( .A(round_reg[1447]), .B(n52034), .Z(n48261) );
  ANDN U52878 ( .B(n51881), .A(n50208), .Z(n52343) );
  XNOR U52879 ( .A(n52344), .B(n48252), .Z(n43900) );
  XNOR U52880 ( .A(round_reg[1508]), .B(n51561), .Z(n48252) );
  IV U52881 ( .A(n51104), .Z(n51561) );
  XOR U52882 ( .A(n52293), .B(n52345), .Z(n51104) );
  XOR U52883 ( .A(n52346), .B(n52347), .Z(n52293) );
  XNOR U52884 ( .A(round_reg[1572]), .B(round_reg[1252]), .Z(n52347) );
  XOR U52885 ( .A(round_reg[292]), .B(n52348), .Z(n52346) );
  XOR U52886 ( .A(round_reg[932]), .B(round_reg[612]), .Z(n52348) );
  NOR U52887 ( .A(n50201), .B(n51879), .Z(n52344) );
  XOR U52888 ( .A(round_reg[1119]), .B(n52025), .Z(n51879) );
  XNOR U52889 ( .A(round_reg[716]), .B(n50999), .Z(n50201) );
  IV U52890 ( .A(n51007), .Z(n50999) );
  XOR U52891 ( .A(n52349), .B(n52350), .Z(n51007) );
  XNOR U52892 ( .A(n52351), .B(n52352), .Z(n48694) );
  XNOR U52893 ( .A(n47106), .B(n44782), .Z(n52352) );
  XOR U52894 ( .A(n52353), .B(n52163), .Z(n44782) );
  XOR U52895 ( .A(round_reg[701]), .B(n52354), .Z(n52163) );
  ANDN U52896 ( .B(n48710), .A(n48711), .Z(n52353) );
  XNOR U52897 ( .A(round_reg[635]), .B(n49897), .Z(n48710) );
  XOR U52898 ( .A(n52355), .B(n51890), .Z(n47106) );
  ANDN U52899 ( .B(n48067), .A(n48068), .Z(n52355) );
  XOR U52900 ( .A(round_reg[348]), .B(n48965), .Z(n48067) );
  XOR U52901 ( .A(n52356), .B(n52337), .Z(n48965) );
  XNOR U52902 ( .A(n52357), .B(n52358), .Z(n52337) );
  XNOR U52903 ( .A(round_reg[1563]), .B(round_reg[1243]), .Z(n52358) );
  XOR U52904 ( .A(round_reg[283]), .B(n52359), .Z(n52357) );
  XOR U52905 ( .A(round_reg[923]), .B(round_reg[603]), .Z(n52359) );
  XOR U52906 ( .A(n46624), .B(n52360), .Z(n52351) );
  XOR U52907 ( .A(n43603), .B(n45251), .Z(n52360) );
  XOR U52908 ( .A(n52361), .B(n51900), .Z(n45251) );
  XOR U52909 ( .A(round_reg[929]), .B(n52265), .Z(n51900) );
  IV U52910 ( .A(n50501), .Z(n52265) );
  XOR U52911 ( .A(n52362), .B(n52363), .Z(n50501) );
  ANDN U52912 ( .B(n48073), .A(n48074), .Z(n52361) );
  XNOR U52913 ( .A(round_reg[567]), .B(n51626), .Z(n48073) );
  XNOR U52914 ( .A(n52364), .B(n51894), .Z(n43603) );
  XOR U52915 ( .A(round_reg[825]), .B(n50449), .Z(n51894) );
  IV U52916 ( .A(n51253), .Z(n50449) );
  XOR U52917 ( .A(n52365), .B(n52297), .Z(n51253) );
  XNOR U52918 ( .A(n52366), .B(n52367), .Z(n52297) );
  XNOR U52919 ( .A(round_reg[120]), .B(round_reg[1080]), .Z(n52367) );
  XOR U52920 ( .A(round_reg[1400]), .B(n52368), .Z(n52366) );
  XOR U52921 ( .A(round_reg[760]), .B(round_reg[440]), .Z(n52368) );
  XOR U52922 ( .A(round_reg[399]), .B(n48553), .Z(n48063) );
  XNOR U52923 ( .A(n52239), .B(n52369), .Z(n48553) );
  XOR U52924 ( .A(n52370), .B(n52371), .Z(n52239) );
  XNOR U52925 ( .A(round_reg[14]), .B(round_reg[1294]), .Z(n52371) );
  XOR U52926 ( .A(round_reg[334]), .B(n52372), .Z(n52370) );
  XOR U52927 ( .A(round_reg[974]), .B(round_reg[654]), .Z(n52372) );
  XNOR U52928 ( .A(n52373), .B(n51897), .Z(n46624) );
  XOR U52929 ( .A(round_reg[858]), .B(n50814), .Z(n51897) );
  ANDN U52930 ( .B(n48077), .A(n48078), .Z(n52373) );
  XOR U52931 ( .A(round_reg[469]), .B(n50232), .Z(n48077) );
  XNOR U52932 ( .A(n52374), .B(n51881), .Z(n52007) );
  XOR U52933 ( .A(round_reg[1070]), .B(n51997), .Z(n51881) );
  AND U52934 ( .A(n48260), .B(n50208), .Z(n52374) );
  XNOR U52935 ( .A(round_reg[702]), .B(n50516), .Z(n50208) );
  XOR U52936 ( .A(round_reg[636]), .B(n52375), .Z(n48260) );
  XOR U52937 ( .A(n41888), .B(n47503), .Z(n41415) );
  XNOR U52938 ( .A(n52376), .B(n47865), .Z(n47503) );
  ANDN U52939 ( .B(n49782), .A(n49781), .Z(n52376) );
  XOR U52940 ( .A(round_reg[884]), .B(n51246), .Z(n49782) );
  IV U52941 ( .A(n51227), .Z(n51246) );
  XOR U52942 ( .A(n52377), .B(n52378), .Z(n51227) );
  IV U52943 ( .A(n47140), .Z(n41888) );
  XNOR U52944 ( .A(n51833), .B(n47689), .Z(n47140) );
  XNOR U52945 ( .A(n52379), .B(n52380), .Z(n47689) );
  XOR U52946 ( .A(n41877), .B(n45715), .Z(n52380) );
  XOR U52947 ( .A(n52381), .B(n49084), .Z(n45715) );
  XOR U52948 ( .A(round_reg[1001]), .B(n51006), .Z(n49084) );
  XOR U52949 ( .A(n52382), .B(n52383), .Z(n51006) );
  XOR U52950 ( .A(round_reg[954]), .B(n52384), .Z(n47014) );
  XOR U52951 ( .A(round_reg[528]), .B(n51516), .Z(n46858) );
  XNOR U52952 ( .A(n52385), .B(n47877), .Z(n41877) );
  XOR U52953 ( .A(round_reg[1169]), .B(n49898), .Z(n47877) );
  XNOR U52954 ( .A(n52386), .B(n52208), .Z(n49898) );
  XNOR U52955 ( .A(n52387), .B(n52388), .Z(n52208) );
  XNOR U52956 ( .A(round_reg[1424]), .B(round_reg[1104]), .Z(n52388) );
  XOR U52957 ( .A(round_reg[144]), .B(n52389), .Z(n52387) );
  XOR U52958 ( .A(round_reg[784]), .B(round_reg[464]), .Z(n52389) );
  AND U52959 ( .A(n46864), .B(n47016), .Z(n52385) );
  XOR U52960 ( .A(round_reg[786]), .B(n51100), .Z(n47016) );
  XOR U52961 ( .A(round_reg[424]), .B(n51016), .Z(n46864) );
  IV U52962 ( .A(n51042), .Z(n51016) );
  XOR U52963 ( .A(n52390), .B(n52391), .Z(n51042) );
  XOR U52964 ( .A(n45600), .B(n52392), .Z(n52379) );
  XOR U52965 ( .A(n44166), .B(n45269), .Z(n52392) );
  XNOR U52966 ( .A(n52393), .B(n47880), .Z(n45269) );
  XOR U52967 ( .A(round_reg[1241]), .B(n50434), .Z(n47880) );
  NOR U52968 ( .A(n47881), .B(n47001), .Z(n52393) );
  XNOR U52969 ( .A(round_reg[494]), .B(n51525), .Z(n47001) );
  IV U52970 ( .A(n50394), .Z(n51525) );
  XOR U52971 ( .A(n52394), .B(n52395), .Z(n50394) );
  XOR U52972 ( .A(round_reg[883]), .B(n50966), .Z(n47881) );
  XNOR U52973 ( .A(n52396), .B(n52397), .Z(n50966) );
  XNOR U52974 ( .A(n52398), .B(n47883), .Z(n44166) );
  XNOR U52975 ( .A(round_reg[1030]), .B(n49271), .Z(n47883) );
  AND U52976 ( .A(n46868), .B(n47691), .Z(n52398) );
  XOR U52977 ( .A(round_reg[596]), .B(n51984), .Z(n46868) );
  IV U52978 ( .A(n51332), .Z(n51984) );
  XNOR U52979 ( .A(n52401), .B(n47885), .Z(n45600) );
  XOR U52980 ( .A(round_reg[1143]), .B(n50523), .Z(n47885) );
  XOR U52981 ( .A(n52402), .B(n52403), .Z(n50523) );
  XNOR U52982 ( .A(round_reg[373]), .B(n51195), .Z(n46854) );
  XOR U52983 ( .A(round_reg[740]), .B(n51816), .Z(n47008) );
  IV U52984 ( .A(n52304), .Z(n51816) );
  XOR U52985 ( .A(n52404), .B(n52405), .Z(n51833) );
  XNOR U52986 ( .A(n45805), .B(n43780), .Z(n52405) );
  XNOR U52987 ( .A(n52406), .B(n47864), .Z(n43780) );
  XNOR U52988 ( .A(round_reg[70]), .B(n49271), .Z(n47864) );
  XOR U52989 ( .A(n52407), .B(n52278), .Z(n49271) );
  XNOR U52990 ( .A(n52408), .B(n52409), .Z(n52278) );
  XNOR U52991 ( .A(round_reg[134]), .B(round_reg[1094]), .Z(n52409) );
  XOR U52992 ( .A(round_reg[1414]), .B(n52410), .Z(n52408) );
  XOR U52993 ( .A(round_reg[774]), .B(round_reg[454]), .Z(n52410) );
  XOR U52994 ( .A(round_reg[1242]), .B(n49625), .Z(n49781) );
  XOR U52995 ( .A(round_reg[1315]), .B(n51179), .Z(n47865) );
  IV U52996 ( .A(n51533), .Z(n51179) );
  XNOR U52997 ( .A(n52411), .B(n52412), .Z(n51533) );
  XNOR U52998 ( .A(n52413), .B(n47857), .Z(n45805) );
  XNOR U52999 ( .A(round_reg[300]), .B(n50749), .Z(n47857) );
  AND U53000 ( .A(n47501), .B(n47500), .Z(n52413) );
  XNOR U53001 ( .A(round_reg[1533]), .B(n50837), .Z(n47500) );
  XOR U53002 ( .A(round_reg[1144]), .B(n51907), .Z(n47501) );
  XOR U53003 ( .A(n45365), .B(n52414), .Z(n52404) );
  XNOR U53004 ( .A(n47852), .B(n45967), .Z(n52414) );
  XNOR U53005 ( .A(n52415), .B(n47868), .Z(n45967) );
  XOR U53006 ( .A(round_reg[48]), .B(n49856), .Z(n47868) );
  XNOR U53007 ( .A(n52416), .B(n52417), .Z(n49856) );
  ANDN U53008 ( .B(n47496), .A(n47498), .Z(n52415) );
  XOR U53009 ( .A(round_reg[1170]), .B(n52418), .Z(n47498) );
  XNOR U53010 ( .A(round_reg[1598]), .B(n50777), .Z(n47496) );
  IV U53011 ( .A(n52090), .Z(n50777) );
  XOR U53012 ( .A(n52419), .B(n52420), .Z(n52090) );
  XOR U53013 ( .A(n52421), .B(n47871), .Z(n47852) );
  XOR U53014 ( .A(round_reg[252]), .B(n50522), .Z(n47871) );
  ANDN U53015 ( .B(n47506), .A(n47508), .Z(n52421) );
  XOR U53016 ( .A(round_reg[1031]), .B(n51847), .Z(n47508) );
  IV U53017 ( .A(n48706), .Z(n51847) );
  XOR U53018 ( .A(round_reg[1408]), .B(n49083), .Z(n47506) );
  XNOR U53019 ( .A(n52422), .B(n52423), .Z(n49083) );
  XNOR U53020 ( .A(n52424), .B(n47860), .Z(n45365) );
  XNOR U53021 ( .A(round_reg[129]), .B(n50127), .Z(n47860) );
  XOR U53022 ( .A(n52121), .B(n52425), .Z(n50127) );
  XNOR U53023 ( .A(n52426), .B(n52427), .Z(n52121) );
  XNOR U53024 ( .A(round_reg[1473]), .B(round_reg[1153]), .Z(n52427) );
  XOR U53025 ( .A(round_reg[193]), .B(n52428), .Z(n52426) );
  XOR U53026 ( .A(round_reg[833]), .B(round_reg[513]), .Z(n52428) );
  ANDN U53027 ( .B(n47510), .A(n47511), .Z(n52424) );
  XOR U53028 ( .A(round_reg[1002]), .B(n51464), .Z(n47511) );
  XNOR U53029 ( .A(round_reg[1378]), .B(n50745), .Z(n47510) );
  XNOR U53030 ( .A(n52431), .B(n44097), .Z(n37074) );
  XOR U53031 ( .A(n43769), .B(n48635), .Z(n44097) );
  XNOR U53032 ( .A(n52432), .B(n48490), .Z(n48635) );
  NOR U53033 ( .A(n52433), .B(n51357), .Z(n52432) );
  XOR U53034 ( .A(round_reg[1485]), .B(n51343), .Z(n51357) );
  XNOR U53035 ( .A(n52349), .B(n52434), .Z(n51343) );
  XOR U53036 ( .A(n52435), .B(n52436), .Z(n52349) );
  XNOR U53037 ( .A(round_reg[140]), .B(round_reg[1100]), .Z(n52436) );
  XOR U53038 ( .A(round_reg[1420]), .B(n52437), .Z(n52435) );
  XOR U53039 ( .A(round_reg[780]), .B(round_reg[460]), .Z(n52437) );
  IV U53040 ( .A(n44929), .Z(n43769) );
  XNOR U53041 ( .A(n47143), .B(n51153), .Z(n44929) );
  XOR U53042 ( .A(n52438), .B(n52439), .Z(n51153) );
  XNOR U53043 ( .A(n43529), .B(n49131), .Z(n52439) );
  XOR U53044 ( .A(n52440), .B(n48477), .Z(n49131) );
  XOR U53045 ( .A(round_reg[144]), .B(n51143), .Z(n48477) );
  IV U53046 ( .A(n50735), .Z(n51143) );
  ANDN U53047 ( .B(n48658), .A(n48659), .Z(n52440) );
  XNOR U53048 ( .A(round_reg[1017]), .B(n50828), .Z(n48659) );
  XNOR U53049 ( .A(n52441), .B(n52333), .Z(n50828) );
  XNOR U53050 ( .A(n52442), .B(n52443), .Z(n52333) );
  XNOR U53051 ( .A(round_reg[121]), .B(round_reg[1081]), .Z(n52443) );
  XOR U53052 ( .A(round_reg[1401]), .B(n52444), .Z(n52442) );
  XOR U53053 ( .A(round_reg[761]), .B(round_reg[441]), .Z(n52444) );
  XOR U53054 ( .A(round_reg[1393]), .B(n50514), .Z(n48658) );
  XNOR U53055 ( .A(n52445), .B(n48482), .Z(n43529) );
  XOR U53056 ( .A(round_reg[315]), .B(n49897), .Z(n48482) );
  ANDN U53057 ( .B(n48647), .A(n48648), .Z(n52445) );
  XNOR U53058 ( .A(round_reg[1095]), .B(n50158), .Z(n48648) );
  XOR U53059 ( .A(n52446), .B(n52447), .Z(n50158) );
  XNOR U53060 ( .A(round_reg[1484]), .B(n51140), .Z(n48647) );
  XOR U53061 ( .A(n50525), .B(n52448), .Z(n52438) );
  XNOR U53062 ( .A(n46129), .B(n45758), .Z(n52448) );
  XNOR U53063 ( .A(n52449), .B(n48486), .Z(n45758) );
  XOR U53064 ( .A(round_reg[63]), .B(n50841), .Z(n48486) );
  IV U53065 ( .A(n48879), .Z(n50841) );
  XNOR U53066 ( .A(n52451), .B(n52452), .Z(n52423) );
  XNOR U53067 ( .A(round_reg[127]), .B(round_reg[1087]), .Z(n52452) );
  XOR U53068 ( .A(round_reg[1407]), .B(n52453), .Z(n52451) );
  XOR U53069 ( .A(round_reg[767]), .B(round_reg[447]), .Z(n52453) );
  ANDN U53070 ( .B(n48651), .A(n48652), .Z(n52449) );
  XOR U53071 ( .A(round_reg[1185]), .B(n51478), .Z(n48652) );
  XOR U53072 ( .A(round_reg[1549]), .B(n51093), .Z(n48651) );
  XNOR U53073 ( .A(n52454), .B(n48693), .Z(n46129) );
  XOR U53074 ( .A(round_reg[85]), .B(n48948), .Z(n48693) );
  ANDN U53075 ( .B(n48656), .A(n48654), .Z(n52454) );
  XOR U53076 ( .A(round_reg[1330]), .B(n50404), .Z(n48654) );
  XOR U53077 ( .A(n52455), .B(n52456), .Z(n50404) );
  XOR U53078 ( .A(round_reg[1257]), .B(n51520), .Z(n48656) );
  XNOR U53079 ( .A(n52457), .B(n49539), .Z(n50525) );
  XOR U53080 ( .A(round_reg[203]), .B(n51726), .Z(n49539) );
  XNOR U53081 ( .A(n52458), .B(n52459), .Z(n51726) );
  AND U53082 ( .A(n51166), .B(n50530), .Z(n52457) );
  XNOR U53083 ( .A(round_reg[1423]), .B(n50859), .Z(n50530) );
  XOR U53084 ( .A(round_reg[1046]), .B(n51183), .Z(n51166) );
  XOR U53085 ( .A(n52460), .B(n52461), .Z(n47143) );
  XOR U53086 ( .A(n48222), .B(n46175), .Z(n52461) );
  XOR U53087 ( .A(n52462), .B(n48241), .Z(n46175) );
  XNOR U53088 ( .A(round_reg[907]), .B(n51647), .Z(n48241) );
  NOR U53089 ( .A(n48631), .B(n48633), .Z(n52462) );
  XOR U53090 ( .A(round_reg[145]), .B(n51342), .Z(n48633) );
  XNOR U53091 ( .A(round_reg[545]), .B(n51478), .Z(n48631) );
  XNOR U53092 ( .A(n52463), .B(n52464), .Z(n51478) );
  XNOR U53093 ( .A(n52465), .B(n48234), .Z(n48222) );
  XOR U53094 ( .A(round_reg[803]), .B(n51459), .Z(n48234) );
  XNOR U53095 ( .A(n52466), .B(n52467), .Z(n51459) );
  XNOR U53096 ( .A(round_reg[441]), .B(n51177), .Z(n48233) );
  XOR U53097 ( .A(round_reg[0]), .B(n50457), .Z(n48642) );
  XOR U53098 ( .A(n47846), .B(n52468), .Z(n52460) );
  XOR U53099 ( .A(n45897), .B(n47438), .Z(n52468) );
  XNOR U53100 ( .A(n52469), .B(n48237), .Z(n47438) );
  XNOR U53101 ( .A(round_reg[836]), .B(n50505), .Z(n48237) );
  XNOR U53102 ( .A(n52470), .B(n51591), .Z(n50505) );
  XNOR U53103 ( .A(n52471), .B(n52472), .Z(n51591) );
  XNOR U53104 ( .A(round_reg[1540]), .B(round_reg[1220]), .Z(n52472) );
  XOR U53105 ( .A(round_reg[260]), .B(n52473), .Z(n52471) );
  XOR U53106 ( .A(round_reg[900]), .B(round_reg[580]), .Z(n52473) );
  NOR U53107 ( .A(n48637), .B(n48638), .Z(n52469) );
  XNOR U53108 ( .A(round_reg[86]), .B(n51183), .Z(n48638) );
  XNOR U53109 ( .A(round_reg[511]), .B(n49081), .Z(n48637) );
  XOR U53110 ( .A(n52474), .B(n48228), .Z(n45897) );
  XOR U53111 ( .A(round_reg[679]), .B(n50732), .Z(n48228) );
  ANDN U53112 ( .B(n48229), .A(n48628), .Z(n52474) );
  XNOR U53113 ( .A(round_reg[204]), .B(n51140), .Z(n48628) );
  XOR U53114 ( .A(round_reg[613]), .B(n52332), .Z(n48229) );
  XNOR U53115 ( .A(n52477), .B(n48491), .Z(n47846) );
  XNOR U53116 ( .A(round_reg[757]), .B(n52032), .Z(n48491) );
  IV U53117 ( .A(n51526), .Z(n52032) );
  NOR U53118 ( .A(n51611), .B(n48490), .Z(n52477) );
  XNOR U53119 ( .A(round_reg[326]), .B(n50643), .Z(n48490) );
  XOR U53120 ( .A(n51937), .B(n52446), .Z(n50643) );
  XNOR U53121 ( .A(n52478), .B(n52479), .Z(n52446) );
  XNOR U53122 ( .A(round_reg[1350]), .B(round_reg[1030]), .Z(n52479) );
  XOR U53123 ( .A(round_reg[390]), .B(n52480), .Z(n52478) );
  XOR U53124 ( .A(round_reg[710]), .B(round_reg[70]), .Z(n52480) );
  XOR U53125 ( .A(n52481), .B(n52482), .Z(n51937) );
  XNOR U53126 ( .A(round_reg[1541]), .B(round_reg[1221]), .Z(n52482) );
  XOR U53127 ( .A(round_reg[261]), .B(n52483), .Z(n52481) );
  XOR U53128 ( .A(round_reg[901]), .B(round_reg[581]), .Z(n52483) );
  IV U53129 ( .A(n52433), .Z(n51611) );
  XOR U53130 ( .A(round_reg[316]), .B(n52375), .Z(n52433) );
  IV U53131 ( .A(n50719), .Z(n52375) );
  XNOR U53132 ( .A(n52484), .B(n52270), .Z(n50719) );
  XOR U53133 ( .A(n52485), .B(n52486), .Z(n52270) );
  XNOR U53134 ( .A(round_reg[1531]), .B(round_reg[1211]), .Z(n52486) );
  XOR U53135 ( .A(round_reg[251]), .B(n52487), .Z(n52485) );
  XOR U53136 ( .A(round_reg[891]), .B(round_reg[571]), .Z(n52487) );
  ANDN U53137 ( .B(n41404), .A(n44465), .Z(n52431) );
  IV U53138 ( .A(n41405), .Z(n44465) );
  XOR U53139 ( .A(n50056), .B(n47809), .Z(n41405) );
  XOR U53140 ( .A(n46291), .B(n47258), .Z(n47809) );
  XNOR U53141 ( .A(n52488), .B(n52489), .Z(n47258) );
  XNOR U53142 ( .A(n45722), .B(n46303), .Z(n52489) );
  XOR U53143 ( .A(n52490), .B(n50762), .Z(n46303) );
  XOR U53144 ( .A(round_reg[7]), .B(n51699), .Z(n50762) );
  IV U53145 ( .A(n51349), .Z(n51699) );
  XNOR U53146 ( .A(n52492), .B(n52493), .Z(n51455) );
  XNOR U53147 ( .A(round_reg[1542]), .B(round_reg[1222]), .Z(n52493) );
  XOR U53148 ( .A(round_reg[262]), .B(n52494), .Z(n52492) );
  XOR U53149 ( .A(round_reg[902]), .B(round_reg[582]), .Z(n52494) );
  ANDN U53150 ( .B(n50058), .A(n47753), .Z(n52490) );
  XNOR U53151 ( .A(round_reg[1193]), .B(n48368), .Z(n47753) );
  IV U53152 ( .A(n50942), .Z(n48368) );
  XOR U53153 ( .A(n52390), .B(n52430), .Z(n50942) );
  XNOR U53154 ( .A(n52495), .B(n52496), .Z(n52430) );
  XNOR U53155 ( .A(round_reg[1577]), .B(round_reg[1257]), .Z(n52496) );
  XOR U53156 ( .A(round_reg[297]), .B(n52497), .Z(n52495) );
  XOR U53157 ( .A(round_reg[937]), .B(round_reg[617]), .Z(n52497) );
  XOR U53158 ( .A(n52498), .B(n52499), .Z(n52390) );
  XNOR U53159 ( .A(round_reg[1448]), .B(round_reg[1128]), .Z(n52499) );
  XOR U53160 ( .A(round_reg[168]), .B(n52500), .Z(n52498) );
  XOR U53161 ( .A(round_reg[808]), .B(round_reg[488]), .Z(n52500) );
  XOR U53162 ( .A(round_reg[1557]), .B(n52501), .Z(n50058) );
  XNOR U53163 ( .A(n52502), .B(n50169), .Z(n45722) );
  XNOR U53164 ( .A(round_reg[152]), .B(n51145), .Z(n50169) );
  NOR U53165 ( .A(n50170), .B(n50062), .Z(n52502) );
  XOR U53166 ( .A(round_reg[961]), .B(n51347), .Z(n50062) );
  XNOR U53167 ( .A(n52268), .B(n52300), .Z(n51347) );
  XNOR U53168 ( .A(n52503), .B(n52504), .Z(n52300) );
  XNOR U53169 ( .A(round_reg[1345]), .B(round_reg[1025]), .Z(n52504) );
  XOR U53170 ( .A(round_reg[385]), .B(n52505), .Z(n52503) );
  XOR U53171 ( .A(round_reg[705]), .B(round_reg[65]), .Z(n52505) );
  XNOR U53172 ( .A(n52506), .B(n52507), .Z(n52268) );
  XNOR U53173 ( .A(round_reg[1536]), .B(round_reg[1216]), .Z(n52507) );
  XOR U53174 ( .A(round_reg[256]), .B(n52508), .Z(n52506) );
  XOR U53175 ( .A(round_reg[896]), .B(round_reg[576]), .Z(n52508) );
  XNOR U53176 ( .A(round_reg[1401]), .B(n51177), .Z(n50170) );
  XOR U53177 ( .A(n44534), .B(n52509), .Z(n52488) );
  XOR U53178 ( .A(n45164), .B(n47413), .Z(n52509) );
  XNOR U53179 ( .A(n52510), .B(n50163), .Z(n47413) );
  XNOR U53180 ( .A(round_reg[93]), .B(n51781), .Z(n50163) );
  ANDN U53181 ( .B(n50065), .A(n49803), .Z(n52510) );
  XOR U53182 ( .A(round_reg[1265]), .B(n48935), .Z(n49803) );
  XNOR U53183 ( .A(n52511), .B(n52512), .Z(n48935) );
  XOR U53184 ( .A(round_reg[1338]), .B(n51609), .Z(n50065) );
  IV U53185 ( .A(n50110), .Z(n51609) );
  XNOR U53186 ( .A(n52513), .B(n52514), .Z(n52271) );
  XNOR U53187 ( .A(round_reg[122]), .B(round_reg[1082]), .Z(n52514) );
  XOR U53188 ( .A(round_reg[1402]), .B(n52515), .Z(n52513) );
  XOR U53189 ( .A(round_reg[762]), .B(round_reg[442]), .Z(n52515) );
  XNOR U53190 ( .A(n52517), .B(n50166), .Z(n45164) );
  XOR U53191 ( .A(round_reg[211]), .B(n52123), .Z(n50166) );
  IV U53192 ( .A(n52303), .Z(n52123) );
  NOR U53193 ( .A(n50165), .B(n48313), .Z(n52517) );
  XNOR U53194 ( .A(n52518), .B(n50172), .Z(n44534) );
  XOR U53195 ( .A(round_reg[259]), .B(n48514), .Z(n50172) );
  XNOR U53196 ( .A(n52519), .B(n52301), .Z(n48514) );
  XOR U53197 ( .A(n52520), .B(n52521), .Z(n52301) );
  XNOR U53198 ( .A(round_reg[1474]), .B(round_reg[1154]), .Z(n52521) );
  XOR U53199 ( .A(round_reg[194]), .B(n52522), .Z(n52520) );
  XOR U53200 ( .A(round_reg[834]), .B(round_reg[514]), .Z(n52522) );
  ANDN U53201 ( .B(n50067), .A(n47746), .Z(n52518) );
  XNOR U53202 ( .A(round_reg[1103]), .B(n50859), .Z(n47746) );
  IV U53203 ( .A(n52523), .Z(n50859) );
  XOR U53204 ( .A(round_reg[1492]), .B(n50231), .Z(n50067) );
  IV U53205 ( .A(n49608), .Z(n50231) );
  XOR U53206 ( .A(n52524), .B(n52525), .Z(n46291) );
  XOR U53207 ( .A(n43852), .B(n46028), .Z(n52525) );
  XOR U53208 ( .A(n52526), .B(n52119), .Z(n46028) );
  XNOR U53209 ( .A(round_reg[1053]), .B(n51781), .Z(n52119) );
  IV U53210 ( .A(n51456), .Z(n51781) );
  XOR U53211 ( .A(n52527), .B(n52528), .Z(n51456) );
  AND U53212 ( .A(n48609), .B(n50048), .Z(n52526) );
  XOR U53213 ( .A(round_reg[685]), .B(n52089), .Z(n50048) );
  XNOR U53214 ( .A(round_reg[619]), .B(n48452), .Z(n48609) );
  XNOR U53215 ( .A(n52529), .B(n52530), .Z(n48452) );
  XNOR U53216 ( .A(n52531), .B(n47429), .Z(n43852) );
  XNOR U53217 ( .A(round_reg[1102]), .B(n50853), .Z(n47429) );
  ANDN U53218 ( .B(n47430), .A(n48617), .Z(n52531) );
  XNOR U53219 ( .A(round_reg[332]), .B(n50933), .Z(n48617) );
  IV U53220 ( .A(n52176), .Z(n50933) );
  XOR U53221 ( .A(n52532), .B(n52533), .Z(n52458) );
  XNOR U53222 ( .A(round_reg[1547]), .B(round_reg[1227]), .Z(n52533) );
  XOR U53223 ( .A(round_reg[267]), .B(n52534), .Z(n52532) );
  XOR U53224 ( .A(round_reg[907]), .B(round_reg[587]), .Z(n52534) );
  XOR U53225 ( .A(n43107), .B(n52536), .Z(n52524) );
  XOR U53226 ( .A(n43292), .B(n46130), .Z(n52536) );
  XNOR U53227 ( .A(n52537), .B(n47420), .Z(n46130) );
  XNOR U53228 ( .A(round_reg[1192]), .B(n52538), .Z(n47420) );
  XOR U53229 ( .A(round_reg[447]), .B(n51703), .Z(n48620) );
  XOR U53230 ( .A(round_reg[809]), .B(n52181), .Z(n47421) );
  IV U53231 ( .A(n49947), .Z(n52181) );
  XOR U53232 ( .A(n52539), .B(n52540), .Z(n49947) );
  XNOR U53233 ( .A(n52541), .B(n47433), .Z(n43292) );
  XNOR U53234 ( .A(round_reg[1264]), .B(n51953), .Z(n47433) );
  ANDN U53235 ( .B(n47434), .A(n48606), .Z(n52541) );
  XNOR U53236 ( .A(round_reg[453]), .B(n51293), .Z(n48606) );
  IV U53237 ( .A(n50998), .Z(n51293) );
  XOR U53238 ( .A(n52542), .B(n52543), .Z(n50998) );
  XOR U53239 ( .A(round_reg[842]), .B(n50852), .Z(n47434) );
  XNOR U53240 ( .A(n52544), .B(n52342), .Z(n50852) );
  XOR U53241 ( .A(n52545), .B(n52546), .Z(n52342) );
  XNOR U53242 ( .A(round_reg[137]), .B(round_reg[1097]), .Z(n52546) );
  XOR U53243 ( .A(round_reg[1417]), .B(n52547), .Z(n52545) );
  XOR U53244 ( .A(round_reg[777]), .B(round_reg[457]), .Z(n52547) );
  XNOR U53245 ( .A(n52548), .B(n47425), .Z(n43107) );
  XNOR U53246 ( .A(round_reg[960]), .B(n50457), .Z(n47425) );
  IV U53247 ( .A(n51026), .Z(n50457) );
  XOR U53248 ( .A(n52325), .B(n52425), .Z(n51026) );
  XNOR U53249 ( .A(n52549), .B(n52550), .Z(n52425) );
  XNOR U53250 ( .A(round_reg[1344]), .B(round_reg[1024]), .Z(n52550) );
  XOR U53251 ( .A(round_reg[384]), .B(n52551), .Z(n52549) );
  XOR U53252 ( .A(round_reg[704]), .B(round_reg[64]), .Z(n52551) );
  XOR U53253 ( .A(n52552), .B(n52553), .Z(n52325) );
  XNOR U53254 ( .A(round_reg[1599]), .B(round_reg[1279]), .Z(n52553) );
  XOR U53255 ( .A(round_reg[319]), .B(n52554), .Z(n52552) );
  XOR U53256 ( .A(round_reg[959]), .B(round_reg[639]), .Z(n52554) );
  XNOR U53257 ( .A(round_reg[551]), .B(n51947), .Z(n48614) );
  XOR U53258 ( .A(round_reg[913]), .B(n52148), .Z(n47426) );
  XNOR U53259 ( .A(n52555), .B(n50165), .Z(n50056) );
  XNOR U53260 ( .A(round_reg[1431]), .B(n49833), .Z(n50165) );
  IV U53261 ( .A(n52113), .Z(n49833) );
  ANDN U53262 ( .B(n48313), .A(n48315), .Z(n52555) );
  XOR U53263 ( .A(round_reg[686]), .B(n50718), .Z(n48315) );
  XNOR U53264 ( .A(n52556), .B(n52038), .Z(n50718) );
  XNOR U53265 ( .A(n52557), .B(n52558), .Z(n52038) );
  XNOR U53266 ( .A(round_reg[110]), .B(round_reg[1070]), .Z(n52558) );
  XOR U53267 ( .A(round_reg[1390]), .B(n52559), .Z(n52557) );
  XOR U53268 ( .A(round_reg[750]), .B(round_reg[430]), .Z(n52559) );
  XOR U53269 ( .A(round_reg[1054]), .B(n49606), .Z(n48313) );
  XOR U53270 ( .A(n51125), .B(n44859), .Z(n41404) );
  XOR U53271 ( .A(n52127), .B(n51151), .Z(n44859) );
  XNOR U53272 ( .A(n52560), .B(n52561), .Z(n51151) );
  XNOR U53273 ( .A(n47386), .B(n47628), .Z(n52561) );
  XNOR U53274 ( .A(n52562), .B(n48854), .Z(n47628) );
  XNOR U53275 ( .A(round_reg[1346]), .B(n49989), .Z(n48854) );
  XOR U53276 ( .A(round_reg[970]), .B(n52336), .Z(n49150) );
  XNOR U53277 ( .A(round_reg[923]), .B(n51009), .Z(n49282) );
  XNOR U53278 ( .A(n52117), .B(n52563), .Z(n51009) );
  XNOR U53279 ( .A(n52564), .B(n52565), .Z(n52117) );
  XNOR U53280 ( .A(round_reg[27]), .B(round_reg[1307]), .Z(n52565) );
  XOR U53281 ( .A(round_reg[347]), .B(n52566), .Z(n52564) );
  XOR U53282 ( .A(round_reg[987]), .B(round_reg[667]), .Z(n52566) );
  XOR U53283 ( .A(n52567), .B(n48850), .Z(n47386) );
  XOR U53284 ( .A(round_reg[1566]), .B(n51486), .Z(n48850) );
  IV U53285 ( .A(n50835), .Z(n51486) );
  NOR U53286 ( .A(n50178), .B(n49140), .Z(n52567) );
  XNOR U53287 ( .A(round_reg[1202]), .B(n51466), .Z(n49140) );
  XOR U53288 ( .A(round_reg[819]), .B(n48942), .Z(n50178) );
  XOR U53289 ( .A(n52455), .B(n52570), .Z(n48942) );
  XOR U53290 ( .A(n52571), .B(n52572), .Z(n52455) );
  XNOR U53291 ( .A(round_reg[114]), .B(round_reg[1074]), .Z(n52572) );
  XOR U53292 ( .A(round_reg[1394]), .B(n52573), .Z(n52571) );
  XOR U53293 ( .A(round_reg[754]), .B(round_reg[434]), .Z(n52573) );
  XOR U53294 ( .A(n49136), .B(n52574), .Z(n52560) );
  XOR U53295 ( .A(n44873), .B(n46402), .Z(n52574) );
  XNOR U53296 ( .A(n52575), .B(n48842), .Z(n46402) );
  IV U53297 ( .A(n49143), .Z(n48842) );
  XOR U53298 ( .A(round_reg[1440]), .B(n52000), .Z(n49143) );
  NOR U53299 ( .A(n51111), .B(n49142), .Z(n52575) );
  XNOR U53300 ( .A(round_reg[1063]), .B(n50224), .Z(n49142) );
  XOR U53301 ( .A(round_reg[695]), .B(n50507), .Z(n51111) );
  XOR U53302 ( .A(n52576), .B(n48845), .Z(n44873) );
  XOR U53303 ( .A(round_reg[1283]), .B(n51985), .Z(n48845) );
  NOR U53304 ( .A(n49279), .B(n49148), .Z(n52576) );
  XNOR U53305 ( .A(round_reg[1274]), .B(n52384), .Z(n49148) );
  IV U53306 ( .A(n51117), .Z(n49279) );
  XOR U53307 ( .A(round_reg[852]), .B(n49608), .Z(n51117) );
  XOR U53308 ( .A(n52579), .B(n48858), .Z(n49136) );
  XOR U53309 ( .A(round_reg[1501]), .B(n51032), .Z(n48858) );
  NOR U53310 ( .A(n49426), .B(n49146), .Z(n52579) );
  XOR U53311 ( .A(round_reg[1112]), .B(n51145), .Z(n49146) );
  XOR U53312 ( .A(n52580), .B(n52581), .Z(n51145) );
  IV U53313 ( .A(n51113), .Z(n49426) );
  XOR U53314 ( .A(round_reg[709]), .B(n49074), .Z(n51113) );
  XOR U53315 ( .A(n52582), .B(n52583), .Z(n52127) );
  XNOR U53316 ( .A(n48286), .B(n43643), .Z(n52583) );
  XNOR U53317 ( .A(n52584), .B(n48300), .Z(n43643) );
  XOR U53318 ( .A(round_reg[464]), .B(n50735), .Z(n48300) );
  ANDN U53319 ( .B(n49267), .A(n48299), .Z(n52584) );
  XOR U53320 ( .A(n52587), .B(n48688), .Z(n48286) );
  XOR U53321 ( .A(round_reg[630]), .B(n50106), .Z(n48688) );
  ANDN U53322 ( .B(n48689), .A(n49264), .Z(n52587) );
  XNOR U53323 ( .A(round_reg[1441]), .B(n49175), .Z(n49264) );
  XNOR U53324 ( .A(n52588), .B(n52589), .Z(n49175) );
  XNOR U53325 ( .A(round_reg[221]), .B(n51032), .Z(n48689) );
  XNOR U53326 ( .A(n52116), .B(n51779), .Z(n51032) );
  XNOR U53327 ( .A(n52590), .B(n52591), .Z(n51779) );
  XNOR U53328 ( .A(round_reg[1565]), .B(round_reg[1245]), .Z(n52591) );
  XOR U53329 ( .A(round_reg[285]), .B(n52592), .Z(n52590) );
  XOR U53330 ( .A(round_reg[925]), .B(round_reg[605]), .Z(n52592) );
  XOR U53331 ( .A(n52593), .B(n52594), .Z(n52116) );
  XNOR U53332 ( .A(round_reg[1436]), .B(round_reg[1116]), .Z(n52594) );
  XOR U53333 ( .A(round_reg[156]), .B(n52595), .Z(n52593) );
  XOR U53334 ( .A(round_reg[796]), .B(round_reg[476]), .Z(n52595) );
  XNOR U53335 ( .A(n44548), .B(n52596), .Z(n52582) );
  XOR U53336 ( .A(n44109), .B(n46723), .Z(n52596) );
  XOR U53337 ( .A(n52597), .B(n48294), .Z(n46723) );
  XOR U53338 ( .A(round_reg[343]), .B(n48554), .Z(n48294) );
  XNOR U53339 ( .A(n52598), .B(n52580), .Z(n48554) );
  XOR U53340 ( .A(n52599), .B(n52600), .Z(n52580) );
  XNOR U53341 ( .A(round_reg[1367]), .B(round_reg[1047]), .Z(n52600) );
  XOR U53342 ( .A(round_reg[407]), .B(n52601), .Z(n52599) );
  XOR U53343 ( .A(round_reg[87]), .B(round_reg[727]), .Z(n52601) );
  NOR U53344 ( .A(n49270), .B(n48293), .Z(n52597) );
  XNOR U53345 ( .A(round_reg[269]), .B(n51093), .Z(n48293) );
  XNOR U53346 ( .A(n52602), .B(n52603), .Z(n51093) );
  XOR U53347 ( .A(round_reg[1502]), .B(n51050), .Z(n49270) );
  XNOR U53348 ( .A(n52604), .B(n48304), .Z(n44109) );
  XNOR U53349 ( .A(round_reg[562]), .B(n51466), .Z(n48304) );
  ANDN U53350 ( .B(n48303), .A(n51128), .Z(n52604) );
  XOR U53351 ( .A(round_reg[1347]), .B(n52605), .Z(n51128) );
  XOR U53352 ( .A(round_reg[162]), .B(n51051), .Z(n48303) );
  IV U53353 ( .A(n51595), .Z(n51051) );
  XOR U53354 ( .A(n52607), .B(n52608), .Z(n51916) );
  XNOR U53355 ( .A(round_reg[1506]), .B(round_reg[1186]), .Z(n52608) );
  XOR U53356 ( .A(round_reg[226]), .B(n52609), .Z(n52607) );
  XOR U53357 ( .A(round_reg[866]), .B(round_reg[546]), .Z(n52609) );
  XOR U53358 ( .A(n52610), .B(n48862), .Z(n44548) );
  XOR U53359 ( .A(round_reg[394]), .B(n52004), .Z(n48862) );
  NOR U53360 ( .A(n51122), .B(n51106), .Z(n52610) );
  XNOR U53361 ( .A(round_reg[1567]), .B(n50453), .Z(n51106) );
  XNOR U53362 ( .A(n52611), .B(n52612), .Z(n50453) );
  XNOR U53363 ( .A(round_reg[17]), .B(n51325), .Z(n51122) );
  XOR U53364 ( .A(n52613), .B(n48299), .Z(n51125) );
  XOR U53365 ( .A(round_reg[103]), .B(n52614), .Z(n48299) );
  ANDN U53366 ( .B(n49245), .A(n49267), .Z(n52613) );
  XOR U53367 ( .A(round_reg[1284]), .B(n51538), .Z(n49267) );
  XOR U53368 ( .A(round_reg[1275]), .B(n49897), .Z(n49245) );
  IV U53369 ( .A(n52615), .Z(n49897) );
  XNOR U53370 ( .A(n42783), .B(n52616), .Z(n52287) );
  XNOR U53371 ( .A(n36363), .B(n38660), .Z(n52616) );
  XNOR U53372 ( .A(n52617), .B(n44244), .Z(n38660) );
  XOR U53373 ( .A(n46630), .B(n46758), .Z(n44244) );
  IV U53374 ( .A(n47674), .Z(n46758) );
  XOR U53375 ( .A(n47573), .B(n49070), .Z(n47674) );
  XNOR U53376 ( .A(n52618), .B(n52619), .Z(n49070) );
  XNOR U53377 ( .A(n45725), .B(n41736), .Z(n52619) );
  XOR U53378 ( .A(n52620), .B(n45870), .Z(n41736) );
  XOR U53379 ( .A(round_reg[1168]), .B(n52621), .Z(n45870) );
  ANDN U53380 ( .B(n45871), .A(n47677), .Z(n52620) );
  XNOR U53381 ( .A(round_reg[423]), .B(n52614), .Z(n47677) );
  IV U53382 ( .A(n50224), .Z(n52614) );
  XNOR U53383 ( .A(n52622), .B(n52623), .Z(n50224) );
  XOR U53384 ( .A(round_reg[785]), .B(n51342), .Z(n45871) );
  XOR U53385 ( .A(n52624), .B(n52625), .Z(n51342) );
  XOR U53386 ( .A(n52626), .B(n50716), .Z(n45725) );
  XOR U53387 ( .A(round_reg[1240]), .B(n48962), .Z(n50716) );
  ANDN U53388 ( .B(n45884), .A(n48186), .Z(n52626) );
  XNOR U53389 ( .A(round_reg[493]), .B(n51467), .Z(n48186) );
  IV U53390 ( .A(n48558), .Z(n51467) );
  XOR U53391 ( .A(n52627), .B(n52628), .Z(n51466) );
  XNOR U53392 ( .A(n44268), .B(n52629), .Z(n52618) );
  XOR U53393 ( .A(n44853), .B(n42538), .Z(n52629) );
  XOR U53394 ( .A(n52630), .B(n45876), .Z(n42538) );
  XOR U53395 ( .A(round_reg[1029]), .B(n51437), .Z(n45876) );
  IV U53396 ( .A(n49074), .Z(n51437) );
  XNOR U53397 ( .A(n51454), .B(n52190), .Z(n49074) );
  XNOR U53398 ( .A(n52631), .B(n52632), .Z(n52190) );
  XNOR U53399 ( .A(round_reg[324]), .B(round_reg[1284]), .Z(n52632) );
  XOR U53400 ( .A(round_reg[4]), .B(n52633), .Z(n52631) );
  XOR U53401 ( .A(round_reg[964]), .B(round_reg[644]), .Z(n52633) );
  XOR U53402 ( .A(n52634), .B(n52635), .Z(n51454) );
  XNOR U53403 ( .A(round_reg[133]), .B(round_reg[1093]), .Z(n52635) );
  XOR U53404 ( .A(round_reg[1413]), .B(n52636), .Z(n52634) );
  XOR U53405 ( .A(round_reg[773]), .B(round_reg[453]), .Z(n52636) );
  ANDN U53406 ( .B(n45875), .A(n46760), .Z(n52630) );
  XOR U53407 ( .A(round_reg[595]), .B(n50480), .Z(n46760) );
  XOR U53408 ( .A(n52637), .B(n52638), .Z(n50480) );
  XNOR U53409 ( .A(round_reg[661]), .B(n51961), .Z(n45875) );
  XOR U53410 ( .A(n52639), .B(n50725), .Z(n44853) );
  XOR U53411 ( .A(round_reg[1142]), .B(n49795), .Z(n50725) );
  ANDN U53412 ( .B(n45880), .A(n49573), .Z(n52639) );
  XOR U53413 ( .A(n52642), .B(n50722), .Z(n44268) );
  IV U53414 ( .A(n50710), .Z(n50722) );
  XOR U53415 ( .A(round_reg[1000]), .B(n48442), .Z(n50710) );
  XNOR U53416 ( .A(n52540), .B(n52643), .Z(n48442) );
  XOR U53417 ( .A(n52644), .B(n52645), .Z(n52540) );
  XNOR U53418 ( .A(round_reg[1064]), .B(round_reg[104]), .Z(n52645) );
  XOR U53419 ( .A(round_reg[1384]), .B(n52646), .Z(n52644) );
  XOR U53420 ( .A(round_reg[744]), .B(round_reg[424]), .Z(n52646) );
  ANDN U53421 ( .B(n47636), .A(n47638), .Z(n52642) );
  XOR U53422 ( .A(round_reg[527]), .B(n50401), .Z(n47638) );
  XNOR U53423 ( .A(round_reg[953]), .B(n51672), .Z(n47636) );
  XOR U53424 ( .A(n52647), .B(n52648), .Z(n47573) );
  XOR U53425 ( .A(n46177), .B(n48370), .Z(n52648) );
  XOR U53426 ( .A(n52649), .B(n48384), .Z(n48370) );
  XOR U53427 ( .A(round_reg[422]), .B(n49280), .Z(n48384) );
  ANDN U53428 ( .B(n46903), .A(n46904), .Z(n52649) );
  XOR U53429 ( .A(round_reg[1595]), .B(n52615), .Z(n46904) );
  XOR U53430 ( .A(n52334), .B(n52650), .Z(n52615) );
  XOR U53431 ( .A(n52651), .B(n52652), .Z(n52334) );
  XNOR U53432 ( .A(round_reg[1530]), .B(round_reg[1210]), .Z(n52652) );
  XOR U53433 ( .A(round_reg[250]), .B(n52653), .Z(n52651) );
  XOR U53434 ( .A(round_reg[890]), .B(round_reg[570]), .Z(n52653) );
  XNOR U53435 ( .A(round_reg[45]), .B(n50120), .Z(n46903) );
  IV U53436 ( .A(n52089), .Z(n50120) );
  XNOR U53437 ( .A(n52655), .B(n52656), .Z(n52395) );
  XNOR U53438 ( .A(round_reg[109]), .B(round_reg[1069]), .Z(n52656) );
  XOR U53439 ( .A(round_reg[1389]), .B(n52657), .Z(n52655) );
  XOR U53440 ( .A(round_reg[749]), .B(round_reg[429]), .Z(n52657) );
  XNOR U53441 ( .A(n52658), .B(n48378), .Z(n46177) );
  XOR U53442 ( .A(round_reg[371]), .B(n50136), .Z(n48378) );
  XOR U53443 ( .A(n52659), .B(n52660), .Z(n52627) );
  XNOR U53444 ( .A(round_reg[1586]), .B(round_reg[1266]), .Z(n52660) );
  XOR U53445 ( .A(round_reg[306]), .B(n52661), .Z(n52659) );
  XOR U53446 ( .A(round_reg[946]), .B(round_reg[626]), .Z(n52661) );
  ANDN U53447 ( .B(n46897), .A(n46898), .Z(n52658) );
  XOR U53448 ( .A(round_reg[1530]), .B(n50727), .Z(n46898) );
  IV U53449 ( .A(n49861), .Z(n50727) );
  XOR U53450 ( .A(n52663), .B(n52284), .Z(n49861) );
  XNOR U53451 ( .A(n52664), .B(n52665), .Z(n52284) );
  XNOR U53452 ( .A(round_reg[1594]), .B(round_reg[1274]), .Z(n52665) );
  XOR U53453 ( .A(round_reg[314]), .B(n52666), .Z(n52664) );
  XOR U53454 ( .A(round_reg[954]), .B(round_reg[634]), .Z(n52666) );
  XNOR U53455 ( .A(round_reg[297]), .B(n51520), .Z(n46897) );
  XOR U53456 ( .A(n47326), .B(n52667), .Z(n52647) );
  XOR U53457 ( .A(n47157), .B(n43545), .Z(n52667) );
  XNOR U53458 ( .A(n52668), .B(n48375), .Z(n43545) );
  XOR U53459 ( .A(round_reg[594]), .B(n50755), .Z(n48375) );
  ANDN U53460 ( .B(n46907), .A(n46908), .Z(n52668) );
  XOR U53461 ( .A(round_reg[1469]), .B(n49992), .Z(n46908) );
  XNOR U53462 ( .A(n52419), .B(n52669), .Z(n49992) );
  XOR U53463 ( .A(n52670), .B(n52671), .Z(n52419) );
  XNOR U53464 ( .A(round_reg[1533]), .B(round_reg[1213]), .Z(n52671) );
  XOR U53465 ( .A(round_reg[253]), .B(n52672), .Z(n52670) );
  XOR U53466 ( .A(round_reg[893]), .B(round_reg[573]), .Z(n52672) );
  XOR U53467 ( .A(round_reg[249]), .B(n49836), .Z(n46907) );
  XNOR U53468 ( .A(n52673), .B(n49433), .Z(n47157) );
  XOR U53469 ( .A(round_reg[492]), .B(n48365), .Z(n49433) );
  ANDN U53470 ( .B(n47570), .A(n47571), .Z(n52673) );
  XOR U53471 ( .A(round_reg[1312]), .B(n50834), .Z(n47571) );
  XOR U53472 ( .A(round_reg[67]), .B(n52605), .Z(n47570) );
  XNOR U53473 ( .A(n52674), .B(n49994), .Z(n47326) );
  XNOR U53474 ( .A(round_reg[526]), .B(n50772), .Z(n49994) );
  ANDN U53475 ( .B(n47101), .A(n47102), .Z(n52674) );
  XOR U53476 ( .A(round_reg[1375]), .B(n52675), .Z(n47102) );
  XNOR U53477 ( .A(round_reg[190]), .B(n50728), .Z(n47101) );
  XNOR U53478 ( .A(n52676), .B(n52677), .Z(n50728) );
  XNOR U53479 ( .A(n52678), .B(n45880), .Z(n46630) );
  XOR U53480 ( .A(round_reg[739]), .B(n51624), .Z(n45880) );
  XNOR U53481 ( .A(n52679), .B(n52680), .Z(n52345) );
  XNOR U53482 ( .A(round_reg[1443]), .B(round_reg[1123]), .Z(n52680) );
  XOR U53483 ( .A(round_reg[163]), .B(n52681), .Z(n52679) );
  XOR U53484 ( .A(round_reg[803]), .B(round_reg[483]), .Z(n52681) );
  AND U53485 ( .A(n49574), .B(n49573), .Z(n52678) );
  XOR U53486 ( .A(round_reg[372]), .B(n50440), .Z(n49573) );
  XOR U53487 ( .A(n52132), .B(n52397), .Z(n50440) );
  XNOR U53488 ( .A(n52683), .B(n52684), .Z(n52397) );
  XNOR U53489 ( .A(round_reg[1587]), .B(round_reg[1267]), .Z(n52684) );
  XOR U53490 ( .A(round_reg[307]), .B(n52685), .Z(n52683) );
  XOR U53491 ( .A(round_reg[947]), .B(round_reg[627]), .Z(n52685) );
  XOR U53492 ( .A(n52686), .B(n52687), .Z(n52132) );
  XNOR U53493 ( .A(round_reg[116]), .B(round_reg[1076]), .Z(n52687) );
  XOR U53494 ( .A(round_reg[1396]), .B(n52688), .Z(n52686) );
  XOR U53495 ( .A(round_reg[756]), .B(round_reg[436]), .Z(n52688) );
  XNOR U53496 ( .A(round_reg[298]), .B(n48356), .Z(n49574) );
  XOR U53497 ( .A(n52539), .B(n52306), .Z(n48356) );
  XNOR U53498 ( .A(n52689), .B(n52690), .Z(n52306) );
  XNOR U53499 ( .A(round_reg[1322]), .B(round_reg[1002]), .Z(n52690) );
  XOR U53500 ( .A(round_reg[362]), .B(n52691), .Z(n52689) );
  XOR U53501 ( .A(round_reg[682]), .B(round_reg[42]), .Z(n52691) );
  XOR U53502 ( .A(n52692), .B(n52693), .Z(n52539) );
  XNOR U53503 ( .A(round_reg[1513]), .B(round_reg[1193]), .Z(n52693) );
  XOR U53504 ( .A(round_reg[233]), .B(n52694), .Z(n52692) );
  XOR U53505 ( .A(round_reg[873]), .B(round_reg[553]), .Z(n52694) );
  ANDN U53506 ( .B(n43068), .A(n43066), .Z(n52617) );
  XOR U53507 ( .A(n45621), .B(n52247), .Z(n43066) );
  XNOR U53508 ( .A(n52695), .B(n49107), .Z(n52247) );
  XOR U53509 ( .A(round_reg[1335]), .B(n50507), .Z(n50464) );
  XOR U53510 ( .A(n46691), .B(n48802), .Z(n45621) );
  XNOR U53511 ( .A(n52698), .B(n52699), .Z(n48802) );
  XOR U53512 ( .A(n43320), .B(n43873), .Z(n52699) );
  XOR U53513 ( .A(n52700), .B(n49097), .Z(n43873) );
  XOR U53514 ( .A(round_reg[683]), .B(n50823), .Z(n49097) );
  ANDN U53515 ( .B(n49098), .A(n51574), .Z(n52700) );
  XNOR U53516 ( .A(round_reg[208]), .B(n51516), .Z(n51574) );
  XOR U53517 ( .A(round_reg[617]), .B(n52701), .Z(n49098) );
  XNOR U53518 ( .A(n52702), .B(n50268), .Z(n43320) );
  XOR U53519 ( .A(round_reg[761]), .B(n51177), .Z(n50268) );
  XOR U53520 ( .A(n52703), .B(n52663), .Z(n51177) );
  XNOR U53521 ( .A(n52704), .B(n52705), .Z(n52663) );
  XNOR U53522 ( .A(round_reg[1465]), .B(round_reg[1145]), .Z(n52705) );
  XOR U53523 ( .A(round_reg[185]), .B(n52706), .Z(n52704) );
  XOR U53524 ( .A(round_reg[825]), .B(round_reg[505]), .Z(n52706) );
  ANDN U53525 ( .B(n50269), .A(n51578), .Z(n52702) );
  XOR U53526 ( .A(round_reg[256]), .B(n51199), .Z(n51578) );
  XOR U53527 ( .A(round_reg[330]), .B(n52336), .Z(n50269) );
  XOR U53528 ( .A(n52707), .B(n52708), .Z(n52336) );
  XOR U53529 ( .A(n48435), .B(n52709), .Z(n52698) );
  XOR U53530 ( .A(n49090), .B(n47164), .Z(n52709) );
  XNOR U53531 ( .A(n52710), .B(n49102), .Z(n47164) );
  XNOR U53532 ( .A(round_reg[807]), .B(n52034), .Z(n49102) );
  NOR U53533 ( .A(n49103), .B(n51571), .Z(n52710) );
  XNOR U53534 ( .A(round_reg[4]), .B(n51538), .Z(n51571) );
  XOR U53535 ( .A(round_reg[445]), .B(n50949), .Z(n49103) );
  XNOR U53536 ( .A(n52711), .B(n49106), .Z(n49090) );
  XOR U53537 ( .A(round_reg[840]), .B(n50947), .Z(n49106) );
  ANDN U53538 ( .B(n49107), .A(n51581), .Z(n52711) );
  XOR U53539 ( .A(round_reg[90]), .B(n51468), .Z(n51581) );
  XOR U53540 ( .A(round_reg[451]), .B(n50421), .Z(n49107) );
  IV U53541 ( .A(n52028), .Z(n50421) );
  XNOR U53542 ( .A(n52712), .B(n52713), .Z(n52191) );
  XNOR U53543 ( .A(round_reg[1475]), .B(round_reg[1155]), .Z(n52713) );
  XOR U53544 ( .A(round_reg[195]), .B(n52714), .Z(n52712) );
  XOR U53545 ( .A(round_reg[835]), .B(round_reg[515]), .Z(n52714) );
  XNOR U53546 ( .A(n52716), .B(n49110), .Z(n48435) );
  XOR U53547 ( .A(round_reg[911]), .B(n51346), .Z(n49110) );
  XNOR U53548 ( .A(n52717), .B(n52207), .Z(n51346) );
  XOR U53549 ( .A(n52718), .B(n52719), .Z(n52207) );
  XNOR U53550 ( .A(round_reg[15]), .B(round_reg[1295]), .Z(n52719) );
  XOR U53551 ( .A(round_reg[335]), .B(n52720), .Z(n52718) );
  XOR U53552 ( .A(round_reg[975]), .B(round_reg[655]), .Z(n52720) );
  ANDN U53553 ( .B(n49111), .A(n52252), .Z(n52716) );
  XOR U53554 ( .A(round_reg[149]), .B(n50232), .Z(n52252) );
  XOR U53555 ( .A(n52721), .B(n52722), .Z(n50232) );
  XNOR U53556 ( .A(round_reg[549]), .B(n52001), .Z(n49111) );
  XNOR U53557 ( .A(n52723), .B(n52724), .Z(n46691) );
  XNOR U53558 ( .A(n47464), .B(n46241), .Z(n52724) );
  XOR U53559 ( .A(n52725), .B(n50782), .Z(n46241) );
  XOR U53560 ( .A(round_reg[89]), .B(n51656), .Z(n50782) );
  IV U53561 ( .A(n51101), .Z(n51656) );
  XOR U53562 ( .A(n52726), .B(n52727), .Z(n51101) );
  ANDN U53563 ( .B(n51079), .A(n51563), .Z(n52725) );
  XOR U53564 ( .A(round_reg[1261]), .B(n51839), .Z(n51563) );
  IV U53565 ( .A(n50153), .Z(n51839) );
  XOR U53566 ( .A(n52728), .B(n52729), .Z(n50153) );
  XOR U53567 ( .A(round_reg[1334]), .B(n51020), .Z(n51079) );
  IV U53568 ( .A(n49902), .Z(n51020) );
  XOR U53569 ( .A(n52730), .B(n50264), .Z(n47464) );
  XNOR U53570 ( .A(round_reg[148]), .B(n51789), .Z(n50264) );
  ANDN U53571 ( .B(n51084), .A(n51560), .Z(n52730) );
  XNOR U53572 ( .A(round_reg[1021]), .B(n49800), .Z(n51560) );
  XOR U53573 ( .A(round_reg[1397]), .B(n51526), .Z(n51084) );
  XOR U53574 ( .A(n52731), .B(n52732), .Z(n51526) );
  XOR U53575 ( .A(n51075), .B(n52733), .Z(n52723) );
  XOR U53576 ( .A(n45396), .B(n46714), .Z(n52733) );
  XNOR U53577 ( .A(n52734), .B(n50261), .Z(n46714) );
  XNOR U53578 ( .A(round_reg[319]), .B(n52065), .Z(n50261) );
  IV U53579 ( .A(n52313), .Z(n52065) );
  ANDN U53580 ( .B(n51088), .A(n51556), .Z(n52734) );
  XNOR U53581 ( .A(round_reg[1099]), .B(n50138), .Z(n51556) );
  IV U53582 ( .A(n51434), .Z(n50138) );
  XNOR U53583 ( .A(n52735), .B(n52736), .Z(n51921) );
  XNOR U53584 ( .A(round_reg[1483]), .B(round_reg[1163]), .Z(n52736) );
  XOR U53585 ( .A(round_reg[203]), .B(n52737), .Z(n52735) );
  XOR U53586 ( .A(round_reg[843]), .B(round_reg[523]), .Z(n52737) );
  XNOR U53587 ( .A(n52738), .B(n52739), .Z(n52708) );
  XNOR U53588 ( .A(round_reg[1354]), .B(round_reg[1034]), .Z(n52739) );
  XOR U53589 ( .A(round_reg[394]), .B(n52740), .Z(n52738) );
  XOR U53590 ( .A(round_reg[74]), .B(round_reg[714]), .Z(n52740) );
  XOR U53591 ( .A(round_reg[1488]), .B(n52621), .Z(n51088) );
  IV U53592 ( .A(n51516), .Z(n52621) );
  XOR U53593 ( .A(n52369), .B(n52741), .Z(n51516) );
  XOR U53594 ( .A(n52742), .B(n52743), .Z(n52369) );
  XNOR U53595 ( .A(round_reg[1423]), .B(round_reg[1103]), .Z(n52743) );
  XOR U53596 ( .A(round_reg[143]), .B(n52744), .Z(n52742) );
  XOR U53597 ( .A(round_reg[783]), .B(round_reg[463]), .Z(n52744) );
  XNOR U53598 ( .A(n52745), .B(n50250), .Z(n45396) );
  XNOR U53599 ( .A(round_reg[3]), .B(n51985), .Z(n50250) );
  NOR U53600 ( .A(n51081), .B(n51566), .Z(n52745) );
  XNOR U53601 ( .A(round_reg[1189]), .B(n52001), .Z(n51566) );
  IV U53602 ( .A(n52746), .Z(n52001) );
  XOR U53603 ( .A(round_reg[1553]), .B(n51664), .Z(n51081) );
  IV U53604 ( .A(n52148), .Z(n51664) );
  XOR U53605 ( .A(n52747), .B(n52585), .Z(n52148) );
  XNOR U53606 ( .A(n52748), .B(n52749), .Z(n52585) );
  XNOR U53607 ( .A(round_reg[1488]), .B(round_reg[1168]), .Z(n52749) );
  XOR U53608 ( .A(round_reg[208]), .B(n52750), .Z(n52748) );
  XOR U53609 ( .A(round_reg[848]), .B(round_reg[528]), .Z(n52750) );
  XOR U53610 ( .A(n52751), .B(n50254), .Z(n51075) );
  XNOR U53611 ( .A(round_reg[207]), .B(n50401), .Z(n50254) );
  XOR U53612 ( .A(n52752), .B(n52753), .Z(n50401) );
  ANDN U53613 ( .B(n51086), .A(n51554), .Z(n52751) );
  XOR U53614 ( .A(round_reg[1050]), .B(n51468), .Z(n51554) );
  XOR U53615 ( .A(round_reg[1427]), .B(n51698), .Z(n51086) );
  XOR U53616 ( .A(n52754), .B(n52400), .Z(n51698) );
  XNOR U53617 ( .A(n52755), .B(n52756), .Z(n52400) );
  XNOR U53618 ( .A(round_reg[1491]), .B(round_reg[1171]), .Z(n52756) );
  XOR U53619 ( .A(round_reg[211]), .B(n52757), .Z(n52755) );
  XOR U53620 ( .A(round_reg[851]), .B(round_reg[531]), .Z(n52757) );
  XOR U53621 ( .A(n51416), .B(n45308), .Z(n43068) );
  XNOR U53622 ( .A(n46268), .B(n50787), .Z(n45308) );
  XNOR U53623 ( .A(n52758), .B(n52759), .Z(n50787) );
  XNOR U53624 ( .A(n46668), .B(n42330), .Z(n52759) );
  XNOR U53625 ( .A(n52760), .B(n48579), .Z(n42330) );
  XNOR U53626 ( .A(round_reg[624]), .B(n51953), .Z(n48579) );
  IV U53627 ( .A(n50939), .Z(n51953) );
  XNOR U53628 ( .A(n52037), .B(n52761), .Z(n50939) );
  XOR U53629 ( .A(n52762), .B(n52763), .Z(n52037) );
  XNOR U53630 ( .A(round_reg[1519]), .B(round_reg[1199]), .Z(n52763) );
  XOR U53631 ( .A(round_reg[239]), .B(n52764), .Z(n52762) );
  XOR U53632 ( .A(round_reg[879]), .B(round_reg[559]), .Z(n52764) );
  ANDN U53633 ( .B(n48580), .A(n50403), .Z(n52760) );
  XNOR U53634 ( .A(n52765), .B(n48596), .Z(n46668) );
  XNOR U53635 ( .A(round_reg[388]), .B(n50714), .Z(n48596) );
  XNOR U53636 ( .A(round_reg[1561]), .B(n50434), .Z(n50393) );
  XNOR U53637 ( .A(round_reg[11]), .B(n51127), .Z(n48597) );
  IV U53638 ( .A(n51461), .Z(n51127) );
  XOR U53639 ( .A(n52544), .B(n52766), .Z(n51461) );
  XOR U53640 ( .A(n52767), .B(n52768), .Z(n52544) );
  XNOR U53641 ( .A(round_reg[1546]), .B(round_reg[1226]), .Z(n52768) );
  XOR U53642 ( .A(round_reg[266]), .B(n52769), .Z(n52767) );
  XOR U53643 ( .A(round_reg[906]), .B(round_reg[586]), .Z(n52769) );
  XOR U53644 ( .A(n47354), .B(n52770), .Z(n52758) );
  XOR U53645 ( .A(n45617), .B(n47163), .Z(n52770) );
  XNOR U53646 ( .A(n52771), .B(n48588), .Z(n47163) );
  XOR U53647 ( .A(round_reg[556]), .B(n51911), .Z(n48588) );
  AND U53648 ( .A(n50396), .B(n48589), .Z(n52771) );
  XNOR U53649 ( .A(round_reg[156]), .B(n51544), .Z(n48589) );
  IV U53650 ( .A(n50827), .Z(n51544) );
  XOR U53651 ( .A(n52772), .B(n52773), .Z(n50827) );
  XOR U53652 ( .A(round_reg[1405]), .B(n50949), .Z(n50396) );
  XOR U53653 ( .A(n52484), .B(n52774), .Z(n50949) );
  XOR U53654 ( .A(n52775), .B(n52776), .Z(n52484) );
  XNOR U53655 ( .A(round_reg[1340]), .B(round_reg[1020]), .Z(n52776) );
  XOR U53656 ( .A(round_reg[380]), .B(n52777), .Z(n52775) );
  XOR U53657 ( .A(round_reg[700]), .B(round_reg[60]), .Z(n52777) );
  XNOR U53658 ( .A(n52778), .B(n48592), .Z(n45617) );
  XOR U53659 ( .A(round_reg[458]), .B(n50117), .Z(n48592) );
  XNOR U53660 ( .A(n52779), .B(n52780), .Z(n50117) );
  ANDN U53661 ( .B(n48593), .A(n50400), .Z(n52778) );
  XOR U53662 ( .A(round_reg[1342]), .B(n52255), .Z(n50400) );
  IV U53663 ( .A(n50516), .Z(n52255) );
  XNOR U53664 ( .A(n52781), .B(n52782), .Z(n50516) );
  XOR U53665 ( .A(round_reg[97]), .B(n52783), .Z(n48593) );
  XNOR U53666 ( .A(n52784), .B(n48583), .Z(n47354) );
  XOR U53667 ( .A(round_reg[337]), .B(n51325), .Z(n48583) );
  XOR U53668 ( .A(n52741), .B(n52785), .Z(n51325) );
  XOR U53669 ( .A(n52786), .B(n52787), .Z(n52741) );
  XNOR U53670 ( .A(round_reg[1552]), .B(round_reg[1232]), .Z(n52787) );
  XOR U53671 ( .A(round_reg[272]), .B(n52788), .Z(n52786) );
  XOR U53672 ( .A(round_reg[912]), .B(round_reg[592]), .Z(n52788) );
  ANDN U53673 ( .B(n48584), .A(n50406), .Z(n52784) );
  IV U53674 ( .A(n51420), .Z(n50406) );
  XNOR U53675 ( .A(round_reg[1496]), .B(n49789), .Z(n51420) );
  XOR U53676 ( .A(n52171), .B(n51605), .Z(n49789) );
  XNOR U53677 ( .A(n52789), .B(n52790), .Z(n51605) );
  XNOR U53678 ( .A(round_reg[1431]), .B(round_reg[1111]), .Z(n52790) );
  XOR U53679 ( .A(round_reg[151]), .B(n52791), .Z(n52789) );
  XOR U53680 ( .A(round_reg[791]), .B(round_reg[471]), .Z(n52791) );
  XOR U53681 ( .A(n52792), .B(n52793), .Z(n52171) );
  XNOR U53682 ( .A(round_reg[1560]), .B(round_reg[1240]), .Z(n52793) );
  XOR U53683 ( .A(round_reg[280]), .B(n52794), .Z(n52792) );
  XOR U53684 ( .A(round_reg[920]), .B(round_reg[600]), .Z(n52794) );
  XNOR U53685 ( .A(round_reg[263]), .B(n50132), .Z(n48584) );
  XNOR U53686 ( .A(n52795), .B(n51939), .Z(n50132) );
  XNOR U53687 ( .A(n52796), .B(n52797), .Z(n51939) );
  XNOR U53688 ( .A(round_reg[1478]), .B(round_reg[1158]), .Z(n52797) );
  XOR U53689 ( .A(round_reg[198]), .B(n52798), .Z(n52796) );
  XOR U53690 ( .A(round_reg[838]), .B(round_reg[518]), .Z(n52798) );
  XOR U53691 ( .A(n52799), .B(n52800), .Z(n46268) );
  XNOR U53692 ( .A(n44318), .B(n45081), .Z(n52800) );
  XOR U53693 ( .A(n52801), .B(n50597), .Z(n45081) );
  XOR U53694 ( .A(round_reg[1560]), .B(n48962), .Z(n50597) );
  IV U53695 ( .A(n51812), .Z(n48962) );
  XNOR U53696 ( .A(n52726), .B(n52802), .Z(n51812) );
  XOR U53697 ( .A(n52803), .B(n52804), .Z(n52726) );
  XNOR U53698 ( .A(round_reg[24]), .B(round_reg[1304]), .Z(n52804) );
  XOR U53699 ( .A(round_reg[344]), .B(n52805), .Z(n52803) );
  XOR U53700 ( .A(round_reg[984]), .B(round_reg[664]), .Z(n52805) );
  NOR U53701 ( .A(n50387), .B(n50596), .Z(n52801) );
  XNOR U53702 ( .A(n52806), .B(n51971), .Z(n44318) );
  XOR U53703 ( .A(round_reg[1434]), .B(n52807), .Z(n51971) );
  NOR U53704 ( .A(n50373), .B(n51970), .Z(n52806) );
  XNOR U53705 ( .A(n43286), .B(n52808), .Z(n52799) );
  XOR U53706 ( .A(n50591), .B(n44526), .Z(n52808) );
  XOR U53707 ( .A(n52809), .B(n50605), .Z(n44526) );
  XOR U53708 ( .A(round_reg[1404]), .B(n51567), .Z(n50605) );
  XNOR U53709 ( .A(n52811), .B(n52812), .Z(n52650) );
  XNOR U53710 ( .A(round_reg[1339]), .B(round_reg[1019]), .Z(n52812) );
  XOR U53711 ( .A(round_reg[379]), .B(n52813), .Z(n52811) );
  XOR U53712 ( .A(round_reg[699]), .B(round_reg[59]), .Z(n52813) );
  ANDN U53713 ( .B(n50604), .A(n50383), .Z(n52809) );
  XOR U53714 ( .A(n52814), .B(n50602), .Z(n50591) );
  ANDN U53715 ( .B(n50377), .A(n50601), .Z(n52814) );
  XOR U53716 ( .A(n52815), .B(n50810), .Z(n43286) );
  XOR U53717 ( .A(round_reg[1341]), .B(n52354), .Z(n50810) );
  ANDN U53718 ( .B(n50809), .A(n52816), .Z(n52815) );
  XNOR U53719 ( .A(n52817), .B(n48580), .Z(n51416) );
  XNOR U53720 ( .A(round_reg[215]), .B(n50995), .Z(n48580) );
  XOR U53721 ( .A(n52322), .B(n52818), .Z(n50995) );
  XNOR U53722 ( .A(n52819), .B(n52820), .Z(n52322) );
  XNOR U53723 ( .A(round_reg[1559]), .B(round_reg[1239]), .Z(n52820) );
  XOR U53724 ( .A(round_reg[279]), .B(n52821), .Z(n52819) );
  XOR U53725 ( .A(round_reg[919]), .B(round_reg[599]), .Z(n52821) );
  XOR U53726 ( .A(round_reg[1435]), .B(n51694), .Z(n50403) );
  XOR U53727 ( .A(round_reg[1058]), .B(n50745), .Z(n50369) );
  XNOR U53728 ( .A(n52822), .B(n52823), .Z(n52363) );
  XNOR U53729 ( .A(round_reg[33]), .B(round_reg[1313]), .Z(n52823) );
  XOR U53730 ( .A(round_reg[353]), .B(n52824), .Z(n52822) );
  XOR U53731 ( .A(round_reg[993]), .B(round_reg[673]), .Z(n52824) );
  XNOR U53732 ( .A(n52826), .B(n44091), .Z(n36363) );
  XNOR U53733 ( .A(n49420), .B(n49153), .Z(n44091) );
  XNOR U53734 ( .A(n52827), .B(n50913), .Z(n49153) );
  ANDN U53735 ( .B(n51389), .A(n51388), .Z(n52827) );
  XNOR U53736 ( .A(round_reg[341]), .B(n52153), .Z(n51389) );
  IV U53737 ( .A(n51961), .Z(n52153) );
  XOR U53738 ( .A(n52125), .B(n52578), .Z(n51961) );
  XOR U53739 ( .A(n52828), .B(n52829), .Z(n52578) );
  XNOR U53740 ( .A(round_reg[1556]), .B(round_reg[1236]), .Z(n52829) );
  XOR U53741 ( .A(round_reg[276]), .B(n52830), .Z(n52828) );
  XOR U53742 ( .A(round_reg[916]), .B(round_reg[596]), .Z(n52830) );
  XOR U53743 ( .A(n52831), .B(n52832), .Z(n52125) );
  XNOR U53744 ( .A(round_reg[1365]), .B(round_reg[1045]), .Z(n52832) );
  XOR U53745 ( .A(round_reg[405]), .B(n52833), .Z(n52831) );
  XOR U53746 ( .A(round_reg[85]), .B(round_reg[725]), .Z(n52833) );
  IV U53747 ( .A(n47396), .Z(n49420) );
  XOR U53748 ( .A(n47215), .B(n47520), .Z(n47396) );
  XOR U53749 ( .A(n52834), .B(n52835), .Z(n47520) );
  XNOR U53750 ( .A(n48797), .B(n49821), .Z(n52835) );
  XNOR U53751 ( .A(n52836), .B(n50632), .Z(n49821) );
  XNOR U53752 ( .A(round_reg[1345]), .B(n51512), .Z(n50632) );
  ANDN U53753 ( .B(n49424), .A(n49422), .Z(n52836) );
  XOR U53754 ( .A(round_reg[969]), .B(n51408), .Z(n49422) );
  XOR U53755 ( .A(round_reg[922]), .B(n49625), .Z(n49424) );
  XNOR U53756 ( .A(n51951), .B(n52837), .Z(n49625) );
  XOR U53757 ( .A(n52838), .B(n52839), .Z(n51951) );
  XNOR U53758 ( .A(round_reg[26]), .B(round_reg[1306]), .Z(n52839) );
  XOR U53759 ( .A(round_reg[346]), .B(n52840), .Z(n52838) );
  XOR U53760 ( .A(round_reg[986]), .B(round_reg[666]), .Z(n52840) );
  XNOR U53761 ( .A(n52841), .B(n50629), .Z(n48797) );
  XOR U53762 ( .A(round_reg[1565]), .B(n50520), .Z(n50629) );
  ANDN U53763 ( .B(n49159), .A(n51392), .Z(n52841) );
  IV U53764 ( .A(n49161), .Z(n51392) );
  XOR U53765 ( .A(round_reg[818]), .B(n52086), .Z(n49161) );
  XOR U53766 ( .A(round_reg[1201]), .B(n50739), .Z(n49159) );
  XNOR U53767 ( .A(n52842), .B(n52843), .Z(n52227) );
  XNOR U53768 ( .A(round_reg[1456]), .B(round_reg[1136]), .Z(n52843) );
  XOR U53769 ( .A(round_reg[176]), .B(n52844), .Z(n52842) );
  XOR U53770 ( .A(round_reg[816]), .B(round_reg[496]), .Z(n52844) );
  XOR U53771 ( .A(n52845), .B(n52846), .Z(n52456) );
  XNOR U53772 ( .A(round_reg[1585]), .B(round_reg[1265]), .Z(n52846) );
  XOR U53773 ( .A(round_reg[305]), .B(n52847), .Z(n52845) );
  XOR U53774 ( .A(round_reg[945]), .B(round_reg[625]), .Z(n52847) );
  XOR U53775 ( .A(n50903), .B(n52848), .Z(n52834) );
  XOR U53776 ( .A(n46354), .B(n43766), .Z(n52848) );
  XNOR U53777 ( .A(n52849), .B(n50620), .Z(n43766) );
  XOR U53778 ( .A(round_reg[1282]), .B(n50775), .Z(n50620) );
  XNOR U53779 ( .A(n52850), .B(n52715), .Z(n50775) );
  XOR U53780 ( .A(n52851), .B(n52852), .Z(n52715) );
  XNOR U53781 ( .A(round_reg[1346]), .B(round_reg[1026]), .Z(n52852) );
  XOR U53782 ( .A(round_reg[386]), .B(n52853), .Z(n52851) );
  XOR U53783 ( .A(round_reg[706]), .B(round_reg[66]), .Z(n52853) );
  ANDN U53784 ( .B(n49529), .A(n49528), .Z(n52849) );
  XOR U53785 ( .A(round_reg[1273]), .B(n51672), .Z(n49528) );
  XOR U53786 ( .A(round_reg[851]), .B(n52303), .Z(n49529) );
  XNOR U53787 ( .A(n52856), .B(n50624), .Z(n46354) );
  XNOR U53788 ( .A(round_reg[1439]), .B(n52025), .Z(n50624) );
  AND U53789 ( .A(n51037), .B(n50908), .Z(n52856) );
  XOR U53790 ( .A(round_reg[1062]), .B(n49280), .Z(n50908) );
  XOR U53791 ( .A(n52857), .B(n52475), .Z(n49280) );
  XNOR U53792 ( .A(n52858), .B(n52859), .Z(n52475) );
  XNOR U53793 ( .A(round_reg[357]), .B(round_reg[1317]), .Z(n52859) );
  XOR U53794 ( .A(round_reg[37]), .B(n52860), .Z(n52858) );
  XOR U53795 ( .A(round_reg[997]), .B(round_reg[677]), .Z(n52860) );
  XOR U53796 ( .A(round_reg[694]), .B(n49902), .Z(n51037) );
  XNOR U53797 ( .A(n52861), .B(n50912), .Z(n50903) );
  XNOR U53798 ( .A(round_reg[1500]), .B(n50635), .Z(n50912) );
  XOR U53799 ( .A(n52009), .B(n51952), .Z(n50635) );
  XOR U53800 ( .A(n52862), .B(n52863), .Z(n51952) );
  XNOR U53801 ( .A(round_reg[1435]), .B(round_reg[1115]), .Z(n52863) );
  XOR U53802 ( .A(round_reg[155]), .B(n52864), .Z(n52862) );
  XOR U53803 ( .A(round_reg[795]), .B(round_reg[475]), .Z(n52864) );
  XOR U53804 ( .A(n52865), .B(n52866), .Z(n52009) );
  XNOR U53805 ( .A(round_reg[1564]), .B(round_reg[1244]), .Z(n52866) );
  XOR U53806 ( .A(round_reg[284]), .B(n52867), .Z(n52865) );
  XOR U53807 ( .A(round_reg[924]), .B(round_reg[604]), .Z(n52867) );
  ANDN U53808 ( .B(n51388), .A(n50913), .Z(n52861) );
  XOR U53809 ( .A(round_reg[1111]), .B(n52113), .Z(n50913) );
  XNOR U53810 ( .A(n52868), .B(n52869), .Z(n52802) );
  XNOR U53811 ( .A(round_reg[1495]), .B(round_reg[1175]), .Z(n52869) );
  XOR U53812 ( .A(round_reg[215]), .B(n52870), .Z(n52868) );
  XOR U53813 ( .A(round_reg[855]), .B(round_reg[535]), .Z(n52870) );
  XOR U53814 ( .A(round_reg[708]), .B(n50714), .Z(n51388) );
  IV U53815 ( .A(n50741), .Z(n50714) );
  XOR U53816 ( .A(n52872), .B(n52873), .Z(n52519) );
  XNOR U53817 ( .A(round_reg[323]), .B(round_reg[1283]), .Z(n52873) );
  XOR U53818 ( .A(round_reg[3]), .B(n52874), .Z(n52872) );
  XOR U53819 ( .A(round_reg[963]), .B(round_reg[643]), .Z(n52874) );
  XOR U53820 ( .A(n52875), .B(n52876), .Z(n51938) );
  XNOR U53821 ( .A(round_reg[132]), .B(round_reg[1092]), .Z(n52876) );
  XOR U53822 ( .A(round_reg[1412]), .B(n52877), .Z(n52875) );
  XOR U53823 ( .A(round_reg[772]), .B(round_reg[452]), .Z(n52877) );
  XOR U53824 ( .A(n52878), .B(n52879), .Z(n47215) );
  XNOR U53825 ( .A(n45603), .B(n45970), .Z(n52879) );
  XNOR U53826 ( .A(n52880), .B(n48902), .Z(n45970) );
  XNOR U53827 ( .A(round_reg[693]), .B(n51195), .Z(n48902) );
  IV U53828 ( .A(n51097), .Z(n51195) );
  XOR U53829 ( .A(n52640), .B(n52378), .Z(n51097) );
  XNOR U53830 ( .A(n52881), .B(n52882), .Z(n52378) );
  XNOR U53831 ( .A(round_reg[1588]), .B(round_reg[1268]), .Z(n52882) );
  XOR U53832 ( .A(round_reg[308]), .B(n52883), .Z(n52881) );
  XOR U53833 ( .A(round_reg[948]), .B(round_reg[628]), .Z(n52883) );
  XOR U53834 ( .A(n52884), .B(n52885), .Z(n52640) );
  XNOR U53835 ( .A(round_reg[117]), .B(round_reg[1077]), .Z(n52885) );
  XOR U53836 ( .A(round_reg[1397]), .B(n52886), .Z(n52884) );
  XOR U53837 ( .A(round_reg[757]), .B(round_reg[437]), .Z(n52886) );
  ANDN U53838 ( .B(n50924), .A(n51823), .Z(n52880) );
  XOR U53839 ( .A(round_reg[218]), .B(n50814), .Z(n51823) );
  XOR U53840 ( .A(n52887), .B(n52727), .Z(n50814) );
  XNOR U53841 ( .A(n52888), .B(n52889), .Z(n52727) );
  XNOR U53842 ( .A(round_reg[1433]), .B(round_reg[1113]), .Z(n52889) );
  XOR U53843 ( .A(round_reg[153]), .B(n52890), .Z(n52888) );
  XOR U53844 ( .A(round_reg[793]), .B(round_reg[473]), .Z(n52890) );
  XNOR U53845 ( .A(round_reg[627]), .B(n50504), .Z(n50924) );
  IV U53846 ( .A(n51990), .Z(n50504) );
  XNOR U53847 ( .A(n52891), .B(n51751), .Z(n51990) );
  XNOR U53848 ( .A(n52892), .B(n52893), .Z(n51751) );
  XNOR U53849 ( .A(round_reg[1331]), .B(round_reg[1011]), .Z(n52893) );
  XOR U53850 ( .A(round_reg[371]), .B(n52894), .Z(n52892) );
  XOR U53851 ( .A(round_reg[691]), .B(round_reg[51]), .Z(n52894) );
  XNOR U53852 ( .A(n52895), .B(n48906), .Z(n45603) );
  XOR U53853 ( .A(round_reg[707]), .B(n52605), .Z(n48906) );
  NOR U53854 ( .A(n50919), .B(n51383), .Z(n52895) );
  XOR U53855 ( .A(round_reg[266]), .B(n50934), .Z(n51383) );
  XOR U53856 ( .A(round_reg[340]), .B(n50742), .Z(n50919) );
  IV U53857 ( .A(n51676), .Z(n50742) );
  XOR U53858 ( .A(n52722), .B(n52854), .Z(n51676) );
  XNOR U53859 ( .A(n52896), .B(n52897), .Z(n52854) );
  XNOR U53860 ( .A(round_reg[1555]), .B(round_reg[1235]), .Z(n52897) );
  XOR U53861 ( .A(round_reg[275]), .B(n52898), .Z(n52896) );
  XOR U53862 ( .A(round_reg[915]), .B(round_reg[595]), .Z(n52898) );
  XOR U53863 ( .A(n52899), .B(n52900), .Z(n52722) );
  XNOR U53864 ( .A(round_reg[1364]), .B(round_reg[1044]), .Z(n52900) );
  XOR U53865 ( .A(round_reg[404]), .B(n52901), .Z(n52899) );
  XOR U53866 ( .A(round_reg[84]), .B(round_reg[724]), .Z(n52901) );
  XNOR U53867 ( .A(n46271), .B(n52902), .Z(n52878) );
  XNOR U53868 ( .A(n42688), .B(n45444), .Z(n52902) );
  XNOR U53869 ( .A(n52903), .B(n48897), .Z(n45444) );
  XOR U53870 ( .A(round_reg[850]), .B(n50475), .Z(n48897) );
  IV U53871 ( .A(n52418), .Z(n50475) );
  XOR U53872 ( .A(n52904), .B(n52905), .Z(n52418) );
  ANDN U53873 ( .B(n50921), .A(n51381), .Z(n52903) );
  XNOR U53874 ( .A(round_reg[100]), .B(n52304), .Z(n51381) );
  XOR U53875 ( .A(round_reg[461]), .B(n51330), .Z(n50921) );
  XNOR U53876 ( .A(n52906), .B(n48893), .Z(n42688) );
  XOR U53877 ( .A(round_reg[921]), .B(n50434), .Z(n48893) );
  XOR U53878 ( .A(n52908), .B(n52909), .Z(n52581) );
  XNOR U53879 ( .A(round_reg[1496]), .B(round_reg[1176]), .Z(n52909) );
  XOR U53880 ( .A(round_reg[216]), .B(n52910), .Z(n52908) );
  XOR U53881 ( .A(round_reg[856]), .B(round_reg[536]), .Z(n52910) );
  ANDN U53882 ( .B(n50926), .A(n51376), .Z(n52906) );
  XNOR U53883 ( .A(n51778), .B(n52911), .Z(n52025) );
  XOR U53884 ( .A(n52912), .B(n52913), .Z(n51778) );
  XNOR U53885 ( .A(round_reg[1374]), .B(round_reg[1054]), .Z(n52913) );
  XOR U53886 ( .A(round_reg[414]), .B(n52914), .Z(n52912) );
  XOR U53887 ( .A(round_reg[94]), .B(round_reg[734]), .Z(n52914) );
  XOR U53888 ( .A(round_reg[559]), .B(n51172), .Z(n50926) );
  XOR U53889 ( .A(n52915), .B(n50329), .Z(n46271) );
  XOR U53890 ( .A(round_reg[817]), .B(n51708), .Z(n50329) );
  ANDN U53891 ( .B(n51826), .A(n50928), .Z(n52915) );
  XOR U53892 ( .A(round_reg[391]), .B(n48706), .Z(n50928) );
  XOR U53893 ( .A(n52916), .B(n52917), .Z(n48706) );
  XNOR U53894 ( .A(round_reg[14]), .B(n51491), .Z(n51826) );
  ANDN U53895 ( .B(n41408), .A(n44458), .Z(n52826) );
  IV U53896 ( .A(n41409), .Z(n44458) );
  XOR U53897 ( .A(n51865), .B(n45902), .Z(n41409) );
  XNOR U53898 ( .A(n48308), .B(n50331), .Z(n45902) );
  XNOR U53899 ( .A(n52918), .B(n52919), .Z(n50331) );
  XNOR U53900 ( .A(n45935), .B(n45399), .Z(n52919) );
  XOR U53901 ( .A(n52920), .B(n49668), .Z(n45399) );
  XOR U53902 ( .A(round_reg[648]), .B(n51377), .Z(n49668) );
  XOR U53903 ( .A(n52921), .B(n52277), .Z(n51377) );
  XNOR U53904 ( .A(n52922), .B(n52923), .Z(n52277) );
  XNOR U53905 ( .A(round_reg[1543]), .B(round_reg[1223]), .Z(n52923) );
  XOR U53906 ( .A(round_reg[263]), .B(n52924), .Z(n52922) );
  XOR U53907 ( .A(round_reg[903]), .B(round_reg[583]), .Z(n52924) );
  ANDN U53908 ( .B(n49669), .A(n49949), .Z(n52920) );
  XOR U53909 ( .A(n52925), .B(n49672), .Z(n45935) );
  XOR U53910 ( .A(round_reg[726]), .B(n51542), .Z(n49672) );
  IV U53911 ( .A(n51183), .Z(n51542) );
  XNOR U53912 ( .A(n52926), .B(n52818), .Z(n51183) );
  XNOR U53913 ( .A(n52927), .B(n52928), .Z(n52818) );
  XNOR U53914 ( .A(round_reg[1430]), .B(round_reg[1110]), .Z(n52928) );
  XOR U53915 ( .A(round_reg[150]), .B(n52929), .Z(n52927) );
  XOR U53916 ( .A(round_reg[790]), .B(round_reg[470]), .Z(n52929) );
  ANDN U53917 ( .B(n49671), .A(n49946), .Z(n52925) );
  XOR U53918 ( .A(round_reg[285]), .B(n50520), .Z(n49946) );
  XNOR U53919 ( .A(n52930), .B(n52931), .Z(n52772) );
  XNOR U53920 ( .A(round_reg[1500]), .B(round_reg[1180]), .Z(n52931) );
  XOR U53921 ( .A(round_reg[220]), .B(n52932), .Z(n52930) );
  XOR U53922 ( .A(round_reg[860]), .B(round_reg[540]), .Z(n52932) );
  XNOR U53923 ( .A(round_reg[359]), .B(n50732), .Z(n49671) );
  IV U53924 ( .A(n51927), .Z(n50732) );
  XNOR U53925 ( .A(n52229), .B(n52934), .Z(n51927) );
  XNOR U53926 ( .A(n52935), .B(n52936), .Z(n52229) );
  XNOR U53927 ( .A(round_reg[1574]), .B(round_reg[1254]), .Z(n52936) );
  XOR U53928 ( .A(round_reg[294]), .B(n52937), .Z(n52935) );
  XOR U53929 ( .A(round_reg[934]), .B(round_reg[614]), .Z(n52937) );
  XNOR U53930 ( .A(n46704), .B(n52938), .Z(n52918) );
  XNOR U53931 ( .A(n44192), .B(n42401), .Z(n52938) );
  XOR U53932 ( .A(n52939), .B(n48675), .Z(n42401) );
  XOR U53933 ( .A(round_reg[772]), .B(n52076), .Z(n48675) );
  IV U53934 ( .A(n50419), .Z(n52076) );
  ANDN U53935 ( .B(n49662), .A(n49957), .Z(n52939) );
  XOR U53936 ( .A(round_reg[33]), .B(n50715), .Z(n49957) );
  IV U53937 ( .A(n50452), .Z(n50715) );
  XOR U53938 ( .A(round_reg[410]), .B(n51468), .Z(n49662) );
  XNOR U53939 ( .A(n52940), .B(n52941), .Z(n52907) );
  XNOR U53940 ( .A(round_reg[25]), .B(round_reg[1305]), .Z(n52941) );
  XOR U53941 ( .A(round_reg[345]), .B(n52942), .Z(n52940) );
  XOR U53942 ( .A(round_reg[985]), .B(round_reg[665]), .Z(n52942) );
  XOR U53943 ( .A(n52943), .B(n52944), .Z(n52338) );
  XNOR U53944 ( .A(round_reg[1434]), .B(round_reg[1114]), .Z(n52944) );
  XOR U53945 ( .A(round_reg[154]), .B(n52945), .Z(n52943) );
  XOR U53946 ( .A(round_reg[794]), .B(round_reg[474]), .Z(n52945) );
  XNOR U53947 ( .A(n52946), .B(n48681), .Z(n44192) );
  XOR U53948 ( .A(round_reg[869]), .B(n52746), .Z(n48681) );
  XNOR U53949 ( .A(n52947), .B(n52948), .Z(n52746) );
  ANDN U53950 ( .B(n49665), .A(n51867), .Z(n52946) );
  XNOR U53951 ( .A(round_reg[119]), .B(n50483), .Z(n51867) );
  IV U53952 ( .A(n52949), .Z(n50483) );
  XOR U53953 ( .A(round_reg[480]), .B(n51397), .Z(n49665) );
  XOR U53954 ( .A(n52950), .B(n48671), .Z(n46704) );
  XOR U53955 ( .A(round_reg[940]), .B(n51098), .Z(n48671) );
  IV U53956 ( .A(n50749), .Z(n51098) );
  XOR U53957 ( .A(n52951), .B(n52952), .Z(n50749) );
  ANDN U53958 ( .B(n49660), .A(n49954), .Z(n52950) );
  XOR U53959 ( .A(round_reg[178]), .B(n51327), .Z(n49954) );
  IV U53960 ( .A(n52086), .Z(n51327) );
  XNOR U53961 ( .A(n52953), .B(n52891), .Z(n52086) );
  XNOR U53962 ( .A(n52954), .B(n52955), .Z(n52891) );
  XNOR U53963 ( .A(round_reg[1522]), .B(round_reg[1202]), .Z(n52955) );
  XOR U53964 ( .A(round_reg[242]), .B(n52956), .Z(n52954) );
  XOR U53965 ( .A(round_reg[882]), .B(round_reg[562]), .Z(n52956) );
  XNOR U53966 ( .A(round_reg[514]), .B(n51001), .Z(n49660) );
  IV U53967 ( .A(n51010), .Z(n51001) );
  XOR U53968 ( .A(n52957), .B(n52958), .Z(n48308) );
  XNOR U53969 ( .A(n47599), .B(n44970), .Z(n52958) );
  XNOR U53970 ( .A(n52959), .B(n49361), .Z(n44970) );
  XNOR U53971 ( .A(round_reg[284]), .B(n49261), .Z(n49361) );
  IV U53972 ( .A(n49798), .Z(n49261) );
  XOR U53973 ( .A(n52960), .B(n52528), .Z(n49798) );
  XNOR U53974 ( .A(n52961), .B(n52962), .Z(n52528) );
  XNOR U53975 ( .A(round_reg[28]), .B(round_reg[1308]), .Z(n52962) );
  XOR U53976 ( .A(round_reg[348]), .B(n52963), .Z(n52961) );
  XOR U53977 ( .A(round_reg[988]), .B(round_reg[668]), .Z(n52963) );
  ANDN U53978 ( .B(n49362), .A(n49974), .Z(n52959) );
  XOR U53979 ( .A(round_reg[1128]), .B(n51317), .Z(n49974) );
  IV U53980 ( .A(n51883), .Z(n51317) );
  XOR U53981 ( .A(n52964), .B(n52934), .Z(n51883) );
  XNOR U53982 ( .A(n52965), .B(n52966), .Z(n52934) );
  XNOR U53983 ( .A(round_reg[1063]), .B(round_reg[103]), .Z(n52966) );
  XOR U53984 ( .A(round_reg[1383]), .B(n52967), .Z(n52965) );
  XOR U53985 ( .A(round_reg[743]), .B(round_reg[423]), .Z(n52967) );
  XOR U53986 ( .A(round_reg[1517]), .B(n50693), .Z(n49362) );
  XNOR U53987 ( .A(n52968), .B(n49372), .Z(n47599) );
  XOR U53988 ( .A(round_reg[177]), .B(n51708), .Z(n49372) );
  ANDN U53989 ( .B(n49373), .A(n49971), .Z(n52968) );
  XOR U53990 ( .A(round_reg[986]), .B(n51663), .Z(n49971) );
  IV U53991 ( .A(n52081), .Z(n51663) );
  XOR U53992 ( .A(round_reg[1362]), .B(n51532), .Z(n49373) );
  XNOR U53993 ( .A(n49356), .B(n52971), .Z(n52957) );
  XOR U53994 ( .A(n46663), .B(n43968), .Z(n52971) );
  XNOR U53995 ( .A(n52972), .B(n52021), .Z(n43968) );
  XOR U53996 ( .A(round_reg[236]), .B(n51911), .Z(n52021) );
  ANDN U53997 ( .B(n51857), .A(n49965), .Z(n52972) );
  XOR U53998 ( .A(round_reg[1079]), .B(n52949), .Z(n49965) );
  XNOR U53999 ( .A(n52973), .B(n52974), .Z(n52949) );
  XNOR U54000 ( .A(round_reg[1456]), .B(n51818), .Z(n51857) );
  XNOR U54001 ( .A(n52512), .B(n52975), .Z(n51818) );
  XNOR U54002 ( .A(n52976), .B(n52977), .Z(n52512) );
  XNOR U54003 ( .A(round_reg[1520]), .B(round_reg[1200]), .Z(n52977) );
  XOR U54004 ( .A(round_reg[240]), .B(n52978), .Z(n52976) );
  XOR U54005 ( .A(round_reg[880]), .B(round_reg[560]), .Z(n52978) );
  XNOR U54006 ( .A(n52979), .B(n49365), .Z(n46663) );
  XNOR U54007 ( .A(round_reg[118]), .B(n48445), .Z(n49365) );
  ANDN U54008 ( .B(n49366), .A(n50637), .Z(n52979) );
  XOR U54009 ( .A(round_reg[1226]), .B(n50934), .Z(n50637) );
  XOR U54010 ( .A(round_reg[1299]), .B(n49181), .Z(n49366) );
  XNOR U54011 ( .A(n52980), .B(n49533), .Z(n49356) );
  XOR U54012 ( .A(round_reg[32]), .B(n50957), .Z(n49533) );
  IV U54013 ( .A(n50834), .Z(n50957) );
  XNOR U54014 ( .A(n52981), .B(n52982), .Z(n52589) );
  XNOR U54015 ( .A(round_reg[1376]), .B(round_reg[1056]), .Z(n52982) );
  XOR U54016 ( .A(round_reg[416]), .B(n52983), .Z(n52981) );
  XOR U54017 ( .A(round_reg[96]), .B(round_reg[736]), .Z(n52983) );
  XNOR U54018 ( .A(n52984), .B(n52985), .Z(n52202) );
  XNOR U54019 ( .A(round_reg[1567]), .B(round_reg[1247]), .Z(n52985) );
  XOR U54020 ( .A(round_reg[287]), .B(n52986), .Z(n52984) );
  XOR U54021 ( .A(round_reg[927]), .B(round_reg[607]), .Z(n52986) );
  ANDN U54022 ( .B(n49534), .A(n49962), .Z(n52980) );
  XOR U54023 ( .A(round_reg[1154]), .B(n51010), .Z(n49962) );
  XOR U54024 ( .A(n52987), .B(n52988), .Z(n51010) );
  XOR U54025 ( .A(round_reg[1582]), .B(n51582), .Z(n49534) );
  XNOR U54026 ( .A(n52989), .B(n49669), .Z(n51865) );
  XNOR U54027 ( .A(round_reg[582]), .B(n50815), .Z(n49669) );
  ANDN U54028 ( .B(n49949), .A(n49950), .Z(n52989) );
  XOR U54029 ( .A(round_reg[1457]), .B(n51708), .Z(n49950) );
  XNOR U54030 ( .A(n52990), .B(n52991), .Z(n52417) );
  XNOR U54031 ( .A(round_reg[112]), .B(round_reg[1072]), .Z(n52991) );
  XOR U54032 ( .A(round_reg[1392]), .B(n52992), .Z(n52990) );
  XOR U54033 ( .A(round_reg[752]), .B(round_reg[432]), .Z(n52992) );
  XOR U54034 ( .A(n52993), .B(n52994), .Z(n51924) );
  XNOR U54035 ( .A(round_reg[1521]), .B(round_reg[1201]), .Z(n52994) );
  XOR U54036 ( .A(round_reg[241]), .B(n52995), .Z(n52993) );
  XOR U54037 ( .A(round_reg[881]), .B(round_reg[561]), .Z(n52995) );
  XOR U54038 ( .A(round_reg[237]), .B(n50693), .Z(n49949) );
  XOR U54039 ( .A(n52996), .B(n52556), .Z(n50693) );
  XNOR U54040 ( .A(n52997), .B(n52998), .Z(n52556) );
  XNOR U54041 ( .A(round_reg[1581]), .B(round_reg[1261]), .Z(n52998) );
  XOR U54042 ( .A(round_reg[301]), .B(n52999), .Z(n52997) );
  XOR U54043 ( .A(round_reg[941]), .B(round_reg[621]), .Z(n52999) );
  XNOR U54044 ( .A(n50381), .B(n46027), .Z(n41408) );
  IV U54045 ( .A(n45922), .Z(n46027) );
  XOR U54046 ( .A(n51131), .B(n50102), .Z(n45922) );
  XOR U54047 ( .A(n53000), .B(n53001), .Z(n50102) );
  XOR U54048 ( .A(n42680), .B(n46267), .Z(n53001) );
  XNOR U54049 ( .A(n53002), .B(n51970), .Z(n46267) );
  XOR U54050 ( .A(round_reg[1057]), .B(n49089), .Z(n51970) );
  IV U54051 ( .A(n52783), .Z(n49089) );
  ANDN U54052 ( .B(n50373), .A(n50374), .Z(n53002) );
  XOR U54053 ( .A(round_reg[623]), .B(n50414), .Z(n50374) );
  XOR U54054 ( .A(n52394), .B(n52226), .Z(n50414) );
  XNOR U54055 ( .A(n53003), .B(n53004), .Z(n52226) );
  XNOR U54056 ( .A(round_reg[1327]), .B(round_reg[1007]), .Z(n53004) );
  XOR U54057 ( .A(round_reg[367]), .B(n53005), .Z(n53003) );
  XOR U54058 ( .A(round_reg[687]), .B(round_reg[47]), .Z(n53005) );
  XOR U54059 ( .A(n53006), .B(n53007), .Z(n52394) );
  XNOR U54060 ( .A(round_reg[1518]), .B(round_reg[1198]), .Z(n53007) );
  XOR U54061 ( .A(round_reg[238]), .B(n53008), .Z(n53006) );
  XOR U54062 ( .A(round_reg[878]), .B(round_reg[558]), .Z(n53008) );
  XOR U54063 ( .A(round_reg[689]), .B(n50498), .Z(n50373) );
  XOR U54064 ( .A(n53009), .B(n50601), .Z(n42680) );
  XNOR U54065 ( .A(round_reg[1106]), .B(n51100), .Z(n50601) );
  XNOR U54066 ( .A(n52785), .B(n52638), .Z(n51100) );
  XNOR U54067 ( .A(n53010), .B(n53011), .Z(n52638) );
  XNOR U54068 ( .A(round_reg[1490]), .B(round_reg[1170]), .Z(n53011) );
  XOR U54069 ( .A(round_reg[210]), .B(n53012), .Z(n53010) );
  XOR U54070 ( .A(round_reg[850]), .B(round_reg[530]), .Z(n53012) );
  XNOR U54071 ( .A(n53013), .B(n53014), .Z(n52785) );
  XNOR U54072 ( .A(round_reg[1361]), .B(round_reg[1041]), .Z(n53014) );
  XOR U54073 ( .A(round_reg[401]), .B(n53015), .Z(n53013) );
  XOR U54074 ( .A(round_reg[81]), .B(round_reg[721]), .Z(n53015) );
  NOR U54075 ( .A(n50377), .B(n50378), .Z(n53009) );
  XOR U54076 ( .A(round_reg[336]), .B(n48561), .Z(n50378) );
  XNOR U54077 ( .A(round_reg[767]), .B(n51703), .Z(n50377) );
  XOR U54078 ( .A(n52267), .B(n52420), .Z(n51703) );
  XNOR U54079 ( .A(n53016), .B(n53017), .Z(n52420) );
  XNOR U54080 ( .A(round_reg[1342]), .B(round_reg[1022]), .Z(n53017) );
  XOR U54081 ( .A(round_reg[382]), .B(n53018), .Z(n53016) );
  XOR U54082 ( .A(round_reg[702]), .B(round_reg[62]), .Z(n53018) );
  XOR U54083 ( .A(n53019), .B(n53020), .Z(n52267) );
  XNOR U54084 ( .A(round_reg[1471]), .B(round_reg[1151]), .Z(n53020) );
  XOR U54085 ( .A(round_reg[191]), .B(n53021), .Z(n53019) );
  XOR U54086 ( .A(round_reg[831]), .B(round_reg[511]), .Z(n53021) );
  XOR U54087 ( .A(n45990), .B(n53022), .Z(n53000) );
  XOR U54088 ( .A(n43724), .B(n45963), .Z(n53022) );
  XOR U54089 ( .A(n53023), .B(n50596), .Z(n45963) );
  XNOR U54090 ( .A(round_reg[1196]), .B(n51911), .Z(n50596) );
  XNOR U54091 ( .A(n52654), .B(n52307), .Z(n51911) );
  XNOR U54092 ( .A(n53024), .B(n53025), .Z(n52307) );
  XNOR U54093 ( .A(round_reg[1451]), .B(round_reg[1131]), .Z(n53025) );
  XOR U54094 ( .A(round_reg[171]), .B(n53026), .Z(n53024) );
  XOR U54095 ( .A(round_reg[811]), .B(round_reg[491]), .Z(n53026) );
  XNOR U54096 ( .A(n53027), .B(n53028), .Z(n52654) );
  XNOR U54097 ( .A(round_reg[1580]), .B(round_reg[1260]), .Z(n53028) );
  XOR U54098 ( .A(round_reg[300]), .B(n53029), .Z(n53027) );
  XOR U54099 ( .A(round_reg[940]), .B(round_reg[620]), .Z(n53029) );
  XOR U54100 ( .A(round_reg[387]), .B(n52605), .Z(n50388) );
  XOR U54101 ( .A(round_reg[813]), .B(n48558), .Z(n50387) );
  XOR U54102 ( .A(n52096), .B(n53030), .Z(n48558) );
  XOR U54103 ( .A(n53031), .B(n53032), .Z(n52096) );
  XNOR U54104 ( .A(round_reg[108]), .B(round_reg[1068]), .Z(n53032) );
  XOR U54105 ( .A(round_reg[1388]), .B(n53033), .Z(n53031) );
  XOR U54106 ( .A(round_reg[748]), .B(round_reg[428]), .Z(n53033) );
  XNOR U54107 ( .A(n53034), .B(n50809), .Z(n43724) );
  XOR U54108 ( .A(round_reg[1268]), .B(n50299), .Z(n50809) );
  XNOR U54109 ( .A(n52570), .B(n52732), .Z(n50299) );
  XNOR U54110 ( .A(n53035), .B(n53036), .Z(n52732) );
  XNOR U54111 ( .A(round_reg[1332]), .B(round_reg[1012]), .Z(n53036) );
  XOR U54112 ( .A(round_reg[372]), .B(n53037), .Z(n53035) );
  XOR U54113 ( .A(round_reg[692]), .B(round_reg[52]), .Z(n53037) );
  XNOR U54114 ( .A(n53038), .B(n53039), .Z(n52570) );
  XNOR U54115 ( .A(round_reg[1523]), .B(round_reg[1203]), .Z(n53039) );
  XOR U54116 ( .A(round_reg[243]), .B(n53040), .Z(n53038) );
  XOR U54117 ( .A(round_reg[883]), .B(round_reg[563]), .Z(n53040) );
  ANDN U54118 ( .B(n52816), .A(n51975), .Z(n53034) );
  XNOR U54119 ( .A(n53041), .B(n50604), .Z(n45990) );
  XNOR U54120 ( .A(round_reg[964]), .B(n51538), .Z(n50604) );
  IV U54121 ( .A(n51158), .Z(n51538) );
  XOR U54122 ( .A(n51964), .B(n52543), .Z(n51158) );
  XNOR U54123 ( .A(n53042), .B(n53043), .Z(n52543) );
  XNOR U54124 ( .A(round_reg[1348]), .B(round_reg[1028]), .Z(n53043) );
  XOR U54125 ( .A(round_reg[388]), .B(n53044), .Z(n53042) );
  XOR U54126 ( .A(round_reg[708]), .B(round_reg[68]), .Z(n53044) );
  XOR U54127 ( .A(n53045), .B(n53046), .Z(n51964) );
  XNOR U54128 ( .A(round_reg[1539]), .B(round_reg[1219]), .Z(n53046) );
  XOR U54129 ( .A(round_reg[259]), .B(n53047), .Z(n53045) );
  XOR U54130 ( .A(round_reg[899]), .B(round_reg[579]), .Z(n53047) );
  ANDN U54131 ( .B(n50383), .A(n50384), .Z(n53041) );
  XOR U54132 ( .A(round_reg[555]), .B(n51528), .Z(n50384) );
  XNOR U54133 ( .A(n52097), .B(n51844), .Z(n51528) );
  XNOR U54134 ( .A(n53048), .B(n53049), .Z(n51844) );
  XNOR U54135 ( .A(round_reg[1450]), .B(round_reg[1130]), .Z(n53049) );
  XOR U54136 ( .A(round_reg[170]), .B(n53050), .Z(n53048) );
  XOR U54137 ( .A(round_reg[810]), .B(round_reg[490]), .Z(n53050) );
  XNOR U54138 ( .A(n53051), .B(n53052), .Z(n52097) );
  XNOR U54139 ( .A(round_reg[1579]), .B(round_reg[1259]), .Z(n53052) );
  XOR U54140 ( .A(round_reg[299]), .B(n53053), .Z(n53051) );
  XOR U54141 ( .A(round_reg[939]), .B(round_reg[619]), .Z(n53053) );
  XOR U54142 ( .A(round_reg[917]), .B(n52501), .Z(n50383) );
  IV U54143 ( .A(n49907), .Z(n52501) );
  XOR U54144 ( .A(n52926), .B(n53054), .Z(n49907) );
  XOR U54145 ( .A(n53055), .B(n53056), .Z(n52926) );
  XNOR U54146 ( .A(round_reg[21]), .B(round_reg[1301]), .Z(n53056) );
  XOR U54147 ( .A(round_reg[341]), .B(n53057), .Z(n53055) );
  XOR U54148 ( .A(round_reg[981]), .B(round_reg[661]), .Z(n53057) );
  XOR U54149 ( .A(n53058), .B(n53059), .Z(n51131) );
  XNOR U54150 ( .A(n43871), .B(n44005), .Z(n53059) );
  XNOR U54151 ( .A(n53060), .B(n47532), .Z(n44005) );
  XOR U54152 ( .A(round_reg[456]), .B(n50497), .Z(n47532) );
  XNOR U54153 ( .A(n52491), .B(n52285), .Z(n50497) );
  XNOR U54154 ( .A(n53061), .B(n53062), .Z(n52285) );
  XNOR U54155 ( .A(round_reg[1480]), .B(round_reg[1160]), .Z(n53062) );
  XOR U54156 ( .A(round_reg[200]), .B(n53063), .Z(n53061) );
  XOR U54157 ( .A(round_reg[840]), .B(round_reg[520]), .Z(n53063) );
  XNOR U54158 ( .A(n53064), .B(n53065), .Z(n52491) );
  XNOR U54159 ( .A(round_reg[1351]), .B(round_reg[1031]), .Z(n53065) );
  XOR U54160 ( .A(round_reg[391]), .B(n53066), .Z(n53064) );
  XOR U54161 ( .A(round_reg[71]), .B(round_reg[711]), .Z(n53066) );
  ANDN U54162 ( .B(n47533), .A(n51149), .Z(n53060) );
  XNOR U54163 ( .A(round_reg[1340]), .B(n51013), .Z(n51149) );
  XNOR U54164 ( .A(round_reg[95]), .B(n51147), .Z(n47533) );
  IV U54165 ( .A(n52675), .Z(n51147) );
  XOR U54166 ( .A(n52568), .B(n53067), .Z(n52675) );
  XOR U54167 ( .A(n53068), .B(n53069), .Z(n52568) );
  XNOR U54168 ( .A(round_reg[30]), .B(round_reg[1310]), .Z(n53069) );
  XOR U54169 ( .A(round_reg[350]), .B(n53070), .Z(n53068) );
  XOR U54170 ( .A(round_reg[990]), .B(round_reg[670]), .Z(n53070) );
  XNOR U54171 ( .A(n53071), .B(n46785), .Z(n43871) );
  XOR U54172 ( .A(round_reg[622]), .B(n51582), .Z(n46785) );
  XNOR U54173 ( .A(n53072), .B(n53073), .Z(n52178) );
  XNOR U54174 ( .A(round_reg[1326]), .B(round_reg[1006]), .Z(n53073) );
  XOR U54175 ( .A(round_reg[366]), .B(n53074), .Z(n53072) );
  XOR U54176 ( .A(round_reg[686]), .B(round_reg[46]), .Z(n53074) );
  XNOR U54177 ( .A(n53075), .B(n53076), .Z(n53030) );
  XNOR U54178 ( .A(round_reg[1517]), .B(round_reg[1197]), .Z(n53076) );
  XOR U54179 ( .A(round_reg[237]), .B(n53077), .Z(n53075) );
  XOR U54180 ( .A(round_reg[877]), .B(round_reg[557]), .Z(n53077) );
  ANDN U54181 ( .B(n46786), .A(n48325), .Z(n53071) );
  XNOR U54182 ( .A(round_reg[1433]), .B(n49854), .Z(n48325) );
  IV U54183 ( .A(n50148), .Z(n49854) );
  XOR U54184 ( .A(n52321), .B(n52837), .Z(n50148) );
  XNOR U54185 ( .A(n53078), .B(n53079), .Z(n52837) );
  XNOR U54186 ( .A(round_reg[1497]), .B(round_reg[1177]), .Z(n53079) );
  XOR U54187 ( .A(round_reg[217]), .B(n53080), .Z(n53078) );
  XOR U54188 ( .A(round_reg[857]), .B(round_reg[537]), .Z(n53080) );
  XOR U54189 ( .A(n53081), .B(n53082), .Z(n52321) );
  XNOR U54190 ( .A(round_reg[1368]), .B(round_reg[1048]), .Z(n53082) );
  XOR U54191 ( .A(round_reg[408]), .B(n53083), .Z(n53081) );
  XOR U54192 ( .A(round_reg[88]), .B(round_reg[728]), .Z(n53083) );
  XNOR U54193 ( .A(round_reg[213]), .B(n50430), .Z(n46786) );
  IV U54194 ( .A(n49268), .Z(n50430) );
  XOR U54195 ( .A(n53084), .B(n53085), .Z(n49268) );
  XOR U54196 ( .A(n43549), .B(n53086), .Z(n53058) );
  XOR U54197 ( .A(n46401), .B(n46771), .Z(n53086) );
  XNOR U54198 ( .A(n53087), .B(n48910), .Z(n46771) );
  XOR U54199 ( .A(round_reg[554]), .B(n48564), .Z(n48910) );
  XOR U54200 ( .A(n52138), .B(n53088), .Z(n48564) );
  XOR U54201 ( .A(n53089), .B(n53090), .Z(n52138) );
  XNOR U54202 ( .A(round_reg[1449]), .B(round_reg[1129]), .Z(n53090) );
  XOR U54203 ( .A(round_reg[169]), .B(n53091), .Z(n53089) );
  XOR U54204 ( .A(round_reg[809]), .B(round_reg[489]), .Z(n53091) );
  ANDN U54205 ( .B(n48332), .A(n48333), .Z(n53087) );
  XNOR U54206 ( .A(round_reg[1403]), .B(n50984), .Z(n48333) );
  XNOR U54207 ( .A(round_reg[154]), .B(n52807), .Z(n48332) );
  XNOR U54208 ( .A(n53094), .B(n49601), .Z(n46401) );
  XOR U54209 ( .A(round_reg[335]), .B(n48362), .Z(n49601) );
  ANDN U54210 ( .B(n48336), .A(n48337), .Z(n53094) );
  XOR U54211 ( .A(round_reg[1494]), .B(n51200), .Z(n48337) );
  XOR U54212 ( .A(n52598), .B(n53095), .Z(n51200) );
  XOR U54213 ( .A(n53096), .B(n53097), .Z(n52598) );
  XNOR U54214 ( .A(round_reg[1558]), .B(round_reg[1238]), .Z(n53097) );
  XOR U54215 ( .A(round_reg[278]), .B(n53098), .Z(n53096) );
  XOR U54216 ( .A(round_reg[918]), .B(round_reg[598]), .Z(n53098) );
  XOR U54217 ( .A(round_reg[261]), .B(n50441), .Z(n48336) );
  XNOR U54218 ( .A(n53099), .B(n52407), .Z(n50441) );
  XNOR U54219 ( .A(n53100), .B(n53101), .Z(n52407) );
  XNOR U54220 ( .A(round_reg[325]), .B(round_reg[1285]), .Z(n53101) );
  XOR U54221 ( .A(round_reg[5]), .B(n53102), .Z(n53100) );
  XOR U54222 ( .A(round_reg[965]), .B(round_reg[645]), .Z(n53102) );
  XNOR U54223 ( .A(n53103), .B(n46778), .Z(n43549) );
  XNOR U54224 ( .A(round_reg[386]), .B(n49989), .Z(n46778) );
  IV U54225 ( .A(n51630), .Z(n49989) );
  XOR U54226 ( .A(n51963), .B(n53104), .Z(n51630) );
  XOR U54227 ( .A(n53105), .B(n53106), .Z(n51963) );
  XNOR U54228 ( .A(round_reg[130]), .B(round_reg[1090]), .Z(n53106) );
  XOR U54229 ( .A(round_reg[1410]), .B(n53107), .Z(n53105) );
  XOR U54230 ( .A(round_reg[770]), .B(round_reg[450]), .Z(n53107) );
  ANDN U54231 ( .B(n46779), .A(n48329), .Z(n53103) );
  XOR U54232 ( .A(round_reg[1559]), .B(n50738), .Z(n48329) );
  XNOR U54233 ( .A(round_reg[9]), .B(n51408), .Z(n46779) );
  XOR U54234 ( .A(n53108), .B(n52816), .Z(n50381) );
  XOR U54235 ( .A(round_reg[846]), .B(n53109), .Z(n52816) );
  ANDN U54236 ( .B(n51975), .A(n50808), .Z(n53108) );
  XNOR U54237 ( .A(round_reg[96]), .B(n51928), .Z(n50808) );
  XNOR U54238 ( .A(round_reg[457]), .B(n50124), .Z(n51975) );
  IV U54239 ( .A(n51364), .Z(n50124) );
  XOR U54240 ( .A(n52921), .B(n53110), .Z(n51364) );
  XOR U54241 ( .A(n53111), .B(n53112), .Z(n52921) );
  XNOR U54242 ( .A(round_reg[1352]), .B(round_reg[1032]), .Z(n53112) );
  XOR U54243 ( .A(round_reg[392]), .B(n53113), .Z(n53111) );
  XOR U54244 ( .A(round_reg[72]), .B(round_reg[712]), .Z(n53113) );
  XNOR U54245 ( .A(n53114), .B(n44086), .Z(n42783) );
  XNOR U54246 ( .A(n52158), .B(n46877), .Z(n44086) );
  XNOR U54247 ( .A(n53115), .B(n53116), .Z(n50197) );
  XNOR U54248 ( .A(n43464), .B(n44017), .Z(n53116) );
  XNOR U54249 ( .A(n53117), .B(n48078), .Z(n44017) );
  XOR U54250 ( .A(round_reg[108]), .B(n49801), .Z(n48078) );
  ANDN U54251 ( .B(n48079), .A(n51896), .Z(n53117) );
  XOR U54252 ( .A(round_reg[1216]), .B(n51199), .Z(n51896) );
  XOR U54253 ( .A(round_reg[1289]), .B(n51557), .Z(n48079) );
  IV U54254 ( .A(n51408), .Z(n51557) );
  XNOR U54255 ( .A(n53118), .B(n52779), .Z(n51408) );
  XNOR U54256 ( .A(n53119), .B(n53120), .Z(n52779) );
  XNOR U54257 ( .A(round_reg[1353]), .B(round_reg[1033]), .Z(n53120) );
  XOR U54258 ( .A(round_reg[393]), .B(n53121), .Z(n53119) );
  XOR U54259 ( .A(round_reg[73]), .B(round_reg[713]), .Z(n53121) );
  XNOR U54260 ( .A(n53122), .B(n48711), .Z(n43464) );
  XNOR U54261 ( .A(round_reg[226]), .B(n48708), .Z(n48711) );
  IV U54262 ( .A(n51352), .Z(n48708) );
  XNOR U54263 ( .A(n52411), .B(n53123), .Z(n51352) );
  XOR U54264 ( .A(n53124), .B(n53125), .Z(n52411) );
  XNOR U54265 ( .A(round_reg[1570]), .B(round_reg[1250]), .Z(n53125) );
  XOR U54266 ( .A(round_reg[290]), .B(n53126), .Z(n53124) );
  XOR U54267 ( .A(round_reg[930]), .B(round_reg[610]), .Z(n53126) );
  ANDN U54268 ( .B(n48712), .A(n52162), .Z(n53122) );
  XOR U54269 ( .A(round_reg[1069]), .B(n50432), .Z(n52162) );
  XOR U54270 ( .A(n51958), .B(n52951), .Z(n50432) );
  XNOR U54271 ( .A(n53127), .B(n53128), .Z(n52951) );
  XNOR U54272 ( .A(round_reg[1324]), .B(round_reg[1004]), .Z(n53128) );
  XOR U54273 ( .A(round_reg[364]), .B(n53129), .Z(n53127) );
  XOR U54274 ( .A(round_reg[684]), .B(round_reg[44]), .Z(n53129) );
  XOR U54275 ( .A(n53130), .B(n53131), .Z(n51958) );
  XNOR U54276 ( .A(round_reg[1453]), .B(round_reg[1133]), .Z(n53131) );
  XOR U54277 ( .A(round_reg[173]), .B(n53132), .Z(n53130) );
  XOR U54278 ( .A(round_reg[813]), .B(round_reg[493]), .Z(n53132) );
  XOR U54279 ( .A(round_reg[1446]), .B(n51547), .Z(n48712) );
  XNOR U54280 ( .A(n53134), .B(n53135), .Z(n52294) );
  XNOR U54281 ( .A(round_reg[1061]), .B(round_reg[101]), .Z(n53135) );
  XOR U54282 ( .A(round_reg[1381]), .B(n53136), .Z(n53134) );
  XOR U54283 ( .A(round_reg[741]), .B(round_reg[421]), .Z(n53136) );
  XOR U54284 ( .A(n46728), .B(n53137), .Z(n53115) );
  XOR U54285 ( .A(n44668), .B(n48040), .Z(n53137) );
  XNOR U54286 ( .A(n53138), .B(n48068), .Z(n48040) );
  XOR U54287 ( .A(round_reg[274]), .B(n50755), .Z(n48068) );
  XNOR U54288 ( .A(n53139), .B(n52624), .Z(n50755) );
  XOR U54289 ( .A(n53140), .B(n53141), .Z(n52624) );
  XNOR U54290 ( .A(round_reg[1489]), .B(round_reg[1169]), .Z(n53141) );
  XOR U54291 ( .A(round_reg[209]), .B(n53142), .Z(n53140) );
  XOR U54292 ( .A(round_reg[849]), .B(round_reg[529]), .Z(n53142) );
  ANDN U54293 ( .B(n48069), .A(n51889), .Z(n53138) );
  XNOR U54294 ( .A(n53143), .B(n48064), .Z(n44668) );
  XNOR U54295 ( .A(round_reg[22]), .B(n48945), .Z(n48064) );
  ANDN U54296 ( .B(n48065), .A(n51893), .Z(n53143) );
  XNOR U54297 ( .A(round_reg[1208]), .B(n50427), .Z(n51893) );
  IV U54298 ( .A(n52015), .Z(n50427) );
  XNOR U54299 ( .A(n52973), .B(n52441), .Z(n52015) );
  XOR U54300 ( .A(n53144), .B(n53145), .Z(n52441) );
  XNOR U54301 ( .A(round_reg[1592]), .B(round_reg[1272]), .Z(n53145) );
  XOR U54302 ( .A(round_reg[312]), .B(n53146), .Z(n53144) );
  XOR U54303 ( .A(round_reg[952]), .B(round_reg[632]), .Z(n53146) );
  XOR U54304 ( .A(n53147), .B(n53148), .Z(n52973) );
  XNOR U54305 ( .A(round_reg[1463]), .B(round_reg[1143]), .Z(n53148) );
  XOR U54306 ( .A(round_reg[183]), .B(n53149), .Z(n53147) );
  XOR U54307 ( .A(round_reg[823]), .B(round_reg[503]), .Z(n53149) );
  XNOR U54308 ( .A(round_reg[1572]), .B(n51250), .Z(n48065) );
  XOR U54309 ( .A(n52466), .B(n51764), .Z(n51250) );
  XOR U54310 ( .A(n53150), .B(n53151), .Z(n51764) );
  XNOR U54311 ( .A(round_reg[356]), .B(round_reg[1316]), .Z(n53151) );
  XOR U54312 ( .A(round_reg[36]), .B(n53152), .Z(n53150) );
  XOR U54313 ( .A(round_reg[996]), .B(round_reg[676]), .Z(n53152) );
  XOR U54314 ( .A(n53153), .B(n53154), .Z(n52466) );
  XNOR U54315 ( .A(round_reg[1507]), .B(round_reg[1187]), .Z(n53154) );
  XOR U54316 ( .A(round_reg[227]), .B(n53155), .Z(n53153) );
  XOR U54317 ( .A(round_reg[867]), .B(round_reg[547]), .Z(n53155) );
  XNOR U54318 ( .A(n53156), .B(n48074), .Z(n46728) );
  XNOR U54319 ( .A(round_reg[167]), .B(n52034), .Z(n48074) );
  IV U54320 ( .A(n51723), .Z(n52034) );
  XOR U54321 ( .A(n53157), .B(n52212), .Z(n51723) );
  XNOR U54322 ( .A(n53158), .B(n53159), .Z(n52212) );
  XNOR U54323 ( .A(round_reg[1511]), .B(round_reg[1191]), .Z(n53159) );
  XOR U54324 ( .A(round_reg[231]), .B(n53160), .Z(n53158) );
  XOR U54325 ( .A(round_reg[871]), .B(round_reg[551]), .Z(n53160) );
  ANDN U54326 ( .B(n48075), .A(n51899), .Z(n53156) );
  XOR U54327 ( .A(round_reg[976]), .B(n48561), .Z(n51899) );
  XNOR U54328 ( .A(n52625), .B(n52752), .Z(n48561) );
  XNOR U54329 ( .A(n53161), .B(n53162), .Z(n52752) );
  XNOR U54330 ( .A(round_reg[1551]), .B(round_reg[1231]), .Z(n53162) );
  XOR U54331 ( .A(round_reg[271]), .B(n53163), .Z(n53161) );
  XOR U54332 ( .A(round_reg[911]), .B(round_reg[591]), .Z(n53163) );
  XNOR U54333 ( .A(n53164), .B(n53165), .Z(n52625) );
  XNOR U54334 ( .A(round_reg[1360]), .B(round_reg[1040]), .Z(n53165) );
  XOR U54335 ( .A(round_reg[400]), .B(n53166), .Z(n53164) );
  XOR U54336 ( .A(round_reg[80]), .B(round_reg[720]), .Z(n53166) );
  XOR U54337 ( .A(round_reg[1352]), .B(n51393), .Z(n48075) );
  XOR U54338 ( .A(n52795), .B(n53167), .Z(n51393) );
  XOR U54339 ( .A(n53168), .B(n53169), .Z(n52795) );
  XNOR U54340 ( .A(round_reg[327]), .B(round_reg[1287]), .Z(n53169) );
  XOR U54341 ( .A(round_reg[647]), .B(n53170), .Z(n53168) );
  XOR U54342 ( .A(round_reg[967]), .B(round_reg[7]), .Z(n53170) );
  XOR U54343 ( .A(n53171), .B(n53172), .Z(n49326) );
  XNOR U54344 ( .A(n45666), .B(n47452), .Z(n53172) );
  XOR U54345 ( .A(n53173), .B(n48056), .Z(n47452) );
  XOR U54346 ( .A(round_reg[1068]), .B(n50139), .Z(n48056) );
  IV U54347 ( .A(n49801), .Z(n50139) );
  XOR U54348 ( .A(n52996), .B(n52530), .Z(n49801) );
  XNOR U54349 ( .A(n53174), .B(n53175), .Z(n52530) );
  XNOR U54350 ( .A(round_reg[1323]), .B(round_reg[1003]), .Z(n53175) );
  XOR U54351 ( .A(round_reg[363]), .B(n53176), .Z(n53174) );
  XOR U54352 ( .A(round_reg[683]), .B(round_reg[43]), .Z(n53176) );
  XOR U54353 ( .A(n53177), .B(n53178), .Z(n52996) );
  XNOR U54354 ( .A(round_reg[1452]), .B(round_reg[1132]), .Z(n53178) );
  XOR U54355 ( .A(round_reg[172]), .B(n53179), .Z(n53177) );
  XOR U54356 ( .A(round_reg[812]), .B(round_reg[492]), .Z(n53179) );
  NOR U54357 ( .A(n50584), .B(n48055), .Z(n53173) );
  XNOR U54358 ( .A(round_reg[700]), .B(n51094), .Z(n48055) );
  XOR U54359 ( .A(round_reg[634]), .B(n52384), .Z(n50584) );
  IV U54360 ( .A(n50857), .Z(n52384) );
  XOR U54361 ( .A(n53180), .B(n48059), .Z(n45666) );
  XOR U54362 ( .A(round_reg[1117]), .B(n48517), .Z(n48059) );
  XOR U54363 ( .A(n52356), .B(n52569), .Z(n48517) );
  XOR U54364 ( .A(n53181), .B(n53182), .Z(n52569) );
  XNOR U54365 ( .A(round_reg[1501]), .B(round_reg[1181]), .Z(n53182) );
  XOR U54366 ( .A(round_reg[221]), .B(n53183), .Z(n53181) );
  XOR U54367 ( .A(round_reg[861]), .B(round_reg[541]), .Z(n53183) );
  XOR U54368 ( .A(n53184), .B(n53185), .Z(n52356) );
  XNOR U54369 ( .A(round_reg[1372]), .B(round_reg[1052]), .Z(n53185) );
  XOR U54370 ( .A(round_reg[412]), .B(n53186), .Z(n53184) );
  XOR U54371 ( .A(round_reg[92]), .B(round_reg[732]), .Z(n53186) );
  NOR U54372 ( .A(n47207), .B(n48058), .Z(n53180) );
  XNOR U54373 ( .A(round_reg[714]), .B(n52004), .Z(n48058) );
  XOR U54374 ( .A(n52459), .B(n52286), .Z(n52004) );
  XNOR U54375 ( .A(n53187), .B(n53188), .Z(n52286) );
  XNOR U54376 ( .A(round_reg[329]), .B(round_reg[1289]), .Z(n53188) );
  XOR U54377 ( .A(round_reg[649]), .B(n53189), .Z(n53187) );
  XOR U54378 ( .A(round_reg[9]), .B(round_reg[969]), .Z(n53189) );
  XOR U54379 ( .A(n53190), .B(n53191), .Z(n52459) );
  XNOR U54380 ( .A(round_reg[138]), .B(round_reg[1098]), .Z(n53191) );
  XOR U54381 ( .A(round_reg[1418]), .B(n53192), .Z(n53190) );
  XOR U54382 ( .A(round_reg[778]), .B(round_reg[458]), .Z(n53192) );
  XOR U54383 ( .A(round_reg[347]), .B(n49955), .Z(n47207) );
  XOR U54384 ( .A(n47109), .B(n53193), .Z(n53171) );
  XOR U54385 ( .A(n47146), .B(n45134), .Z(n53193) );
  XOR U54386 ( .A(n53194), .B(n48048), .Z(n45134) );
  XOR U54387 ( .A(round_reg[1207]), .B(n51626), .Z(n48048) );
  NOR U54388 ( .A(n47203), .B(n48047), .Z(n53194) );
  XOR U54389 ( .A(round_reg[824]), .B(n51907), .Z(n48047) );
  XOR U54390 ( .A(n53195), .B(n52697), .Z(n51907) );
  XOR U54391 ( .A(n53196), .B(n53197), .Z(n52697) );
  XNOR U54392 ( .A(round_reg[119]), .B(round_reg[1079]), .Z(n53197) );
  XOR U54393 ( .A(round_reg[1399]), .B(n53198), .Z(n53196) );
  XOR U54394 ( .A(round_reg[759]), .B(round_reg[439]), .Z(n53198) );
  XNOR U54395 ( .A(round_reg[398]), .B(n48957), .Z(n47203) );
  XNOR U54396 ( .A(n52753), .B(n52602), .Z(n48957) );
  XNOR U54397 ( .A(n53199), .B(n53200), .Z(n52602) );
  XNOR U54398 ( .A(round_reg[13]), .B(round_reg[1293]), .Z(n53200) );
  XOR U54399 ( .A(round_reg[333]), .B(n53201), .Z(n53199) );
  XOR U54400 ( .A(round_reg[973]), .B(round_reg[653]), .Z(n53201) );
  XOR U54401 ( .A(n53202), .B(n53203), .Z(n52753) );
  XNOR U54402 ( .A(round_reg[1422]), .B(round_reg[1102]), .Z(n53203) );
  XOR U54403 ( .A(round_reg[142]), .B(n53204), .Z(n53202) );
  XOR U54404 ( .A(round_reg[782]), .B(round_reg[462]), .Z(n53204) );
  XNOR U54405 ( .A(n53205), .B(n48051), .Z(n47146) );
  XOR U54406 ( .A(round_reg[1279]), .B(n52313), .Z(n48051) );
  XOR U54407 ( .A(n53206), .B(n53207), .Z(n52676) );
  XNOR U54408 ( .A(round_reg[1534]), .B(round_reg[1214]), .Z(n53207) );
  XOR U54409 ( .A(round_reg[254]), .B(n53208), .Z(n53206) );
  XOR U54410 ( .A(round_reg[894]), .B(round_reg[574]), .Z(n53208) );
  XOR U54411 ( .A(n53209), .B(n53210), .Z(n51830) );
  XNOR U54412 ( .A(round_reg[1343]), .B(round_reg[1023]), .Z(n53210) );
  XOR U54413 ( .A(round_reg[383]), .B(n53211), .Z(n53209) );
  XOR U54414 ( .A(round_reg[703]), .B(round_reg[63]), .Z(n53211) );
  ANDN U54415 ( .B(n48052), .A(n47198), .Z(n53205) );
  XOR U54416 ( .A(round_reg[468]), .B(n51789), .Z(n47198) );
  XOR U54417 ( .A(n53213), .B(n53214), .Z(n53054) );
  XNOR U54418 ( .A(round_reg[1492]), .B(round_reg[1172]), .Z(n53214) );
  XOR U54419 ( .A(round_reg[212]), .B(n53215), .Z(n53213) );
  XOR U54420 ( .A(round_reg[852]), .B(round_reg[532]), .Z(n53215) );
  XOR U54421 ( .A(round_reg[857]), .B(n51790), .Z(n48052) );
  IV U54422 ( .A(n50508), .Z(n51790) );
  XNOR U54423 ( .A(n52969), .B(n51944), .Z(n50508) );
  XNOR U54424 ( .A(n53216), .B(n53217), .Z(n51944) );
  XNOR U54425 ( .A(round_reg[1432]), .B(round_reg[1112]), .Z(n53217) );
  XOR U54426 ( .A(round_reg[152]), .B(n53218), .Z(n53216) );
  XOR U54427 ( .A(round_reg[792]), .B(round_reg[472]), .Z(n53218) );
  XOR U54428 ( .A(n53219), .B(n53220), .Z(n52969) );
  XNOR U54429 ( .A(round_reg[1561]), .B(round_reg[1241]), .Z(n53220) );
  XOR U54430 ( .A(round_reg[281]), .B(n53221), .Z(n53219) );
  XOR U54431 ( .A(round_reg[921]), .B(round_reg[601]), .Z(n53221) );
  XNOR U54432 ( .A(n53222), .B(n48044), .Z(n47109) );
  XOR U54433 ( .A(round_reg[975]), .B(n48362), .Z(n48044) );
  XNOR U54434 ( .A(n53223), .B(n52586), .Z(n48362) );
  XOR U54435 ( .A(n53224), .B(n53225), .Z(n52586) );
  XNOR U54436 ( .A(round_reg[1359]), .B(round_reg[1039]), .Z(n53225) );
  XOR U54437 ( .A(round_reg[399]), .B(n53226), .Z(n53224) );
  XOR U54438 ( .A(round_reg[79]), .B(round_reg[719]), .Z(n53226) );
  ANDN U54439 ( .B(n48045), .A(n47211), .Z(n53222) );
  XOR U54440 ( .A(round_reg[566]), .B(n50234), .Z(n47211) );
  XNOR U54441 ( .A(n52696), .B(n52731), .Z(n50234) );
  XOR U54442 ( .A(n53227), .B(n53228), .Z(n52731) );
  XNOR U54443 ( .A(round_reg[1461]), .B(round_reg[1141]), .Z(n53228) );
  XOR U54444 ( .A(round_reg[181]), .B(n53229), .Z(n53227) );
  XOR U54445 ( .A(round_reg[821]), .B(round_reg[501]), .Z(n53229) );
  XOR U54446 ( .A(n53230), .B(n53231), .Z(n52696) );
  XNOR U54447 ( .A(round_reg[1590]), .B(round_reg[1270]), .Z(n53231) );
  XOR U54448 ( .A(round_reg[310]), .B(n53232), .Z(n53230) );
  XOR U54449 ( .A(round_reg[950]), .B(round_reg[630]), .Z(n53232) );
  XOR U54450 ( .A(round_reg[928]), .B(n49860), .Z(n48045) );
  XNOR U54451 ( .A(n52911), .B(n53233), .Z(n49860) );
  XNOR U54452 ( .A(n53234), .B(n53235), .Z(n52911) );
  XNOR U54453 ( .A(round_reg[1503]), .B(round_reg[1183]), .Z(n53235) );
  XOR U54454 ( .A(round_reg[223]), .B(n53236), .Z(n53234) );
  XOR U54455 ( .A(round_reg[863]), .B(round_reg[543]), .Z(n53236) );
  XOR U54456 ( .A(n53237), .B(n48069), .Z(n52158) );
  XOR U54457 ( .A(round_reg[1507]), .B(n48450), .Z(n48069) );
  XNOR U54458 ( .A(n53238), .B(n52825), .Z(n48450) );
  XOR U54459 ( .A(n53239), .B(n53240), .Z(n52825) );
  XNOR U54460 ( .A(round_reg[1442]), .B(round_reg[1122]), .Z(n53240) );
  XOR U54461 ( .A(round_reg[162]), .B(n53241), .Z(n53239) );
  XOR U54462 ( .A(round_reg[802]), .B(round_reg[482]), .Z(n53241) );
  ANDN U54463 ( .B(n51889), .A(n51890), .Z(n53237) );
  XNOR U54464 ( .A(round_reg[715]), .B(n51205), .Z(n51890) );
  XNOR U54465 ( .A(round_reg[1118]), .B(n50650), .Z(n51889) );
  XNOR U54466 ( .A(n53244), .B(n53245), .Z(n52612) );
  XNOR U54467 ( .A(round_reg[1502]), .B(round_reg[1182]), .Z(n53245) );
  XOR U54468 ( .A(round_reg[222]), .B(n53246), .Z(n53244) );
  XOR U54469 ( .A(round_reg[862]), .B(round_reg[542]), .Z(n53246) );
  XOR U54470 ( .A(n53247), .B(n53248), .Z(n52010) );
  XNOR U54471 ( .A(round_reg[1373]), .B(round_reg[1053]), .Z(n53248) );
  XOR U54472 ( .A(round_reg[413]), .B(n53249), .Z(n53247) );
  XOR U54473 ( .A(round_reg[93]), .B(round_reg[733]), .Z(n53249) );
  XOR U54474 ( .A(n53250), .B(n44248), .Z(n41411) );
  XOR U54475 ( .A(n51766), .B(n43958), .Z(n44248) );
  XOR U54476 ( .A(n47574), .B(n47252), .Z(n43958) );
  XNOR U54477 ( .A(n53251), .B(n53252), .Z(n47252) );
  XOR U54478 ( .A(n45829), .B(n46651), .Z(n53252) );
  XNOR U54479 ( .A(n53253), .B(n49678), .Z(n46651) );
  XNOR U54480 ( .A(round_reg[658]), .B(n51053), .Z(n49678) );
  IV U54481 ( .A(n51428), .Z(n51053) );
  XOR U54482 ( .A(n52754), .B(n52386), .Z(n51428) );
  XNOR U54483 ( .A(n53254), .B(n53255), .Z(n52386) );
  XNOR U54484 ( .A(round_reg[1553]), .B(round_reg[1233]), .Z(n53255) );
  XOR U54485 ( .A(round_reg[273]), .B(n53256), .Z(n53254) );
  XOR U54486 ( .A(round_reg[913]), .B(round_reg[593]), .Z(n53256) );
  XOR U54487 ( .A(n53257), .B(n53258), .Z(n52754) );
  XNOR U54488 ( .A(round_reg[1362]), .B(round_reg[1042]), .Z(n53258) );
  XOR U54489 ( .A(round_reg[402]), .B(n53259), .Z(n53257) );
  XOR U54490 ( .A(round_reg[82]), .B(round_reg[722]), .Z(n53259) );
  ANDN U54491 ( .B(n48824), .A(n51631), .Z(n53253) );
  XOR U54492 ( .A(round_reg[592]), .B(n50955), .Z(n51631) );
  IV U54493 ( .A(n51103), .Z(n50955) );
  XOR U54494 ( .A(n53260), .B(n53261), .Z(n51103) );
  XNOR U54495 ( .A(round_reg[247]), .B(n52087), .Z(n48824) );
  IV U54496 ( .A(n51626), .Z(n52087) );
  XOR U54497 ( .A(n52296), .B(n53262), .Z(n51626) );
  XOR U54498 ( .A(n53263), .B(n53264), .Z(n52296) );
  XNOR U54499 ( .A(round_reg[1591]), .B(round_reg[1271]), .Z(n53264) );
  XOR U54500 ( .A(round_reg[311]), .B(n53265), .Z(n53263) );
  XOR U54501 ( .A(round_reg[951]), .B(round_reg[631]), .Z(n53265) );
  XNOR U54502 ( .A(n53266), .B(n49681), .Z(n45829) );
  XOR U54503 ( .A(round_reg[736]), .B(n51928), .Z(n49681) );
  XNOR U54504 ( .A(n52611), .B(n52463), .Z(n51928) );
  XNOR U54505 ( .A(n53267), .B(n53268), .Z(n52463) );
  XNOR U54506 ( .A(round_reg[1440]), .B(round_reg[1120]), .Z(n53268) );
  XOR U54507 ( .A(round_reg[160]), .B(n53269), .Z(n53267) );
  XOR U54508 ( .A(round_reg[800]), .B(round_reg[480]), .Z(n53269) );
  XOR U54509 ( .A(n53270), .B(n53271), .Z(n52611) );
  XNOR U54510 ( .A(round_reg[31]), .B(round_reg[1311]), .Z(n53271) );
  XOR U54511 ( .A(round_reg[351]), .B(n53272), .Z(n53270) );
  XOR U54512 ( .A(round_reg[991]), .B(round_reg[671]), .Z(n53272) );
  ANDN U54513 ( .B(n50696), .A(n51633), .Z(n53266) );
  XNOR U54514 ( .A(round_reg[369]), .B(n50498), .Z(n51633) );
  XNOR U54515 ( .A(n52953), .B(n53273), .Z(n50498) );
  XOR U54516 ( .A(n53274), .B(n53275), .Z(n52953) );
  XNOR U54517 ( .A(round_reg[113]), .B(round_reg[1073]), .Z(n53275) );
  XOR U54518 ( .A(round_reg[1393]), .B(n53276), .Z(n53274) );
  XOR U54519 ( .A(round_reg[753]), .B(round_reg[433]), .Z(n53276) );
  XNOR U54520 ( .A(round_reg[295]), .B(n52170), .Z(n50696) );
  XOR U54521 ( .A(n46518), .B(n53277), .Z(n53251) );
  XNOR U54522 ( .A(n51613), .B(n44682), .Z(n53277) );
  XOR U54523 ( .A(n53278), .B(n49689), .Z(n44682) );
  XOR U54524 ( .A(round_reg[950]), .B(n50106), .Z(n49689) );
  XNOR U54525 ( .A(n52974), .B(n52133), .Z(n50106) );
  XOR U54526 ( .A(n53279), .B(n53280), .Z(n52133) );
  XNOR U54527 ( .A(round_reg[1525]), .B(round_reg[1205]), .Z(n53280) );
  XOR U54528 ( .A(round_reg[245]), .B(n53281), .Z(n53279) );
  XOR U54529 ( .A(round_reg[885]), .B(round_reg[565]), .Z(n53281) );
  XOR U54530 ( .A(n53282), .B(n53283), .Z(n52974) );
  XNOR U54531 ( .A(round_reg[1334]), .B(round_reg[1014]), .Z(n53283) );
  XOR U54532 ( .A(round_reg[374]), .B(n53284), .Z(n53282) );
  XOR U54533 ( .A(round_reg[694]), .B(round_reg[54]), .Z(n53284) );
  ANDN U54534 ( .B(n48832), .A(n51641), .Z(n53278) );
  XOR U54535 ( .A(round_reg[524]), .B(n51140), .Z(n51641) );
  XOR U54536 ( .A(n52224), .B(n53243), .Z(n51140) );
  XOR U54537 ( .A(n53285), .B(n53286), .Z(n53243) );
  XNOR U54538 ( .A(round_reg[139]), .B(round_reg[1099]), .Z(n53286) );
  XOR U54539 ( .A(round_reg[1419]), .B(n53287), .Z(n53285) );
  XOR U54540 ( .A(round_reg[779]), .B(round_reg[459]), .Z(n53287) );
  XOR U54541 ( .A(n53288), .B(n53289), .Z(n52224) );
  XNOR U54542 ( .A(round_reg[1548]), .B(round_reg[1228]), .Z(n53289) );
  XOR U54543 ( .A(round_reg[268]), .B(n53290), .Z(n53288) );
  XOR U54544 ( .A(round_reg[908]), .B(round_reg[588]), .Z(n53290) );
  XNOR U54545 ( .A(round_reg[188]), .B(n51030), .Z(n48832) );
  IV U54546 ( .A(n52072), .Z(n51030) );
  XNOR U54547 ( .A(n53291), .B(n49691), .Z(n51613) );
  XNOR U54548 ( .A(round_reg[782]), .B(n50853), .Z(n49691) );
  ANDN U54549 ( .B(n48828), .A(n51636), .Z(n53291) );
  XOR U54550 ( .A(round_reg[420]), .B(n52304), .Z(n51636) );
  XOR U54551 ( .A(n52948), .B(n51917), .Z(n52304) );
  XOR U54552 ( .A(n53292), .B(n53293), .Z(n51917) );
  XNOR U54553 ( .A(round_reg[355]), .B(round_reg[1315]), .Z(n53293) );
  XOR U54554 ( .A(round_reg[35]), .B(n53294), .Z(n53292) );
  XOR U54555 ( .A(round_reg[995]), .B(round_reg[675]), .Z(n53294) );
  XOR U54556 ( .A(n53295), .B(n53296), .Z(n52948) );
  XNOR U54557 ( .A(round_reg[1444]), .B(round_reg[1124]), .Z(n53296) );
  XOR U54558 ( .A(round_reg[164]), .B(n53297), .Z(n53295) );
  XOR U54559 ( .A(round_reg[804]), .B(round_reg[484]), .Z(n53297) );
  XNOR U54560 ( .A(round_reg[43]), .B(n50823), .Z(n48828) );
  XNOR U54561 ( .A(n53298), .B(n53088), .Z(n50823) );
  XNOR U54562 ( .A(n53299), .B(n53300), .Z(n53088) );
  XNOR U54563 ( .A(round_reg[1578]), .B(round_reg[1258]), .Z(n53300) );
  XOR U54564 ( .A(round_reg[298]), .B(n53301), .Z(n53299) );
  XOR U54565 ( .A(round_reg[938]), .B(round_reg[618]), .Z(n53301) );
  XOR U54566 ( .A(n53302), .B(n49686), .Z(n46518) );
  XNOR U54567 ( .A(round_reg[879]), .B(n51172), .Z(n49686) );
  XOR U54568 ( .A(n53303), .B(n52416), .Z(n51172) );
  XNOR U54569 ( .A(n53304), .B(n53305), .Z(n52416) );
  XNOR U54570 ( .A(round_reg[1583]), .B(round_reg[1263]), .Z(n53305) );
  XOR U54571 ( .A(round_reg[303]), .B(n53306), .Z(n53304) );
  XOR U54572 ( .A(round_reg[943]), .B(round_reg[623]), .Z(n53306) );
  XOR U54573 ( .A(round_reg[490]), .B(n50761), .Z(n51638) );
  XOR U54574 ( .A(n52382), .B(n52529), .Z(n50761) );
  XNOR U54575 ( .A(n53307), .B(n53308), .Z(n52529) );
  XNOR U54576 ( .A(round_reg[1514]), .B(round_reg[1194]), .Z(n53308) );
  XOR U54577 ( .A(round_reg[234]), .B(n53309), .Z(n53307) );
  XOR U54578 ( .A(round_reg[874]), .B(round_reg[554]), .Z(n53309) );
  XOR U54579 ( .A(n53310), .B(n53311), .Z(n52382) );
  XNOR U54580 ( .A(round_reg[1065]), .B(round_reg[105]), .Z(n53311) );
  XOR U54581 ( .A(round_reg[1385]), .B(n53312), .Z(n53310) );
  XOR U54582 ( .A(round_reg[745]), .B(round_reg[425]), .Z(n53312) );
  XNOR U54583 ( .A(round_reg[65]), .B(n50156), .Z(n48819) );
  IV U54584 ( .A(n51512), .Z(n50156) );
  XOR U54585 ( .A(n52987), .B(n53313), .Z(n51512) );
  XOR U54586 ( .A(n53314), .B(n53315), .Z(n52987) );
  XNOR U54587 ( .A(round_reg[129]), .B(round_reg[1089]), .Z(n53315) );
  XOR U54588 ( .A(round_reg[1409]), .B(n53316), .Z(n53314) );
  XOR U54589 ( .A(round_reg[769]), .B(round_reg[449]), .Z(n53316) );
  XOR U54590 ( .A(n53317), .B(n53318), .Z(n47574) );
  XNOR U54591 ( .A(n43345), .B(n47993), .Z(n53318) );
  XNOR U54592 ( .A(n53319), .B(n48395), .Z(n47993) );
  XNOR U54593 ( .A(round_reg[1468]), .B(n52072), .Z(n48395) );
  AND U54594 ( .A(n51758), .B(n48396), .Z(n53319) );
  XOR U54595 ( .A(round_reg[1027]), .B(n52605), .Z(n48396) );
  XNOR U54596 ( .A(n52470), .B(n52122), .Z(n52605) );
  XOR U54597 ( .A(n53320), .B(n53321), .Z(n52122) );
  XNOR U54598 ( .A(round_reg[2]), .B(round_reg[1282]), .Z(n53321) );
  XOR U54599 ( .A(round_reg[322]), .B(n53322), .Z(n53320) );
  XOR U54600 ( .A(round_reg[962]), .B(round_reg[642]), .Z(n53322) );
  XOR U54601 ( .A(n53323), .B(n53324), .Z(n52470) );
  XNOR U54602 ( .A(round_reg[131]), .B(round_reg[1091]), .Z(n53324) );
  XOR U54603 ( .A(round_reg[1411]), .B(n53325), .Z(n53323) );
  XOR U54604 ( .A(round_reg[771]), .B(round_reg[451]), .Z(n53325) );
  XNOR U54605 ( .A(round_reg[659]), .B(n49181), .Z(n51758) );
  XOR U54606 ( .A(n52904), .B(n53212), .Z(n49181) );
  XNOR U54607 ( .A(n53326), .B(n53327), .Z(n53212) );
  XNOR U54608 ( .A(round_reg[1363]), .B(round_reg[1043]), .Z(n53327) );
  XOR U54609 ( .A(round_reg[403]), .B(n53328), .Z(n53326) );
  XOR U54610 ( .A(round_reg[83]), .B(round_reg[723]), .Z(n53328) );
  XOR U54611 ( .A(n53329), .B(n53330), .Z(n52904) );
  XNOR U54612 ( .A(round_reg[1554]), .B(round_reg[1234]), .Z(n53330) );
  XOR U54613 ( .A(round_reg[274]), .B(n53331), .Z(n53329) );
  XOR U54614 ( .A(round_reg[914]), .B(round_reg[594]), .Z(n53331) );
  XNOR U54615 ( .A(n53332), .B(n48983), .Z(n43345) );
  XOR U54616 ( .A(round_reg[1529]), .B(n49836), .Z(n48983) );
  XNOR U54617 ( .A(n52236), .B(n52516), .Z(n49836) );
  XOR U54618 ( .A(n53333), .B(n53334), .Z(n52516) );
  XNOR U54619 ( .A(round_reg[1593]), .B(round_reg[1273]), .Z(n53334) );
  XOR U54620 ( .A(round_reg[313]), .B(n53335), .Z(n53333) );
  XOR U54621 ( .A(round_reg[953]), .B(round_reg[633]), .Z(n53335) );
  XOR U54622 ( .A(n53336), .B(n53337), .Z(n52236) );
  XNOR U54623 ( .A(round_reg[1464]), .B(round_reg[1144]), .Z(n53337) );
  XOR U54624 ( .A(round_reg[184]), .B(n53338), .Z(n53336) );
  XOR U54625 ( .A(round_reg[824]), .B(round_reg[504]), .Z(n53338) );
  ANDN U54626 ( .B(n48984), .A(n51769), .Z(n53332) );
  XOR U54627 ( .A(round_reg[737]), .B(n52783), .Z(n51769) );
  XOR U54628 ( .A(n53123), .B(n53233), .Z(n52783) );
  XNOR U54629 ( .A(n53339), .B(n53340), .Z(n53233) );
  XNOR U54630 ( .A(round_reg[32]), .B(round_reg[1312]), .Z(n53340) );
  XOR U54631 ( .A(round_reg[352]), .B(n53341), .Z(n53339) );
  XOR U54632 ( .A(round_reg[992]), .B(round_reg[672]), .Z(n53341) );
  XOR U54633 ( .A(n53342), .B(n53343), .Z(n53123) );
  XNOR U54634 ( .A(round_reg[1441]), .B(round_reg[1121]), .Z(n53343) );
  XOR U54635 ( .A(round_reg[161]), .B(n53344), .Z(n53342) );
  XOR U54636 ( .A(round_reg[801]), .B(round_reg[481]), .Z(n53344) );
  XNOR U54637 ( .A(round_reg[1140]), .B(n51185), .Z(n48984) );
  XOR U54638 ( .A(n51658), .B(n52662), .Z(n51185) );
  XOR U54639 ( .A(n53345), .B(n53346), .Z(n52662) );
  XNOR U54640 ( .A(round_reg[115]), .B(round_reg[1075]), .Z(n53346) );
  XOR U54641 ( .A(round_reg[1395]), .B(n53347), .Z(n53345) );
  XOR U54642 ( .A(round_reg[755]), .B(round_reg[435]), .Z(n53347) );
  XOR U54643 ( .A(n53348), .B(n53349), .Z(n51658) );
  XNOR U54644 ( .A(round_reg[1524]), .B(round_reg[1204]), .Z(n53349) );
  XOR U54645 ( .A(round_reg[244]), .B(n53350), .Z(n53348) );
  XOR U54646 ( .A(round_reg[884]), .B(round_reg[564]), .Z(n53350) );
  XNOR U54647 ( .A(n47684), .B(n53351), .Z(n53317) );
  XNOR U54648 ( .A(n45141), .B(n47401), .Z(n53351) );
  XNOR U54649 ( .A(n53352), .B(n48398), .Z(n47401) );
  IV U54650 ( .A(n49991), .Z(n48398) );
  XOR U54651 ( .A(round_reg[1374]), .B(n49606), .Z(n49991) );
  XNOR U54652 ( .A(n52201), .B(n52933), .Z(n49606) );
  XOR U54653 ( .A(n53353), .B(n53354), .Z(n52933) );
  XNOR U54654 ( .A(round_reg[29]), .B(round_reg[1309]), .Z(n53354) );
  XOR U54655 ( .A(round_reg[349]), .B(n53355), .Z(n53353) );
  XOR U54656 ( .A(round_reg[989]), .B(round_reg[669]), .Z(n53355) );
  XOR U54657 ( .A(n53356), .B(n53357), .Z(n52201) );
  XNOR U54658 ( .A(round_reg[1438]), .B(round_reg[1118]), .Z(n53357) );
  XOR U54659 ( .A(round_reg[158]), .B(n53358), .Z(n53356) );
  XOR U54660 ( .A(round_reg[798]), .B(round_reg[478]), .Z(n53358) );
  ANDN U54661 ( .B(n48399), .A(n47049), .Z(n53352) );
  XOR U54662 ( .A(round_reg[951]), .B(n51810), .Z(n47049) );
  XOR U54663 ( .A(n52237), .B(n52641), .Z(n51810) );
  XOR U54664 ( .A(n53359), .B(n53360), .Z(n52641) );
  XNOR U54665 ( .A(round_reg[1526]), .B(round_reg[1206]), .Z(n53360) );
  XOR U54666 ( .A(round_reg[246]), .B(n53361), .Z(n53359) );
  XOR U54667 ( .A(round_reg[886]), .B(round_reg[566]), .Z(n53361) );
  XNOR U54668 ( .A(n53362), .B(n53363), .Z(n52237) );
  XNOR U54669 ( .A(round_reg[1335]), .B(round_reg[1015]), .Z(n53363) );
  XOR U54670 ( .A(round_reg[375]), .B(n53364), .Z(n53362) );
  XOR U54671 ( .A(round_reg[695]), .B(round_reg[55]), .Z(n53364) );
  XNOR U54672 ( .A(round_reg[998]), .B(n50412), .Z(n48399) );
  IV U54673 ( .A(n51589), .Z(n50412) );
  XNOR U54674 ( .A(n52947), .B(n53157), .Z(n51589) );
  XOR U54675 ( .A(n53365), .B(n53366), .Z(n53157) );
  XNOR U54676 ( .A(round_reg[1062]), .B(round_reg[102]), .Z(n53366) );
  XOR U54677 ( .A(round_reg[1382]), .B(n53367), .Z(n53365) );
  XOR U54678 ( .A(round_reg[742]), .B(round_reg[422]), .Z(n53367) );
  XOR U54679 ( .A(n53368), .B(n53369), .Z(n52947) );
  XNOR U54680 ( .A(round_reg[1573]), .B(round_reg[1253]), .Z(n53369) );
  XOR U54681 ( .A(round_reg[293]), .B(n53370), .Z(n53368) );
  XOR U54682 ( .A(round_reg[933]), .B(round_reg[613]), .Z(n53370) );
  XNOR U54683 ( .A(n53371), .B(n49693), .Z(n45141) );
  XNOR U54684 ( .A(round_reg[1311]), .B(n52041), .Z(n49693) );
  IV U54685 ( .A(n50519), .Z(n52041) );
  XOR U54686 ( .A(n53372), .B(n53373), .Z(n50519) );
  ANDN U54687 ( .B(n49694), .A(n47043), .Z(n53371) );
  XOR U54688 ( .A(n53374), .B(n48391), .Z(n47684) );
  XNOR U54689 ( .A(round_reg[1594]), .B(n50857), .Z(n48391) );
  XOR U54690 ( .A(n52365), .B(n53093), .Z(n50857) );
  XOR U54691 ( .A(n53375), .B(n53376), .Z(n53093) );
  XNOR U54692 ( .A(round_reg[1338]), .B(round_reg[1018]), .Z(n53376) );
  XOR U54693 ( .A(round_reg[378]), .B(n53377), .Z(n53375) );
  XOR U54694 ( .A(round_reg[698]), .B(round_reg[58]), .Z(n53377) );
  XOR U54695 ( .A(n53378), .B(n53379), .Z(n52365) );
  XNOR U54696 ( .A(round_reg[1529]), .B(round_reg[1209]), .Z(n53379) );
  XOR U54697 ( .A(round_reg[249]), .B(n53380), .Z(n53378) );
  XOR U54698 ( .A(round_reg[889]), .B(round_reg[569]), .Z(n53380) );
  AND U54699 ( .A(n47053), .B(n48392), .Z(n53374) );
  XNOR U54700 ( .A(round_reg[1166]), .B(n50772), .Z(n48392) );
  IV U54701 ( .A(n53109), .Z(n50772) );
  XNOR U54702 ( .A(n53381), .B(n53223), .Z(n53109) );
  XOR U54703 ( .A(n53382), .B(n53383), .Z(n53223) );
  XNOR U54704 ( .A(round_reg[1550]), .B(round_reg[1230]), .Z(n53383) );
  XOR U54705 ( .A(round_reg[270]), .B(n53384), .Z(n53382) );
  XOR U54706 ( .A(round_reg[910]), .B(round_reg[590]), .Z(n53384) );
  XNOR U54707 ( .A(round_reg[783]), .B(n52523), .Z(n47053) );
  XNOR U54708 ( .A(n53386), .B(n53387), .Z(n53261) );
  XNOR U54709 ( .A(round_reg[1487]), .B(round_reg[1167]), .Z(n53387) );
  XOR U54710 ( .A(round_reg[207]), .B(n53388), .Z(n53386) );
  XOR U54711 ( .A(round_reg[847]), .B(round_reg[527]), .Z(n53388) );
  XNOR U54712 ( .A(n53389), .B(n49694), .Z(n51766) );
  XOR U54713 ( .A(round_reg[1238]), .B(n50397), .Z(n49694) );
  XOR U54714 ( .A(n51604), .B(n52721), .Z(n50397) );
  XNOR U54715 ( .A(n53390), .B(n53391), .Z(n52721) );
  XNOR U54716 ( .A(round_reg[1493]), .B(round_reg[1173]), .Z(n53391) );
  XOR U54717 ( .A(round_reg[213]), .B(n53392), .Z(n53390) );
  XOR U54718 ( .A(round_reg[853]), .B(round_reg[533]), .Z(n53392) );
  XOR U54719 ( .A(n53393), .B(n53394), .Z(n51604) );
  XNOR U54720 ( .A(round_reg[22]), .B(round_reg[1302]), .Z(n53394) );
  XOR U54721 ( .A(round_reg[342]), .B(n53395), .Z(n53393) );
  XOR U54722 ( .A(round_reg[982]), .B(round_reg[662]), .Z(n53395) );
  ANDN U54723 ( .B(n47043), .A(n47044), .Z(n53389) );
  XOR U54724 ( .A(round_reg[491]), .B(n51135), .Z(n47044) );
  XOR U54725 ( .A(n53273), .B(n52177), .Z(n48938) );
  XOR U54726 ( .A(n53396), .B(n53397), .Z(n52177) );
  XNOR U54727 ( .A(round_reg[1455]), .B(round_reg[1135]), .Z(n53397) );
  XOR U54728 ( .A(round_reg[175]), .B(n53398), .Z(n53396) );
  XOR U54729 ( .A(round_reg[815]), .B(round_reg[495]), .Z(n53398) );
  XOR U54730 ( .A(n53399), .B(n53400), .Z(n53273) );
  XNOR U54731 ( .A(round_reg[1584]), .B(round_reg[1264]), .Z(n53400) );
  XOR U54732 ( .A(round_reg[304]), .B(n53401), .Z(n53399) );
  XOR U54733 ( .A(round_reg[944]), .B(round_reg[624]), .Z(n53401) );
  NOR U54734 ( .A(n44475), .B(n44085), .Z(n53250) );
  XOR U54735 ( .A(n52050), .B(n45814), .Z(n44085) );
  XOR U54736 ( .A(n47839), .B(n49581), .Z(n45814) );
  XNOR U54737 ( .A(n53402), .B(n53403), .Z(n49581) );
  XNOR U54738 ( .A(n47474), .B(n46996), .Z(n53403) );
  XOR U54739 ( .A(n53404), .B(n51275), .Z(n46996) );
  IV U54740 ( .A(n52269), .Z(n51275) );
  XOR U54741 ( .A(round_reg[82]), .B(n51532), .Z(n52269) );
  XNOR U54742 ( .A(n52747), .B(n52855), .Z(n51532) );
  XOR U54743 ( .A(n53405), .B(n53406), .Z(n52855) );
  XNOR U54744 ( .A(round_reg[1426]), .B(round_reg[1106]), .Z(n53406) );
  XOR U54745 ( .A(round_reg[146]), .B(n53407), .Z(n53405) );
  XOR U54746 ( .A(round_reg[786]), .B(round_reg[466]), .Z(n53407) );
  XOR U54747 ( .A(n53408), .B(n53409), .Z(n52747) );
  XNOR U54748 ( .A(round_reg[17]), .B(round_reg[1297]), .Z(n53409) );
  XOR U54749 ( .A(round_reg[337]), .B(n53410), .Z(n53408) );
  XOR U54750 ( .A(round_reg[977]), .B(round_reg[657]), .Z(n53410) );
  NOR U54751 ( .A(n51744), .B(n51274), .Z(n53404) );
  XNOR U54752 ( .A(round_reg[1327]), .B(n51146), .Z(n51274) );
  XOR U54753 ( .A(n52975), .B(n51959), .Z(n51146) );
  XNOR U54754 ( .A(n53411), .B(n53412), .Z(n51959) );
  XNOR U54755 ( .A(round_reg[1582]), .B(round_reg[1262]), .Z(n53412) );
  XOR U54756 ( .A(round_reg[302]), .B(n53413), .Z(n53411) );
  XOR U54757 ( .A(round_reg[942]), .B(round_reg[622]), .Z(n53413) );
  XOR U54758 ( .A(n53414), .B(n53415), .Z(n52975) );
  XNOR U54759 ( .A(round_reg[111]), .B(round_reg[1071]), .Z(n53415) );
  XOR U54760 ( .A(round_reg[1391]), .B(n53416), .Z(n53414) );
  XOR U54761 ( .A(round_reg[751]), .B(round_reg[431]), .Z(n53416) );
  XOR U54762 ( .A(round_reg[1254]), .B(n51341), .Z(n51744) );
  XNOR U54763 ( .A(n52623), .B(n51681), .Z(n51341) );
  XOR U54764 ( .A(n53417), .B(n53418), .Z(n51681) );
  XNOR U54765 ( .A(round_reg[1509]), .B(round_reg[1189]), .Z(n53418) );
  XOR U54766 ( .A(round_reg[229]), .B(n53419), .Z(n53417) );
  XOR U54767 ( .A(round_reg[869]), .B(round_reg[549]), .Z(n53419) );
  XOR U54768 ( .A(n53420), .B(n53421), .Z(n52623) );
  XNOR U54769 ( .A(round_reg[358]), .B(round_reg[1318]), .Z(n53421) );
  XOR U54770 ( .A(round_reg[38]), .B(n53422), .Z(n53420) );
  XOR U54771 ( .A(round_reg[998]), .B(round_reg[678]), .Z(n53422) );
  XOR U54772 ( .A(n53423), .B(n52258), .Z(n47474) );
  XOR U54773 ( .A(round_reg[60]), .B(n51013), .Z(n52258) );
  IV U54774 ( .A(n51094), .Z(n51013) );
  XNOR U54775 ( .A(n53424), .B(n53425), .Z(n52222) );
  XNOR U54776 ( .A(round_reg[1595]), .B(round_reg[1275]), .Z(n53425) );
  XOR U54777 ( .A(round_reg[315]), .B(n53426), .Z(n53424) );
  XOR U54778 ( .A(round_reg[955]), .B(round_reg[635]), .Z(n53426) );
  XOR U54779 ( .A(n53427), .B(n53428), .Z(n52669) );
  XNOR U54780 ( .A(round_reg[124]), .B(round_reg[1084]), .Z(n53428) );
  XOR U54781 ( .A(round_reg[1404]), .B(n53429), .Z(n53427) );
  XOR U54782 ( .A(round_reg[764]), .B(round_reg[444]), .Z(n53429) );
  ANDN U54783 ( .B(n46843), .A(n52257), .Z(n53423) );
  IV U54784 ( .A(n52058), .Z(n52257) );
  XOR U54785 ( .A(round_reg[1546]), .B(n50934), .Z(n52058) );
  IV U54786 ( .A(n51599), .Z(n50934) );
  XOR U54787 ( .A(n53242), .B(n53110), .Z(n51599) );
  XNOR U54788 ( .A(n53430), .B(n53431), .Z(n53110) );
  XNOR U54789 ( .A(round_reg[1481]), .B(round_reg[1161]), .Z(n53431) );
  XOR U54790 ( .A(round_reg[201]), .B(n53432), .Z(n53430) );
  XOR U54791 ( .A(round_reg[841]), .B(round_reg[521]), .Z(n53432) );
  XNOR U54792 ( .A(n53433), .B(n53434), .Z(n53242) );
  XNOR U54793 ( .A(round_reg[1290]), .B(round_reg[10]), .Z(n53434) );
  XOR U54794 ( .A(round_reg[330]), .B(n53435), .Z(n53433) );
  XOR U54795 ( .A(round_reg[970]), .B(round_reg[650]), .Z(n53435) );
  XNOR U54796 ( .A(round_reg[1182]), .B(n51050), .Z(n46843) );
  XOR U54797 ( .A(n47168), .B(n53436), .Z(n53402) );
  XOR U54798 ( .A(n47405), .B(n45079), .Z(n53436) );
  XNOR U54799 ( .A(n53437), .B(n51278), .Z(n45079) );
  XOR U54800 ( .A(round_reg[200]), .B(n50947), .Z(n51278) );
  XOR U54801 ( .A(n53118), .B(n52916), .Z(n50947) );
  XNOR U54802 ( .A(n53438), .B(n53439), .Z(n52916) );
  XNOR U54803 ( .A(round_reg[135]), .B(round_reg[1095]), .Z(n53439) );
  XOR U54804 ( .A(round_reg[1415]), .B(n53440), .Z(n53438) );
  XOR U54805 ( .A(round_reg[775]), .B(round_reg[455]), .Z(n53440) );
  XOR U54806 ( .A(n53441), .B(n53442), .Z(n53118) );
  XNOR U54807 ( .A(round_reg[1544]), .B(round_reg[1224]), .Z(n53442) );
  XOR U54808 ( .A(round_reg[264]), .B(n53443), .Z(n53441) );
  XOR U54809 ( .A(round_reg[904]), .B(round_reg[584]), .Z(n53443) );
  ANDN U54810 ( .B(n47952), .A(n51277), .Z(n53437) );
  XOR U54811 ( .A(round_reg[1420]), .B(n51727), .Z(n51277) );
  IV U54812 ( .A(n51579), .Z(n51727) );
  XNOR U54813 ( .A(n53444), .B(n53445), .Z(n52603) );
  XNOR U54814 ( .A(round_reg[1484]), .B(round_reg[1164]), .Z(n53445) );
  XOR U54815 ( .A(round_reg[204]), .B(n53446), .Z(n53444) );
  XOR U54816 ( .A(round_reg[844]), .B(round_reg[524]), .Z(n53446) );
  XNOR U54817 ( .A(n53447), .B(n53448), .Z(n52766) );
  XNOR U54818 ( .A(round_reg[1355]), .B(round_reg[1035]), .Z(n53448) );
  XOR U54819 ( .A(round_reg[395]), .B(n53449), .Z(n53447) );
  XOR U54820 ( .A(round_reg[75]), .B(round_reg[715]), .Z(n53449) );
  XOR U54821 ( .A(round_reg[1043]), .B(n52166), .Z(n47952) );
  XNOR U54822 ( .A(n53450), .B(n51286), .Z(n47405) );
  XOR U54823 ( .A(round_reg[141]), .B(n51330), .Z(n51286) );
  XNOR U54824 ( .A(n52240), .B(n52535), .Z(n51330) );
  XOR U54825 ( .A(n53451), .B(n53452), .Z(n52535) );
  XNOR U54826 ( .A(round_reg[1356]), .B(round_reg[1036]), .Z(n53452) );
  XOR U54827 ( .A(round_reg[396]), .B(n53453), .Z(n53451) );
  XOR U54828 ( .A(round_reg[76]), .B(round_reg[716]), .Z(n53453) );
  XOR U54829 ( .A(n53454), .B(n53455), .Z(n52240) );
  XNOR U54830 ( .A(round_reg[1485]), .B(round_reg[1165]), .Z(n53455) );
  XOR U54831 ( .A(round_reg[205]), .B(n53456), .Z(n53454) );
  XOR U54832 ( .A(round_reg[845]), .B(round_reg[525]), .Z(n53456) );
  ANDN U54833 ( .B(n51287), .A(n51304), .Z(n53450) );
  XNOR U54834 ( .A(round_reg[1014]), .B(n49902), .Z(n51304) );
  XOR U54835 ( .A(n52316), .B(n52403), .Z(n49902) );
  XNOR U54836 ( .A(n53457), .B(n53458), .Z(n52403) );
  XNOR U54837 ( .A(round_reg[118]), .B(round_reg[1078]), .Z(n53458) );
  XOR U54838 ( .A(round_reg[1398]), .B(n53459), .Z(n53457) );
  XOR U54839 ( .A(round_reg[758]), .B(round_reg[438]), .Z(n53459) );
  XNOR U54840 ( .A(n53460), .B(n53461), .Z(n52316) );
  XNOR U54841 ( .A(round_reg[1589]), .B(round_reg[1269]), .Z(n53461) );
  XOR U54842 ( .A(round_reg[309]), .B(n53462), .Z(n53460) );
  XOR U54843 ( .A(round_reg[949]), .B(round_reg[629]), .Z(n53462) );
  XOR U54844 ( .A(round_reg[1390]), .B(n51997), .Z(n51287) );
  IV U54845 ( .A(n50831), .Z(n51997) );
  XNOR U54846 ( .A(n53303), .B(n52728), .Z(n50831) );
  XNOR U54847 ( .A(n53463), .B(n53464), .Z(n52728) );
  XNOR U54848 ( .A(round_reg[1325]), .B(round_reg[1005]), .Z(n53464) );
  XOR U54849 ( .A(round_reg[365]), .B(n53465), .Z(n53463) );
  XOR U54850 ( .A(round_reg[685]), .B(round_reg[45]), .Z(n53465) );
  XOR U54851 ( .A(n53466), .B(n53467), .Z(n53303) );
  XNOR U54852 ( .A(round_reg[1454]), .B(round_reg[1134]), .Z(n53467) );
  XOR U54853 ( .A(round_reg[174]), .B(n53468), .Z(n53466) );
  XOR U54854 ( .A(round_reg[814]), .B(round_reg[494]), .Z(n53468) );
  XOR U54855 ( .A(n53469), .B(n51283), .Z(n47168) );
  XOR U54856 ( .A(round_reg[312]), .B(n50733), .Z(n51283) );
  IV U54857 ( .A(n51224), .Z(n50733) );
  XNOR U54858 ( .A(n52703), .B(n52402), .Z(n51224) );
  XOR U54859 ( .A(n53470), .B(n53471), .Z(n52402) );
  XNOR U54860 ( .A(round_reg[1527]), .B(round_reg[1207]), .Z(n53471) );
  XOR U54861 ( .A(round_reg[247]), .B(n53472), .Z(n53470) );
  XOR U54862 ( .A(round_reg[887]), .B(round_reg[567]), .Z(n53472) );
  XOR U54863 ( .A(n53473), .B(n53474), .Z(n52703) );
  XNOR U54864 ( .A(round_reg[1336]), .B(round_reg[1016]), .Z(n53474) );
  XOR U54865 ( .A(round_reg[376]), .B(n53475), .Z(n53473) );
  XOR U54866 ( .A(round_reg[696]), .B(round_reg[56]), .Z(n53475) );
  XNOR U54867 ( .A(round_reg[1481]), .B(n51660), .Z(n51282) );
  XOR U54868 ( .A(round_reg[1092]), .B(n50419), .Z(n46836) );
  XNOR U54869 ( .A(n53476), .B(n53099), .Z(n50419) );
  XNOR U54870 ( .A(n53477), .B(n53478), .Z(n53099) );
  XNOR U54871 ( .A(round_reg[1476]), .B(round_reg[1156]), .Z(n53478) );
  XOR U54872 ( .A(round_reg[196]), .B(n53479), .Z(n53477) );
  XOR U54873 ( .A(round_reg[836]), .B(round_reg[516]), .Z(n53479) );
  XOR U54874 ( .A(n53480), .B(n53481), .Z(n47839) );
  XOR U54875 ( .A(n46523), .B(n42505), .Z(n53481) );
  XNOR U54876 ( .A(n53482), .B(n50863), .Z(n42505) );
  IV U54877 ( .A(n51300), .Z(n50863) );
  XOR U54878 ( .A(round_reg[904]), .B(n50111), .Z(n51300) );
  IV U54879 ( .A(n51788), .Z(n50111) );
  XOR U54880 ( .A(n52341), .B(n52447), .Z(n51788) );
  XNOR U54881 ( .A(n53483), .B(n53484), .Z(n52447) );
  XNOR U54882 ( .A(round_reg[1479]), .B(round_reg[1159]), .Z(n53484) );
  XOR U54883 ( .A(round_reg[199]), .B(n53485), .Z(n53483) );
  XOR U54884 ( .A(round_reg[839]), .B(round_reg[519]), .Z(n53485) );
  XOR U54885 ( .A(n53486), .B(n53487), .Z(n52341) );
  XNOR U54886 ( .A(round_reg[328]), .B(round_reg[1288]), .Z(n53487) );
  XOR U54887 ( .A(round_reg[648]), .B(n53488), .Z(n53486) );
  XOR U54888 ( .A(round_reg[968]), .B(round_reg[8]), .Z(n53488) );
  ANDN U54889 ( .B(n49047), .A(n51299), .Z(n53482) );
  XNOR U54890 ( .A(round_reg[542]), .B(n51050), .Z(n51299) );
  XNOR U54891 ( .A(n53372), .B(n52527), .Z(n51050) );
  XOR U54892 ( .A(n53489), .B(n53490), .Z(n52527) );
  XNOR U54893 ( .A(round_reg[1437]), .B(round_reg[1117]), .Z(n53490) );
  XOR U54894 ( .A(round_reg[157]), .B(n53491), .Z(n53489) );
  XOR U54895 ( .A(round_reg[797]), .B(round_reg[477]), .Z(n53491) );
  XOR U54896 ( .A(n53492), .B(n53493), .Z(n53372) );
  XNOR U54897 ( .A(round_reg[1566]), .B(round_reg[1246]), .Z(n53493) );
  XOR U54898 ( .A(round_reg[286]), .B(n53494), .Z(n53492) );
  XOR U54899 ( .A(round_reg[926]), .B(round_reg[606]), .Z(n53494) );
  XNOR U54900 ( .A(round_reg[142]), .B(n51395), .Z(n49047) );
  IV U54901 ( .A(n50853), .Z(n51395) );
  XOR U54902 ( .A(n52717), .B(n52225), .Z(n50853) );
  XOR U54903 ( .A(n53495), .B(n53496), .Z(n52225) );
  XNOR U54904 ( .A(round_reg[1357]), .B(round_reg[1037]), .Z(n53496) );
  XOR U54905 ( .A(round_reg[397]), .B(n53497), .Z(n53495) );
  XOR U54906 ( .A(round_reg[77]), .B(round_reg[717]), .Z(n53497) );
  XOR U54907 ( .A(n53498), .B(n53499), .Z(n52717) );
  XNOR U54908 ( .A(round_reg[1486]), .B(round_reg[1166]), .Z(n53499) );
  XOR U54909 ( .A(round_reg[206]), .B(n53500), .Z(n53498) );
  XOR U54910 ( .A(round_reg[846]), .B(round_reg[526]), .Z(n53500) );
  XNOR U54911 ( .A(n53501), .B(n50872), .Z(n46523) );
  XOR U54912 ( .A(round_reg[676]), .B(n50888), .Z(n50872) );
  IV U54913 ( .A(n51335), .Z(n50888) );
  XOR U54914 ( .A(n53238), .B(n51680), .Z(n51335) );
  XNOR U54915 ( .A(n53502), .B(n53503), .Z(n51680) );
  XNOR U54916 ( .A(round_reg[1060]), .B(round_reg[100]), .Z(n53503) );
  XOR U54917 ( .A(round_reg[1380]), .B(n53504), .Z(n53502) );
  XOR U54918 ( .A(round_reg[740]), .B(round_reg[420]), .Z(n53504) );
  XOR U54919 ( .A(n53505), .B(n53506), .Z(n53238) );
  XNOR U54920 ( .A(round_reg[1571]), .B(round_reg[1251]), .Z(n53506) );
  XOR U54921 ( .A(round_reg[291]), .B(n53507), .Z(n53505) );
  XOR U54922 ( .A(round_reg[931]), .B(round_reg[611]), .Z(n53507) );
  ANDN U54923 ( .B(n49056), .A(n51291), .Z(n53501) );
  XOR U54924 ( .A(round_reg[610]), .B(n50822), .Z(n51291) );
  XOR U54925 ( .A(n52588), .B(n52682), .Z(n50822) );
  XOR U54926 ( .A(n53508), .B(n53509), .Z(n52682) );
  XNOR U54927 ( .A(round_reg[34]), .B(round_reg[1314]), .Z(n53509) );
  XOR U54928 ( .A(round_reg[354]), .B(n53510), .Z(n53508) );
  XOR U54929 ( .A(round_reg[994]), .B(round_reg[674]), .Z(n53510) );
  XOR U54930 ( .A(n53511), .B(n53512), .Z(n52588) );
  XNOR U54931 ( .A(round_reg[1505]), .B(round_reg[1185]), .Z(n53512) );
  XOR U54932 ( .A(round_reg[225]), .B(n53513), .Z(n53511) );
  XOR U54933 ( .A(round_reg[865]), .B(round_reg[545]), .Z(n53513) );
  XNOR U54934 ( .A(round_reg[201]), .B(n51660), .Z(n49056) );
  IV U54935 ( .A(n51721), .Z(n51660) );
  XOR U54936 ( .A(n53514), .B(n53515), .Z(n52707) );
  XNOR U54937 ( .A(round_reg[1545]), .B(round_reg[1225]), .Z(n53515) );
  XOR U54938 ( .A(round_reg[265]), .B(n53516), .Z(n53514) );
  XOR U54939 ( .A(round_reg[905]), .B(round_reg[585]), .Z(n53516) );
  XNOR U54940 ( .A(n53517), .B(n53518), .Z(n53167) );
  XNOR U54941 ( .A(round_reg[136]), .B(round_reg[1096]), .Z(n53518) );
  XOR U54942 ( .A(round_reg[1416]), .B(n53519), .Z(n53517) );
  XOR U54943 ( .A(round_reg[776]), .B(round_reg[456]), .Z(n53519) );
  XNOR U54944 ( .A(n45974), .B(n53520), .Z(n53480) );
  XNOR U54945 ( .A(n51269), .B(n49415), .Z(n53520) );
  XNOR U54946 ( .A(n53521), .B(n50866), .Z(n49415) );
  XNOR U54947 ( .A(round_reg[800]), .B(n52000), .Z(n50866) );
  IV U54948 ( .A(n51397), .Z(n52000) );
  XNOR U54949 ( .A(n53522), .B(n53523), .Z(n52362) );
  XNOR U54950 ( .A(round_reg[1504]), .B(round_reg[1184]), .Z(n53523) );
  XOR U54951 ( .A(round_reg[224]), .B(n53524), .Z(n53522) );
  XOR U54952 ( .A(round_reg[864]), .B(round_reg[544]), .Z(n53524) );
  XNOR U54953 ( .A(n53525), .B(n53526), .Z(n53373) );
  XNOR U54954 ( .A(round_reg[1375]), .B(round_reg[1055]), .Z(n53526) );
  XOR U54955 ( .A(round_reg[415]), .B(n53527), .Z(n53525) );
  XOR U54956 ( .A(round_reg[95]), .B(round_reg[735]), .Z(n53527) );
  ANDN U54957 ( .B(n52044), .A(n53528), .Z(n53521) );
  XNOR U54958 ( .A(n53529), .B(n50874), .Z(n51269) );
  XOR U54959 ( .A(round_reg[754]), .B(n50829), .Z(n50874) );
  XNOR U54960 ( .A(n52396), .B(n52511), .Z(n50829) );
  XNOR U54961 ( .A(n53530), .B(n53531), .Z(n52511) );
  XNOR U54962 ( .A(round_reg[1329]), .B(round_reg[1009]), .Z(n53531) );
  XOR U54963 ( .A(round_reg[369]), .B(n53532), .Z(n53530) );
  XOR U54964 ( .A(round_reg[689]), .B(round_reg[49]), .Z(n53532) );
  XOR U54965 ( .A(n53533), .B(n53534), .Z(n52396) );
  XNOR U54966 ( .A(round_reg[1458]), .B(round_reg[1138]), .Z(n53534) );
  XOR U54967 ( .A(round_reg[178]), .B(n53535), .Z(n53533) );
  XOR U54968 ( .A(round_reg[818]), .B(round_reg[498]), .Z(n53535) );
  XOR U54969 ( .A(round_reg[313]), .B(n51672), .Z(n49060) );
  IV U54970 ( .A(n51773), .Z(n51672) );
  XOR U54971 ( .A(n53195), .B(n52100), .Z(n51773) );
  XNOR U54972 ( .A(n53536), .B(n53537), .Z(n52100) );
  XNOR U54973 ( .A(round_reg[1337]), .B(round_reg[1017]), .Z(n53537) );
  XOR U54974 ( .A(round_reg[377]), .B(n53538), .Z(n53536) );
  XOR U54975 ( .A(round_reg[697]), .B(round_reg[57]), .Z(n53538) );
  XOR U54976 ( .A(n53539), .B(n53540), .Z(n53195) );
  XNOR U54977 ( .A(round_reg[1528]), .B(round_reg[1208]), .Z(n53540) );
  XOR U54978 ( .A(round_reg[248]), .B(n53541), .Z(n53539) );
  XOR U54979 ( .A(round_reg[888]), .B(round_reg[568]), .Z(n53541) );
  XNOR U54980 ( .A(round_reg[323]), .B(n51985), .Z(n51294) );
  XNOR U54981 ( .A(n53542), .B(n50870), .Z(n45974) );
  XOR U54982 ( .A(round_reg[833]), .B(n51203), .Z(n50870) );
  IV U54983 ( .A(n52073), .Z(n51203) );
  XNOR U54984 ( .A(n51829), .B(n52850), .Z(n52073) );
  XOR U54985 ( .A(n53543), .B(n53544), .Z(n52850) );
  XNOR U54986 ( .A(round_reg[1537]), .B(round_reg[1217]), .Z(n53544) );
  XOR U54987 ( .A(round_reg[257]), .B(n53545), .Z(n53543) );
  XOR U54988 ( .A(round_reg[897]), .B(round_reg[577]), .Z(n53545) );
  XOR U54989 ( .A(n53546), .B(n53547), .Z(n51829) );
  XNOR U54990 ( .A(round_reg[128]), .B(round_reg[1088]), .Z(n53547) );
  XOR U54991 ( .A(round_reg[1408]), .B(n53548), .Z(n53546) );
  XOR U54992 ( .A(round_reg[768]), .B(round_reg[448]), .Z(n53548) );
  NOR U54993 ( .A(n51297), .B(n49052), .Z(n53542) );
  XOR U54994 ( .A(round_reg[83]), .B(n51548), .Z(n49052) );
  IV U54995 ( .A(n52166), .Z(n51548) );
  XNOR U54996 ( .A(n53139), .B(n52577), .Z(n52166) );
  XNOR U54997 ( .A(n53549), .B(n53550), .Z(n52577) );
  XNOR U54998 ( .A(round_reg[1427]), .B(round_reg[1107]), .Z(n53550) );
  XOR U54999 ( .A(round_reg[147]), .B(n53551), .Z(n53549) );
  XOR U55000 ( .A(round_reg[787]), .B(round_reg[467]), .Z(n53551) );
  XOR U55001 ( .A(n53552), .B(n53553), .Z(n53139) );
  XNOR U55002 ( .A(round_reg[18]), .B(round_reg[1298]), .Z(n53553) );
  XOR U55003 ( .A(round_reg[338]), .B(n53554), .Z(n53552) );
  XOR U55004 ( .A(round_reg[978]), .B(round_reg[658]), .Z(n53554) );
  XOR U55005 ( .A(round_reg[508]), .B(n52072), .Z(n51297) );
  XNOR U55006 ( .A(n51691), .B(n52283), .Z(n52072) );
  XNOR U55007 ( .A(n53555), .B(n53556), .Z(n52283) );
  XNOR U55008 ( .A(round_reg[123]), .B(round_reg[1083]), .Z(n53556) );
  XOR U55009 ( .A(round_reg[1403]), .B(n53557), .Z(n53555) );
  XOR U55010 ( .A(round_reg[763]), .B(round_reg[443]), .Z(n53557) );
  XOR U55011 ( .A(n53558), .B(n53559), .Z(n51691) );
  XNOR U55012 ( .A(round_reg[1532]), .B(round_reg[1212]), .Z(n53559) );
  XOR U55013 ( .A(round_reg[252]), .B(n53560), .Z(n53558) );
  XOR U55014 ( .A(round_reg[892]), .B(round_reg[572]), .Z(n53560) );
  XNOR U55015 ( .A(n53561), .B(n51302), .Z(n52050) );
  IV U55016 ( .A(n53528), .Z(n51302) );
  XOR U55017 ( .A(round_reg[438]), .B(n48445), .Z(n53528) );
  XNOR U55018 ( .A(n53562), .B(n53563), .Z(n51659) );
  XNOR U55019 ( .A(round_reg[1333]), .B(round_reg[1013]), .Z(n53563) );
  XOR U55020 ( .A(round_reg[373]), .B(n53564), .Z(n53562) );
  XOR U55021 ( .A(round_reg[693]), .B(round_reg[53]), .Z(n53564) );
  XOR U55022 ( .A(n53565), .B(n53566), .Z(n53262) );
  XNOR U55023 ( .A(round_reg[1462]), .B(round_reg[1142]), .Z(n53566) );
  XOR U55024 ( .A(round_reg[182]), .B(n53567), .Z(n53565) );
  XOR U55025 ( .A(round_reg[822]), .B(round_reg[502]), .Z(n53567) );
  ANDN U55026 ( .B(n50865), .A(n52044), .Z(n53561) );
  XNOR U55027 ( .A(round_reg[61]), .B(n52354), .Z(n52044) );
  IV U55028 ( .A(n49800), .Z(n52354) );
  XOR U55029 ( .A(n52677), .B(n53568), .Z(n49800) );
  XNOR U55030 ( .A(n53569), .B(n53570), .Z(n52677) );
  XNOR U55031 ( .A(round_reg[125]), .B(round_reg[1085]), .Z(n53570) );
  XOR U55032 ( .A(round_reg[1405]), .B(n53571), .Z(n53569) );
  XOR U55033 ( .A(round_reg[765]), .B(round_reg[445]), .Z(n53571) );
  XOR U55034 ( .A(round_reg[1547]), .B(n51647), .Z(n50865) );
  IV U55035 ( .A(n51399), .Z(n51647) );
  XNOR U55036 ( .A(n53572), .B(n53573), .Z(n52780) );
  XNOR U55037 ( .A(round_reg[1482]), .B(round_reg[1162]), .Z(n53573) );
  XOR U55038 ( .A(round_reg[202]), .B(n53574), .Z(n53572) );
  XOR U55039 ( .A(round_reg[842]), .B(round_reg[522]), .Z(n53574) );
  XNOR U55040 ( .A(n53575), .B(n53576), .Z(n52350) );
  XNOR U55041 ( .A(round_reg[1291]), .B(round_reg[11]), .Z(n53576) );
  XOR U55042 ( .A(round_reg[331]), .B(n53577), .Z(n53575) );
  XOR U55043 ( .A(round_reg[971]), .B(round_reg[651]), .Z(n53577) );
  XOR U55044 ( .A(n48960), .B(n44986), .Z(n44475) );
  XOR U55045 ( .A(n51728), .B(n47094), .Z(n44986) );
  XOR U55046 ( .A(n53578), .B(n53579), .Z(n47094) );
  XNOR U55047 ( .A(n46646), .B(n45406), .Z(n53579) );
  XOR U55048 ( .A(n53580), .B(n46820), .Z(n45406) );
  XOR U55049 ( .A(round_reg[1075]), .B(n51545), .Z(n46820) );
  IV U55050 ( .A(n50444), .Z(n51545) );
  XOR U55051 ( .A(n52377), .B(n51925), .Z(n50444) );
  XOR U55052 ( .A(n53581), .B(n53582), .Z(n51925) );
  XNOR U55053 ( .A(round_reg[1330]), .B(round_reg[1010]), .Z(n53582) );
  XOR U55054 ( .A(round_reg[370]), .B(n53583), .Z(n53581) );
  XOR U55055 ( .A(round_reg[690]), .B(round_reg[50]), .Z(n53583) );
  XOR U55056 ( .A(n53584), .B(n53585), .Z(n52377) );
  XNOR U55057 ( .A(round_reg[1459]), .B(round_reg[1139]), .Z(n53585) );
  XOR U55058 ( .A(round_reg[179]), .B(n53586), .Z(n53584) );
  XOR U55059 ( .A(round_reg[819]), .B(round_reg[499]), .Z(n53586) );
  ANDN U55060 ( .B(n48366), .A(n46484), .Z(n53580) );
  XNOR U55061 ( .A(n53587), .B(n46818), .Z(n46646) );
  XOR U55062 ( .A(round_reg[1124]), .B(n48449), .Z(n46818) );
  XOR U55063 ( .A(n52412), .B(n52476), .Z(n48449) );
  XNOR U55064 ( .A(n53588), .B(n53589), .Z(n52476) );
  XNOR U55065 ( .A(round_reg[1508]), .B(round_reg[1188]), .Z(n53589) );
  XOR U55066 ( .A(round_reg[228]), .B(n53590), .Z(n53588) );
  XOR U55067 ( .A(round_reg[868]), .B(round_reg[548]), .Z(n53590) );
  XNOR U55068 ( .A(n53591), .B(n53592), .Z(n52412) );
  XNOR U55069 ( .A(round_reg[1379]), .B(round_reg[1059]), .Z(n53592) );
  XOR U55070 ( .A(round_reg[419]), .B(n53593), .Z(n53591) );
  XOR U55071 ( .A(round_reg[99]), .B(round_reg[739]), .Z(n53593) );
  ANDN U55072 ( .B(n48369), .A(n46475), .Z(n53587) );
  XNOR U55073 ( .A(round_reg[354]), .B(n49075), .Z(n46475) );
  IV U55074 ( .A(n51954), .Z(n49075) );
  XOR U55075 ( .A(n52467), .B(n52464), .Z(n51954) );
  XNOR U55076 ( .A(n53594), .B(n53595), .Z(n52464) );
  XNOR U55077 ( .A(round_reg[1569]), .B(round_reg[1249]), .Z(n53595) );
  XOR U55078 ( .A(round_reg[289]), .B(n53596), .Z(n53594) );
  XOR U55079 ( .A(round_reg[929]), .B(round_reg[609]), .Z(n53596) );
  XOR U55080 ( .A(n53597), .B(n53598), .Z(n52467) );
  XNOR U55081 ( .A(round_reg[1378]), .B(round_reg[1058]), .Z(n53598) );
  XOR U55082 ( .A(round_reg[418]), .B(n53599), .Z(n53597) );
  XOR U55083 ( .A(round_reg[98]), .B(round_reg[738]), .Z(n53599) );
  XNOR U55084 ( .A(round_reg[721]), .B(n50451), .Z(n48369) );
  XNOR U55085 ( .A(n53260), .B(n52905), .Z(n50451) );
  XNOR U55086 ( .A(n53600), .B(n53601), .Z(n52905) );
  XNOR U55087 ( .A(round_reg[1425]), .B(round_reg[1105]), .Z(n53601) );
  XOR U55088 ( .A(round_reg[145]), .B(n53602), .Z(n53600) );
  XOR U55089 ( .A(round_reg[785]), .B(round_reg[465]), .Z(n53602) );
  XOR U55090 ( .A(n53603), .B(n53604), .Z(n53260) );
  XNOR U55091 ( .A(round_reg[16]), .B(round_reg[1296]), .Z(n53604) );
  XOR U55092 ( .A(round_reg[336]), .B(n53605), .Z(n53603) );
  XOR U55093 ( .A(round_reg[976]), .B(round_reg[656]), .Z(n53605) );
  XOR U55094 ( .A(n44105), .B(n53606), .Z(n53578) );
  XOR U55095 ( .A(n48351), .B(n45290), .Z(n53606) );
  XNOR U55096 ( .A(n53607), .B(n46813), .Z(n45290) );
  XOR U55097 ( .A(round_reg[1214]), .B(n50448), .Z(n46813) );
  XNOR U55098 ( .A(n53608), .B(n53609), .Z(n52450) );
  XNOR U55099 ( .A(round_reg[1598]), .B(round_reg[1278]), .Z(n53609) );
  XOR U55100 ( .A(round_reg[318]), .B(n53610), .Z(n53608) );
  XOR U55101 ( .A(round_reg[958]), .B(round_reg[638]), .Z(n53610) );
  XOR U55102 ( .A(n53611), .B(n53612), .Z(n52774) );
  XNOR U55103 ( .A(round_reg[1469]), .B(round_reg[1149]), .Z(n53612) );
  XOR U55104 ( .A(round_reg[189]), .B(n53613), .Z(n53611) );
  XOR U55105 ( .A(round_reg[829]), .B(round_reg[509]), .Z(n53613) );
  ANDN U55106 ( .B(n48357), .A(n46480), .Z(n53607) );
  XOR U55107 ( .A(round_reg[405]), .B(n48948), .Z(n46480) );
  XNOR U55108 ( .A(n53095), .B(n52399), .Z(n48948) );
  XNOR U55109 ( .A(n53614), .B(n53615), .Z(n52399) );
  XNOR U55110 ( .A(round_reg[20]), .B(round_reg[1300]), .Z(n53615) );
  XOR U55111 ( .A(round_reg[340]), .B(n53616), .Z(n53614) );
  XOR U55112 ( .A(round_reg[980]), .B(round_reg[660]), .Z(n53616) );
  XNOR U55113 ( .A(n53617), .B(n53618), .Z(n53095) );
  XNOR U55114 ( .A(round_reg[1429]), .B(round_reg[1109]), .Z(n53618) );
  XOR U55115 ( .A(round_reg[149]), .B(n53619), .Z(n53617) );
  XOR U55116 ( .A(round_reg[789]), .B(round_reg[469]), .Z(n53619) );
  XOR U55117 ( .A(round_reg[831]), .B(n49081), .Z(n48357) );
  XNOR U55118 ( .A(n52782), .B(n53620), .Z(n49081) );
  XNOR U55119 ( .A(n53621), .B(n53622), .Z(n52782) );
  XNOR U55120 ( .A(round_reg[126]), .B(round_reg[1086]), .Z(n53622) );
  XOR U55121 ( .A(round_reg[1406]), .B(n53623), .Z(n53621) );
  XOR U55122 ( .A(round_reg[766]), .B(round_reg[446]), .Z(n53623) );
  XNOR U55123 ( .A(n53624), .B(n46816), .Z(n48351) );
  XNOR U55124 ( .A(round_reg[1222]), .B(n50815), .Z(n46816) );
  XOR U55125 ( .A(n53625), .B(n53626), .Z(n52542) );
  XNOR U55126 ( .A(round_reg[1477]), .B(round_reg[1157]), .Z(n53626) );
  XOR U55127 ( .A(round_reg[197]), .B(n53627), .Z(n53625) );
  XOR U55128 ( .A(round_reg[837]), .B(round_reg[517]), .Z(n53627) );
  XNOR U55129 ( .A(n53628), .B(n53629), .Z(n52917) );
  XNOR U55130 ( .A(round_reg[326]), .B(round_reg[1286]), .Z(n53629) );
  XOR U55131 ( .A(round_reg[646]), .B(n53630), .Z(n53628) );
  XOR U55132 ( .A(round_reg[966]), .B(round_reg[6]), .Z(n53630) );
  ANDN U55133 ( .B(n48363), .A(n46488), .Z(n53624) );
  XNOR U55134 ( .A(round_reg[475]), .B(n50513), .Z(n46488) );
  IV U55135 ( .A(n51694), .Z(n50513) );
  XOR U55136 ( .A(n52960), .B(n52970), .Z(n51694) );
  XNOR U55137 ( .A(n53631), .B(n53632), .Z(n52970) );
  XNOR U55138 ( .A(round_reg[1370]), .B(round_reg[1050]), .Z(n53632) );
  XOR U55139 ( .A(round_reg[410]), .B(n53633), .Z(n53631) );
  XOR U55140 ( .A(round_reg[90]), .B(round_reg[730]), .Z(n53633) );
  XOR U55141 ( .A(n53634), .B(n53635), .Z(n52960) );
  XNOR U55142 ( .A(round_reg[1499]), .B(round_reg[1179]), .Z(n53635) );
  XOR U55143 ( .A(round_reg[219]), .B(n53636), .Z(n53634) );
  XOR U55144 ( .A(round_reg[859]), .B(round_reg[539]), .Z(n53636) );
  XNOR U55145 ( .A(round_reg[864]), .B(n51161), .Z(n48363) );
  IV U55146 ( .A(n51671), .Z(n51161) );
  XOR U55147 ( .A(n53637), .B(n53067), .Z(n51671) );
  XNOR U55148 ( .A(n53638), .B(n53639), .Z(n53067) );
  XNOR U55149 ( .A(round_reg[1439]), .B(round_reg[1119]), .Z(n53639) );
  XOR U55150 ( .A(round_reg[159]), .B(n53640), .Z(n53638) );
  XOR U55151 ( .A(round_reg[799]), .B(round_reg[479]), .Z(n53640) );
  XNOR U55152 ( .A(n53641), .B(n46810), .Z(n44105) );
  XNOR U55153 ( .A(round_reg[982]), .B(n48945), .Z(n46810) );
  XOR U55154 ( .A(n53084), .B(n52871), .Z(n48945) );
  XOR U55155 ( .A(n53642), .B(n53643), .Z(n52871) );
  XNOR U55156 ( .A(round_reg[1366]), .B(round_reg[1046]), .Z(n53643) );
  XOR U55157 ( .A(round_reg[406]), .B(n53644), .Z(n53642) );
  XOR U55158 ( .A(round_reg[86]), .B(round_reg[726]), .Z(n53644) );
  XOR U55159 ( .A(n53645), .B(n53646), .Z(n53084) );
  XNOR U55160 ( .A(round_reg[1557]), .B(round_reg[1237]), .Z(n53646) );
  XOR U55161 ( .A(round_reg[277]), .B(n53647), .Z(n53645) );
  XOR U55162 ( .A(round_reg[917]), .B(round_reg[597]), .Z(n53647) );
  ANDN U55163 ( .B(n48359), .A(n48956), .Z(n53641) );
  XNOR U55164 ( .A(round_reg[573]), .B(n50837), .Z(n48956) );
  IV U55165 ( .A(n51837), .Z(n50837) );
  XOR U55166 ( .A(n52781), .B(n52810), .Z(n51837) );
  XNOR U55167 ( .A(n53648), .B(n53649), .Z(n52810) );
  XNOR U55168 ( .A(round_reg[1468]), .B(round_reg[1148]), .Z(n53649) );
  XOR U55169 ( .A(round_reg[188]), .B(n53650), .Z(n53648) );
  XOR U55170 ( .A(round_reg[828]), .B(round_reg[508]), .Z(n53650) );
  XOR U55171 ( .A(n53651), .B(n53652), .Z(n52781) );
  XNOR U55172 ( .A(round_reg[1597]), .B(round_reg[1277]), .Z(n53652) );
  XOR U55173 ( .A(round_reg[317]), .B(n53653), .Z(n53651) );
  XOR U55174 ( .A(round_reg[957]), .B(round_reg[637]), .Z(n53653) );
  XNOR U55175 ( .A(round_reg[935]), .B(n50988), .Z(n48359) );
  IV U55176 ( .A(n52170), .Z(n50988) );
  XNOR U55177 ( .A(n53133), .B(n52391), .Z(n52170) );
  XNOR U55178 ( .A(n53654), .B(n53655), .Z(n52391) );
  XNOR U55179 ( .A(round_reg[359]), .B(round_reg[1319]), .Z(n53655) );
  XOR U55180 ( .A(round_reg[39]), .B(n53656), .Z(n53654) );
  XOR U55181 ( .A(round_reg[999]), .B(round_reg[679]), .Z(n53656) );
  XNOR U55182 ( .A(n53657), .B(n53658), .Z(n53133) );
  XNOR U55183 ( .A(round_reg[1510]), .B(round_reg[1190]), .Z(n53658) );
  XOR U55184 ( .A(round_reg[230]), .B(n53659), .Z(n53657) );
  XOR U55185 ( .A(round_reg[870]), .B(round_reg[550]), .Z(n53659) );
  XNOR U55186 ( .A(n53660), .B(n53661), .Z(n51728) );
  XOR U55187 ( .A(n49635), .B(n44923), .Z(n53661) );
  XNOR U55188 ( .A(n53662), .B(n50670), .Z(n44923) );
  XNOR U55189 ( .A(round_reg[404]), .B(n50849), .Z(n50670) );
  XNOR U55190 ( .A(n52637), .B(n53085), .Z(n50849) );
  XNOR U55191 ( .A(n53663), .B(n53664), .Z(n53085) );
  XNOR U55192 ( .A(round_reg[1428]), .B(round_reg[1108]), .Z(n53664) );
  XOR U55193 ( .A(round_reg[148]), .B(n53665), .Z(n53663) );
  XOR U55194 ( .A(round_reg[788]), .B(round_reg[468]), .Z(n53665) );
  XOR U55195 ( .A(n53666), .B(n53667), .Z(n52637) );
  XNOR U55196 ( .A(round_reg[19]), .B(round_reg[1299]), .Z(n53667) );
  XOR U55197 ( .A(round_reg[339]), .B(n53668), .Z(n53666) );
  XOR U55198 ( .A(round_reg[979]), .B(round_reg[659]), .Z(n53668) );
  ANDN U55199 ( .B(n48972), .A(n46607), .Z(n53662) );
  XOR U55200 ( .A(round_reg[1577]), .B(n52701), .Z(n46607) );
  IV U55201 ( .A(n51520), .Z(n52701) );
  XNOR U55202 ( .A(n51843), .B(n52964), .Z(n51520) );
  XNOR U55203 ( .A(n53669), .B(n53670), .Z(n52964) );
  XNOR U55204 ( .A(round_reg[1512]), .B(round_reg[1192]), .Z(n53670) );
  XOR U55205 ( .A(round_reg[232]), .B(n53671), .Z(n53669) );
  XOR U55206 ( .A(round_reg[872]), .B(round_reg[552]), .Z(n53671) );
  XOR U55207 ( .A(n53672), .B(n53673), .Z(n51843) );
  XNOR U55208 ( .A(round_reg[1321]), .B(round_reg[1001]), .Z(n53673) );
  XOR U55209 ( .A(round_reg[361]), .B(n53674), .Z(n53672) );
  XOR U55210 ( .A(round_reg[681]), .B(round_reg[41]), .Z(n53674) );
  XOR U55211 ( .A(round_reg[27]), .B(n49955), .Z(n48972) );
  XOR U55212 ( .A(n53675), .B(n53676), .Z(n52887) );
  XNOR U55213 ( .A(round_reg[1562]), .B(round_reg[1242]), .Z(n53676) );
  XOR U55214 ( .A(round_reg[282]), .B(n53677), .Z(n53675) );
  XOR U55215 ( .A(round_reg[922]), .B(round_reg[602]), .Z(n53677) );
  XOR U55216 ( .A(n53678), .B(n53679), .Z(n52773) );
  XNOR U55217 ( .A(round_reg[1371]), .B(round_reg[1051]), .Z(n53679) );
  XOR U55218 ( .A(round_reg[411]), .B(n53680), .Z(n53678) );
  XOR U55219 ( .A(round_reg[91]), .B(round_reg[731]), .Z(n53680) );
  XOR U55220 ( .A(n53681), .B(n50663), .Z(n49635) );
  XNOR U55221 ( .A(round_reg[353]), .B(n50452), .Z(n50663) );
  XNOR U55222 ( .A(n53637), .B(n52606), .Z(n50452) );
  XNOR U55223 ( .A(n53682), .B(n53683), .Z(n52606) );
  XNOR U55224 ( .A(round_reg[1377]), .B(round_reg[1057]), .Z(n53683) );
  XOR U55225 ( .A(round_reg[417]), .B(n53684), .Z(n53682) );
  XOR U55226 ( .A(round_reg[97]), .B(round_reg[737]), .Z(n53684) );
  XOR U55227 ( .A(n53685), .B(n53686), .Z(n53637) );
  XNOR U55228 ( .A(round_reg[1568]), .B(round_reg[1248]), .Z(n53686) );
  XOR U55229 ( .A(round_reg[288]), .B(n53687), .Z(n53685) );
  XOR U55230 ( .A(round_reg[928]), .B(round_reg[608]), .Z(n53687) );
  XNOR U55231 ( .A(round_reg[1512]), .B(n52538), .Z(n46621) );
  XOR U55232 ( .A(round_reg[279]), .B(n50738), .Z(n48980) );
  XNOR U55233 ( .A(n53688), .B(n53689), .Z(n51945) );
  XNOR U55234 ( .A(round_reg[23]), .B(round_reg[1303]), .Z(n53689) );
  XOR U55235 ( .A(round_reg[343]), .B(n53690), .Z(n53688) );
  XOR U55236 ( .A(round_reg[983]), .B(round_reg[663]), .Z(n53690) );
  XOR U55237 ( .A(n53691), .B(n53692), .Z(n52126) );
  XNOR U55238 ( .A(round_reg[1494]), .B(round_reg[1174]), .Z(n53692) );
  XOR U55239 ( .A(round_reg[214]), .B(n53693), .Z(n53691) );
  XOR U55240 ( .A(round_reg[854]), .B(round_reg[534]), .Z(n53693) );
  XOR U55241 ( .A(n42661), .B(n53694), .Z(n53660) );
  XOR U55242 ( .A(n44185), .B(n50658), .Z(n53694) );
  XNOR U55243 ( .A(n53695), .B(n50668), .Z(n50658) );
  XOR U55244 ( .A(round_reg[572]), .B(n49077), .Z(n50668) );
  IV U55245 ( .A(n50522), .Z(n49077) );
  XNOR U55246 ( .A(n53092), .B(n53568), .Z(n50522) );
  XNOR U55247 ( .A(n53696), .B(n53697), .Z(n53568) );
  XNOR U55248 ( .A(round_reg[1596]), .B(round_reg[1276]), .Z(n53697) );
  XOR U55249 ( .A(round_reg[316]), .B(n53698), .Z(n53696) );
  XOR U55250 ( .A(round_reg[956]), .B(round_reg[636]), .Z(n53698) );
  XNOR U55251 ( .A(n53699), .B(n53700), .Z(n53092) );
  XNOR U55252 ( .A(round_reg[1467]), .B(round_reg[1147]), .Z(n53700) );
  XOR U55253 ( .A(round_reg[187]), .B(n53701), .Z(n53699) );
  XOR U55254 ( .A(round_reg[827]), .B(round_reg[507]), .Z(n53701) );
  ANDN U55255 ( .B(n48974), .A(n46611), .Z(n53695) );
  XOR U55256 ( .A(round_reg[1357]), .B(n49863), .Z(n46611) );
  IV U55257 ( .A(n48869), .Z(n49863) );
  XOR U55258 ( .A(n53381), .B(n51922), .Z(n48869) );
  XOR U55259 ( .A(n53702), .B(n53703), .Z(n51922) );
  XNOR U55260 ( .A(round_reg[12]), .B(round_reg[1292]), .Z(n53703) );
  XOR U55261 ( .A(round_reg[332]), .B(n53704), .Z(n53702) );
  XOR U55262 ( .A(round_reg[972]), .B(round_reg[652]), .Z(n53704) );
  XOR U55263 ( .A(n53705), .B(n53706), .Z(n53381) );
  XNOR U55264 ( .A(round_reg[141]), .B(round_reg[1101]), .Z(n53706) );
  XOR U55265 ( .A(round_reg[1421]), .B(n53707), .Z(n53705) );
  XOR U55266 ( .A(round_reg[781]), .B(round_reg[461]), .Z(n53707) );
  XOR U55267 ( .A(round_reg[172]), .B(n48365), .Z(n48974) );
  XNOR U55268 ( .A(n53708), .B(n53709), .Z(n53298) );
  XNOR U55269 ( .A(round_reg[107]), .B(round_reg[1067]), .Z(n53709) );
  XOR U55270 ( .A(round_reg[1387]), .B(n53710), .Z(n53708) );
  XOR U55271 ( .A(round_reg[747]), .B(round_reg[427]), .Z(n53710) );
  XNOR U55272 ( .A(n53711), .B(n53712), .Z(n52729) );
  XNOR U55273 ( .A(round_reg[1516]), .B(round_reg[1196]), .Z(n53712) );
  XOR U55274 ( .A(round_reg[236]), .B(n53713), .Z(n53711) );
  XOR U55275 ( .A(round_reg[876]), .B(round_reg[556]), .Z(n53713) );
  XNOR U55276 ( .A(n53714), .B(n50666), .Z(n44185) );
  XOR U55277 ( .A(round_reg[474]), .B(n52807), .Z(n50666) );
  IV U55278 ( .A(n49792), .Z(n52807) );
  XNOR U55279 ( .A(n52563), .B(n52172), .Z(n49792) );
  XNOR U55280 ( .A(n53715), .B(n53716), .Z(n52172) );
  XNOR U55281 ( .A(round_reg[1369]), .B(round_reg[1049]), .Z(n53716) );
  XOR U55282 ( .A(round_reg[409]), .B(n53717), .Z(n53715) );
  XOR U55283 ( .A(round_reg[89]), .B(round_reg[729]), .Z(n53717) );
  XNOR U55284 ( .A(n53718), .B(n53719), .Z(n52563) );
  XNOR U55285 ( .A(round_reg[1498]), .B(round_reg[1178]), .Z(n53719) );
  XOR U55286 ( .A(round_reg[218]), .B(n53720), .Z(n53718) );
  XOR U55287 ( .A(round_reg[858]), .B(round_reg[538]), .Z(n53720) );
  ANDN U55288 ( .B(n48978), .A(n46950), .Z(n53714) );
  XNOR U55289 ( .A(round_reg[1294]), .B(n50765), .Z(n46950) );
  IV U55290 ( .A(n51491), .Z(n50765) );
  XOR U55291 ( .A(n52434), .B(n53385), .Z(n51491) );
  XNOR U55292 ( .A(n53721), .B(n53722), .Z(n53385) );
  XNOR U55293 ( .A(round_reg[1358]), .B(round_reg[1038]), .Z(n53722) );
  XOR U55294 ( .A(round_reg[398]), .B(n53723), .Z(n53721) );
  XOR U55295 ( .A(round_reg[78]), .B(round_reg[718]), .Z(n53723) );
  XOR U55296 ( .A(n53724), .B(n53725), .Z(n52434) );
  XNOR U55297 ( .A(round_reg[1549]), .B(round_reg[1229]), .Z(n53725) );
  XOR U55298 ( .A(round_reg[269]), .B(n53726), .Z(n53724) );
  XOR U55299 ( .A(round_reg[909]), .B(round_reg[589]), .Z(n53726) );
  XOR U55300 ( .A(round_reg[113]), .B(n50514), .Z(n48978) );
  XOR U55301 ( .A(n52761), .B(n52628), .Z(n50514) );
  XNOR U55302 ( .A(n53727), .B(n53728), .Z(n52628) );
  XNOR U55303 ( .A(round_reg[1457]), .B(round_reg[1137]), .Z(n53728) );
  XOR U55304 ( .A(round_reg[177]), .B(n53729), .Z(n53727) );
  XOR U55305 ( .A(round_reg[817]), .B(round_reg[497]), .Z(n53729) );
  XOR U55306 ( .A(n53730), .B(n53731), .Z(n52761) );
  XNOR U55307 ( .A(round_reg[1328]), .B(round_reg[1008]), .Z(n53731) );
  XOR U55308 ( .A(round_reg[368]), .B(n53732), .Z(n53730) );
  XOR U55309 ( .A(round_reg[688]), .B(round_reg[48]), .Z(n53732) );
  XNOR U55310 ( .A(n53733), .B(n52196), .Z(n42661) );
  XOR U55311 ( .A(round_reg[576]), .B(n51199), .Z(n52196) );
  XNOR U55312 ( .A(n53734), .B(n53735), .Z(n53620) );
  XNOR U55313 ( .A(round_reg[1535]), .B(round_reg[1215]), .Z(n53735) );
  XOR U55314 ( .A(round_reg[255]), .B(n53736), .Z(n53734) );
  XOR U55315 ( .A(round_reg[895]), .B(round_reg[575]), .Z(n53736) );
  XOR U55316 ( .A(n53737), .B(n53738), .Z(n53313) );
  XNOR U55317 ( .A(round_reg[1280]), .B(round_reg[0]), .Z(n53738) );
  XOR U55318 ( .A(round_reg[320]), .B(n53739), .Z(n53737) );
  XOR U55319 ( .A(round_reg[960]), .B(round_reg[640]), .Z(n53739) );
  ANDN U55320 ( .B(n51740), .A(n46617), .Z(n53733) );
  XOR U55321 ( .A(round_reg[1451]), .B(n51135), .Z(n46617) );
  XNOR U55322 ( .A(n52952), .B(n52429), .Z(n51135) );
  XNOR U55323 ( .A(n53740), .B(n53741), .Z(n52429) );
  XNOR U55324 ( .A(round_reg[106]), .B(round_reg[1066]), .Z(n53741) );
  XOR U55325 ( .A(round_reg[1386]), .B(n53742), .Z(n53740) );
  XOR U55326 ( .A(round_reg[746]), .B(round_reg[426]), .Z(n53742) );
  XNOR U55327 ( .A(n53743), .B(n53744), .Z(n52952) );
  XNOR U55328 ( .A(round_reg[1515]), .B(round_reg[1195]), .Z(n53744) );
  XOR U55329 ( .A(round_reg[235]), .B(n53745), .Z(n53743) );
  XOR U55330 ( .A(round_reg[875]), .B(round_reg[555]), .Z(n53745) );
  XNOR U55331 ( .A(round_reg[231]), .B(n51947), .Z(n51740) );
  XNOR U55332 ( .A(n52857), .B(n52643), .Z(n51947) );
  XNOR U55333 ( .A(n53746), .B(n53747), .Z(n52643) );
  XNOR U55334 ( .A(round_reg[1575]), .B(round_reg[1255]), .Z(n53747) );
  XOR U55335 ( .A(round_reg[295]), .B(n53748), .Z(n53746) );
  XOR U55336 ( .A(round_reg[935]), .B(round_reg[615]), .Z(n53748) );
  XOR U55337 ( .A(n53749), .B(n53750), .Z(n52857) );
  XNOR U55338 ( .A(round_reg[1446]), .B(round_reg[1126]), .Z(n53750) );
  XOR U55339 ( .A(round_reg[166]), .B(n53751), .Z(n53749) );
  XOR U55340 ( .A(round_reg[806]), .B(round_reg[486]), .Z(n53751) );
  XOR U55341 ( .A(n53752), .B(n48366), .Z(n48960) );
  XNOR U55342 ( .A(round_reg[643]), .B(n51985), .Z(n48366) );
  XNOR U55343 ( .A(n53476), .B(n52988), .Z(n51985) );
  XNOR U55344 ( .A(n53753), .B(n53754), .Z(n52988) );
  XNOR U55345 ( .A(round_reg[1538]), .B(round_reg[1218]), .Z(n53754) );
  XOR U55346 ( .A(round_reg[258]), .B(n53755), .Z(n53753) );
  XOR U55347 ( .A(round_reg[898]), .B(round_reg[578]), .Z(n53755) );
  XOR U55348 ( .A(n53756), .B(n53757), .Z(n53476) );
  XNOR U55349 ( .A(round_reg[1347]), .B(round_reg[1027]), .Z(n53757) );
  XOR U55350 ( .A(round_reg[387]), .B(n53758), .Z(n53756) );
  XOR U55351 ( .A(round_reg[707]), .B(round_reg[67]), .Z(n53758) );
  ANDN U55352 ( .B(n46484), .A(n46486), .Z(n53752) );
  XOR U55353 ( .A(round_reg[232]), .B(n50756), .Z(n46486) );
  IV U55354 ( .A(n52538), .Z(n50756) );
  XNOR U55355 ( .A(n52622), .B(n52383), .Z(n52538) );
  XNOR U55356 ( .A(n53759), .B(n53760), .Z(n52383) );
  XNOR U55357 ( .A(round_reg[1576]), .B(round_reg[1256]), .Z(n53760) );
  XOR U55358 ( .A(round_reg[296]), .B(n53761), .Z(n53759) );
  XOR U55359 ( .A(round_reg[936]), .B(round_reg[616]), .Z(n53761) );
  XOR U55360 ( .A(n53762), .B(n53763), .Z(n52622) );
  XNOR U55361 ( .A(round_reg[1447]), .B(round_reg[1127]), .Z(n53763) );
  XOR U55362 ( .A(round_reg[167]), .B(n53764), .Z(n53762) );
  XOR U55363 ( .A(round_reg[807]), .B(round_reg[487]), .Z(n53764) );
  XOR U55364 ( .A(round_reg[577]), .B(n49857), .Z(n46484) );
  XNOR U55365 ( .A(n53765), .B(n53766), .Z(n52422) );
  XNOR U55366 ( .A(round_reg[1472]), .B(round_reg[1152]), .Z(n53766) );
  XOR U55367 ( .A(round_reg[192]), .B(n53767), .Z(n53765) );
  XOR U55368 ( .A(round_reg[832]), .B(round_reg[512]), .Z(n53767) );
  XNOR U55369 ( .A(n53768), .B(n53769), .Z(n53104) );
  XNOR U55370 ( .A(round_reg[1]), .B(round_reg[1281]), .Z(n53769) );
  XOR U55371 ( .A(round_reg[321]), .B(n53770), .Z(n53768) );
  XOR U55372 ( .A(round_reg[961]), .B(round_reg[641]), .Z(n53770) );
  IV U55373 ( .A(init), .Z(n1029) );
endmodule

