
module mult_N64_CC64 ( clk, rst, a, b, c );
  input [63:0] a;
  input [0:0] b;
  output [127:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378;
  wire   [127:0] sreg;

  DFF \sreg_reg[126]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(sreg[126]) );
  DFF \sreg_reg[125]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(sreg[125]) );
  DFF \sreg_reg[124]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(sreg[124]) );
  DFF \sreg_reg[123]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(sreg[123]) );
  DFF \sreg_reg[122]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(sreg[122]) );
  DFF \sreg_reg[121]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(sreg[121]) );
  DFF \sreg_reg[120]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(sreg[120]) );
  DFF \sreg_reg[119]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(sreg[119]) );
  DFF \sreg_reg[118]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(sreg[118]) );
  DFF \sreg_reg[117]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(sreg[117]) );
  DFF \sreg_reg[116]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(sreg[116]) );
  DFF \sreg_reg[115]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(sreg[115]) );
  DFF \sreg_reg[114]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(sreg[114]) );
  DFF \sreg_reg[113]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(sreg[113]) );
  DFF \sreg_reg[112]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(sreg[112]) );
  DFF \sreg_reg[111]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(sreg[111]) );
  DFF \sreg_reg[110]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(sreg[110]) );
  DFF \sreg_reg[109]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(sreg[109]) );
  DFF \sreg_reg[108]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(sreg[108]) );
  DFF \sreg_reg[107]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(sreg[107]) );
  DFF \sreg_reg[106]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(sreg[106]) );
  DFF \sreg_reg[105]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(sreg[105]) );
  DFF \sreg_reg[104]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(sreg[104]) );
  DFF \sreg_reg[103]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(sreg[103]) );
  DFF \sreg_reg[102]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(sreg[102]) );
  DFF \sreg_reg[101]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(sreg[101]) );
  DFF \sreg_reg[100]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(sreg[100]) );
  DFF \sreg_reg[99]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(sreg[99]) );
  DFF \sreg_reg[98]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(sreg[98]) );
  DFF \sreg_reg[97]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(sreg[97]) );
  DFF \sreg_reg[96]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(sreg[96]) );
  DFF \sreg_reg[95]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(sreg[95]) );
  DFF \sreg_reg[94]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(sreg[94]) );
  DFF \sreg_reg[93]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(sreg[93]) );
  DFF \sreg_reg[92]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(sreg[92]) );
  DFF \sreg_reg[91]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(sreg[91]) );
  DFF \sreg_reg[90]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(sreg[90]) );
  DFF \sreg_reg[89]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(sreg[89]) );
  DFF \sreg_reg[88]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(sreg[88]) );
  DFF \sreg_reg[87]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(sreg[87]) );
  DFF \sreg_reg[86]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(sreg[86]) );
  DFF \sreg_reg[85]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(sreg[85]) );
  DFF \sreg_reg[84]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(sreg[84]) );
  DFF \sreg_reg[83]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(sreg[83]) );
  DFF \sreg_reg[82]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(sreg[82]) );
  DFF \sreg_reg[81]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(sreg[81]) );
  DFF \sreg_reg[80]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(sreg[80]) );
  DFF \sreg_reg[79]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(sreg[79]) );
  DFF \sreg_reg[78]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(sreg[78]) );
  DFF \sreg_reg[77]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(sreg[77]) );
  DFF \sreg_reg[76]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(sreg[76]) );
  DFF \sreg_reg[75]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(sreg[75]) );
  DFF \sreg_reg[74]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(sreg[74]) );
  DFF \sreg_reg[73]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(sreg[73]) );
  DFF \sreg_reg[72]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(sreg[72]) );
  DFF \sreg_reg[71]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(sreg[71]) );
  DFF \sreg_reg[70]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(sreg[70]) );
  DFF \sreg_reg[69]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(sreg[69]) );
  DFF \sreg_reg[68]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(sreg[68]) );
  DFF \sreg_reg[67]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(sreg[67]) );
  DFF \sreg_reg[66]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(sreg[66]) );
  DFF \sreg_reg[65]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(sreg[65]) );
  DFF \sreg_reg[64]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(sreg[64]) );
  DFF \sreg_reg[63]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(sreg[63]) );
  DFF \sreg_reg[62]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[61]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[7]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[6]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[5]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[4]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[3]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[2]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[1]), .CLK(clk), .RST(rst), .Q(c[0]) );
  XOR U4 ( .A(sreg[66]), .B(n195), .Z(n1) );
  NANDN U5 ( .A(n196), .B(n1), .Z(n2) );
  NAND U6 ( .A(sreg[66]), .B(n195), .Z(n3) );
  AND U7 ( .A(n2), .B(n3), .Z(n199) );
  XOR U8 ( .A(sreg[69]), .B(n204), .Z(n4) );
  NANDN U9 ( .A(n205), .B(n4), .Z(n5) );
  NAND U10 ( .A(sreg[69]), .B(n204), .Z(n6) );
  AND U11 ( .A(n5), .B(n6), .Z(n208) );
  XOR U12 ( .A(sreg[72]), .B(n213), .Z(n7) );
  NANDN U13 ( .A(n214), .B(n7), .Z(n8) );
  NAND U14 ( .A(sreg[72]), .B(n213), .Z(n9) );
  AND U15 ( .A(n8), .B(n9), .Z(n217) );
  XOR U16 ( .A(sreg[75]), .B(n222), .Z(n10) );
  NANDN U17 ( .A(n223), .B(n10), .Z(n11) );
  NAND U18 ( .A(sreg[75]), .B(n222), .Z(n12) );
  AND U19 ( .A(n11), .B(n12), .Z(n226) );
  XOR U20 ( .A(sreg[78]), .B(n231), .Z(n13) );
  NANDN U21 ( .A(n232), .B(n13), .Z(n14) );
  NAND U22 ( .A(sreg[78]), .B(n231), .Z(n15) );
  AND U23 ( .A(n14), .B(n15), .Z(n235) );
  XOR U24 ( .A(sreg[81]), .B(n240), .Z(n16) );
  NANDN U25 ( .A(n241), .B(n16), .Z(n17) );
  NAND U26 ( .A(sreg[81]), .B(n240), .Z(n18) );
  AND U27 ( .A(n17), .B(n18), .Z(n244) );
  XOR U28 ( .A(sreg[84]), .B(n249), .Z(n19) );
  NANDN U29 ( .A(n250), .B(n19), .Z(n20) );
  NAND U30 ( .A(sreg[84]), .B(n249), .Z(n21) );
  AND U31 ( .A(n20), .B(n21), .Z(n253) );
  XOR U32 ( .A(sreg[87]), .B(n258), .Z(n22) );
  NANDN U33 ( .A(n259), .B(n22), .Z(n23) );
  NAND U34 ( .A(sreg[87]), .B(n258), .Z(n24) );
  AND U35 ( .A(n23), .B(n24), .Z(n262) );
  XOR U36 ( .A(sreg[90]), .B(n267), .Z(n25) );
  NANDN U37 ( .A(n268), .B(n25), .Z(n26) );
  NAND U38 ( .A(sreg[90]), .B(n267), .Z(n27) );
  AND U39 ( .A(n26), .B(n27), .Z(n271) );
  XOR U40 ( .A(sreg[93]), .B(n276), .Z(n28) );
  NANDN U41 ( .A(n277), .B(n28), .Z(n29) );
  NAND U42 ( .A(sreg[93]), .B(n276), .Z(n30) );
  AND U43 ( .A(n29), .B(n30), .Z(n280) );
  XOR U44 ( .A(sreg[96]), .B(n285), .Z(n31) );
  NANDN U45 ( .A(n286), .B(n31), .Z(n32) );
  NAND U46 ( .A(sreg[96]), .B(n285), .Z(n33) );
  AND U47 ( .A(n32), .B(n33), .Z(n289) );
  XOR U48 ( .A(sreg[99]), .B(n294), .Z(n34) );
  NANDN U49 ( .A(n295), .B(n34), .Z(n35) );
  NAND U50 ( .A(sreg[99]), .B(n294), .Z(n36) );
  AND U51 ( .A(n35), .B(n36), .Z(n298) );
  XOR U52 ( .A(sreg[102]), .B(n303), .Z(n37) );
  NANDN U53 ( .A(n304), .B(n37), .Z(n38) );
  NAND U54 ( .A(sreg[102]), .B(n303), .Z(n39) );
  AND U55 ( .A(n38), .B(n39), .Z(n307) );
  XOR U56 ( .A(sreg[105]), .B(n312), .Z(n40) );
  NANDN U57 ( .A(n313), .B(n40), .Z(n41) );
  NAND U58 ( .A(sreg[105]), .B(n312), .Z(n42) );
  AND U59 ( .A(n41), .B(n42), .Z(n316) );
  XOR U60 ( .A(sreg[108]), .B(n321), .Z(n43) );
  NANDN U61 ( .A(n322), .B(n43), .Z(n44) );
  NAND U62 ( .A(sreg[108]), .B(n321), .Z(n45) );
  AND U63 ( .A(n44), .B(n45), .Z(n325) );
  XOR U64 ( .A(sreg[111]), .B(n330), .Z(n46) );
  NANDN U65 ( .A(n331), .B(n46), .Z(n47) );
  NAND U66 ( .A(sreg[111]), .B(n330), .Z(n48) );
  AND U67 ( .A(n47), .B(n48), .Z(n334) );
  XOR U68 ( .A(sreg[114]), .B(n339), .Z(n49) );
  NANDN U69 ( .A(n340), .B(n49), .Z(n50) );
  NAND U70 ( .A(sreg[114]), .B(n339), .Z(n51) );
  AND U71 ( .A(n50), .B(n51), .Z(n343) );
  XOR U72 ( .A(sreg[117]), .B(n348), .Z(n52) );
  NANDN U73 ( .A(n349), .B(n52), .Z(n53) );
  NAND U74 ( .A(sreg[117]), .B(n348), .Z(n54) );
  AND U75 ( .A(n53), .B(n54), .Z(n352) );
  XOR U76 ( .A(sreg[120]), .B(n357), .Z(n55) );
  NANDN U77 ( .A(n358), .B(n55), .Z(n56) );
  NAND U78 ( .A(sreg[120]), .B(n357), .Z(n57) );
  AND U79 ( .A(n56), .B(n57), .Z(n361) );
  XOR U80 ( .A(sreg[123]), .B(n366), .Z(n58) );
  NANDN U81 ( .A(n367), .B(n58), .Z(n59) );
  NAND U82 ( .A(sreg[123]), .B(n366), .Z(n60) );
  AND U83 ( .A(n59), .B(n60), .Z(n370) );
  XOR U84 ( .A(n189), .B(sreg[64]), .Z(n61) );
  NANDN U85 ( .A(n190), .B(n61), .Z(n62) );
  NAND U86 ( .A(n189), .B(sreg[64]), .Z(n63) );
  AND U87 ( .A(n62), .B(n63), .Z(n193) );
  XOR U88 ( .A(sreg[67]), .B(n198), .Z(n64) );
  NANDN U89 ( .A(n199), .B(n64), .Z(n65) );
  NAND U90 ( .A(sreg[67]), .B(n198), .Z(n66) );
  AND U91 ( .A(n65), .B(n66), .Z(n202) );
  XOR U92 ( .A(sreg[70]), .B(n207), .Z(n67) );
  NANDN U93 ( .A(n208), .B(n67), .Z(n68) );
  NAND U94 ( .A(sreg[70]), .B(n207), .Z(n69) );
  AND U95 ( .A(n68), .B(n69), .Z(n211) );
  XOR U96 ( .A(sreg[73]), .B(n216), .Z(n70) );
  NANDN U97 ( .A(n217), .B(n70), .Z(n71) );
  NAND U98 ( .A(sreg[73]), .B(n216), .Z(n72) );
  AND U99 ( .A(n71), .B(n72), .Z(n220) );
  XOR U100 ( .A(sreg[76]), .B(n225), .Z(n73) );
  NANDN U101 ( .A(n226), .B(n73), .Z(n74) );
  NAND U102 ( .A(sreg[76]), .B(n225), .Z(n75) );
  AND U103 ( .A(n74), .B(n75), .Z(n229) );
  XOR U104 ( .A(sreg[79]), .B(n234), .Z(n76) );
  NANDN U105 ( .A(n235), .B(n76), .Z(n77) );
  NAND U106 ( .A(sreg[79]), .B(n234), .Z(n78) );
  AND U107 ( .A(n77), .B(n78), .Z(n238) );
  XOR U108 ( .A(sreg[82]), .B(n243), .Z(n79) );
  NANDN U109 ( .A(n244), .B(n79), .Z(n80) );
  NAND U110 ( .A(sreg[82]), .B(n243), .Z(n81) );
  AND U111 ( .A(n80), .B(n81), .Z(n247) );
  XOR U112 ( .A(sreg[85]), .B(n252), .Z(n82) );
  NANDN U113 ( .A(n253), .B(n82), .Z(n83) );
  NAND U114 ( .A(sreg[85]), .B(n252), .Z(n84) );
  AND U115 ( .A(n83), .B(n84), .Z(n256) );
  XOR U116 ( .A(sreg[88]), .B(n261), .Z(n85) );
  NANDN U117 ( .A(n262), .B(n85), .Z(n86) );
  NAND U118 ( .A(sreg[88]), .B(n261), .Z(n87) );
  AND U119 ( .A(n86), .B(n87), .Z(n265) );
  XOR U120 ( .A(sreg[91]), .B(n270), .Z(n88) );
  NANDN U121 ( .A(n271), .B(n88), .Z(n89) );
  NAND U122 ( .A(sreg[91]), .B(n270), .Z(n90) );
  AND U123 ( .A(n89), .B(n90), .Z(n274) );
  XOR U124 ( .A(sreg[94]), .B(n279), .Z(n91) );
  NANDN U125 ( .A(n280), .B(n91), .Z(n92) );
  NAND U126 ( .A(sreg[94]), .B(n279), .Z(n93) );
  AND U127 ( .A(n92), .B(n93), .Z(n283) );
  XOR U128 ( .A(sreg[97]), .B(n288), .Z(n94) );
  NANDN U129 ( .A(n289), .B(n94), .Z(n95) );
  NAND U130 ( .A(sreg[97]), .B(n288), .Z(n96) );
  AND U131 ( .A(n95), .B(n96), .Z(n292) );
  XOR U132 ( .A(sreg[100]), .B(n297), .Z(n97) );
  NANDN U133 ( .A(n298), .B(n97), .Z(n98) );
  NAND U134 ( .A(sreg[100]), .B(n297), .Z(n99) );
  AND U135 ( .A(n98), .B(n99), .Z(n301) );
  XOR U136 ( .A(sreg[103]), .B(n306), .Z(n100) );
  NANDN U137 ( .A(n307), .B(n100), .Z(n101) );
  NAND U138 ( .A(sreg[103]), .B(n306), .Z(n102) );
  AND U139 ( .A(n101), .B(n102), .Z(n310) );
  XOR U140 ( .A(sreg[106]), .B(n315), .Z(n103) );
  NANDN U141 ( .A(n316), .B(n103), .Z(n104) );
  NAND U142 ( .A(sreg[106]), .B(n315), .Z(n105) );
  AND U143 ( .A(n104), .B(n105), .Z(n319) );
  XOR U144 ( .A(sreg[109]), .B(n324), .Z(n106) );
  NANDN U145 ( .A(n325), .B(n106), .Z(n107) );
  NAND U146 ( .A(sreg[109]), .B(n324), .Z(n108) );
  AND U147 ( .A(n107), .B(n108), .Z(n328) );
  XOR U148 ( .A(sreg[112]), .B(n333), .Z(n109) );
  NANDN U149 ( .A(n334), .B(n109), .Z(n110) );
  NAND U150 ( .A(sreg[112]), .B(n333), .Z(n111) );
  AND U151 ( .A(n110), .B(n111), .Z(n337) );
  XOR U152 ( .A(sreg[115]), .B(n342), .Z(n112) );
  NANDN U153 ( .A(n343), .B(n112), .Z(n113) );
  NAND U154 ( .A(sreg[115]), .B(n342), .Z(n114) );
  AND U155 ( .A(n113), .B(n114), .Z(n346) );
  XOR U156 ( .A(sreg[118]), .B(n351), .Z(n115) );
  NANDN U157 ( .A(n352), .B(n115), .Z(n116) );
  NAND U158 ( .A(sreg[118]), .B(n351), .Z(n117) );
  AND U159 ( .A(n116), .B(n117), .Z(n355) );
  XOR U160 ( .A(sreg[121]), .B(n360), .Z(n118) );
  NANDN U161 ( .A(n361), .B(n118), .Z(n119) );
  NAND U162 ( .A(sreg[121]), .B(n360), .Z(n120) );
  AND U163 ( .A(n119), .B(n120), .Z(n364) );
  XOR U164 ( .A(sreg[124]), .B(n369), .Z(n121) );
  NANDN U165 ( .A(n370), .B(n121), .Z(n122) );
  NAND U166 ( .A(sreg[124]), .B(n369), .Z(n123) );
  AND U167 ( .A(n122), .B(n123), .Z(n373) );
  XOR U168 ( .A(sreg[65]), .B(n192), .Z(n124) );
  NANDN U169 ( .A(n193), .B(n124), .Z(n125) );
  NAND U170 ( .A(sreg[65]), .B(n192), .Z(n126) );
  AND U171 ( .A(n125), .B(n126), .Z(n196) );
  XOR U172 ( .A(sreg[68]), .B(n201), .Z(n127) );
  NANDN U173 ( .A(n202), .B(n127), .Z(n128) );
  NAND U174 ( .A(sreg[68]), .B(n201), .Z(n129) );
  AND U175 ( .A(n128), .B(n129), .Z(n205) );
  XOR U176 ( .A(sreg[71]), .B(n210), .Z(n130) );
  NANDN U177 ( .A(n211), .B(n130), .Z(n131) );
  NAND U178 ( .A(sreg[71]), .B(n210), .Z(n132) );
  AND U179 ( .A(n131), .B(n132), .Z(n214) );
  XOR U180 ( .A(sreg[74]), .B(n219), .Z(n133) );
  NANDN U181 ( .A(n220), .B(n133), .Z(n134) );
  NAND U182 ( .A(sreg[74]), .B(n219), .Z(n135) );
  AND U183 ( .A(n134), .B(n135), .Z(n223) );
  XOR U184 ( .A(sreg[77]), .B(n228), .Z(n136) );
  NANDN U185 ( .A(n229), .B(n136), .Z(n137) );
  NAND U186 ( .A(sreg[77]), .B(n228), .Z(n138) );
  AND U187 ( .A(n137), .B(n138), .Z(n232) );
  XOR U188 ( .A(sreg[80]), .B(n237), .Z(n139) );
  NANDN U189 ( .A(n238), .B(n139), .Z(n140) );
  NAND U190 ( .A(sreg[80]), .B(n237), .Z(n141) );
  AND U191 ( .A(n140), .B(n141), .Z(n241) );
  XOR U192 ( .A(sreg[83]), .B(n246), .Z(n142) );
  NANDN U193 ( .A(n247), .B(n142), .Z(n143) );
  NAND U194 ( .A(sreg[83]), .B(n246), .Z(n144) );
  AND U195 ( .A(n143), .B(n144), .Z(n250) );
  XOR U196 ( .A(sreg[86]), .B(n255), .Z(n145) );
  NANDN U197 ( .A(n256), .B(n145), .Z(n146) );
  NAND U198 ( .A(sreg[86]), .B(n255), .Z(n147) );
  AND U199 ( .A(n146), .B(n147), .Z(n259) );
  XOR U200 ( .A(sreg[89]), .B(n264), .Z(n148) );
  NANDN U201 ( .A(n265), .B(n148), .Z(n149) );
  NAND U202 ( .A(sreg[89]), .B(n264), .Z(n150) );
  AND U203 ( .A(n149), .B(n150), .Z(n268) );
  XOR U204 ( .A(sreg[92]), .B(n273), .Z(n151) );
  NANDN U205 ( .A(n274), .B(n151), .Z(n152) );
  NAND U206 ( .A(sreg[92]), .B(n273), .Z(n153) );
  AND U207 ( .A(n152), .B(n153), .Z(n277) );
  XOR U208 ( .A(sreg[95]), .B(n282), .Z(n154) );
  NANDN U209 ( .A(n283), .B(n154), .Z(n155) );
  NAND U210 ( .A(sreg[95]), .B(n282), .Z(n156) );
  AND U211 ( .A(n155), .B(n156), .Z(n286) );
  XOR U212 ( .A(sreg[98]), .B(n291), .Z(n157) );
  NANDN U213 ( .A(n292), .B(n157), .Z(n158) );
  NAND U214 ( .A(sreg[98]), .B(n291), .Z(n159) );
  AND U215 ( .A(n158), .B(n159), .Z(n295) );
  XOR U216 ( .A(sreg[101]), .B(n300), .Z(n160) );
  NANDN U217 ( .A(n301), .B(n160), .Z(n161) );
  NAND U218 ( .A(sreg[101]), .B(n300), .Z(n162) );
  AND U219 ( .A(n161), .B(n162), .Z(n304) );
  XOR U220 ( .A(sreg[104]), .B(n309), .Z(n163) );
  NANDN U221 ( .A(n310), .B(n163), .Z(n164) );
  NAND U222 ( .A(sreg[104]), .B(n309), .Z(n165) );
  AND U223 ( .A(n164), .B(n165), .Z(n313) );
  XOR U224 ( .A(sreg[107]), .B(n318), .Z(n166) );
  NANDN U225 ( .A(n319), .B(n166), .Z(n167) );
  NAND U226 ( .A(sreg[107]), .B(n318), .Z(n168) );
  AND U227 ( .A(n167), .B(n168), .Z(n322) );
  XOR U228 ( .A(sreg[110]), .B(n327), .Z(n169) );
  NANDN U229 ( .A(n328), .B(n169), .Z(n170) );
  NAND U230 ( .A(sreg[110]), .B(n327), .Z(n171) );
  AND U231 ( .A(n170), .B(n171), .Z(n331) );
  XOR U232 ( .A(sreg[113]), .B(n336), .Z(n172) );
  NANDN U233 ( .A(n337), .B(n172), .Z(n173) );
  NAND U234 ( .A(sreg[113]), .B(n336), .Z(n174) );
  AND U235 ( .A(n173), .B(n174), .Z(n340) );
  XOR U236 ( .A(sreg[116]), .B(n345), .Z(n175) );
  NANDN U237 ( .A(n346), .B(n175), .Z(n176) );
  NAND U238 ( .A(sreg[116]), .B(n345), .Z(n177) );
  AND U239 ( .A(n176), .B(n177), .Z(n349) );
  XOR U240 ( .A(sreg[119]), .B(n354), .Z(n178) );
  NANDN U241 ( .A(n355), .B(n178), .Z(n179) );
  NAND U242 ( .A(sreg[119]), .B(n354), .Z(n180) );
  AND U243 ( .A(n179), .B(n180), .Z(n358) );
  XOR U244 ( .A(sreg[122]), .B(n363), .Z(n181) );
  NANDN U245 ( .A(n364), .B(n181), .Z(n182) );
  NAND U246 ( .A(sreg[122]), .B(n363), .Z(n183) );
  AND U247 ( .A(n182), .B(n183), .Z(n367) );
  XOR U248 ( .A(sreg[125]), .B(n372), .Z(n184) );
  NANDN U249 ( .A(n373), .B(n184), .Z(n185) );
  NAND U250 ( .A(sreg[125]), .B(n372), .Z(n186) );
  AND U251 ( .A(n185), .B(n186), .Z(n376) );
  AND U252 ( .A(b[0]), .B(a[0]), .Z(n187) );
  XOR U253 ( .A(n187), .B(sreg[63]), .Z(c[63]) );
  NAND U254 ( .A(b[0]), .B(a[1]), .Z(n190) );
  AND U255 ( .A(n187), .B(sreg[63]), .Z(n189) );
  XOR U256 ( .A(sreg[64]), .B(n189), .Z(n188) );
  XNOR U257 ( .A(n190), .B(n188), .Z(c[64]) );
  AND U258 ( .A(b[0]), .B(a[2]), .Z(n192) );
  XNOR U259 ( .A(n193), .B(sreg[65]), .Z(n191) );
  XOR U260 ( .A(n192), .B(n191), .Z(c[65]) );
  AND U261 ( .A(b[0]), .B(a[3]), .Z(n195) );
  XNOR U262 ( .A(n196), .B(sreg[66]), .Z(n194) );
  XOR U263 ( .A(n195), .B(n194), .Z(c[66]) );
  AND U264 ( .A(b[0]), .B(a[4]), .Z(n198) );
  XNOR U265 ( .A(n199), .B(sreg[67]), .Z(n197) );
  XOR U266 ( .A(n198), .B(n197), .Z(c[67]) );
  AND U267 ( .A(b[0]), .B(a[5]), .Z(n201) );
  XNOR U268 ( .A(n202), .B(sreg[68]), .Z(n200) );
  XOR U269 ( .A(n201), .B(n200), .Z(c[68]) );
  AND U270 ( .A(b[0]), .B(a[6]), .Z(n204) );
  XNOR U271 ( .A(n205), .B(sreg[69]), .Z(n203) );
  XOR U272 ( .A(n204), .B(n203), .Z(c[69]) );
  AND U273 ( .A(b[0]), .B(a[7]), .Z(n207) );
  XNOR U274 ( .A(n208), .B(sreg[70]), .Z(n206) );
  XOR U275 ( .A(n207), .B(n206), .Z(c[70]) );
  AND U276 ( .A(b[0]), .B(a[8]), .Z(n210) );
  XNOR U277 ( .A(n211), .B(sreg[71]), .Z(n209) );
  XOR U278 ( .A(n210), .B(n209), .Z(c[71]) );
  AND U279 ( .A(b[0]), .B(a[9]), .Z(n213) );
  XNOR U280 ( .A(n214), .B(sreg[72]), .Z(n212) );
  XOR U281 ( .A(n213), .B(n212), .Z(c[72]) );
  AND U282 ( .A(b[0]), .B(a[10]), .Z(n216) );
  XNOR U283 ( .A(n217), .B(sreg[73]), .Z(n215) );
  XOR U284 ( .A(n216), .B(n215), .Z(c[73]) );
  AND U285 ( .A(b[0]), .B(a[11]), .Z(n219) );
  XNOR U286 ( .A(n220), .B(sreg[74]), .Z(n218) );
  XOR U287 ( .A(n219), .B(n218), .Z(c[74]) );
  AND U288 ( .A(b[0]), .B(a[12]), .Z(n222) );
  XNOR U289 ( .A(n223), .B(sreg[75]), .Z(n221) );
  XOR U290 ( .A(n222), .B(n221), .Z(c[75]) );
  AND U291 ( .A(b[0]), .B(a[13]), .Z(n225) );
  XNOR U292 ( .A(n226), .B(sreg[76]), .Z(n224) );
  XOR U293 ( .A(n225), .B(n224), .Z(c[76]) );
  AND U294 ( .A(b[0]), .B(a[14]), .Z(n228) );
  XNOR U295 ( .A(n229), .B(sreg[77]), .Z(n227) );
  XOR U296 ( .A(n228), .B(n227), .Z(c[77]) );
  AND U297 ( .A(b[0]), .B(a[15]), .Z(n231) );
  XNOR U298 ( .A(n232), .B(sreg[78]), .Z(n230) );
  XOR U299 ( .A(n231), .B(n230), .Z(c[78]) );
  AND U300 ( .A(b[0]), .B(a[16]), .Z(n234) );
  XNOR U301 ( .A(n235), .B(sreg[79]), .Z(n233) );
  XOR U302 ( .A(n234), .B(n233), .Z(c[79]) );
  AND U303 ( .A(b[0]), .B(a[17]), .Z(n237) );
  XNOR U304 ( .A(n238), .B(sreg[80]), .Z(n236) );
  XOR U305 ( .A(n237), .B(n236), .Z(c[80]) );
  AND U306 ( .A(b[0]), .B(a[18]), .Z(n240) );
  XNOR U307 ( .A(n241), .B(sreg[81]), .Z(n239) );
  XOR U308 ( .A(n240), .B(n239), .Z(c[81]) );
  AND U309 ( .A(b[0]), .B(a[19]), .Z(n243) );
  XNOR U310 ( .A(n244), .B(sreg[82]), .Z(n242) );
  XOR U311 ( .A(n243), .B(n242), .Z(c[82]) );
  AND U312 ( .A(b[0]), .B(a[20]), .Z(n246) );
  XNOR U313 ( .A(n247), .B(sreg[83]), .Z(n245) );
  XOR U314 ( .A(n246), .B(n245), .Z(c[83]) );
  AND U315 ( .A(b[0]), .B(a[21]), .Z(n249) );
  XNOR U316 ( .A(n250), .B(sreg[84]), .Z(n248) );
  XOR U317 ( .A(n249), .B(n248), .Z(c[84]) );
  AND U318 ( .A(b[0]), .B(a[22]), .Z(n252) );
  XNOR U319 ( .A(n253), .B(sreg[85]), .Z(n251) );
  XOR U320 ( .A(n252), .B(n251), .Z(c[85]) );
  AND U321 ( .A(b[0]), .B(a[23]), .Z(n255) );
  XNOR U322 ( .A(n256), .B(sreg[86]), .Z(n254) );
  XOR U323 ( .A(n255), .B(n254), .Z(c[86]) );
  AND U324 ( .A(b[0]), .B(a[24]), .Z(n258) );
  XNOR U325 ( .A(n259), .B(sreg[87]), .Z(n257) );
  XOR U326 ( .A(n258), .B(n257), .Z(c[87]) );
  AND U327 ( .A(b[0]), .B(a[25]), .Z(n261) );
  XNOR U328 ( .A(n262), .B(sreg[88]), .Z(n260) );
  XOR U329 ( .A(n261), .B(n260), .Z(c[88]) );
  AND U330 ( .A(b[0]), .B(a[26]), .Z(n264) );
  XNOR U331 ( .A(n265), .B(sreg[89]), .Z(n263) );
  XOR U332 ( .A(n264), .B(n263), .Z(c[89]) );
  AND U333 ( .A(b[0]), .B(a[27]), .Z(n267) );
  XNOR U334 ( .A(n268), .B(sreg[90]), .Z(n266) );
  XOR U335 ( .A(n267), .B(n266), .Z(c[90]) );
  AND U336 ( .A(b[0]), .B(a[28]), .Z(n270) );
  XNOR U337 ( .A(n271), .B(sreg[91]), .Z(n269) );
  XOR U338 ( .A(n270), .B(n269), .Z(c[91]) );
  AND U339 ( .A(b[0]), .B(a[29]), .Z(n273) );
  XNOR U340 ( .A(n274), .B(sreg[92]), .Z(n272) );
  XOR U341 ( .A(n273), .B(n272), .Z(c[92]) );
  AND U342 ( .A(b[0]), .B(a[30]), .Z(n276) );
  XNOR U343 ( .A(n277), .B(sreg[93]), .Z(n275) );
  XOR U344 ( .A(n276), .B(n275), .Z(c[93]) );
  AND U345 ( .A(b[0]), .B(a[31]), .Z(n279) );
  XNOR U346 ( .A(n280), .B(sreg[94]), .Z(n278) );
  XOR U347 ( .A(n279), .B(n278), .Z(c[94]) );
  AND U348 ( .A(b[0]), .B(a[32]), .Z(n282) );
  XNOR U349 ( .A(n283), .B(sreg[95]), .Z(n281) );
  XOR U350 ( .A(n282), .B(n281), .Z(c[95]) );
  AND U351 ( .A(b[0]), .B(a[33]), .Z(n285) );
  XNOR U352 ( .A(n286), .B(sreg[96]), .Z(n284) );
  XOR U353 ( .A(n285), .B(n284), .Z(c[96]) );
  AND U354 ( .A(b[0]), .B(a[34]), .Z(n288) );
  XNOR U355 ( .A(n289), .B(sreg[97]), .Z(n287) );
  XOR U356 ( .A(n288), .B(n287), .Z(c[97]) );
  AND U357 ( .A(b[0]), .B(a[35]), .Z(n291) );
  XNOR U358 ( .A(n292), .B(sreg[98]), .Z(n290) );
  XOR U359 ( .A(n291), .B(n290), .Z(c[98]) );
  AND U360 ( .A(b[0]), .B(a[36]), .Z(n294) );
  XNOR U361 ( .A(n295), .B(sreg[99]), .Z(n293) );
  XOR U362 ( .A(n294), .B(n293), .Z(c[99]) );
  AND U363 ( .A(b[0]), .B(a[37]), .Z(n297) );
  XNOR U364 ( .A(n298), .B(sreg[100]), .Z(n296) );
  XOR U365 ( .A(n297), .B(n296), .Z(c[100]) );
  AND U366 ( .A(b[0]), .B(a[38]), .Z(n300) );
  XNOR U367 ( .A(n301), .B(sreg[101]), .Z(n299) );
  XOR U368 ( .A(n300), .B(n299), .Z(c[101]) );
  AND U369 ( .A(b[0]), .B(a[39]), .Z(n303) );
  XNOR U370 ( .A(n304), .B(sreg[102]), .Z(n302) );
  XOR U371 ( .A(n303), .B(n302), .Z(c[102]) );
  AND U372 ( .A(b[0]), .B(a[40]), .Z(n306) );
  XNOR U373 ( .A(n307), .B(sreg[103]), .Z(n305) );
  XOR U374 ( .A(n306), .B(n305), .Z(c[103]) );
  AND U375 ( .A(b[0]), .B(a[41]), .Z(n309) );
  XNOR U376 ( .A(n310), .B(sreg[104]), .Z(n308) );
  XOR U377 ( .A(n309), .B(n308), .Z(c[104]) );
  AND U378 ( .A(b[0]), .B(a[42]), .Z(n312) );
  XNOR U379 ( .A(n313), .B(sreg[105]), .Z(n311) );
  XOR U380 ( .A(n312), .B(n311), .Z(c[105]) );
  AND U381 ( .A(b[0]), .B(a[43]), .Z(n315) );
  XNOR U382 ( .A(n316), .B(sreg[106]), .Z(n314) );
  XOR U383 ( .A(n315), .B(n314), .Z(c[106]) );
  AND U384 ( .A(b[0]), .B(a[44]), .Z(n318) );
  XNOR U385 ( .A(n319), .B(sreg[107]), .Z(n317) );
  XOR U386 ( .A(n318), .B(n317), .Z(c[107]) );
  AND U387 ( .A(b[0]), .B(a[45]), .Z(n321) );
  XNOR U388 ( .A(n322), .B(sreg[108]), .Z(n320) );
  XOR U389 ( .A(n321), .B(n320), .Z(c[108]) );
  AND U390 ( .A(b[0]), .B(a[46]), .Z(n324) );
  XNOR U391 ( .A(n325), .B(sreg[109]), .Z(n323) );
  XOR U392 ( .A(n324), .B(n323), .Z(c[109]) );
  AND U393 ( .A(b[0]), .B(a[47]), .Z(n327) );
  XNOR U394 ( .A(n328), .B(sreg[110]), .Z(n326) );
  XOR U395 ( .A(n327), .B(n326), .Z(c[110]) );
  AND U396 ( .A(b[0]), .B(a[48]), .Z(n330) );
  XNOR U397 ( .A(n331), .B(sreg[111]), .Z(n329) );
  XOR U398 ( .A(n330), .B(n329), .Z(c[111]) );
  AND U399 ( .A(b[0]), .B(a[49]), .Z(n333) );
  XNOR U400 ( .A(n334), .B(sreg[112]), .Z(n332) );
  XOR U401 ( .A(n333), .B(n332), .Z(c[112]) );
  AND U402 ( .A(b[0]), .B(a[50]), .Z(n336) );
  XNOR U403 ( .A(n337), .B(sreg[113]), .Z(n335) );
  XOR U404 ( .A(n336), .B(n335), .Z(c[113]) );
  AND U405 ( .A(b[0]), .B(a[51]), .Z(n339) );
  XNOR U406 ( .A(n340), .B(sreg[114]), .Z(n338) );
  XOR U407 ( .A(n339), .B(n338), .Z(c[114]) );
  AND U408 ( .A(b[0]), .B(a[52]), .Z(n342) );
  XNOR U409 ( .A(n343), .B(sreg[115]), .Z(n341) );
  XOR U410 ( .A(n342), .B(n341), .Z(c[115]) );
  AND U411 ( .A(b[0]), .B(a[53]), .Z(n345) );
  XNOR U412 ( .A(n346), .B(sreg[116]), .Z(n344) );
  XOR U413 ( .A(n345), .B(n344), .Z(c[116]) );
  AND U414 ( .A(b[0]), .B(a[54]), .Z(n348) );
  XNOR U415 ( .A(n349), .B(sreg[117]), .Z(n347) );
  XOR U416 ( .A(n348), .B(n347), .Z(c[117]) );
  AND U417 ( .A(b[0]), .B(a[55]), .Z(n351) );
  XNOR U418 ( .A(n352), .B(sreg[118]), .Z(n350) );
  XOR U419 ( .A(n351), .B(n350), .Z(c[118]) );
  AND U420 ( .A(b[0]), .B(a[56]), .Z(n354) );
  XNOR U421 ( .A(n355), .B(sreg[119]), .Z(n353) );
  XOR U422 ( .A(n354), .B(n353), .Z(c[119]) );
  AND U423 ( .A(b[0]), .B(a[57]), .Z(n357) );
  XNOR U424 ( .A(n358), .B(sreg[120]), .Z(n356) );
  XOR U425 ( .A(n357), .B(n356), .Z(c[120]) );
  AND U426 ( .A(b[0]), .B(a[58]), .Z(n360) );
  XNOR U427 ( .A(n361), .B(sreg[121]), .Z(n359) );
  XOR U428 ( .A(n360), .B(n359), .Z(c[121]) );
  AND U429 ( .A(b[0]), .B(a[59]), .Z(n363) );
  XNOR U430 ( .A(n364), .B(sreg[122]), .Z(n362) );
  XOR U431 ( .A(n363), .B(n362), .Z(c[122]) );
  AND U432 ( .A(b[0]), .B(a[60]), .Z(n366) );
  XNOR U433 ( .A(n367), .B(sreg[123]), .Z(n365) );
  XOR U434 ( .A(n366), .B(n365), .Z(c[123]) );
  AND U435 ( .A(b[0]), .B(a[61]), .Z(n369) );
  XNOR U436 ( .A(n370), .B(sreg[124]), .Z(n368) );
  XOR U437 ( .A(n369), .B(n368), .Z(c[124]) );
  AND U438 ( .A(b[0]), .B(a[62]), .Z(n372) );
  XNOR U439 ( .A(n373), .B(sreg[125]), .Z(n371) );
  XOR U440 ( .A(n372), .B(n371), .Z(c[125]) );
  NAND U441 ( .A(b[0]), .B(a[63]), .Z(n374) );
  XNOR U442 ( .A(sreg[126]), .B(n376), .Z(n375) );
  XNOR U443 ( .A(n374), .B(n375), .Z(c[126]) );
  NAND U444 ( .A(n375), .B(n374), .Z(n378) );
  NANDN U445 ( .A(sreg[126]), .B(n376), .Z(n377) );
  AND U446 ( .A(n378), .B(n377), .Z(c[127]) );
endmodule

