
module mult_N64_CC4 ( clk, rst, a, b, c );
  input [63:0] a;
  input [15:0] b;
  output [63:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702;
  wire   [63:16] swire;
  wire   [127:64] sreg;

  DFF \sreg_reg[64]  ( .D(swire[16]), .CLK(clk), .RST(rst), .Q(sreg[64]) );
  DFF \sreg_reg[65]  ( .D(swire[17]), .CLK(clk), .RST(rst), .Q(sreg[65]) );
  DFF \sreg_reg[66]  ( .D(swire[18]), .CLK(clk), .RST(rst), .Q(sreg[66]) );
  DFF \sreg_reg[67]  ( .D(swire[19]), .CLK(clk), .RST(rst), .Q(sreg[67]) );
  DFF \sreg_reg[68]  ( .D(swire[20]), .CLK(clk), .RST(rst), .Q(sreg[68]) );
  DFF \sreg_reg[69]  ( .D(swire[21]), .CLK(clk), .RST(rst), .Q(sreg[69]) );
  DFF \sreg_reg[70]  ( .D(swire[22]), .CLK(clk), .RST(rst), .Q(sreg[70]) );
  DFF \sreg_reg[71]  ( .D(swire[23]), .CLK(clk), .RST(rst), .Q(sreg[71]) );
  DFF \sreg_reg[72]  ( .D(swire[24]), .CLK(clk), .RST(rst), .Q(sreg[72]) );
  DFF \sreg_reg[73]  ( .D(swire[25]), .CLK(clk), .RST(rst), .Q(sreg[73]) );
  DFF \sreg_reg[74]  ( .D(swire[26]), .CLK(clk), .RST(rst), .Q(sreg[74]) );
  DFF \sreg_reg[75]  ( .D(swire[27]), .CLK(clk), .RST(rst), .Q(sreg[75]) );
  DFF \sreg_reg[76]  ( .D(swire[28]), .CLK(clk), .RST(rst), .Q(sreg[76]) );
  DFF \sreg_reg[77]  ( .D(swire[29]), .CLK(clk), .RST(rst), .Q(sreg[77]) );
  DFF \sreg_reg[78]  ( .D(swire[30]), .CLK(clk), .RST(rst), .Q(sreg[78]) );
  DFF \sreg_reg[79]  ( .D(swire[31]), .CLK(clk), .RST(rst), .Q(sreg[79]) );
  DFF \sreg_reg[80]  ( .D(swire[32]), .CLK(clk), .RST(rst), .Q(sreg[80]) );
  DFF \sreg_reg[81]  ( .D(swire[33]), .CLK(clk), .RST(rst), .Q(sreg[81]) );
  DFF \sreg_reg[82]  ( .D(swire[34]), .CLK(clk), .RST(rst), .Q(sreg[82]) );
  DFF \sreg_reg[83]  ( .D(swire[35]), .CLK(clk), .RST(rst), .Q(sreg[83]) );
  DFF \sreg_reg[84]  ( .D(swire[36]), .CLK(clk), .RST(rst), .Q(sreg[84]) );
  DFF \sreg_reg[85]  ( .D(swire[37]), .CLK(clk), .RST(rst), .Q(sreg[85]) );
  DFF \sreg_reg[86]  ( .D(swire[38]), .CLK(clk), .RST(rst), .Q(sreg[86]) );
  DFF \sreg_reg[87]  ( .D(swire[39]), .CLK(clk), .RST(rst), .Q(sreg[87]) );
  DFF \sreg_reg[88]  ( .D(swire[40]), .CLK(clk), .RST(rst), .Q(sreg[88]) );
  DFF \sreg_reg[89]  ( .D(swire[41]), .CLK(clk), .RST(rst), .Q(sreg[89]) );
  DFF \sreg_reg[90]  ( .D(swire[42]), .CLK(clk), .RST(rst), .Q(sreg[90]) );
  DFF \sreg_reg[91]  ( .D(swire[43]), .CLK(clk), .RST(rst), .Q(sreg[91]) );
  DFF \sreg_reg[92]  ( .D(swire[44]), .CLK(clk), .RST(rst), .Q(sreg[92]) );
  DFF \sreg_reg[93]  ( .D(swire[45]), .CLK(clk), .RST(rst), .Q(sreg[93]) );
  DFF \sreg_reg[94]  ( .D(swire[46]), .CLK(clk), .RST(rst), .Q(sreg[94]) );
  DFF \sreg_reg[95]  ( .D(swire[47]), .CLK(clk), .RST(rst), .Q(sreg[95]) );
  DFF \sreg_reg[96]  ( .D(swire[48]), .CLK(clk), .RST(rst), .Q(sreg[96]) );
  DFF \sreg_reg[97]  ( .D(swire[49]), .CLK(clk), .RST(rst), .Q(sreg[97]) );
  DFF \sreg_reg[98]  ( .D(swire[50]), .CLK(clk), .RST(rst), .Q(sreg[98]) );
  DFF \sreg_reg[99]  ( .D(swire[51]), .CLK(clk), .RST(rst), .Q(sreg[99]) );
  DFF \sreg_reg[100]  ( .D(swire[52]), .CLK(clk), .RST(rst), .Q(sreg[100]) );
  DFF \sreg_reg[101]  ( .D(swire[53]), .CLK(clk), .RST(rst), .Q(sreg[101]) );
  DFF \sreg_reg[102]  ( .D(swire[54]), .CLK(clk), .RST(rst), .Q(sreg[102]) );
  DFF \sreg_reg[103]  ( .D(swire[55]), .CLK(clk), .RST(rst), .Q(sreg[103]) );
  DFF \sreg_reg[104]  ( .D(swire[56]), .CLK(clk), .RST(rst), .Q(sreg[104]) );
  DFF \sreg_reg[105]  ( .D(swire[57]), .CLK(clk), .RST(rst), .Q(sreg[105]) );
  DFF \sreg_reg[106]  ( .D(swire[58]), .CLK(clk), .RST(rst), .Q(sreg[106]) );
  DFF \sreg_reg[107]  ( .D(swire[59]), .CLK(clk), .RST(rst), .Q(sreg[107]) );
  DFF \sreg_reg[108]  ( .D(swire[60]), .CLK(clk), .RST(rst), .Q(sreg[108]) );
  DFF \sreg_reg[109]  ( .D(swire[61]), .CLK(clk), .RST(rst), .Q(sreg[109]) );
  DFF \sreg_reg[110]  ( .D(swire[62]), .CLK(clk), .RST(rst), .Q(sreg[110]) );
  DFF \sreg_reg[111]  ( .D(swire[63]), .CLK(clk), .RST(rst), .Q(sreg[111]) );
  DFF \sreg_reg[63]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[62]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[61]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[60]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[59]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[58]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[57]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[56]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[55]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[54]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[53]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[52]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[51]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[50]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[49]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[48]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[47]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[46]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[45]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[44]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[43]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[42]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[41]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[40]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[39]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[38]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[37]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[36]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[35]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[34]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[33]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[32]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[31]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[30]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[29]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[28]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[27]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[26]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[25]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[24]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[23]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[22]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[21]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[20]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[19]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[18]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[17]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[16]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[0]) );
  XOR U19 ( .A(n381), .B(n441), .Z(n385) );
  XOR U20 ( .A(n309), .B(n358), .Z(n313) );
  XOR U21 ( .A(n239), .B(n275), .Z(n243) );
  XOR U22 ( .A(n4146), .B(n4215), .Z(n4151) );
  XOR U23 ( .A(n3977), .B(n4045), .Z(n3981) );
  XOR U24 ( .A(n544), .B(n611), .Z(n548) );
  XOR U25 ( .A(n714), .B(n780), .Z(n718) );
  XOR U26 ( .A(n883), .B(n949), .Z(n887) );
  XOR U27 ( .A(n1052), .B(n1118), .Z(n1056) );
  XOR U28 ( .A(n1221), .B(n1293), .Z(n1225) );
  XOR U29 ( .A(n1397), .B(n1465), .Z(n1401) );
  XOR U30 ( .A(n1569), .B(n1637), .Z(n1573) );
  XOR U31 ( .A(n1741), .B(n1809), .Z(n1745) );
  XOR U32 ( .A(n1913), .B(n1981), .Z(n1917) );
  XOR U33 ( .A(n2085), .B(n2153), .Z(n2089) );
  XOR U34 ( .A(n2257), .B(n2325), .Z(n2261) );
  XOR U35 ( .A(n2429), .B(n2497), .Z(n2433) );
  XOR U36 ( .A(n2601), .B(n2669), .Z(n2605) );
  XOR U37 ( .A(n2773), .B(n2841), .Z(n2777) );
  XOR U38 ( .A(n2945), .B(n3013), .Z(n2949) );
  XOR U39 ( .A(n3117), .B(n3185), .Z(n3121) );
  XOR U40 ( .A(n3289), .B(n3357), .Z(n3293) );
  XOR U41 ( .A(n3461), .B(n3529), .Z(n3465) );
  XOR U42 ( .A(n3633), .B(n3701), .Z(n3637) );
  XOR U43 ( .A(n3805), .B(n3873), .Z(n3809) );
  XOR U44 ( .A(n4306), .B(n4356), .Z(n4310) );
  XOR U45 ( .A(n4162), .B(n4212), .Z(n4166) );
  XOR U46 ( .A(n3992), .B(n4042), .Z(n3996) );
  XOR U47 ( .A(n224), .B(n278), .Z(n228) );
  XOR U48 ( .A(n559), .B(n608), .Z(n563) );
  XOR U49 ( .A(n729), .B(n777), .Z(n733) );
  XOR U50 ( .A(n898), .B(n946), .Z(n902) );
  XOR U51 ( .A(n1067), .B(n1115), .Z(n1071) );
  XOR U52 ( .A(n1236), .B(n1290), .Z(n1240) );
  XOR U53 ( .A(n1412), .B(n1462), .Z(n1416) );
  XOR U54 ( .A(n1584), .B(n1634), .Z(n1588) );
  XOR U55 ( .A(n1756), .B(n1806), .Z(n1760) );
  XOR U56 ( .A(n1928), .B(n1978), .Z(n1932) );
  XOR U57 ( .A(n2100), .B(n2150), .Z(n2104) );
  XOR U58 ( .A(n2272), .B(n2322), .Z(n2276) );
  XOR U59 ( .A(n2444), .B(n2494), .Z(n2448) );
  XOR U60 ( .A(n2616), .B(n2666), .Z(n2620) );
  XOR U61 ( .A(n2788), .B(n2838), .Z(n2792) );
  XOR U62 ( .A(n2960), .B(n3010), .Z(n2964) );
  XOR U63 ( .A(n3132), .B(n3182), .Z(n3136) );
  XOR U64 ( .A(n3304), .B(n3354), .Z(n3308) );
  XOR U65 ( .A(n3476), .B(n3526), .Z(n3480) );
  XOR U66 ( .A(n3648), .B(n3698), .Z(n3652) );
  XOR U67 ( .A(n3820), .B(n3870), .Z(n3824) );
  XOR U68 ( .A(n401), .B(n437), .Z(n405) );
  XOR U69 ( .A(n4536), .B(n4569), .Z(n4541) );
  XOR U70 ( .A(n4441), .B(n4473), .Z(n4445) );
  XOR U71 ( .A(n4321), .B(n4353), .Z(n4325) );
  XOR U72 ( .A(n4177), .B(n4209), .Z(n4181) );
  XOR U73 ( .A(n4007), .B(n4039), .Z(n4011) );
  XOR U74 ( .A(n244), .B(n274), .Z(n248) );
  XOR U75 ( .A(n574), .B(n605), .Z(n578) );
  XOR U76 ( .A(n744), .B(n774), .Z(n748) );
  XOR U77 ( .A(n913), .B(n943), .Z(n917) );
  XOR U78 ( .A(n1082), .B(n1112), .Z(n1086) );
  XOR U79 ( .A(n1251), .B(n1287), .Z(n1255) );
  XOR U80 ( .A(n1427), .B(n1459), .Z(n1431) );
  XOR U81 ( .A(n1599), .B(n1631), .Z(n1603) );
  XOR U82 ( .A(n1771), .B(n1803), .Z(n1775) );
  XOR U83 ( .A(n1943), .B(n1975), .Z(n1947) );
  XOR U84 ( .A(n2115), .B(n2147), .Z(n2119) );
  XOR U85 ( .A(n2287), .B(n2319), .Z(n2291) );
  XOR U86 ( .A(n2459), .B(n2491), .Z(n2463) );
  XOR U87 ( .A(n2631), .B(n2663), .Z(n2635) );
  XOR U88 ( .A(n2803), .B(n2835), .Z(n2807) );
  XOR U89 ( .A(n2975), .B(n3007), .Z(n2979) );
  XOR U90 ( .A(n3147), .B(n3179), .Z(n3151) );
  XOR U91 ( .A(n3319), .B(n3351), .Z(n3323) );
  XOR U92 ( .A(n3491), .B(n3523), .Z(n3495) );
  XOR U93 ( .A(n3663), .B(n3695), .Z(n3667) );
  XOR U94 ( .A(n3835), .B(n3867), .Z(n3839) );
  XOR U95 ( .A(n4063), .B(n4131), .Z(n4067) );
  XOR U96 ( .A(n293), .B(n362), .Z(n298) );
  XOR U97 ( .A(n455), .B(n523), .Z(n460) );
  XOR U98 ( .A(n629), .B(n696), .Z(n633) );
  XOR U99 ( .A(n798), .B(n865), .Z(n802) );
  XOR U100 ( .A(n967), .B(n1034), .Z(n971) );
  XOR U101 ( .A(n1136), .B(n1203), .Z(n1140) );
  XOR U102 ( .A(n1311), .B(n1379), .Z(n1315) );
  XOR U103 ( .A(n1483), .B(n1551), .Z(n1487) );
  XOR U104 ( .A(n1655), .B(n1723), .Z(n1659) );
  XOR U105 ( .A(n1827), .B(n1895), .Z(n1831) );
  XOR U106 ( .A(n1999), .B(n2067), .Z(n2003) );
  XOR U107 ( .A(n2171), .B(n2239), .Z(n2175) );
  XOR U108 ( .A(n2343), .B(n2411), .Z(n2347) );
  XOR U109 ( .A(n2515), .B(n2583), .Z(n2519) );
  XOR U110 ( .A(n2687), .B(n2755), .Z(n2691) );
  XOR U111 ( .A(n2859), .B(n2927), .Z(n2863) );
  XOR U112 ( .A(n3031), .B(n3099), .Z(n3035) );
  XOR U113 ( .A(n3203), .B(n3271), .Z(n3207) );
  XOR U114 ( .A(n3375), .B(n3443), .Z(n3379) );
  XOR U115 ( .A(n3547), .B(n3615), .Z(n3551) );
  XOR U116 ( .A(n3719), .B(n3787), .Z(n3723) );
  XOR U117 ( .A(n3891), .B(n3959), .Z(n3895) );
  XOR U118 ( .A(n4368), .B(n4419), .Z(n4373) );
  XOR U119 ( .A(n4237), .B(n4287), .Z(n4241) );
  XOR U120 ( .A(n4078), .B(n4128), .Z(n4082) );
  XOR U121 ( .A(n471), .B(n520), .Z(n475) );
  XOR U122 ( .A(n644), .B(n693), .Z(n648) );
  XOR U123 ( .A(n813), .B(n862), .Z(n817) );
  XOR U124 ( .A(n982), .B(n1031), .Z(n986) );
  XOR U125 ( .A(n1151), .B(n1200), .Z(n1155) );
  XOR U126 ( .A(n1326), .B(n1376), .Z(n1330) );
  XOR U127 ( .A(n1498), .B(n1548), .Z(n1502) );
  XOR U128 ( .A(n1670), .B(n1720), .Z(n1674) );
  XOR U129 ( .A(n1842), .B(n1892), .Z(n1846) );
  XOR U130 ( .A(n2014), .B(n2064), .Z(n2018) );
  XOR U131 ( .A(n2186), .B(n2236), .Z(n2190) );
  XOR U132 ( .A(n2358), .B(n2408), .Z(n2362) );
  XOR U133 ( .A(n2530), .B(n2580), .Z(n2534) );
  XOR U134 ( .A(n2702), .B(n2752), .Z(n2706) );
  XOR U135 ( .A(n2874), .B(n2924), .Z(n2878) );
  XOR U136 ( .A(n3046), .B(n3096), .Z(n3050) );
  XOR U137 ( .A(n3218), .B(n3268), .Z(n3222) );
  XOR U138 ( .A(n3390), .B(n3440), .Z(n3394) );
  XOR U139 ( .A(n3562), .B(n3612), .Z(n3566) );
  XOR U140 ( .A(n3734), .B(n3784), .Z(n3738) );
  XOR U141 ( .A(n3906), .B(n3956), .Z(n3910) );
  XOR U142 ( .A(n396), .B(n438), .Z(n400) );
  XOR U143 ( .A(n4492), .B(n4524), .Z(n4496) );
  XOR U144 ( .A(n4384), .B(n4416), .Z(n4388) );
  XOR U145 ( .A(n4252), .B(n4284), .Z(n4256) );
  XOR U146 ( .A(n4093), .B(n4125), .Z(n4097) );
  XOR U147 ( .A(n164), .B(n194), .Z(n168) );
  XOR U148 ( .A(n324), .B(n355), .Z(n328) );
  XOR U149 ( .A(n659), .B(n690), .Z(n663) );
  XOR U150 ( .A(n828), .B(n859), .Z(n832) );
  XOR U151 ( .A(n997), .B(n1028), .Z(n1001) );
  XOR U152 ( .A(n1166), .B(n1197), .Z(n1170) );
  XOR U153 ( .A(n1341), .B(n1373), .Z(n1345) );
  XOR U154 ( .A(n1513), .B(n1545), .Z(n1517) );
  XOR U155 ( .A(n1685), .B(n1717), .Z(n1689) );
  XOR U156 ( .A(n1857), .B(n1889), .Z(n1861) );
  XOR U157 ( .A(n2029), .B(n2061), .Z(n2033) );
  XOR U158 ( .A(n2201), .B(n2233), .Z(n2205) );
  XOR U159 ( .A(n2373), .B(n2405), .Z(n2377) );
  XOR U160 ( .A(n2545), .B(n2577), .Z(n2549) );
  XOR U161 ( .A(n2717), .B(n2749), .Z(n2721) );
  XOR U162 ( .A(n2889), .B(n2921), .Z(n2893) );
  XOR U163 ( .A(n3061), .B(n3093), .Z(n3065) );
  XOR U164 ( .A(n3233), .B(n3265), .Z(n3237) );
  XOR U165 ( .A(n3405), .B(n3437), .Z(n3409) );
  XOR U166 ( .A(n3577), .B(n3609), .Z(n3581) );
  XOR U167 ( .A(n3749), .B(n3781), .Z(n3753) );
  XOR U168 ( .A(n3921), .B(n3953), .Z(n3925) );
  XOR U169 ( .A(n491), .B(n516), .Z(n495) );
  XOR U170 ( .A(n375), .B(n442), .Z(n380) );
  XOR U171 ( .A(n4152), .B(n4214), .Z(n4156) );
  XOR U172 ( .A(n3982), .B(n4044), .Z(n3986) );
  XOR U173 ( .A(n549), .B(n610), .Z(n553) );
  XOR U174 ( .A(n719), .B(n779), .Z(n723) );
  XOR U175 ( .A(n888), .B(n948), .Z(n892) );
  XOR U176 ( .A(n1057), .B(n1117), .Z(n1061) );
  XOR U177 ( .A(n1226), .B(n1292), .Z(n1230) );
  XOR U178 ( .A(n1402), .B(n1464), .Z(n1406) );
  XOR U179 ( .A(n1574), .B(n1636), .Z(n1578) );
  XOR U180 ( .A(n1746), .B(n1808), .Z(n1750) );
  XOR U181 ( .A(n1918), .B(n1980), .Z(n1922) );
  XOR U182 ( .A(n2090), .B(n2152), .Z(n2094) );
  XOR U183 ( .A(n2262), .B(n2324), .Z(n2266) );
  XOR U184 ( .A(n2434), .B(n2496), .Z(n2438) );
  XOR U185 ( .A(n2606), .B(n2668), .Z(n2610) );
  XOR U186 ( .A(n2778), .B(n2840), .Z(n2782) );
  XOR U187 ( .A(n2950), .B(n3012), .Z(n2954) );
  XOR U188 ( .A(n3122), .B(n3184), .Z(n3126) );
  XOR U189 ( .A(n3294), .B(n3356), .Z(n3298) );
  XOR U190 ( .A(n3466), .B(n3528), .Z(n3470) );
  XOR U191 ( .A(n3638), .B(n3700), .Z(n3642) );
  XOR U192 ( .A(n3810), .B(n3872), .Z(n3814) );
  XOR U193 ( .A(n391), .B(n439), .Z(n395) );
  XOR U194 ( .A(n4430), .B(n4475), .Z(n4435) );
  XOR U195 ( .A(n4311), .B(n4355), .Z(n4315) );
  XOR U196 ( .A(n4167), .B(n4211), .Z(n4171) );
  XOR U197 ( .A(n3997), .B(n4041), .Z(n4001) );
  XOR U198 ( .A(n229), .B(n277), .Z(n233) );
  XOR U199 ( .A(n154), .B(n196), .Z(n158) );
  XOR U200 ( .A(n564), .B(n607), .Z(n568) );
  XOR U201 ( .A(n734), .B(n776), .Z(n738) );
  XOR U202 ( .A(n903), .B(n945), .Z(n907) );
  XOR U203 ( .A(n1072), .B(n1114), .Z(n1076) );
  XOR U204 ( .A(n1241), .B(n1289), .Z(n1245) );
  XOR U205 ( .A(n1417), .B(n1461), .Z(n1421) );
  XOR U206 ( .A(n1589), .B(n1633), .Z(n1593) );
  XOR U207 ( .A(n1761), .B(n1805), .Z(n1765) );
  XOR U208 ( .A(n1933), .B(n1977), .Z(n1937) );
  XOR U209 ( .A(n2105), .B(n2149), .Z(n2109) );
  XOR U210 ( .A(n2277), .B(n2321), .Z(n2281) );
  XOR U211 ( .A(n2449), .B(n2493), .Z(n2453) );
  XOR U212 ( .A(n2621), .B(n2665), .Z(n2625) );
  XOR U213 ( .A(n2793), .B(n2837), .Z(n2797) );
  XOR U214 ( .A(n2965), .B(n3009), .Z(n2969) );
  XOR U215 ( .A(n3137), .B(n3181), .Z(n3141) );
  XOR U216 ( .A(n3309), .B(n3353), .Z(n3313) );
  XOR U217 ( .A(n3481), .B(n3525), .Z(n3485) );
  XOR U218 ( .A(n3653), .B(n3697), .Z(n3657) );
  XOR U219 ( .A(n3825), .B(n3869), .Z(n3829) );
  XOR U220 ( .A(n406), .B(n436), .Z(n410) );
  XOR U221 ( .A(n4542), .B(n4568), .Z(n4546) );
  XOR U222 ( .A(n4446), .B(n4472), .Z(n4450) );
  XOR U223 ( .A(n4326), .B(n4352), .Z(n4330) );
  XOR U224 ( .A(n4182), .B(n4208), .Z(n4186) );
  XOR U225 ( .A(n4012), .B(n4038), .Z(n4016) );
  XOR U226 ( .A(n169), .B(n193), .Z(n173) );
  XOR U227 ( .A(n329), .B(n354), .Z(n333) );
  XOR U228 ( .A(n579), .B(n604), .Z(n583) );
  XOR U229 ( .A(n749), .B(n773), .Z(n753) );
  XOR U230 ( .A(n918), .B(n942), .Z(n922) );
  XOR U231 ( .A(n1087), .B(n1111), .Z(n1091) );
  XOR U232 ( .A(n1256), .B(n1286), .Z(n1260) );
  XOR U233 ( .A(n1432), .B(n1458), .Z(n1436) );
  XOR U234 ( .A(n1604), .B(n1630), .Z(n1608) );
  XOR U235 ( .A(n1776), .B(n1802), .Z(n1780) );
  XOR U236 ( .A(n1948), .B(n1974), .Z(n1952) );
  XOR U237 ( .A(n2120), .B(n2146), .Z(n2124) );
  XOR U238 ( .A(n2292), .B(n2318), .Z(n2296) );
  XOR U239 ( .A(n2464), .B(n2490), .Z(n2468) );
  XOR U240 ( .A(n2636), .B(n2662), .Z(n2640) );
  XOR U241 ( .A(n2808), .B(n2834), .Z(n2812) );
  XOR U242 ( .A(n2980), .B(n3006), .Z(n2984) );
  XOR U243 ( .A(n3152), .B(n3178), .Z(n3156) );
  XOR U244 ( .A(n3324), .B(n3350), .Z(n3328) );
  XOR U245 ( .A(n3496), .B(n3522), .Z(n3500) );
  XOR U246 ( .A(n3668), .B(n3694), .Z(n3672) );
  XOR U247 ( .A(n3840), .B(n3866), .Z(n3844) );
  AND U248 ( .A(n265), .B(n264), .Z(n184) );
  AND U249 ( .A(n595), .B(n594), .Z(n506) );
  AND U250 ( .A(n934), .B(n933), .Z(n848) );
  XOR U251 ( .A(n4226), .B(n4289), .Z(n4231) );
  XOR U252 ( .A(n4068), .B(n4130), .Z(n4072) );
  XOR U253 ( .A(n213), .B(n280), .Z(n218) );
  XOR U254 ( .A(n461), .B(n522), .Z(n465) );
  XOR U255 ( .A(n634), .B(n695), .Z(n638) );
  XOR U256 ( .A(n803), .B(n864), .Z(n807) );
  XOR U257 ( .A(n972), .B(n1033), .Z(n976) );
  XOR U258 ( .A(n1141), .B(n1202), .Z(n1145) );
  XOR U259 ( .A(n1316), .B(n1378), .Z(n1320) );
  XOR U260 ( .A(n1488), .B(n1550), .Z(n1492) );
  XOR U261 ( .A(n1660), .B(n1722), .Z(n1664) );
  XOR U262 ( .A(n1832), .B(n1894), .Z(n1836) );
  XOR U263 ( .A(n2004), .B(n2066), .Z(n2008) );
  XOR U264 ( .A(n2176), .B(n2238), .Z(n2180) );
  XOR U265 ( .A(n2348), .B(n2410), .Z(n2352) );
  XOR U266 ( .A(n2520), .B(n2582), .Z(n2524) );
  XOR U267 ( .A(n2692), .B(n2754), .Z(n2696) );
  XOR U268 ( .A(n2864), .B(n2926), .Z(n2868) );
  XOR U269 ( .A(n3036), .B(n3098), .Z(n3040) );
  XOR U270 ( .A(n3208), .B(n3270), .Z(n3212) );
  XOR U271 ( .A(n3380), .B(n3442), .Z(n3384) );
  XOR U272 ( .A(n3552), .B(n3614), .Z(n3556) );
  XOR U273 ( .A(n3724), .B(n3786), .Z(n3728) );
  XOR U274 ( .A(n3896), .B(n3958), .Z(n3900) );
  XOR U275 ( .A(n4374), .B(n4418), .Z(n4378) );
  XOR U276 ( .A(n4242), .B(n4286), .Z(n4246) );
  XOR U277 ( .A(n4083), .B(n4127), .Z(n4087) );
  XOR U278 ( .A(n139), .B(n199), .Z(n143) );
  XOR U279 ( .A(n476), .B(n519), .Z(n480) );
  XOR U280 ( .A(n649), .B(n692), .Z(n653) );
  XOR U281 ( .A(n818), .B(n861), .Z(n822) );
  XOR U282 ( .A(n987), .B(n1030), .Z(n991) );
  XOR U283 ( .A(n1156), .B(n1199), .Z(n1160) );
  XOR U284 ( .A(n1331), .B(n1375), .Z(n1335) );
  XOR U285 ( .A(n1503), .B(n1547), .Z(n1507) );
  XOR U286 ( .A(n1675), .B(n1719), .Z(n1679) );
  XOR U287 ( .A(n1847), .B(n1891), .Z(n1851) );
  XOR U288 ( .A(n2019), .B(n2063), .Z(n2023) );
  XOR U289 ( .A(n2191), .B(n2235), .Z(n2195) );
  XOR U290 ( .A(n2363), .B(n2407), .Z(n2367) );
  XOR U291 ( .A(n2535), .B(n2579), .Z(n2539) );
  XOR U292 ( .A(n2707), .B(n2751), .Z(n2711) );
  XOR U293 ( .A(n2879), .B(n2923), .Z(n2883) );
  XOR U294 ( .A(n3051), .B(n3095), .Z(n3055) );
  XOR U295 ( .A(n3223), .B(n3267), .Z(n3227) );
  XOR U296 ( .A(n3395), .B(n3439), .Z(n3399) );
  XOR U297 ( .A(n3567), .B(n3611), .Z(n3571) );
  XOR U298 ( .A(n3739), .B(n3783), .Z(n3743) );
  XOR U299 ( .A(n3911), .B(n3955), .Z(n3915) );
  XOR U300 ( .A(n234), .B(n276), .Z(n238) );
  XOR U301 ( .A(n4580), .B(n4607), .Z(n4585) );
  XOR U302 ( .A(n4497), .B(n4523), .Z(n4501) );
  XOR U303 ( .A(n4389), .B(n4415), .Z(n4393) );
  XOR U304 ( .A(n4257), .B(n4283), .Z(n4261) );
  XOR U305 ( .A(n4098), .B(n4124), .Z(n4102) );
  XOR U306 ( .A(n249), .B(n273), .Z(n253) );
  XOR U307 ( .A(n411), .B(n435), .Z(n415) );
  XOR U308 ( .A(n664), .B(n689), .Z(n668) );
  XOR U309 ( .A(n833), .B(n858), .Z(n837) );
  XOR U310 ( .A(n1002), .B(n1027), .Z(n1006) );
  XOR U311 ( .A(n1171), .B(n1196), .Z(n1175) );
  XOR U312 ( .A(n1346), .B(n1372), .Z(n1350) );
  XOR U313 ( .A(n1518), .B(n1544), .Z(n1522) );
  XOR U314 ( .A(n1690), .B(n1716), .Z(n1694) );
  XOR U315 ( .A(n1862), .B(n1888), .Z(n1866) );
  XOR U316 ( .A(n2034), .B(n2060), .Z(n2038) );
  XOR U317 ( .A(n2206), .B(n2232), .Z(n2210) );
  XOR U318 ( .A(n2378), .B(n2404), .Z(n2382) );
  XOR U319 ( .A(n2550), .B(n2576), .Z(n2554) );
  XOR U320 ( .A(n2722), .B(n2748), .Z(n2726) );
  XOR U321 ( .A(n2894), .B(n2920), .Z(n2898) );
  XOR U322 ( .A(n3066), .B(n3092), .Z(n3070) );
  XOR U323 ( .A(n3238), .B(n3264), .Z(n3242) );
  XOR U324 ( .A(n3410), .B(n3436), .Z(n3414) );
  XOR U325 ( .A(n3582), .B(n3608), .Z(n3586) );
  XOR U326 ( .A(n3754), .B(n3780), .Z(n3758) );
  XOR U327 ( .A(n3926), .B(n3952), .Z(n3930) );
  XNOR U328 ( .A(n584), .B(n603), .Z(n592) );
  AND U329 ( .A(n345), .B(n344), .Z(n264) );
  AND U330 ( .A(n680), .B(n679), .Z(n594) );
  AND U331 ( .A(n1018), .B(n1017), .Z(n933) );
  XOR U332 ( .A(n3971), .B(n4046), .Z(n3976) );
  XOR U333 ( .A(n538), .B(n612), .Z(n543) );
  XOR U334 ( .A(n708), .B(n781), .Z(n713) );
  XOR U335 ( .A(n877), .B(n950), .Z(n882) );
  XOR U336 ( .A(n1046), .B(n1119), .Z(n1051) );
  XOR U337 ( .A(n1215), .B(n1294), .Z(n1220) );
  XOR U338 ( .A(n1391), .B(n1466), .Z(n1396) );
  XOR U339 ( .A(n1563), .B(n1638), .Z(n1568) );
  XOR U340 ( .A(n1735), .B(n1810), .Z(n1740) );
  XOR U341 ( .A(n1907), .B(n1982), .Z(n1912) );
  XOR U342 ( .A(n2079), .B(n2154), .Z(n2084) );
  XOR U343 ( .A(n2251), .B(n2326), .Z(n2256) );
  XOR U344 ( .A(n2423), .B(n2498), .Z(n2428) );
  XOR U345 ( .A(n2595), .B(n2670), .Z(n2600) );
  XOR U346 ( .A(n2767), .B(n2842), .Z(n2772) );
  XOR U347 ( .A(n2939), .B(n3014), .Z(n2944) );
  XOR U348 ( .A(n3111), .B(n3186), .Z(n3116) );
  XOR U349 ( .A(n3283), .B(n3358), .Z(n3288) );
  XOR U350 ( .A(n3455), .B(n3530), .Z(n3460) );
  XOR U351 ( .A(n3627), .B(n3702), .Z(n3632) );
  XOR U352 ( .A(n3799), .B(n3874), .Z(n3804) );
  XOR U353 ( .A(n4300), .B(n4357), .Z(n4305) );
  XOR U354 ( .A(n4157), .B(n4213), .Z(n4161) );
  XOR U355 ( .A(n3987), .B(n4043), .Z(n3991) );
  XOR U356 ( .A(n219), .B(n279), .Z(n223) );
  XOR U357 ( .A(n386), .B(n440), .Z(n390) );
  XOR U358 ( .A(n554), .B(n609), .Z(n558) );
  XOR U359 ( .A(n724), .B(n778), .Z(n728) );
  XOR U360 ( .A(n893), .B(n947), .Z(n897) );
  XOR U361 ( .A(n1062), .B(n1116), .Z(n1066) );
  XOR U362 ( .A(n1231), .B(n1291), .Z(n1235) );
  XOR U363 ( .A(n1407), .B(n1463), .Z(n1411) );
  XOR U364 ( .A(n1579), .B(n1635), .Z(n1583) );
  XOR U365 ( .A(n1751), .B(n1807), .Z(n1755) );
  XOR U366 ( .A(n1923), .B(n1979), .Z(n1927) );
  XOR U367 ( .A(n2095), .B(n2151), .Z(n2099) );
  XOR U368 ( .A(n2267), .B(n2323), .Z(n2271) );
  XOR U369 ( .A(n2439), .B(n2495), .Z(n2443) );
  XOR U370 ( .A(n2611), .B(n2667), .Z(n2615) );
  XOR U371 ( .A(n2783), .B(n2839), .Z(n2787) );
  XOR U372 ( .A(n2955), .B(n3011), .Z(n2959) );
  XOR U373 ( .A(n3127), .B(n3183), .Z(n3131) );
  XOR U374 ( .A(n3299), .B(n3355), .Z(n3303) );
  XOR U375 ( .A(n3471), .B(n3527), .Z(n3475) );
  XOR U376 ( .A(n3643), .B(n3699), .Z(n3647) );
  XOR U377 ( .A(n3815), .B(n3871), .Z(n3819) );
  XOR U378 ( .A(n4436), .B(n4474), .Z(n4440) );
  XOR U379 ( .A(n4316), .B(n4354), .Z(n4320) );
  XOR U380 ( .A(n4172), .B(n4210), .Z(n4176) );
  XOR U381 ( .A(n4002), .B(n4040), .Z(n4006) );
  XOR U382 ( .A(n144), .B(n198), .Z(n148) );
  XOR U383 ( .A(n159), .B(n195), .Z(n163) );
  XOR U384 ( .A(n319), .B(n356), .Z(n323) );
  XOR U385 ( .A(n569), .B(n606), .Z(n573) );
  XOR U386 ( .A(n739), .B(n775), .Z(n743) );
  XOR U387 ( .A(n908), .B(n944), .Z(n912) );
  XOR U388 ( .A(n1077), .B(n1113), .Z(n1081) );
  XOR U389 ( .A(n1246), .B(n1288), .Z(n1250) );
  XOR U390 ( .A(n1422), .B(n1460), .Z(n1426) );
  XOR U391 ( .A(n1594), .B(n1632), .Z(n1598) );
  XOR U392 ( .A(n1766), .B(n1804), .Z(n1770) );
  XOR U393 ( .A(n1938), .B(n1976), .Z(n1942) );
  XOR U394 ( .A(n2110), .B(n2148), .Z(n2114) );
  XOR U395 ( .A(n2282), .B(n2320), .Z(n2286) );
  XOR U396 ( .A(n2454), .B(n2492), .Z(n2458) );
  XOR U397 ( .A(n2626), .B(n2664), .Z(n2630) );
  XOR U398 ( .A(n2798), .B(n2836), .Z(n2802) );
  XOR U399 ( .A(n2970), .B(n3008), .Z(n2974) );
  XOR U400 ( .A(n3142), .B(n3180), .Z(n3146) );
  XOR U401 ( .A(n3314), .B(n3352), .Z(n3318) );
  XOR U402 ( .A(n3486), .B(n3524), .Z(n3490) );
  XOR U403 ( .A(n3658), .B(n3696), .Z(n3662) );
  XOR U404 ( .A(n3830), .B(n3868), .Z(n3834) );
  XOR U405 ( .A(n486), .B(n517), .Z(n490) );
  XOR U406 ( .A(n4618), .B(n4639), .Z(n4628) );
  XOR U407 ( .A(n4547), .B(n4567), .Z(n4556) );
  XOR U408 ( .A(n4451), .B(n4471), .Z(n4460) );
  XOR U409 ( .A(n4331), .B(n4351), .Z(n4340) );
  XOR U410 ( .A(n4187), .B(n4207), .Z(n4196) );
  XOR U411 ( .A(n4017), .B(n4037), .Z(n4026) );
  XOR U412 ( .A(n254), .B(n272), .Z(n263) );
  XOR U413 ( .A(n416), .B(n434), .Z(n425) );
  XOR U414 ( .A(n754), .B(n772), .Z(n763) );
  XOR U415 ( .A(n923), .B(n941), .Z(n932) );
  XOR U416 ( .A(n1092), .B(n1110), .Z(n1101) );
  XOR U417 ( .A(n1261), .B(n1285), .Z(n1270) );
  XOR U418 ( .A(n1437), .B(n1457), .Z(n1446) );
  XOR U419 ( .A(n1609), .B(n1629), .Z(n1618) );
  XOR U420 ( .A(n1781), .B(n1801), .Z(n1790) );
  XOR U421 ( .A(n1953), .B(n1973), .Z(n1962) );
  XOR U422 ( .A(n2125), .B(n2145), .Z(n2134) );
  XOR U423 ( .A(n2297), .B(n2317), .Z(n2306) );
  XOR U424 ( .A(n2469), .B(n2489), .Z(n2478) );
  XOR U425 ( .A(n2641), .B(n2661), .Z(n2650) );
  XOR U426 ( .A(n2813), .B(n2833), .Z(n2822) );
  XOR U427 ( .A(n2985), .B(n3005), .Z(n2994) );
  XOR U428 ( .A(n3157), .B(n3177), .Z(n3166) );
  XOR U429 ( .A(n3329), .B(n3349), .Z(n3338) );
  XOR U430 ( .A(n3501), .B(n3521), .Z(n3510) );
  XOR U431 ( .A(n3673), .B(n3693), .Z(n3682) );
  XOR U432 ( .A(n3845), .B(n3865), .Z(n3854) );
  XOR U433 ( .A(n592), .B(n599), .Z(n588) );
  AND U434 ( .A(n427), .B(n426), .Z(n344) );
  AND U435 ( .A(n765), .B(n764), .Z(n679) );
  AND U436 ( .A(n1103), .B(n1102), .Z(n1017) );
  XOR U437 ( .A(n4057), .B(n4132), .Z(n4062) );
  XOR U438 ( .A(n623), .B(n697), .Z(n628) );
  XOR U439 ( .A(n792), .B(n866), .Z(n797) );
  XOR U440 ( .A(n961), .B(n1035), .Z(n966) );
  XOR U441 ( .A(n1130), .B(n1204), .Z(n1135) );
  XOR U442 ( .A(n1305), .B(n1380), .Z(n1310) );
  XOR U443 ( .A(n1477), .B(n1552), .Z(n1482) );
  XOR U444 ( .A(n1649), .B(n1724), .Z(n1654) );
  XOR U445 ( .A(n1821), .B(n1896), .Z(n1826) );
  XOR U446 ( .A(n1993), .B(n2068), .Z(n1998) );
  XOR U447 ( .A(n2165), .B(n2240), .Z(n2170) );
  XOR U448 ( .A(n2337), .B(n2412), .Z(n2342) );
  XOR U449 ( .A(n2509), .B(n2584), .Z(n2514) );
  XOR U450 ( .A(n2681), .B(n2756), .Z(n2686) );
  XOR U451 ( .A(n2853), .B(n2928), .Z(n2858) );
  XOR U452 ( .A(n3025), .B(n3100), .Z(n3030) );
  XOR U453 ( .A(n3197), .B(n3272), .Z(n3202) );
  XOR U454 ( .A(n3369), .B(n3444), .Z(n3374) );
  XOR U455 ( .A(n3541), .B(n3616), .Z(n3546) );
  XOR U456 ( .A(n3713), .B(n3788), .Z(n3718) );
  XOR U457 ( .A(n3885), .B(n3960), .Z(n3890) );
  XOR U458 ( .A(n299), .B(n361), .Z(n303) );
  XOR U459 ( .A(n4232), .B(n4288), .Z(n4236) );
  XOR U460 ( .A(n4073), .B(n4129), .Z(n4077) );
  XOR U461 ( .A(n466), .B(n521), .Z(n470) );
  XOR U462 ( .A(n639), .B(n694), .Z(n643) );
  XOR U463 ( .A(n808), .B(n863), .Z(n812) );
  XOR U464 ( .A(n977), .B(n1032), .Z(n981) );
  XOR U465 ( .A(n1146), .B(n1201), .Z(n1150) );
  XOR U466 ( .A(n1321), .B(n1377), .Z(n1325) );
  XOR U467 ( .A(n1493), .B(n1549), .Z(n1497) );
  XOR U468 ( .A(n1665), .B(n1721), .Z(n1669) );
  XOR U469 ( .A(n1837), .B(n1893), .Z(n1841) );
  XOR U470 ( .A(n2009), .B(n2065), .Z(n2013) );
  XOR U471 ( .A(n2181), .B(n2237), .Z(n2185) );
  XOR U472 ( .A(n2353), .B(n2409), .Z(n2357) );
  XOR U473 ( .A(n2525), .B(n2581), .Z(n2529) );
  XOR U474 ( .A(n2697), .B(n2753), .Z(n2701) );
  XOR U475 ( .A(n2869), .B(n2925), .Z(n2873) );
  XOR U476 ( .A(n3041), .B(n3097), .Z(n3045) );
  XOR U477 ( .A(n3213), .B(n3269), .Z(n3217) );
  XOR U478 ( .A(n3385), .B(n3441), .Z(n3389) );
  XOR U479 ( .A(n3557), .B(n3613), .Z(n3561) );
  XOR U480 ( .A(n3729), .B(n3785), .Z(n3733) );
  XOR U481 ( .A(n3901), .B(n3957), .Z(n3905) );
  XOR U482 ( .A(n133), .B(n200), .Z(n138) );
  XOR U483 ( .A(n314), .B(n357), .Z(n318) );
  XOR U484 ( .A(n4486), .B(n4525), .Z(n4491) );
  XOR U485 ( .A(n4379), .B(n4417), .Z(n4383) );
  XOR U486 ( .A(n4247), .B(n4285), .Z(n4251) );
  XOR U487 ( .A(n4088), .B(n4126), .Z(n4092) );
  XOR U488 ( .A(n481), .B(n518), .Z(n485) );
  XOR U489 ( .A(n654), .B(n691), .Z(n658) );
  XOR U490 ( .A(n823), .B(n860), .Z(n827) );
  XOR U491 ( .A(n992), .B(n1029), .Z(n996) );
  XOR U492 ( .A(n1161), .B(n1198), .Z(n1165) );
  XOR U493 ( .A(n1336), .B(n1374), .Z(n1340) );
  XOR U494 ( .A(n1508), .B(n1546), .Z(n1512) );
  XOR U495 ( .A(n1680), .B(n1718), .Z(n1684) );
  XOR U496 ( .A(n1852), .B(n1890), .Z(n1856) );
  XOR U497 ( .A(n2024), .B(n2062), .Z(n2028) );
  XOR U498 ( .A(n2196), .B(n2234), .Z(n2200) );
  XOR U499 ( .A(n2368), .B(n2406), .Z(n2372) );
  XOR U500 ( .A(n2540), .B(n2578), .Z(n2544) );
  XOR U501 ( .A(n2712), .B(n2750), .Z(n2716) );
  XOR U502 ( .A(n2884), .B(n2922), .Z(n2888) );
  XOR U503 ( .A(n3056), .B(n3094), .Z(n3060) );
  XOR U504 ( .A(n3228), .B(n3266), .Z(n3232) );
  XOR U505 ( .A(n3400), .B(n3438), .Z(n3404) );
  XOR U506 ( .A(n3572), .B(n3610), .Z(n3576) );
  XOR U507 ( .A(n3744), .B(n3782), .Z(n3748) );
  XOR U508 ( .A(n3916), .B(n3954), .Z(n3920) );
  XOR U509 ( .A(n149), .B(n197), .Z(n153) );
  XOR U510 ( .A(n4586), .B(n4606), .Z(n4595) );
  XOR U511 ( .A(n4502), .B(n4522), .Z(n4511) );
  XOR U512 ( .A(n4394), .B(n4414), .Z(n4403) );
  XOR U513 ( .A(n4262), .B(n4282), .Z(n4271) );
  XOR U514 ( .A(n4103), .B(n4123), .Z(n4112) );
  XOR U515 ( .A(n174), .B(n192), .Z(n183) );
  XOR U516 ( .A(n334), .B(n353), .Z(n343) );
  XOR U517 ( .A(n496), .B(n515), .Z(n504) );
  XOR U518 ( .A(n669), .B(n688), .Z(n678) );
  XOR U519 ( .A(n838), .B(n857), .Z(n847) );
  XOR U520 ( .A(n1007), .B(n1026), .Z(n1016) );
  XOR U521 ( .A(n1176), .B(n1195), .Z(n1185) );
  XOR U522 ( .A(n1351), .B(n1371), .Z(n1360) );
  XOR U523 ( .A(n1523), .B(n1543), .Z(n1532) );
  XOR U524 ( .A(n1695), .B(n1715), .Z(n1704) );
  XOR U525 ( .A(n1867), .B(n1887), .Z(n1876) );
  XOR U526 ( .A(n2039), .B(n2059), .Z(n2048) );
  XOR U527 ( .A(n2211), .B(n2231), .Z(n2220) );
  XOR U528 ( .A(n2383), .B(n2403), .Z(n2392) );
  XOR U529 ( .A(n2555), .B(n2575), .Z(n2564) );
  XOR U530 ( .A(n2727), .B(n2747), .Z(n2736) );
  XOR U531 ( .A(n2899), .B(n2919), .Z(n2908) );
  XOR U532 ( .A(n3071), .B(n3091), .Z(n3080) );
  XOR U533 ( .A(n3243), .B(n3263), .Z(n3252) );
  XOR U534 ( .A(n3415), .B(n3435), .Z(n3424) );
  XOR U535 ( .A(n3587), .B(n3607), .Z(n3596) );
  XOR U536 ( .A(n3759), .B(n3779), .Z(n3768) );
  XOR U537 ( .A(n3931), .B(n3951), .Z(n3940) );
  XNOR U538 ( .A(n588), .B(n587), .Z(n514) );
  XOR U539 ( .A(n4685), .B(n4679), .Z(n4692) );
  NANDN U540 ( .A(n185), .B(n184), .Z(n75) );
  AND U541 ( .A(n507), .B(n506), .Z(n426) );
  AND U542 ( .A(n849), .B(n848), .Z(n764) );
  AND U543 ( .A(n1187), .B(n1186), .Z(n1102) );
  XOR U544 ( .A(n1), .B(n2), .Z(swire[63]) );
  XOR U545 ( .A(n3), .B(n4), .Z(n2) );
  AND U546 ( .A(a[62]), .B(b[1]), .Z(n4) );
  AND U547 ( .A(a[61]), .B(b[2]), .Z(n3) );
  XOR U548 ( .A(n5), .B(n6), .Z(n1) );
  XOR U549 ( .A(n7), .B(n8), .Z(n6) );
  XOR U550 ( .A(n9), .B(n10), .Z(n8) );
  AND U551 ( .A(a[63]), .B(b[0]), .Z(n10) );
  AND U552 ( .A(a[60]), .B(b[3]), .Z(n9) );
  XOR U553 ( .A(n11), .B(n12), .Z(n7) );
  XOR U554 ( .A(n13), .B(n14), .Z(n12) );
  XOR U555 ( .A(n15), .B(n16), .Z(n14) );
  AND U556 ( .A(a[59]), .B(b[4]), .Z(n16) );
  AND U557 ( .A(a[54]), .B(b[9]), .Z(n15) );
  XOR U558 ( .A(n17), .B(n18), .Z(n13) );
  AND U559 ( .A(a[53]), .B(b[10]), .Z(n18) );
  AND U560 ( .A(a[52]), .B(b[11]), .Z(n17) );
  XOR U561 ( .A(n19), .B(n20), .Z(n11) );
  XOR U562 ( .A(n21), .B(n22), .Z(n20) );
  AND U563 ( .A(a[51]), .B(b[12]), .Z(n22) );
  AND U564 ( .A(a[50]), .B(b[13]), .Z(n21) );
  XOR U565 ( .A(n23), .B(n24), .Z(n19) );
  AND U566 ( .A(a[49]), .B(b[14]), .Z(n24) );
  AND U567 ( .A(a[48]), .B(b[15]), .Z(n23) );
  XOR U568 ( .A(n25), .B(n26), .Z(n5) );
  XOR U569 ( .A(n27), .B(n28), .Z(n26) );
  AND U570 ( .A(a[58]), .B(b[5]), .Z(n28) );
  AND U571 ( .A(a[57]), .B(b[6]), .Z(n27) );
  XOR U572 ( .A(n29), .B(n30), .Z(n25) );
  AND U573 ( .A(a[56]), .B(b[7]), .Z(n30) );
  AND U574 ( .A(a[55]), .B(b[8]), .Z(n29) );
  XOR U575 ( .A(n31), .B(n32), .Z(swire[62]) );
  XOR U576 ( .A(n33), .B(n34), .Z(n32) );
  XOR U577 ( .A(n35), .B(n36), .Z(n34) );
  XOR U578 ( .A(n37), .B(n38), .Z(n36) );
  XOR U579 ( .A(n39), .B(n40), .Z(n38) );
  XOR U580 ( .A(n41), .B(n42), .Z(n40) );
  AND U581 ( .A(a[59]), .B(b[3]), .Z(n41) );
  XOR U582 ( .A(n43), .B(n44), .Z(n39) );
  XOR U583 ( .A(n45), .B(n46), .Z(n44) );
  XOR U584 ( .A(n47), .B(n48), .Z(n46) );
  XOR U585 ( .A(n49), .B(n47), .Z(n48) );
  AND U586 ( .A(a[53]), .B(b[9]), .Z(n49) );
  XOR U587 ( .A(n50), .B(n51), .Z(n47) );
  ANDN U588 ( .B(n52), .A(n53), .Z(n50) );
  XOR U589 ( .A(n54), .B(n55), .Z(n45) );
  AND U590 ( .A(a[52]), .B(b[10]), .Z(n55) );
  AND U591 ( .A(a[51]), .B(b[11]), .Z(n54) );
  XOR U592 ( .A(n56), .B(n57), .Z(n43) );
  XOR U593 ( .A(n58), .B(n59), .Z(n57) );
  AND U594 ( .A(a[50]), .B(b[12]), .Z(n59) );
  AND U595 ( .A(a[49]), .B(b[13]), .Z(n58) );
  XOR U596 ( .A(n60), .B(n61), .Z(n56) );
  AND U597 ( .A(b[14]), .B(a[48]), .Z(n61) );
  AND U598 ( .A(b[15]), .B(a[47]), .Z(n60) );
  XOR U599 ( .A(n62), .B(n42), .Z(n37) );
  XNOR U600 ( .A(n63), .B(n64), .Z(n42) );
  ANDN U601 ( .B(n65), .A(n66), .Z(n63) );
  AND U602 ( .A(a[58]), .B(b[4]), .Z(n62) );
  XOR U603 ( .A(n67), .B(n68), .Z(n35) );
  XOR U604 ( .A(n69), .B(n70), .Z(n68) );
  AND U605 ( .A(a[57]), .B(b[5]), .Z(n70) );
  AND U606 ( .A(a[56]), .B(b[6]), .Z(n69) );
  XOR U607 ( .A(n71), .B(n72), .Z(n67) );
  AND U608 ( .A(a[55]), .B(b[7]), .Z(n72) );
  AND U609 ( .A(b[8]), .B(a[54]), .Z(n71) );
  AND U610 ( .A(a[62]), .B(b[0]), .Z(n33) );
  XOR U611 ( .A(n73), .B(n74), .Z(n31) );
  AND U612 ( .A(a[61]), .B(b[1]), .Z(n74) );
  AND U613 ( .A(b[2]), .B(a[60]), .Z(n73) );
  XNOR U614 ( .A(n75), .B(n76), .Z(swire[61]) );
  XOR U615 ( .A(n77), .B(n78), .Z(n76) );
  XNOR U616 ( .A(n79), .B(n75), .Z(n78) );
  AND U617 ( .A(a[61]), .B(b[0]), .Z(n79) );
  XOR U618 ( .A(n80), .B(n81), .Z(n77) );
  XNOR U619 ( .A(n82), .B(n83), .Z(n81) );
  AND U620 ( .A(b[1]), .B(a[60]), .Z(n83) );
  XNOR U621 ( .A(n66), .B(n84), .Z(n80) );
  XNOR U622 ( .A(n82), .B(n65), .Z(n84) );
  XNOR U623 ( .A(n85), .B(n64), .Z(n65) );
  AND U624 ( .A(b[2]), .B(a[59]), .Z(n85) );
  OR U625 ( .A(n86), .B(n87), .Z(n82) );
  XOR U626 ( .A(n88), .B(n89), .Z(n66) );
  XNOR U627 ( .A(n64), .B(n90), .Z(n89) );
  XOR U628 ( .A(n91), .B(n92), .Z(n90) );
  XOR U629 ( .A(n93), .B(n94), .Z(n92) );
  XOR U630 ( .A(n95), .B(n96), .Z(n94) );
  XOR U631 ( .A(n97), .B(n98), .Z(n96) );
  XOR U632 ( .A(n99), .B(n100), .Z(n98) );
  XOR U633 ( .A(n101), .B(n102), .Z(n100) );
  XOR U634 ( .A(n103), .B(n104), .Z(n102) );
  XOR U635 ( .A(n105), .B(n106), .Z(n104) );
  XOR U636 ( .A(n52), .B(n107), .Z(n106) );
  XOR U637 ( .A(n108), .B(n53), .Z(n107) );
  XOR U638 ( .A(n109), .B(n110), .Z(n53) );
  XOR U639 ( .A(n51), .B(n111), .Z(n110) );
  XOR U640 ( .A(n112), .B(n113), .Z(n111) );
  XOR U641 ( .A(n114), .B(n115), .Z(n113) );
  XOR U642 ( .A(n116), .B(n117), .Z(n115) );
  XOR U643 ( .A(n118), .B(n119), .Z(n117) );
  XOR U644 ( .A(n120), .B(n121), .Z(n119) );
  XOR U645 ( .A(n122), .B(n123), .Z(n121) );
  XOR U646 ( .A(n124), .B(n125), .Z(n123) );
  XNOR U647 ( .A(n126), .B(n127), .Z(n125) );
  AND U648 ( .A(b[13]), .B(a[48]), .Z(n126) );
  XOR U649 ( .A(n128), .B(n129), .Z(n124) );
  AND U650 ( .A(b[14]), .B(a[47]), .Z(n129) );
  AND U651 ( .A(b[15]), .B(a[46]), .Z(n128) );
  XOR U652 ( .A(n130), .B(n127), .Z(n120) );
  XOR U653 ( .A(n131), .B(n132), .Z(n127) );
  NOR U654 ( .A(n133), .B(n134), .Z(n131) );
  AND U655 ( .A(a[49]), .B(b[12]), .Z(n130) );
  XOR U656 ( .A(n135), .B(n122), .Z(n116) );
  XOR U657 ( .A(n136), .B(n137), .Z(n122) );
  ANDN U658 ( .B(n138), .A(n139), .Z(n136) );
  AND U659 ( .A(a[50]), .B(b[11]), .Z(n135) );
  XOR U660 ( .A(n140), .B(n118), .Z(n112) );
  XOR U661 ( .A(n141), .B(n142), .Z(n118) );
  ANDN U662 ( .B(n143), .A(n144), .Z(n141) );
  AND U663 ( .A(a[51]), .B(b[10]), .Z(n140) );
  XOR U664 ( .A(n145), .B(n114), .Z(n109) );
  XOR U665 ( .A(n146), .B(n147), .Z(n114) );
  ANDN U666 ( .B(n148), .A(n149), .Z(n146) );
  AND U667 ( .A(a[52]), .B(b[9]), .Z(n145) );
  XOR U668 ( .A(n150), .B(n51), .Z(n52) );
  XOR U669 ( .A(n151), .B(n152), .Z(n51) );
  ANDN U670 ( .B(n153), .A(n154), .Z(n151) );
  AND U671 ( .A(b[8]), .B(a[53]), .Z(n150) );
  XOR U672 ( .A(n155), .B(n108), .Z(n103) );
  XOR U673 ( .A(n156), .B(n157), .Z(n108) );
  ANDN U674 ( .B(n158), .A(n159), .Z(n156) );
  AND U675 ( .A(b[7]), .B(a[54]), .Z(n155) );
  XOR U676 ( .A(n160), .B(n105), .Z(n99) );
  XOR U677 ( .A(n161), .B(n162), .Z(n105) );
  ANDN U678 ( .B(n163), .A(n164), .Z(n161) );
  AND U679 ( .A(a[55]), .B(b[6]), .Z(n160) );
  XOR U680 ( .A(n165), .B(n101), .Z(n95) );
  XOR U681 ( .A(n166), .B(n167), .Z(n101) );
  ANDN U682 ( .B(n168), .A(n169), .Z(n166) );
  AND U683 ( .A(a[56]), .B(b[5]), .Z(n165) );
  XOR U684 ( .A(n170), .B(n97), .Z(n91) );
  XOR U685 ( .A(n171), .B(n172), .Z(n97) );
  ANDN U686 ( .B(n173), .A(n174), .Z(n171) );
  AND U687 ( .A(a[57]), .B(b[4]), .Z(n170) );
  XNOR U688 ( .A(n175), .B(n176), .Z(n64) );
  NANDN U689 ( .A(n177), .B(n178), .Z(n176) );
  XOR U690 ( .A(n179), .B(n93), .Z(n88) );
  XNOR U691 ( .A(n180), .B(n181), .Z(n93) );
  AND U692 ( .A(n182), .B(n183), .Z(n180) );
  AND U693 ( .A(a[58]), .B(b[3]), .Z(n179) );
  XOR U694 ( .A(n184), .B(n185), .Z(swire[60]) );
  XOR U695 ( .A(n87), .B(n186), .Z(n185) );
  XOR U696 ( .A(n86), .B(n184), .Z(n186) );
  NAND U697 ( .A(a[60]), .B(b[0]), .Z(n86) );
  XOR U698 ( .A(n177), .B(n178), .Z(n87) );
  XOR U699 ( .A(n175), .B(n187), .Z(n178) );
  NAND U700 ( .A(b[1]), .B(a[59]), .Z(n187) );
  XOR U701 ( .A(n183), .B(n188), .Z(n177) );
  XOR U702 ( .A(n175), .B(n182), .Z(n188) );
  XNOR U703 ( .A(n189), .B(n181), .Z(n182) );
  AND U704 ( .A(b[2]), .B(a[58]), .Z(n189) );
  NANDN U705 ( .A(n190), .B(n191), .Z(n175) );
  XOR U706 ( .A(n181), .B(n173), .Z(n192) );
  XNOR U707 ( .A(n172), .B(n168), .Z(n193) );
  XNOR U708 ( .A(n167), .B(n163), .Z(n194) );
  XNOR U709 ( .A(n162), .B(n158), .Z(n195) );
  XNOR U710 ( .A(n157), .B(n153), .Z(n196) );
  XNOR U711 ( .A(n152), .B(n148), .Z(n197) );
  XNOR U712 ( .A(n147), .B(n143), .Z(n198) );
  XNOR U713 ( .A(n142), .B(n138), .Z(n199) );
  XOR U714 ( .A(n137), .B(n134), .Z(n200) );
  XOR U715 ( .A(n201), .B(n202), .Z(n134) );
  XOR U716 ( .A(n132), .B(n203), .Z(n202) );
  XOR U717 ( .A(n204), .B(n205), .Z(n203) );
  XNOR U718 ( .A(n206), .B(n207), .Z(n205) );
  AND U719 ( .A(b[13]), .B(a[47]), .Z(n206) );
  XOR U720 ( .A(n208), .B(n209), .Z(n204) );
  AND U721 ( .A(b[14]), .B(a[46]), .Z(n209) );
  AND U722 ( .A(b[15]), .B(a[45]), .Z(n208) );
  XOR U723 ( .A(n210), .B(n207), .Z(n201) );
  XOR U724 ( .A(n211), .B(n212), .Z(n207) );
  NOR U725 ( .A(n213), .B(n214), .Z(n211) );
  AND U726 ( .A(b[12]), .B(a[48]), .Z(n210) );
  XNOR U727 ( .A(n215), .B(n132), .Z(n133) );
  XOR U728 ( .A(n216), .B(n217), .Z(n132) );
  ANDN U729 ( .B(n218), .A(n219), .Z(n216) );
  AND U730 ( .A(a[49]), .B(b[11]), .Z(n215) );
  XNOR U731 ( .A(n220), .B(n137), .Z(n139) );
  XOR U732 ( .A(n221), .B(n222), .Z(n137) );
  ANDN U733 ( .B(n223), .A(n224), .Z(n221) );
  AND U734 ( .A(a[50]), .B(b[10]), .Z(n220) );
  XNOR U735 ( .A(n225), .B(n142), .Z(n144) );
  XOR U736 ( .A(n226), .B(n227), .Z(n142) );
  ANDN U737 ( .B(n228), .A(n229), .Z(n226) );
  AND U738 ( .A(a[51]), .B(b[9]), .Z(n225) );
  XNOR U739 ( .A(n230), .B(n147), .Z(n149) );
  XOR U740 ( .A(n231), .B(n232), .Z(n147) );
  ANDN U741 ( .B(n233), .A(n234), .Z(n231) );
  AND U742 ( .A(b[8]), .B(a[52]), .Z(n230) );
  XNOR U743 ( .A(n235), .B(n152), .Z(n154) );
  XOR U744 ( .A(n236), .B(n237), .Z(n152) );
  ANDN U745 ( .B(n238), .A(n239), .Z(n236) );
  AND U746 ( .A(b[7]), .B(a[53]), .Z(n235) );
  XNOR U747 ( .A(n240), .B(n157), .Z(n159) );
  XOR U748 ( .A(n241), .B(n242), .Z(n157) );
  ANDN U749 ( .B(n243), .A(n244), .Z(n241) );
  AND U750 ( .A(b[6]), .B(a[54]), .Z(n240) );
  XNOR U751 ( .A(n245), .B(n162), .Z(n164) );
  XOR U752 ( .A(n246), .B(n247), .Z(n162) );
  ANDN U753 ( .B(n248), .A(n249), .Z(n246) );
  AND U754 ( .A(a[55]), .B(b[5]), .Z(n245) );
  XNOR U755 ( .A(n250), .B(n167), .Z(n169) );
  XOR U756 ( .A(n251), .B(n252), .Z(n167) );
  ANDN U757 ( .B(n253), .A(n254), .Z(n251) );
  AND U758 ( .A(a[56]), .B(b[4]), .Z(n250) );
  XNOR U759 ( .A(n255), .B(n256), .Z(n181) );
  NANDN U760 ( .A(n257), .B(n258), .Z(n256) );
  XNOR U761 ( .A(n259), .B(n172), .Z(n174) );
  XNOR U762 ( .A(n260), .B(n261), .Z(n172) );
  AND U763 ( .A(n262), .B(n263), .Z(n260) );
  AND U764 ( .A(a[57]), .B(b[3]), .Z(n259) );
  XNOR U765 ( .A(n264), .B(n265), .Z(swire[59]) );
  XOR U766 ( .A(n191), .B(n266), .Z(n265) );
  XOR U767 ( .A(n190), .B(n264), .Z(n266) );
  NAND U768 ( .A(a[59]), .B(b[0]), .Z(n190) );
  XNOR U769 ( .A(n257), .B(n258), .Z(n191) );
  XOR U770 ( .A(n255), .B(n267), .Z(n258) );
  NAND U771 ( .A(b[1]), .B(a[58]), .Z(n267) );
  XOR U772 ( .A(n263), .B(n268), .Z(n257) );
  XOR U773 ( .A(n255), .B(n262), .Z(n268) );
  XNOR U774 ( .A(n269), .B(n261), .Z(n262) );
  AND U775 ( .A(b[2]), .B(a[57]), .Z(n269) );
  NANDN U776 ( .A(n270), .B(n271), .Z(n255) );
  XOR U777 ( .A(n261), .B(n253), .Z(n272) );
  XNOR U778 ( .A(n252), .B(n248), .Z(n273) );
  XNOR U779 ( .A(n247), .B(n243), .Z(n274) );
  XNOR U780 ( .A(n242), .B(n238), .Z(n275) );
  XNOR U781 ( .A(n237), .B(n233), .Z(n276) );
  XNOR U782 ( .A(n232), .B(n228), .Z(n277) );
  XNOR U783 ( .A(n227), .B(n223), .Z(n278) );
  XNOR U784 ( .A(n222), .B(n218), .Z(n279) );
  XOR U785 ( .A(n217), .B(n214), .Z(n280) );
  XOR U786 ( .A(n281), .B(n282), .Z(n214) );
  XOR U787 ( .A(n212), .B(n283), .Z(n282) );
  XOR U788 ( .A(n284), .B(n285), .Z(n283) );
  XNOR U789 ( .A(n286), .B(n287), .Z(n285) );
  AND U790 ( .A(b[13]), .B(a[46]), .Z(n286) );
  XOR U791 ( .A(n288), .B(n289), .Z(n284) );
  AND U792 ( .A(b[14]), .B(a[45]), .Z(n289) );
  AND U793 ( .A(b[15]), .B(a[44]), .Z(n288) );
  XOR U794 ( .A(n290), .B(n287), .Z(n281) );
  XOR U795 ( .A(n291), .B(n292), .Z(n287) );
  NOR U796 ( .A(n293), .B(n294), .Z(n291) );
  AND U797 ( .A(b[12]), .B(a[47]), .Z(n290) );
  XNOR U798 ( .A(n295), .B(n212), .Z(n213) );
  XOR U799 ( .A(n296), .B(n297), .Z(n212) );
  ANDN U800 ( .B(n298), .A(n299), .Z(n296) );
  AND U801 ( .A(b[11]), .B(a[48]), .Z(n295) );
  XNOR U802 ( .A(n300), .B(n217), .Z(n219) );
  XOR U803 ( .A(n301), .B(n302), .Z(n217) );
  ANDN U804 ( .B(n303), .A(n304), .Z(n301) );
  AND U805 ( .A(a[49]), .B(b[10]), .Z(n300) );
  XNOR U806 ( .A(n305), .B(n222), .Z(n224) );
  XOR U807 ( .A(n306), .B(n307), .Z(n222) );
  ANDN U808 ( .B(n308), .A(n309), .Z(n306) );
  AND U809 ( .A(a[50]), .B(b[9]), .Z(n305) );
  XNOR U810 ( .A(n310), .B(n227), .Z(n229) );
  XOR U811 ( .A(n311), .B(n312), .Z(n227) );
  ANDN U812 ( .B(n313), .A(n314), .Z(n311) );
  AND U813 ( .A(b[8]), .B(a[51]), .Z(n310) );
  XNOR U814 ( .A(n315), .B(n232), .Z(n234) );
  XOR U815 ( .A(n316), .B(n317), .Z(n232) );
  ANDN U816 ( .B(n318), .A(n319), .Z(n316) );
  AND U817 ( .A(b[7]), .B(a[52]), .Z(n315) );
  XNOR U818 ( .A(n320), .B(n237), .Z(n239) );
  XOR U819 ( .A(n321), .B(n322), .Z(n237) );
  ANDN U820 ( .B(n323), .A(n324), .Z(n321) );
  AND U821 ( .A(b[6]), .B(a[53]), .Z(n320) );
  XNOR U822 ( .A(n325), .B(n242), .Z(n244) );
  XOR U823 ( .A(n326), .B(n327), .Z(n242) );
  ANDN U824 ( .B(n328), .A(n329), .Z(n326) );
  AND U825 ( .A(b[5]), .B(a[54]), .Z(n325) );
  XNOR U826 ( .A(n330), .B(n247), .Z(n249) );
  XOR U827 ( .A(n331), .B(n332), .Z(n247) );
  ANDN U828 ( .B(n333), .A(n334), .Z(n331) );
  AND U829 ( .A(a[55]), .B(b[4]), .Z(n330) );
  XNOR U830 ( .A(n335), .B(n336), .Z(n261) );
  NANDN U831 ( .A(n337), .B(n338), .Z(n336) );
  XNOR U832 ( .A(n339), .B(n252), .Z(n254) );
  XNOR U833 ( .A(n340), .B(n341), .Z(n252) );
  AND U834 ( .A(n342), .B(n343), .Z(n340) );
  AND U835 ( .A(a[56]), .B(b[3]), .Z(n339) );
  XNOR U836 ( .A(n344), .B(n345), .Z(swire[58]) );
  XOR U837 ( .A(n271), .B(n347), .Z(n345) );
  XNOR U838 ( .A(n270), .B(n346), .Z(n347) );
  IV U839 ( .A(n344), .Z(n346) );
  NAND U840 ( .A(a[58]), .B(b[0]), .Z(n270) );
  XNOR U841 ( .A(n337), .B(n338), .Z(n271) );
  XOR U842 ( .A(n335), .B(n348), .Z(n338) );
  NAND U843 ( .A(b[1]), .B(a[57]), .Z(n348) );
  XOR U844 ( .A(n343), .B(n349), .Z(n337) );
  XOR U845 ( .A(n335), .B(n342), .Z(n349) );
  XNOR U846 ( .A(n350), .B(n341), .Z(n342) );
  AND U847 ( .A(b[2]), .B(a[56]), .Z(n350) );
  NANDN U848 ( .A(n351), .B(n352), .Z(n335) );
  XOR U849 ( .A(n341), .B(n333), .Z(n353) );
  XNOR U850 ( .A(n332), .B(n328), .Z(n354) );
  XNOR U851 ( .A(n327), .B(n323), .Z(n355) );
  XNOR U852 ( .A(n322), .B(n318), .Z(n356) );
  XNOR U853 ( .A(n317), .B(n313), .Z(n357) );
  XNOR U854 ( .A(n312), .B(n308), .Z(n358) );
  XNOR U855 ( .A(n359), .B(n360), .Z(n308) );
  XNOR U856 ( .A(n307), .B(n303), .Z(n360) );
  XNOR U857 ( .A(n302), .B(n298), .Z(n361) );
  XOR U858 ( .A(n297), .B(n294), .Z(n362) );
  XOR U859 ( .A(n363), .B(n364), .Z(n294) );
  XOR U860 ( .A(n292), .B(n365), .Z(n364) );
  XOR U861 ( .A(n366), .B(n367), .Z(n365) );
  XNOR U862 ( .A(n368), .B(n369), .Z(n367) );
  AND U863 ( .A(b[13]), .B(a[45]), .Z(n368) );
  XOR U864 ( .A(n370), .B(n371), .Z(n366) );
  AND U865 ( .A(b[14]), .B(a[44]), .Z(n371) );
  AND U866 ( .A(b[15]), .B(a[43]), .Z(n370) );
  XOR U867 ( .A(n372), .B(n369), .Z(n363) );
  XOR U868 ( .A(n373), .B(n374), .Z(n369) );
  NOR U869 ( .A(n375), .B(n376), .Z(n373) );
  AND U870 ( .A(b[12]), .B(a[46]), .Z(n372) );
  XNOR U871 ( .A(n377), .B(n292), .Z(n293) );
  XOR U872 ( .A(n378), .B(n379), .Z(n292) );
  ANDN U873 ( .B(n380), .A(n381), .Z(n378) );
  AND U874 ( .A(b[11]), .B(a[47]), .Z(n377) );
  XNOR U875 ( .A(n382), .B(n297), .Z(n299) );
  XOR U876 ( .A(n383), .B(n384), .Z(n297) );
  ANDN U877 ( .B(n385), .A(n386), .Z(n383) );
  AND U878 ( .A(a[48]), .B(b[10]), .Z(n382) );
  IV U879 ( .A(n304), .Z(n359) );
  XNOR U880 ( .A(n387), .B(n302), .Z(n304) );
  XOR U881 ( .A(n388), .B(n389), .Z(n302) );
  ANDN U882 ( .B(n390), .A(n391), .Z(n388) );
  AND U883 ( .A(a[49]), .B(b[9]), .Z(n387) );
  XNOR U884 ( .A(n392), .B(n307), .Z(n309) );
  XOR U885 ( .A(n393), .B(n394), .Z(n307) );
  ANDN U886 ( .B(n395), .A(n396), .Z(n393) );
  AND U887 ( .A(b[8]), .B(a[50]), .Z(n392) );
  XNOR U888 ( .A(n397), .B(n312), .Z(n314) );
  XOR U889 ( .A(n398), .B(n399), .Z(n312) );
  ANDN U890 ( .B(n400), .A(n401), .Z(n398) );
  AND U891 ( .A(b[7]), .B(a[51]), .Z(n397) );
  XNOR U892 ( .A(n402), .B(n317), .Z(n319) );
  XOR U893 ( .A(n403), .B(n404), .Z(n317) );
  ANDN U894 ( .B(n405), .A(n406), .Z(n403) );
  AND U895 ( .A(b[6]), .B(a[52]), .Z(n402) );
  XNOR U896 ( .A(n407), .B(n322), .Z(n324) );
  XOR U897 ( .A(n408), .B(n409), .Z(n322) );
  ANDN U898 ( .B(n410), .A(n411), .Z(n408) );
  AND U899 ( .A(b[5]), .B(a[53]), .Z(n407) );
  XNOR U900 ( .A(n412), .B(n327), .Z(n329) );
  XOR U901 ( .A(n413), .B(n414), .Z(n327) );
  ANDN U902 ( .B(n415), .A(n416), .Z(n413) );
  AND U903 ( .A(b[4]), .B(a[54]), .Z(n412) );
  XNOR U904 ( .A(n417), .B(n418), .Z(n341) );
  NANDN U905 ( .A(n419), .B(n420), .Z(n418) );
  XNOR U906 ( .A(n421), .B(n332), .Z(n334) );
  XNOR U907 ( .A(n422), .B(n423), .Z(n332) );
  AND U908 ( .A(n424), .B(n425), .Z(n422) );
  AND U909 ( .A(a[55]), .B(b[3]), .Z(n421) );
  XNOR U910 ( .A(n426), .B(n427), .Z(swire[57]) );
  XOR U911 ( .A(n352), .B(n428), .Z(n427) );
  XOR U912 ( .A(n351), .B(n426), .Z(n428) );
  NAND U913 ( .A(a[57]), .B(b[0]), .Z(n351) );
  XNOR U914 ( .A(n419), .B(n420), .Z(n352) );
  XOR U915 ( .A(n417), .B(n429), .Z(n420) );
  NAND U916 ( .A(b[1]), .B(a[56]), .Z(n429) );
  XOR U917 ( .A(n425), .B(n430), .Z(n419) );
  XOR U918 ( .A(n417), .B(n424), .Z(n430) );
  XNOR U919 ( .A(n431), .B(n423), .Z(n424) );
  AND U920 ( .A(b[2]), .B(a[55]), .Z(n431) );
  NANDN U921 ( .A(n432), .B(n433), .Z(n417) );
  XOR U922 ( .A(n423), .B(n415), .Z(n434) );
  XNOR U923 ( .A(n414), .B(n410), .Z(n435) );
  XNOR U924 ( .A(n409), .B(n405), .Z(n436) );
  XNOR U925 ( .A(n404), .B(n400), .Z(n437) );
  XNOR U926 ( .A(n399), .B(n395), .Z(n438) );
  XNOR U927 ( .A(n394), .B(n390), .Z(n439) );
  XNOR U928 ( .A(n389), .B(n385), .Z(n440) );
  XNOR U929 ( .A(n384), .B(n380), .Z(n441) );
  XOR U930 ( .A(n379), .B(n376), .Z(n442) );
  XOR U931 ( .A(n443), .B(n444), .Z(n376) );
  XOR U932 ( .A(n374), .B(n445), .Z(n444) );
  XOR U933 ( .A(n446), .B(n447), .Z(n445) );
  XNOR U934 ( .A(n448), .B(n449), .Z(n447) );
  AND U935 ( .A(b[13]), .B(a[44]), .Z(n448) );
  XOR U936 ( .A(n450), .B(n451), .Z(n446) );
  AND U937 ( .A(b[14]), .B(a[43]), .Z(n451) );
  AND U938 ( .A(b[15]), .B(a[42]), .Z(n450) );
  XOR U939 ( .A(n452), .B(n449), .Z(n443) );
  XOR U940 ( .A(n453), .B(n454), .Z(n449) );
  NOR U941 ( .A(n455), .B(n456), .Z(n453) );
  AND U942 ( .A(b[12]), .B(a[45]), .Z(n452) );
  XNOR U943 ( .A(n457), .B(n374), .Z(n375) );
  XOR U944 ( .A(n458), .B(n459), .Z(n374) );
  ANDN U945 ( .B(n460), .A(n461), .Z(n458) );
  AND U946 ( .A(b[11]), .B(a[46]), .Z(n457) );
  XNOR U947 ( .A(n462), .B(n379), .Z(n381) );
  XOR U948 ( .A(n463), .B(n464), .Z(n379) );
  ANDN U949 ( .B(n465), .A(n466), .Z(n463) );
  AND U950 ( .A(b[10]), .B(a[47]), .Z(n462) );
  XNOR U951 ( .A(n467), .B(n384), .Z(n386) );
  XOR U952 ( .A(n468), .B(n469), .Z(n384) );
  ANDN U953 ( .B(n470), .A(n471), .Z(n468) );
  AND U954 ( .A(a[48]), .B(b[9]), .Z(n467) );
  XNOR U955 ( .A(n472), .B(n389), .Z(n391) );
  XOR U956 ( .A(n473), .B(n474), .Z(n389) );
  ANDN U957 ( .B(n475), .A(n476), .Z(n473) );
  AND U958 ( .A(b[8]), .B(a[49]), .Z(n472) );
  XNOR U959 ( .A(n477), .B(n394), .Z(n396) );
  XOR U960 ( .A(n478), .B(n479), .Z(n394) );
  ANDN U961 ( .B(n480), .A(n481), .Z(n478) );
  AND U962 ( .A(b[7]), .B(a[50]), .Z(n477) );
  XNOR U963 ( .A(n482), .B(n399), .Z(n401) );
  XOR U964 ( .A(n483), .B(n484), .Z(n399) );
  ANDN U965 ( .B(n485), .A(n486), .Z(n483) );
  AND U966 ( .A(b[6]), .B(a[51]), .Z(n482) );
  XNOR U967 ( .A(n487), .B(n404), .Z(n406) );
  XOR U968 ( .A(n488), .B(n489), .Z(n404) );
  ANDN U969 ( .B(n490), .A(n491), .Z(n488) );
  AND U970 ( .A(b[5]), .B(a[52]), .Z(n487) );
  XNOR U971 ( .A(n492), .B(n409), .Z(n411) );
  XOR U972 ( .A(n493), .B(n494), .Z(n409) );
  ANDN U973 ( .B(n495), .A(n496), .Z(n493) );
  AND U974 ( .A(b[4]), .B(a[53]), .Z(n492) );
  XNOR U975 ( .A(n497), .B(n498), .Z(n423) );
  NANDN U976 ( .A(n499), .B(n500), .Z(n498) );
  XNOR U977 ( .A(n501), .B(n414), .Z(n416) );
  XNOR U978 ( .A(n502), .B(n503), .Z(n414) );
  AND U979 ( .A(n504), .B(n505), .Z(n502) );
  AND U980 ( .A(a[54]), .B(b[3]), .Z(n501) );
  XNOR U981 ( .A(n506), .B(n507), .Z(swire[56]) );
  XOR U982 ( .A(n433), .B(n509), .Z(n507) );
  XNOR U983 ( .A(n432), .B(n508), .Z(n509) );
  IV U984 ( .A(n506), .Z(n508) );
  NAND U985 ( .A(a[56]), .B(b[0]), .Z(n432) );
  XNOR U986 ( .A(n499), .B(n500), .Z(n433) );
  XOR U987 ( .A(n497), .B(n510), .Z(n500) );
  NAND U988 ( .A(b[1]), .B(a[55]), .Z(n510) );
  XOR U989 ( .A(n504), .B(n511), .Z(n499) );
  XOR U990 ( .A(n497), .B(n505), .Z(n511) );
  XNOR U991 ( .A(n512), .B(n503), .Z(n505) );
  AND U992 ( .A(b[2]), .B(a[54]), .Z(n512) );
  NANDN U993 ( .A(n513), .B(n514), .Z(n497) );
  XOR U994 ( .A(n503), .B(n495), .Z(n515) );
  XNOR U995 ( .A(n494), .B(n490), .Z(n516) );
  XNOR U996 ( .A(n489), .B(n485), .Z(n517) );
  XNOR U997 ( .A(n484), .B(n480), .Z(n518) );
  XNOR U998 ( .A(n479), .B(n475), .Z(n519) );
  XNOR U999 ( .A(n474), .B(n470), .Z(n520) );
  XNOR U1000 ( .A(n469), .B(n465), .Z(n521) );
  XNOR U1001 ( .A(n464), .B(n460), .Z(n522) );
  XOR U1002 ( .A(n459), .B(n456), .Z(n523) );
  XOR U1003 ( .A(n524), .B(n525), .Z(n456) );
  XOR U1004 ( .A(n454), .B(n526), .Z(n525) );
  XOR U1005 ( .A(n527), .B(n528), .Z(n526) );
  XOR U1006 ( .A(n529), .B(n530), .Z(n528) );
  XOR U1007 ( .A(n531), .B(n532), .Z(n530) );
  XOR U1008 ( .A(n533), .B(n534), .Z(n532) );
  NAND U1009 ( .A(b[14]), .B(a[42]), .Z(n534) );
  AND U1010 ( .A(b[15]), .B(a[41]), .Z(n533) );
  XOR U1011 ( .A(n535), .B(n531), .Z(n527) );
  XOR U1012 ( .A(n536), .B(n537), .Z(n531) );
  NOR U1013 ( .A(n538), .B(n539), .Z(n536) );
  AND U1014 ( .A(b[13]), .B(a[43]), .Z(n535) );
  XOR U1015 ( .A(n540), .B(n529), .Z(n524) );
  XOR U1016 ( .A(n541), .B(n542), .Z(n529) );
  ANDN U1017 ( .B(n543), .A(n544), .Z(n541) );
  AND U1018 ( .A(b[12]), .B(a[44]), .Z(n540) );
  XNOR U1019 ( .A(n545), .B(n454), .Z(n455) );
  XOR U1020 ( .A(n546), .B(n547), .Z(n454) );
  ANDN U1021 ( .B(n548), .A(n549), .Z(n546) );
  AND U1022 ( .A(b[11]), .B(a[45]), .Z(n545) );
  XNOR U1023 ( .A(n550), .B(n459), .Z(n461) );
  XOR U1024 ( .A(n551), .B(n552), .Z(n459) );
  ANDN U1025 ( .B(n553), .A(n554), .Z(n551) );
  AND U1026 ( .A(b[10]), .B(a[46]), .Z(n550) );
  XNOR U1027 ( .A(n555), .B(n464), .Z(n466) );
  XOR U1028 ( .A(n556), .B(n557), .Z(n464) );
  ANDN U1029 ( .B(n558), .A(n559), .Z(n556) );
  AND U1030 ( .A(b[9]), .B(a[47]), .Z(n555) );
  XNOR U1031 ( .A(n560), .B(n469), .Z(n471) );
  XOR U1032 ( .A(n561), .B(n562), .Z(n469) );
  ANDN U1033 ( .B(n563), .A(n564), .Z(n561) );
  AND U1034 ( .A(b[8]), .B(a[48]), .Z(n560) );
  XNOR U1035 ( .A(n565), .B(n474), .Z(n476) );
  XOR U1036 ( .A(n566), .B(n567), .Z(n474) );
  ANDN U1037 ( .B(n568), .A(n569), .Z(n566) );
  AND U1038 ( .A(b[7]), .B(a[49]), .Z(n565) );
  XNOR U1039 ( .A(n570), .B(n479), .Z(n481) );
  XOR U1040 ( .A(n571), .B(n572), .Z(n479) );
  ANDN U1041 ( .B(n573), .A(n574), .Z(n571) );
  AND U1042 ( .A(b[6]), .B(a[50]), .Z(n570) );
  XNOR U1043 ( .A(n575), .B(n484), .Z(n486) );
  XOR U1044 ( .A(n576), .B(n577), .Z(n484) );
  ANDN U1045 ( .B(n578), .A(n579), .Z(n576) );
  AND U1046 ( .A(b[5]), .B(a[51]), .Z(n575) );
  XNOR U1047 ( .A(n580), .B(n489), .Z(n491) );
  XOR U1048 ( .A(n581), .B(n582), .Z(n489) );
  ANDN U1049 ( .B(n583), .A(n584), .Z(n581) );
  AND U1050 ( .A(b[4]), .B(a[52]), .Z(n580) );
  XNOR U1051 ( .A(n585), .B(n586), .Z(n503) );
  NANDN U1052 ( .A(n587), .B(n588), .Z(n586) );
  XNOR U1053 ( .A(n589), .B(n494), .Z(n496) );
  XNOR U1054 ( .A(n590), .B(n591), .Z(n494) );
  NOR U1055 ( .A(n592), .B(n593), .Z(n590) );
  AND U1056 ( .A(a[53]), .B(b[3]), .Z(n589) );
  XNOR U1057 ( .A(n594), .B(n595), .Z(swire[55]) );
  XOR U1058 ( .A(n514), .B(n596), .Z(n595) );
  XOR U1059 ( .A(n513), .B(n594), .Z(n596) );
  NAND U1060 ( .A(a[55]), .B(b[0]), .Z(n513) );
  XOR U1061 ( .A(n597), .B(n598), .Z(n587) );
  NAND U1062 ( .A(b[1]), .B(a[54]), .Z(n598) );
  XOR U1063 ( .A(n597), .B(n593), .Z(n599) );
  XOR U1064 ( .A(n600), .B(n591), .Z(n593) );
  AND U1065 ( .A(b[2]), .B(a[53]), .Z(n600) );
  IV U1066 ( .A(n585), .Z(n597) );
  NANDN U1067 ( .A(n601), .B(n602), .Z(n585) );
  XOR U1068 ( .A(n591), .B(n583), .Z(n603) );
  XNOR U1069 ( .A(n582), .B(n578), .Z(n604) );
  XNOR U1070 ( .A(n577), .B(n573), .Z(n605) );
  XNOR U1071 ( .A(n572), .B(n568), .Z(n606) );
  XNOR U1072 ( .A(n567), .B(n563), .Z(n607) );
  XNOR U1073 ( .A(n562), .B(n558), .Z(n608) );
  XNOR U1074 ( .A(n557), .B(n553), .Z(n609) );
  XNOR U1075 ( .A(n552), .B(n548), .Z(n610) );
  XNOR U1076 ( .A(n547), .B(n543), .Z(n611) );
  XOR U1077 ( .A(n542), .B(n539), .Z(n612) );
  XOR U1078 ( .A(n613), .B(n614), .Z(n539) );
  XOR U1079 ( .A(n537), .B(n615), .Z(n614) );
  XOR U1080 ( .A(n616), .B(n617), .Z(n615) );
  XOR U1081 ( .A(n618), .B(n619), .Z(n617) );
  NAND U1082 ( .A(b[14]), .B(a[41]), .Z(n619) );
  AND U1083 ( .A(b[15]), .B(a[40]), .Z(n618) );
  XOR U1084 ( .A(n620), .B(n616), .Z(n613) );
  XOR U1085 ( .A(n621), .B(n622), .Z(n616) );
  NOR U1086 ( .A(n623), .B(n624), .Z(n621) );
  AND U1087 ( .A(b[13]), .B(a[42]), .Z(n620) );
  XNOR U1088 ( .A(n625), .B(n537), .Z(n538) );
  XOR U1089 ( .A(n626), .B(n627), .Z(n537) );
  ANDN U1090 ( .B(n628), .A(n629), .Z(n626) );
  AND U1091 ( .A(b[12]), .B(a[43]), .Z(n625) );
  XNOR U1092 ( .A(n630), .B(n542), .Z(n544) );
  XOR U1093 ( .A(n631), .B(n632), .Z(n542) );
  ANDN U1094 ( .B(n633), .A(n634), .Z(n631) );
  AND U1095 ( .A(b[11]), .B(a[44]), .Z(n630) );
  XNOR U1096 ( .A(n635), .B(n547), .Z(n549) );
  XOR U1097 ( .A(n636), .B(n637), .Z(n547) );
  ANDN U1098 ( .B(n638), .A(n639), .Z(n636) );
  AND U1099 ( .A(b[10]), .B(a[45]), .Z(n635) );
  XNOR U1100 ( .A(n640), .B(n552), .Z(n554) );
  XOR U1101 ( .A(n641), .B(n642), .Z(n552) );
  ANDN U1102 ( .B(n643), .A(n644), .Z(n641) );
  AND U1103 ( .A(b[9]), .B(a[46]), .Z(n640) );
  XNOR U1104 ( .A(n645), .B(n557), .Z(n559) );
  XOR U1105 ( .A(n646), .B(n647), .Z(n557) );
  ANDN U1106 ( .B(n648), .A(n649), .Z(n646) );
  AND U1107 ( .A(b[8]), .B(a[47]), .Z(n645) );
  XNOR U1108 ( .A(n650), .B(n562), .Z(n564) );
  XOR U1109 ( .A(n651), .B(n652), .Z(n562) );
  ANDN U1110 ( .B(n653), .A(n654), .Z(n651) );
  AND U1111 ( .A(b[7]), .B(a[48]), .Z(n650) );
  XNOR U1112 ( .A(n655), .B(n567), .Z(n569) );
  XOR U1113 ( .A(n656), .B(n657), .Z(n567) );
  ANDN U1114 ( .B(n658), .A(n659), .Z(n656) );
  AND U1115 ( .A(b[6]), .B(a[49]), .Z(n655) );
  XNOR U1116 ( .A(n660), .B(n572), .Z(n574) );
  XOR U1117 ( .A(n661), .B(n662), .Z(n572) );
  ANDN U1118 ( .B(n663), .A(n664), .Z(n661) );
  AND U1119 ( .A(b[5]), .B(a[50]), .Z(n660) );
  XNOR U1120 ( .A(n665), .B(n577), .Z(n579) );
  XOR U1121 ( .A(n666), .B(n667), .Z(n577) );
  ANDN U1122 ( .B(n668), .A(n669), .Z(n666) );
  AND U1123 ( .A(b[4]), .B(a[51]), .Z(n665) );
  XOR U1124 ( .A(n670), .B(n671), .Z(n591) );
  NANDN U1125 ( .A(n672), .B(n673), .Z(n671) );
  XNOR U1126 ( .A(n674), .B(n582), .Z(n584) );
  XNOR U1127 ( .A(n675), .B(n676), .Z(n582) );
  AND U1128 ( .A(n677), .B(n678), .Z(n675) );
  AND U1129 ( .A(a[52]), .B(b[3]), .Z(n674) );
  XNOR U1130 ( .A(n679), .B(n680), .Z(swire[54]) );
  XOR U1131 ( .A(n602), .B(n682), .Z(n680) );
  XNOR U1132 ( .A(n601), .B(n681), .Z(n682) );
  IV U1133 ( .A(n679), .Z(n681) );
  NAND U1134 ( .A(a[54]), .B(b[0]), .Z(n601) );
  XNOR U1135 ( .A(n673), .B(n672), .Z(n602) );
  XOR U1136 ( .A(n670), .B(n683), .Z(n672) );
  NAND U1137 ( .A(b[1]), .B(a[53]), .Z(n683) );
  XNOR U1138 ( .A(n678), .B(n684), .Z(n673) );
  XNOR U1139 ( .A(n670), .B(n677), .Z(n684) );
  XNOR U1140 ( .A(n685), .B(n676), .Z(n677) );
  AND U1141 ( .A(b[2]), .B(a[52]), .Z(n685) );
  ANDN U1142 ( .B(n686), .A(n687), .Z(n670) );
  XOR U1143 ( .A(n676), .B(n668), .Z(n688) );
  XNOR U1144 ( .A(n667), .B(n663), .Z(n689) );
  XNOR U1145 ( .A(n662), .B(n658), .Z(n690) );
  XNOR U1146 ( .A(n657), .B(n653), .Z(n691) );
  XNOR U1147 ( .A(n652), .B(n648), .Z(n692) );
  XNOR U1148 ( .A(n647), .B(n643), .Z(n693) );
  XNOR U1149 ( .A(n642), .B(n638), .Z(n694) );
  XNOR U1150 ( .A(n637), .B(n633), .Z(n695) );
  XNOR U1151 ( .A(n632), .B(n628), .Z(n696) );
  XOR U1152 ( .A(n627), .B(n624), .Z(n697) );
  XOR U1153 ( .A(n698), .B(n699), .Z(n624) );
  XOR U1154 ( .A(n622), .B(n700), .Z(n699) );
  XOR U1155 ( .A(n701), .B(n702), .Z(n700) );
  XOR U1156 ( .A(n703), .B(n704), .Z(n702) );
  NAND U1157 ( .A(b[14]), .B(a[40]), .Z(n704) );
  AND U1158 ( .A(b[15]), .B(a[39]), .Z(n703) );
  XOR U1159 ( .A(n705), .B(n701), .Z(n698) );
  XOR U1160 ( .A(n706), .B(n707), .Z(n701) );
  NOR U1161 ( .A(n708), .B(n709), .Z(n706) );
  AND U1162 ( .A(b[13]), .B(a[41]), .Z(n705) );
  XNOR U1163 ( .A(n710), .B(n622), .Z(n623) );
  XOR U1164 ( .A(n711), .B(n712), .Z(n622) );
  ANDN U1165 ( .B(n713), .A(n714), .Z(n711) );
  AND U1166 ( .A(b[12]), .B(a[42]), .Z(n710) );
  XNOR U1167 ( .A(n715), .B(n627), .Z(n629) );
  XOR U1168 ( .A(n716), .B(n717), .Z(n627) );
  ANDN U1169 ( .B(n718), .A(n719), .Z(n716) );
  AND U1170 ( .A(b[11]), .B(a[43]), .Z(n715) );
  XNOR U1171 ( .A(n720), .B(n632), .Z(n634) );
  XOR U1172 ( .A(n721), .B(n722), .Z(n632) );
  ANDN U1173 ( .B(n723), .A(n724), .Z(n721) );
  AND U1174 ( .A(b[10]), .B(a[44]), .Z(n720) );
  XNOR U1175 ( .A(n725), .B(n637), .Z(n639) );
  XOR U1176 ( .A(n726), .B(n727), .Z(n637) );
  ANDN U1177 ( .B(n728), .A(n729), .Z(n726) );
  AND U1178 ( .A(b[9]), .B(a[45]), .Z(n725) );
  XNOR U1179 ( .A(n730), .B(n642), .Z(n644) );
  XOR U1180 ( .A(n731), .B(n732), .Z(n642) );
  ANDN U1181 ( .B(n733), .A(n734), .Z(n731) );
  AND U1182 ( .A(b[8]), .B(a[46]), .Z(n730) );
  XNOR U1183 ( .A(n735), .B(n647), .Z(n649) );
  XOR U1184 ( .A(n736), .B(n737), .Z(n647) );
  ANDN U1185 ( .B(n738), .A(n739), .Z(n736) );
  AND U1186 ( .A(b[7]), .B(a[47]), .Z(n735) );
  XNOR U1187 ( .A(n740), .B(n652), .Z(n654) );
  XOR U1188 ( .A(n741), .B(n742), .Z(n652) );
  ANDN U1189 ( .B(n743), .A(n744), .Z(n741) );
  AND U1190 ( .A(b[6]), .B(a[48]), .Z(n740) );
  XNOR U1191 ( .A(n745), .B(n657), .Z(n659) );
  XOR U1192 ( .A(n746), .B(n747), .Z(n657) );
  ANDN U1193 ( .B(n748), .A(n749), .Z(n746) );
  AND U1194 ( .A(b[5]), .B(a[49]), .Z(n745) );
  XNOR U1195 ( .A(n750), .B(n662), .Z(n664) );
  XOR U1196 ( .A(n751), .B(n752), .Z(n662) );
  ANDN U1197 ( .B(n753), .A(n754), .Z(n751) );
  AND U1198 ( .A(b[4]), .B(a[50]), .Z(n750) );
  XNOR U1199 ( .A(n755), .B(n756), .Z(n676) );
  NANDN U1200 ( .A(n757), .B(n758), .Z(n756) );
  XNOR U1201 ( .A(n759), .B(n667), .Z(n669) );
  XNOR U1202 ( .A(n760), .B(n761), .Z(n667) );
  AND U1203 ( .A(n762), .B(n763), .Z(n760) );
  AND U1204 ( .A(a[51]), .B(b[3]), .Z(n759) );
  XNOR U1205 ( .A(n764), .B(n765), .Z(swire[53]) );
  XOR U1206 ( .A(n686), .B(n766), .Z(n765) );
  XOR U1207 ( .A(n687), .B(n764), .Z(n766) );
  NAND U1208 ( .A(a[53]), .B(b[0]), .Z(n687) );
  XNOR U1209 ( .A(n757), .B(n758), .Z(n686) );
  XOR U1210 ( .A(n755), .B(n767), .Z(n758) );
  NAND U1211 ( .A(b[1]), .B(a[52]), .Z(n767) );
  XOR U1212 ( .A(n763), .B(n768), .Z(n757) );
  XOR U1213 ( .A(n755), .B(n762), .Z(n768) );
  XNOR U1214 ( .A(n769), .B(n761), .Z(n762) );
  AND U1215 ( .A(b[2]), .B(a[51]), .Z(n769) );
  NANDN U1216 ( .A(n770), .B(n771), .Z(n755) );
  XOR U1217 ( .A(n761), .B(n753), .Z(n772) );
  XNOR U1218 ( .A(n752), .B(n748), .Z(n773) );
  XNOR U1219 ( .A(n747), .B(n743), .Z(n774) );
  XNOR U1220 ( .A(n742), .B(n738), .Z(n775) );
  XNOR U1221 ( .A(n737), .B(n733), .Z(n776) );
  XNOR U1222 ( .A(n732), .B(n728), .Z(n777) );
  XNOR U1223 ( .A(n727), .B(n723), .Z(n778) );
  XNOR U1224 ( .A(n722), .B(n718), .Z(n779) );
  XNOR U1225 ( .A(n717), .B(n713), .Z(n780) );
  XOR U1226 ( .A(n712), .B(n709), .Z(n781) );
  XOR U1227 ( .A(n782), .B(n783), .Z(n709) );
  XOR U1228 ( .A(n707), .B(n784), .Z(n783) );
  XOR U1229 ( .A(n785), .B(n786), .Z(n784) );
  XOR U1230 ( .A(n787), .B(n788), .Z(n786) );
  NAND U1231 ( .A(b[14]), .B(a[39]), .Z(n788) );
  AND U1232 ( .A(b[15]), .B(a[38]), .Z(n787) );
  XOR U1233 ( .A(n789), .B(n785), .Z(n782) );
  XOR U1234 ( .A(n790), .B(n791), .Z(n785) );
  NOR U1235 ( .A(n792), .B(n793), .Z(n790) );
  AND U1236 ( .A(b[13]), .B(a[40]), .Z(n789) );
  XNOR U1237 ( .A(n794), .B(n707), .Z(n708) );
  XOR U1238 ( .A(n795), .B(n796), .Z(n707) );
  ANDN U1239 ( .B(n797), .A(n798), .Z(n795) );
  AND U1240 ( .A(b[12]), .B(a[41]), .Z(n794) );
  XNOR U1241 ( .A(n799), .B(n712), .Z(n714) );
  XOR U1242 ( .A(n800), .B(n801), .Z(n712) );
  ANDN U1243 ( .B(n802), .A(n803), .Z(n800) );
  AND U1244 ( .A(b[11]), .B(a[42]), .Z(n799) );
  XNOR U1245 ( .A(n804), .B(n717), .Z(n719) );
  XOR U1246 ( .A(n805), .B(n806), .Z(n717) );
  ANDN U1247 ( .B(n807), .A(n808), .Z(n805) );
  AND U1248 ( .A(b[10]), .B(a[43]), .Z(n804) );
  XNOR U1249 ( .A(n809), .B(n722), .Z(n724) );
  XOR U1250 ( .A(n810), .B(n811), .Z(n722) );
  ANDN U1251 ( .B(n812), .A(n813), .Z(n810) );
  AND U1252 ( .A(b[9]), .B(a[44]), .Z(n809) );
  XNOR U1253 ( .A(n814), .B(n727), .Z(n729) );
  XOR U1254 ( .A(n815), .B(n816), .Z(n727) );
  ANDN U1255 ( .B(n817), .A(n818), .Z(n815) );
  AND U1256 ( .A(b[8]), .B(a[45]), .Z(n814) );
  XNOR U1257 ( .A(n819), .B(n732), .Z(n734) );
  XOR U1258 ( .A(n820), .B(n821), .Z(n732) );
  ANDN U1259 ( .B(n822), .A(n823), .Z(n820) );
  AND U1260 ( .A(b[7]), .B(a[46]), .Z(n819) );
  XNOR U1261 ( .A(n824), .B(n737), .Z(n739) );
  XOR U1262 ( .A(n825), .B(n826), .Z(n737) );
  ANDN U1263 ( .B(n827), .A(n828), .Z(n825) );
  AND U1264 ( .A(b[6]), .B(a[47]), .Z(n824) );
  XNOR U1265 ( .A(n829), .B(n742), .Z(n744) );
  XOR U1266 ( .A(n830), .B(n831), .Z(n742) );
  ANDN U1267 ( .B(n832), .A(n833), .Z(n830) );
  AND U1268 ( .A(b[5]), .B(a[48]), .Z(n829) );
  XNOR U1269 ( .A(n834), .B(n747), .Z(n749) );
  XOR U1270 ( .A(n835), .B(n836), .Z(n747) );
  ANDN U1271 ( .B(n837), .A(n838), .Z(n835) );
  AND U1272 ( .A(b[4]), .B(a[49]), .Z(n834) );
  XNOR U1273 ( .A(n839), .B(n840), .Z(n761) );
  NANDN U1274 ( .A(n841), .B(n842), .Z(n840) );
  XNOR U1275 ( .A(n843), .B(n752), .Z(n754) );
  XNOR U1276 ( .A(n844), .B(n845), .Z(n752) );
  AND U1277 ( .A(n846), .B(n847), .Z(n844) );
  AND U1278 ( .A(a[50]), .B(b[3]), .Z(n843) );
  XNOR U1279 ( .A(n848), .B(n849), .Z(swire[52]) );
  XOR U1280 ( .A(n771), .B(n851), .Z(n849) );
  XNOR U1281 ( .A(n770), .B(n850), .Z(n851) );
  IV U1282 ( .A(n848), .Z(n850) );
  NAND U1283 ( .A(a[52]), .B(b[0]), .Z(n770) );
  XNOR U1284 ( .A(n841), .B(n842), .Z(n771) );
  XOR U1285 ( .A(n839), .B(n852), .Z(n842) );
  NAND U1286 ( .A(b[1]), .B(a[51]), .Z(n852) );
  XOR U1287 ( .A(n847), .B(n853), .Z(n841) );
  XOR U1288 ( .A(n839), .B(n846), .Z(n853) );
  XNOR U1289 ( .A(n854), .B(n845), .Z(n846) );
  AND U1290 ( .A(b[2]), .B(a[50]), .Z(n854) );
  NANDN U1291 ( .A(n855), .B(n856), .Z(n839) );
  XOR U1292 ( .A(n845), .B(n837), .Z(n857) );
  XNOR U1293 ( .A(n836), .B(n832), .Z(n858) );
  XNOR U1294 ( .A(n831), .B(n827), .Z(n859) );
  XNOR U1295 ( .A(n826), .B(n822), .Z(n860) );
  XNOR U1296 ( .A(n821), .B(n817), .Z(n861) );
  XNOR U1297 ( .A(n816), .B(n812), .Z(n862) );
  XNOR U1298 ( .A(n811), .B(n807), .Z(n863) );
  XNOR U1299 ( .A(n806), .B(n802), .Z(n864) );
  XNOR U1300 ( .A(n801), .B(n797), .Z(n865) );
  XOR U1301 ( .A(n796), .B(n793), .Z(n866) );
  XOR U1302 ( .A(n867), .B(n868), .Z(n793) );
  XOR U1303 ( .A(n791), .B(n869), .Z(n868) );
  XOR U1304 ( .A(n870), .B(n871), .Z(n869) );
  XOR U1305 ( .A(n872), .B(n873), .Z(n871) );
  NAND U1306 ( .A(b[14]), .B(a[38]), .Z(n873) );
  AND U1307 ( .A(b[15]), .B(a[37]), .Z(n872) );
  XOR U1308 ( .A(n874), .B(n870), .Z(n867) );
  XOR U1309 ( .A(n875), .B(n876), .Z(n870) );
  NOR U1310 ( .A(n877), .B(n878), .Z(n875) );
  AND U1311 ( .A(b[13]), .B(a[39]), .Z(n874) );
  XNOR U1312 ( .A(n879), .B(n791), .Z(n792) );
  XOR U1313 ( .A(n880), .B(n881), .Z(n791) );
  ANDN U1314 ( .B(n882), .A(n883), .Z(n880) );
  AND U1315 ( .A(b[12]), .B(a[40]), .Z(n879) );
  XNOR U1316 ( .A(n884), .B(n796), .Z(n798) );
  XOR U1317 ( .A(n885), .B(n886), .Z(n796) );
  ANDN U1318 ( .B(n887), .A(n888), .Z(n885) );
  AND U1319 ( .A(b[11]), .B(a[41]), .Z(n884) );
  XNOR U1320 ( .A(n889), .B(n801), .Z(n803) );
  XOR U1321 ( .A(n890), .B(n891), .Z(n801) );
  ANDN U1322 ( .B(n892), .A(n893), .Z(n890) );
  AND U1323 ( .A(b[10]), .B(a[42]), .Z(n889) );
  XNOR U1324 ( .A(n894), .B(n806), .Z(n808) );
  XOR U1325 ( .A(n895), .B(n896), .Z(n806) );
  ANDN U1326 ( .B(n897), .A(n898), .Z(n895) );
  AND U1327 ( .A(b[9]), .B(a[43]), .Z(n894) );
  XNOR U1328 ( .A(n899), .B(n811), .Z(n813) );
  XOR U1329 ( .A(n900), .B(n901), .Z(n811) );
  ANDN U1330 ( .B(n902), .A(n903), .Z(n900) );
  AND U1331 ( .A(b[8]), .B(a[44]), .Z(n899) );
  XNOR U1332 ( .A(n904), .B(n816), .Z(n818) );
  XOR U1333 ( .A(n905), .B(n906), .Z(n816) );
  ANDN U1334 ( .B(n907), .A(n908), .Z(n905) );
  AND U1335 ( .A(b[7]), .B(a[45]), .Z(n904) );
  XNOR U1336 ( .A(n909), .B(n821), .Z(n823) );
  XOR U1337 ( .A(n910), .B(n911), .Z(n821) );
  ANDN U1338 ( .B(n912), .A(n913), .Z(n910) );
  AND U1339 ( .A(b[6]), .B(a[46]), .Z(n909) );
  XNOR U1340 ( .A(n914), .B(n826), .Z(n828) );
  XOR U1341 ( .A(n915), .B(n916), .Z(n826) );
  ANDN U1342 ( .B(n917), .A(n918), .Z(n915) );
  AND U1343 ( .A(b[5]), .B(a[47]), .Z(n914) );
  XNOR U1344 ( .A(n919), .B(n831), .Z(n833) );
  XOR U1345 ( .A(n920), .B(n921), .Z(n831) );
  ANDN U1346 ( .B(n922), .A(n923), .Z(n920) );
  AND U1347 ( .A(b[4]), .B(a[48]), .Z(n919) );
  XNOR U1348 ( .A(n924), .B(n925), .Z(n845) );
  NANDN U1349 ( .A(n926), .B(n927), .Z(n925) );
  XNOR U1350 ( .A(n928), .B(n836), .Z(n838) );
  XNOR U1351 ( .A(n929), .B(n930), .Z(n836) );
  AND U1352 ( .A(n931), .B(n932), .Z(n929) );
  AND U1353 ( .A(a[49]), .B(b[3]), .Z(n928) );
  XNOR U1354 ( .A(n933), .B(n934), .Z(swire[51]) );
  XOR U1355 ( .A(n856), .B(n935), .Z(n934) );
  XOR U1356 ( .A(n855), .B(n933), .Z(n935) );
  NAND U1357 ( .A(a[51]), .B(b[0]), .Z(n855) );
  XNOR U1358 ( .A(n926), .B(n927), .Z(n856) );
  XOR U1359 ( .A(n924), .B(n936), .Z(n927) );
  NAND U1360 ( .A(b[1]), .B(a[50]), .Z(n936) );
  XOR U1361 ( .A(n932), .B(n937), .Z(n926) );
  XOR U1362 ( .A(n924), .B(n931), .Z(n937) );
  XNOR U1363 ( .A(n938), .B(n930), .Z(n931) );
  AND U1364 ( .A(b[2]), .B(a[49]), .Z(n938) );
  NANDN U1365 ( .A(n939), .B(n940), .Z(n924) );
  XOR U1366 ( .A(n930), .B(n922), .Z(n941) );
  XNOR U1367 ( .A(n921), .B(n917), .Z(n942) );
  XNOR U1368 ( .A(n916), .B(n912), .Z(n943) );
  XNOR U1369 ( .A(n911), .B(n907), .Z(n944) );
  XNOR U1370 ( .A(n906), .B(n902), .Z(n945) );
  XNOR U1371 ( .A(n901), .B(n897), .Z(n946) );
  XNOR U1372 ( .A(n896), .B(n892), .Z(n947) );
  XNOR U1373 ( .A(n891), .B(n887), .Z(n948) );
  XNOR U1374 ( .A(n886), .B(n882), .Z(n949) );
  XOR U1375 ( .A(n881), .B(n878), .Z(n950) );
  XOR U1376 ( .A(n951), .B(n952), .Z(n878) );
  XOR U1377 ( .A(n876), .B(n953), .Z(n952) );
  XOR U1378 ( .A(n954), .B(n955), .Z(n953) );
  XOR U1379 ( .A(n956), .B(n957), .Z(n955) );
  NAND U1380 ( .A(b[14]), .B(a[37]), .Z(n957) );
  AND U1381 ( .A(b[15]), .B(a[36]), .Z(n956) );
  XOR U1382 ( .A(n958), .B(n954), .Z(n951) );
  XOR U1383 ( .A(n959), .B(n960), .Z(n954) );
  NOR U1384 ( .A(n961), .B(n962), .Z(n959) );
  AND U1385 ( .A(b[13]), .B(a[38]), .Z(n958) );
  XNOR U1386 ( .A(n963), .B(n876), .Z(n877) );
  XOR U1387 ( .A(n964), .B(n965), .Z(n876) );
  ANDN U1388 ( .B(n966), .A(n967), .Z(n964) );
  AND U1389 ( .A(b[12]), .B(a[39]), .Z(n963) );
  XNOR U1390 ( .A(n968), .B(n881), .Z(n883) );
  XOR U1391 ( .A(n969), .B(n970), .Z(n881) );
  ANDN U1392 ( .B(n971), .A(n972), .Z(n969) );
  AND U1393 ( .A(b[11]), .B(a[40]), .Z(n968) );
  XNOR U1394 ( .A(n973), .B(n886), .Z(n888) );
  XOR U1395 ( .A(n974), .B(n975), .Z(n886) );
  ANDN U1396 ( .B(n976), .A(n977), .Z(n974) );
  AND U1397 ( .A(b[10]), .B(a[41]), .Z(n973) );
  XNOR U1398 ( .A(n978), .B(n891), .Z(n893) );
  XOR U1399 ( .A(n979), .B(n980), .Z(n891) );
  ANDN U1400 ( .B(n981), .A(n982), .Z(n979) );
  AND U1401 ( .A(b[9]), .B(a[42]), .Z(n978) );
  XNOR U1402 ( .A(n983), .B(n896), .Z(n898) );
  XOR U1403 ( .A(n984), .B(n985), .Z(n896) );
  ANDN U1404 ( .B(n986), .A(n987), .Z(n984) );
  AND U1405 ( .A(b[8]), .B(a[43]), .Z(n983) );
  XNOR U1406 ( .A(n988), .B(n901), .Z(n903) );
  XOR U1407 ( .A(n989), .B(n990), .Z(n901) );
  ANDN U1408 ( .B(n991), .A(n992), .Z(n989) );
  AND U1409 ( .A(b[7]), .B(a[44]), .Z(n988) );
  XNOR U1410 ( .A(n993), .B(n906), .Z(n908) );
  XOR U1411 ( .A(n994), .B(n995), .Z(n906) );
  ANDN U1412 ( .B(n996), .A(n997), .Z(n994) );
  AND U1413 ( .A(b[6]), .B(a[45]), .Z(n993) );
  XNOR U1414 ( .A(n998), .B(n911), .Z(n913) );
  XOR U1415 ( .A(n999), .B(n1000), .Z(n911) );
  ANDN U1416 ( .B(n1001), .A(n1002), .Z(n999) );
  AND U1417 ( .A(b[5]), .B(a[46]), .Z(n998) );
  XNOR U1418 ( .A(n1003), .B(n916), .Z(n918) );
  XOR U1419 ( .A(n1004), .B(n1005), .Z(n916) );
  ANDN U1420 ( .B(n1006), .A(n1007), .Z(n1004) );
  AND U1421 ( .A(b[4]), .B(a[47]), .Z(n1003) );
  XNOR U1422 ( .A(n1008), .B(n1009), .Z(n930) );
  NANDN U1423 ( .A(n1010), .B(n1011), .Z(n1009) );
  XNOR U1424 ( .A(n1012), .B(n921), .Z(n923) );
  XNOR U1425 ( .A(n1013), .B(n1014), .Z(n921) );
  AND U1426 ( .A(n1015), .B(n1016), .Z(n1013) );
  AND U1427 ( .A(a[48]), .B(b[3]), .Z(n1012) );
  XNOR U1428 ( .A(n1017), .B(n1018), .Z(swire[50]) );
  XOR U1429 ( .A(n940), .B(n1020), .Z(n1018) );
  XNOR U1430 ( .A(n939), .B(n1019), .Z(n1020) );
  IV U1431 ( .A(n1017), .Z(n1019) );
  NAND U1432 ( .A(a[50]), .B(b[0]), .Z(n939) );
  XNOR U1433 ( .A(n1010), .B(n1011), .Z(n940) );
  XOR U1434 ( .A(n1008), .B(n1021), .Z(n1011) );
  NAND U1435 ( .A(b[1]), .B(a[49]), .Z(n1021) );
  XOR U1436 ( .A(n1016), .B(n1022), .Z(n1010) );
  XOR U1437 ( .A(n1008), .B(n1015), .Z(n1022) );
  XNOR U1438 ( .A(n1023), .B(n1014), .Z(n1015) );
  AND U1439 ( .A(b[2]), .B(a[48]), .Z(n1023) );
  NANDN U1440 ( .A(n1024), .B(n1025), .Z(n1008) );
  XOR U1441 ( .A(n1014), .B(n1006), .Z(n1026) );
  XNOR U1442 ( .A(n1005), .B(n1001), .Z(n1027) );
  XNOR U1443 ( .A(n1000), .B(n996), .Z(n1028) );
  XNOR U1444 ( .A(n995), .B(n991), .Z(n1029) );
  XNOR U1445 ( .A(n990), .B(n986), .Z(n1030) );
  XNOR U1446 ( .A(n985), .B(n981), .Z(n1031) );
  XNOR U1447 ( .A(n980), .B(n976), .Z(n1032) );
  XNOR U1448 ( .A(n975), .B(n971), .Z(n1033) );
  XNOR U1449 ( .A(n970), .B(n966), .Z(n1034) );
  XOR U1450 ( .A(n965), .B(n962), .Z(n1035) );
  XOR U1451 ( .A(n1036), .B(n1037), .Z(n962) );
  XOR U1452 ( .A(n960), .B(n1038), .Z(n1037) );
  XOR U1453 ( .A(n1039), .B(n1040), .Z(n1038) );
  XOR U1454 ( .A(n1041), .B(n1042), .Z(n1040) );
  NAND U1455 ( .A(b[14]), .B(a[36]), .Z(n1042) );
  AND U1456 ( .A(b[15]), .B(a[35]), .Z(n1041) );
  XOR U1457 ( .A(n1043), .B(n1039), .Z(n1036) );
  XOR U1458 ( .A(n1044), .B(n1045), .Z(n1039) );
  NOR U1459 ( .A(n1046), .B(n1047), .Z(n1044) );
  AND U1460 ( .A(b[13]), .B(a[37]), .Z(n1043) );
  XNOR U1461 ( .A(n1048), .B(n960), .Z(n961) );
  XOR U1462 ( .A(n1049), .B(n1050), .Z(n960) );
  ANDN U1463 ( .B(n1051), .A(n1052), .Z(n1049) );
  AND U1464 ( .A(b[12]), .B(a[38]), .Z(n1048) );
  XNOR U1465 ( .A(n1053), .B(n965), .Z(n967) );
  XOR U1466 ( .A(n1054), .B(n1055), .Z(n965) );
  ANDN U1467 ( .B(n1056), .A(n1057), .Z(n1054) );
  AND U1468 ( .A(b[11]), .B(a[39]), .Z(n1053) );
  XNOR U1469 ( .A(n1058), .B(n970), .Z(n972) );
  XOR U1470 ( .A(n1059), .B(n1060), .Z(n970) );
  ANDN U1471 ( .B(n1061), .A(n1062), .Z(n1059) );
  AND U1472 ( .A(b[10]), .B(a[40]), .Z(n1058) );
  XNOR U1473 ( .A(n1063), .B(n975), .Z(n977) );
  XOR U1474 ( .A(n1064), .B(n1065), .Z(n975) );
  ANDN U1475 ( .B(n1066), .A(n1067), .Z(n1064) );
  AND U1476 ( .A(b[9]), .B(a[41]), .Z(n1063) );
  XNOR U1477 ( .A(n1068), .B(n980), .Z(n982) );
  XOR U1478 ( .A(n1069), .B(n1070), .Z(n980) );
  ANDN U1479 ( .B(n1071), .A(n1072), .Z(n1069) );
  AND U1480 ( .A(b[8]), .B(a[42]), .Z(n1068) );
  XNOR U1481 ( .A(n1073), .B(n985), .Z(n987) );
  XOR U1482 ( .A(n1074), .B(n1075), .Z(n985) );
  ANDN U1483 ( .B(n1076), .A(n1077), .Z(n1074) );
  AND U1484 ( .A(b[7]), .B(a[43]), .Z(n1073) );
  XNOR U1485 ( .A(n1078), .B(n990), .Z(n992) );
  XOR U1486 ( .A(n1079), .B(n1080), .Z(n990) );
  ANDN U1487 ( .B(n1081), .A(n1082), .Z(n1079) );
  AND U1488 ( .A(b[6]), .B(a[44]), .Z(n1078) );
  XNOR U1489 ( .A(n1083), .B(n995), .Z(n997) );
  XOR U1490 ( .A(n1084), .B(n1085), .Z(n995) );
  ANDN U1491 ( .B(n1086), .A(n1087), .Z(n1084) );
  AND U1492 ( .A(b[5]), .B(a[45]), .Z(n1083) );
  XNOR U1493 ( .A(n1088), .B(n1000), .Z(n1002) );
  XOR U1494 ( .A(n1089), .B(n1090), .Z(n1000) );
  ANDN U1495 ( .B(n1091), .A(n1092), .Z(n1089) );
  AND U1496 ( .A(b[4]), .B(a[46]), .Z(n1088) );
  XNOR U1497 ( .A(n1093), .B(n1094), .Z(n1014) );
  NANDN U1498 ( .A(n1095), .B(n1096), .Z(n1094) );
  XNOR U1499 ( .A(n1097), .B(n1005), .Z(n1007) );
  XNOR U1500 ( .A(n1098), .B(n1099), .Z(n1005) );
  AND U1501 ( .A(n1100), .B(n1101), .Z(n1098) );
  AND U1502 ( .A(b[3]), .B(a[47]), .Z(n1097) );
  XNOR U1503 ( .A(n1102), .B(n1103), .Z(swire[49]) );
  XOR U1504 ( .A(n1025), .B(n1104), .Z(n1103) );
  XOR U1505 ( .A(n1024), .B(n1102), .Z(n1104) );
  NAND U1506 ( .A(a[49]), .B(b[0]), .Z(n1024) );
  XNOR U1507 ( .A(n1095), .B(n1096), .Z(n1025) );
  XOR U1508 ( .A(n1093), .B(n1105), .Z(n1096) );
  NAND U1509 ( .A(b[1]), .B(a[48]), .Z(n1105) );
  XOR U1510 ( .A(n1101), .B(n1106), .Z(n1095) );
  XOR U1511 ( .A(n1093), .B(n1100), .Z(n1106) );
  XNOR U1512 ( .A(n1107), .B(n1099), .Z(n1100) );
  AND U1513 ( .A(b[2]), .B(a[47]), .Z(n1107) );
  NANDN U1514 ( .A(n1108), .B(n1109), .Z(n1093) );
  XOR U1515 ( .A(n1099), .B(n1091), .Z(n1110) );
  XNOR U1516 ( .A(n1090), .B(n1086), .Z(n1111) );
  XNOR U1517 ( .A(n1085), .B(n1081), .Z(n1112) );
  XNOR U1518 ( .A(n1080), .B(n1076), .Z(n1113) );
  XNOR U1519 ( .A(n1075), .B(n1071), .Z(n1114) );
  XNOR U1520 ( .A(n1070), .B(n1066), .Z(n1115) );
  XNOR U1521 ( .A(n1065), .B(n1061), .Z(n1116) );
  XNOR U1522 ( .A(n1060), .B(n1056), .Z(n1117) );
  XNOR U1523 ( .A(n1055), .B(n1051), .Z(n1118) );
  XOR U1524 ( .A(n1050), .B(n1047), .Z(n1119) );
  XOR U1525 ( .A(n1120), .B(n1121), .Z(n1047) );
  XOR U1526 ( .A(n1045), .B(n1122), .Z(n1121) );
  XOR U1527 ( .A(n1123), .B(n1124), .Z(n1122) );
  XOR U1528 ( .A(n1125), .B(n1126), .Z(n1124) );
  NAND U1529 ( .A(b[14]), .B(a[35]), .Z(n1126) );
  AND U1530 ( .A(b[15]), .B(a[34]), .Z(n1125) );
  XOR U1531 ( .A(n1127), .B(n1123), .Z(n1120) );
  XOR U1532 ( .A(n1128), .B(n1129), .Z(n1123) );
  NOR U1533 ( .A(n1130), .B(n1131), .Z(n1128) );
  AND U1534 ( .A(b[13]), .B(a[36]), .Z(n1127) );
  XNOR U1535 ( .A(n1132), .B(n1045), .Z(n1046) );
  XOR U1536 ( .A(n1133), .B(n1134), .Z(n1045) );
  ANDN U1537 ( .B(n1135), .A(n1136), .Z(n1133) );
  AND U1538 ( .A(b[12]), .B(a[37]), .Z(n1132) );
  XNOR U1539 ( .A(n1137), .B(n1050), .Z(n1052) );
  XOR U1540 ( .A(n1138), .B(n1139), .Z(n1050) );
  ANDN U1541 ( .B(n1140), .A(n1141), .Z(n1138) );
  AND U1542 ( .A(b[11]), .B(a[38]), .Z(n1137) );
  XNOR U1543 ( .A(n1142), .B(n1055), .Z(n1057) );
  XOR U1544 ( .A(n1143), .B(n1144), .Z(n1055) );
  ANDN U1545 ( .B(n1145), .A(n1146), .Z(n1143) );
  AND U1546 ( .A(b[10]), .B(a[39]), .Z(n1142) );
  XNOR U1547 ( .A(n1147), .B(n1060), .Z(n1062) );
  XOR U1548 ( .A(n1148), .B(n1149), .Z(n1060) );
  ANDN U1549 ( .B(n1150), .A(n1151), .Z(n1148) );
  AND U1550 ( .A(b[9]), .B(a[40]), .Z(n1147) );
  XNOR U1551 ( .A(n1152), .B(n1065), .Z(n1067) );
  XOR U1552 ( .A(n1153), .B(n1154), .Z(n1065) );
  ANDN U1553 ( .B(n1155), .A(n1156), .Z(n1153) );
  AND U1554 ( .A(b[8]), .B(a[41]), .Z(n1152) );
  XNOR U1555 ( .A(n1157), .B(n1070), .Z(n1072) );
  XOR U1556 ( .A(n1158), .B(n1159), .Z(n1070) );
  ANDN U1557 ( .B(n1160), .A(n1161), .Z(n1158) );
  AND U1558 ( .A(b[7]), .B(a[42]), .Z(n1157) );
  XNOR U1559 ( .A(n1162), .B(n1075), .Z(n1077) );
  XOR U1560 ( .A(n1163), .B(n1164), .Z(n1075) );
  ANDN U1561 ( .B(n1165), .A(n1166), .Z(n1163) );
  AND U1562 ( .A(b[6]), .B(a[43]), .Z(n1162) );
  XNOR U1563 ( .A(n1167), .B(n1080), .Z(n1082) );
  XOR U1564 ( .A(n1168), .B(n1169), .Z(n1080) );
  ANDN U1565 ( .B(n1170), .A(n1171), .Z(n1168) );
  AND U1566 ( .A(b[5]), .B(a[44]), .Z(n1167) );
  XNOR U1567 ( .A(n1172), .B(n1085), .Z(n1087) );
  XOR U1568 ( .A(n1173), .B(n1174), .Z(n1085) );
  ANDN U1569 ( .B(n1175), .A(n1176), .Z(n1173) );
  AND U1570 ( .A(b[4]), .B(a[45]), .Z(n1172) );
  XNOR U1571 ( .A(n1177), .B(n1178), .Z(n1099) );
  NANDN U1572 ( .A(n1179), .B(n1180), .Z(n1178) );
  XNOR U1573 ( .A(n1181), .B(n1090), .Z(n1092) );
  XNOR U1574 ( .A(n1182), .B(n1183), .Z(n1090) );
  AND U1575 ( .A(n1184), .B(n1185), .Z(n1182) );
  AND U1576 ( .A(b[3]), .B(a[46]), .Z(n1181) );
  XNOR U1577 ( .A(n1186), .B(n1187), .Z(swire[48]) );
  XOR U1578 ( .A(n1109), .B(n1189), .Z(n1187) );
  XNOR U1579 ( .A(n1108), .B(n1188), .Z(n1189) );
  IV U1580 ( .A(n1186), .Z(n1188) );
  NAND U1581 ( .A(a[48]), .B(b[0]), .Z(n1108) );
  XNOR U1582 ( .A(n1179), .B(n1180), .Z(n1109) );
  XOR U1583 ( .A(n1177), .B(n1190), .Z(n1180) );
  NAND U1584 ( .A(b[1]), .B(a[47]), .Z(n1190) );
  XOR U1585 ( .A(n1185), .B(n1191), .Z(n1179) );
  XOR U1586 ( .A(n1177), .B(n1184), .Z(n1191) );
  XNOR U1587 ( .A(n1192), .B(n1183), .Z(n1184) );
  AND U1588 ( .A(b[2]), .B(a[46]), .Z(n1192) );
  NANDN U1589 ( .A(n1193), .B(n1194), .Z(n1177) );
  XOR U1590 ( .A(n1183), .B(n1175), .Z(n1195) );
  XNOR U1591 ( .A(n1174), .B(n1170), .Z(n1196) );
  XNOR U1592 ( .A(n1169), .B(n1165), .Z(n1197) );
  XNOR U1593 ( .A(n1164), .B(n1160), .Z(n1198) );
  XNOR U1594 ( .A(n1159), .B(n1155), .Z(n1199) );
  XNOR U1595 ( .A(n1154), .B(n1150), .Z(n1200) );
  XNOR U1596 ( .A(n1149), .B(n1145), .Z(n1201) );
  XNOR U1597 ( .A(n1144), .B(n1140), .Z(n1202) );
  XNOR U1598 ( .A(n1139), .B(n1135), .Z(n1203) );
  XOR U1599 ( .A(n1134), .B(n1131), .Z(n1204) );
  XOR U1600 ( .A(n1205), .B(n1206), .Z(n1131) );
  XOR U1601 ( .A(n1129), .B(n1207), .Z(n1206) );
  XOR U1602 ( .A(n1208), .B(n1209), .Z(n1207) );
  XOR U1603 ( .A(n1210), .B(n1211), .Z(n1209) );
  NAND U1604 ( .A(b[14]), .B(a[34]), .Z(n1211) );
  AND U1605 ( .A(b[15]), .B(a[33]), .Z(n1210) );
  XOR U1606 ( .A(n1212), .B(n1208), .Z(n1205) );
  XOR U1607 ( .A(n1213), .B(n1214), .Z(n1208) );
  NOR U1608 ( .A(n1215), .B(n1216), .Z(n1213) );
  AND U1609 ( .A(b[13]), .B(a[35]), .Z(n1212) );
  XNOR U1610 ( .A(n1217), .B(n1129), .Z(n1130) );
  XOR U1611 ( .A(n1218), .B(n1219), .Z(n1129) );
  ANDN U1612 ( .B(n1220), .A(n1221), .Z(n1218) );
  AND U1613 ( .A(b[12]), .B(a[36]), .Z(n1217) );
  XNOR U1614 ( .A(n1222), .B(n1134), .Z(n1136) );
  XOR U1615 ( .A(n1223), .B(n1224), .Z(n1134) );
  ANDN U1616 ( .B(n1225), .A(n1226), .Z(n1223) );
  AND U1617 ( .A(b[11]), .B(a[37]), .Z(n1222) );
  XNOR U1618 ( .A(n1227), .B(n1139), .Z(n1141) );
  XOR U1619 ( .A(n1228), .B(n1229), .Z(n1139) );
  ANDN U1620 ( .B(n1230), .A(n1231), .Z(n1228) );
  AND U1621 ( .A(b[10]), .B(a[38]), .Z(n1227) );
  XNOR U1622 ( .A(n1232), .B(n1144), .Z(n1146) );
  XOR U1623 ( .A(n1233), .B(n1234), .Z(n1144) );
  ANDN U1624 ( .B(n1235), .A(n1236), .Z(n1233) );
  AND U1625 ( .A(b[9]), .B(a[39]), .Z(n1232) );
  XNOR U1626 ( .A(n1237), .B(n1149), .Z(n1151) );
  XOR U1627 ( .A(n1238), .B(n1239), .Z(n1149) );
  ANDN U1628 ( .B(n1240), .A(n1241), .Z(n1238) );
  AND U1629 ( .A(b[8]), .B(a[40]), .Z(n1237) );
  XNOR U1630 ( .A(n1242), .B(n1154), .Z(n1156) );
  XOR U1631 ( .A(n1243), .B(n1244), .Z(n1154) );
  ANDN U1632 ( .B(n1245), .A(n1246), .Z(n1243) );
  AND U1633 ( .A(b[7]), .B(a[41]), .Z(n1242) );
  XNOR U1634 ( .A(n1247), .B(n1159), .Z(n1161) );
  XOR U1635 ( .A(n1248), .B(n1249), .Z(n1159) );
  ANDN U1636 ( .B(n1250), .A(n1251), .Z(n1248) );
  AND U1637 ( .A(b[6]), .B(a[42]), .Z(n1247) );
  XNOR U1638 ( .A(n1252), .B(n1164), .Z(n1166) );
  XOR U1639 ( .A(n1253), .B(n1254), .Z(n1164) );
  ANDN U1640 ( .B(n1255), .A(n1256), .Z(n1253) );
  AND U1641 ( .A(b[5]), .B(a[43]), .Z(n1252) );
  XNOR U1642 ( .A(n1257), .B(n1169), .Z(n1171) );
  XOR U1643 ( .A(n1258), .B(n1259), .Z(n1169) );
  ANDN U1644 ( .B(n1260), .A(n1261), .Z(n1258) );
  AND U1645 ( .A(b[4]), .B(a[44]), .Z(n1257) );
  XNOR U1646 ( .A(n1262), .B(n1263), .Z(n1183) );
  NANDN U1647 ( .A(n1264), .B(n1265), .Z(n1263) );
  XNOR U1648 ( .A(n1266), .B(n1174), .Z(n1176) );
  XNOR U1649 ( .A(n1267), .B(n1268), .Z(n1174) );
  AND U1650 ( .A(n1269), .B(n1270), .Z(n1267) );
  AND U1651 ( .A(b[3]), .B(a[45]), .Z(n1266) );
  XNOR U1652 ( .A(n1271), .B(n1272), .Z(n1186) );
  NOR U1653 ( .A(n1273), .B(n1274), .Z(n1271) );
  XOR U1654 ( .A(n1274), .B(n1273), .Z(swire[47]) );
  XOR U1655 ( .A(sreg[111]), .B(n1272), .Z(n1273) );
  XOR U1656 ( .A(n1194), .B(n1275), .Z(n1274) );
  XNOR U1657 ( .A(n1193), .B(n1272), .Z(n1275) );
  XOR U1658 ( .A(n1276), .B(n1277), .Z(n1272) );
  NOR U1659 ( .A(n1278), .B(n1279), .Z(n1276) );
  NAND U1660 ( .A(a[47]), .B(b[0]), .Z(n1193) );
  XNOR U1661 ( .A(n1264), .B(n1265), .Z(n1194) );
  XOR U1662 ( .A(n1262), .B(n1280), .Z(n1265) );
  NAND U1663 ( .A(b[1]), .B(a[46]), .Z(n1280) );
  XOR U1664 ( .A(n1270), .B(n1281), .Z(n1264) );
  XOR U1665 ( .A(n1262), .B(n1269), .Z(n1281) );
  XNOR U1666 ( .A(n1282), .B(n1268), .Z(n1269) );
  AND U1667 ( .A(b[2]), .B(a[45]), .Z(n1282) );
  NANDN U1668 ( .A(n1283), .B(n1284), .Z(n1262) );
  XOR U1669 ( .A(n1268), .B(n1260), .Z(n1285) );
  XNOR U1670 ( .A(n1259), .B(n1255), .Z(n1286) );
  XNOR U1671 ( .A(n1254), .B(n1250), .Z(n1287) );
  XNOR U1672 ( .A(n1249), .B(n1245), .Z(n1288) );
  XNOR U1673 ( .A(n1244), .B(n1240), .Z(n1289) );
  XNOR U1674 ( .A(n1239), .B(n1235), .Z(n1290) );
  XNOR U1675 ( .A(n1234), .B(n1230), .Z(n1291) );
  XNOR U1676 ( .A(n1229), .B(n1225), .Z(n1292) );
  XNOR U1677 ( .A(n1224), .B(n1220), .Z(n1293) );
  XOR U1678 ( .A(n1219), .B(n1216), .Z(n1294) );
  XOR U1679 ( .A(n1295), .B(n1296), .Z(n1216) );
  XOR U1680 ( .A(n1214), .B(n1297), .Z(n1296) );
  XOR U1681 ( .A(n1298), .B(n1299), .Z(n1297) );
  XOR U1682 ( .A(n1300), .B(n1301), .Z(n1299) );
  NAND U1683 ( .A(b[14]), .B(a[33]), .Z(n1301) );
  AND U1684 ( .A(b[15]), .B(a[32]), .Z(n1300) );
  XOR U1685 ( .A(n1302), .B(n1298), .Z(n1295) );
  XOR U1686 ( .A(n1303), .B(n1304), .Z(n1298) );
  NOR U1687 ( .A(n1305), .B(n1306), .Z(n1303) );
  AND U1688 ( .A(b[13]), .B(a[34]), .Z(n1302) );
  XNOR U1689 ( .A(n1307), .B(n1214), .Z(n1215) );
  XOR U1690 ( .A(n1308), .B(n1309), .Z(n1214) );
  ANDN U1691 ( .B(n1310), .A(n1311), .Z(n1308) );
  AND U1692 ( .A(b[12]), .B(a[35]), .Z(n1307) );
  XNOR U1693 ( .A(n1312), .B(n1219), .Z(n1221) );
  XOR U1694 ( .A(n1313), .B(n1314), .Z(n1219) );
  ANDN U1695 ( .B(n1315), .A(n1316), .Z(n1313) );
  AND U1696 ( .A(b[11]), .B(a[36]), .Z(n1312) );
  XNOR U1697 ( .A(n1317), .B(n1224), .Z(n1226) );
  XOR U1698 ( .A(n1318), .B(n1319), .Z(n1224) );
  ANDN U1699 ( .B(n1320), .A(n1321), .Z(n1318) );
  AND U1700 ( .A(b[10]), .B(a[37]), .Z(n1317) );
  XNOR U1701 ( .A(n1322), .B(n1229), .Z(n1231) );
  XOR U1702 ( .A(n1323), .B(n1324), .Z(n1229) );
  ANDN U1703 ( .B(n1325), .A(n1326), .Z(n1323) );
  AND U1704 ( .A(b[9]), .B(a[38]), .Z(n1322) );
  XNOR U1705 ( .A(n1327), .B(n1234), .Z(n1236) );
  XOR U1706 ( .A(n1328), .B(n1329), .Z(n1234) );
  ANDN U1707 ( .B(n1330), .A(n1331), .Z(n1328) );
  AND U1708 ( .A(b[8]), .B(a[39]), .Z(n1327) );
  XNOR U1709 ( .A(n1332), .B(n1239), .Z(n1241) );
  XOR U1710 ( .A(n1333), .B(n1334), .Z(n1239) );
  ANDN U1711 ( .B(n1335), .A(n1336), .Z(n1333) );
  AND U1712 ( .A(b[7]), .B(a[40]), .Z(n1332) );
  XNOR U1713 ( .A(n1337), .B(n1244), .Z(n1246) );
  XOR U1714 ( .A(n1338), .B(n1339), .Z(n1244) );
  ANDN U1715 ( .B(n1340), .A(n1341), .Z(n1338) );
  AND U1716 ( .A(b[6]), .B(a[41]), .Z(n1337) );
  XNOR U1717 ( .A(n1342), .B(n1249), .Z(n1251) );
  XOR U1718 ( .A(n1343), .B(n1344), .Z(n1249) );
  ANDN U1719 ( .B(n1345), .A(n1346), .Z(n1343) );
  AND U1720 ( .A(b[5]), .B(a[42]), .Z(n1342) );
  XNOR U1721 ( .A(n1347), .B(n1254), .Z(n1256) );
  XOR U1722 ( .A(n1348), .B(n1349), .Z(n1254) );
  ANDN U1723 ( .B(n1350), .A(n1351), .Z(n1348) );
  AND U1724 ( .A(b[4]), .B(a[43]), .Z(n1347) );
  XNOR U1725 ( .A(n1352), .B(n1353), .Z(n1268) );
  NANDN U1726 ( .A(n1354), .B(n1355), .Z(n1353) );
  XNOR U1727 ( .A(n1356), .B(n1259), .Z(n1261) );
  XNOR U1728 ( .A(n1357), .B(n1358), .Z(n1259) );
  AND U1729 ( .A(n1359), .B(n1360), .Z(n1357) );
  AND U1730 ( .A(b[3]), .B(a[44]), .Z(n1356) );
  XOR U1731 ( .A(n1279), .B(n1278), .Z(swire[46]) );
  XOR U1732 ( .A(sreg[110]), .B(n1277), .Z(n1278) );
  XOR U1733 ( .A(n1284), .B(n1361), .Z(n1279) );
  XNOR U1734 ( .A(n1283), .B(n1277), .Z(n1361) );
  XOR U1735 ( .A(n1362), .B(n1363), .Z(n1277) );
  NOR U1736 ( .A(n1364), .B(n1365), .Z(n1362) );
  NAND U1737 ( .A(a[46]), .B(b[0]), .Z(n1283) );
  XNOR U1738 ( .A(n1354), .B(n1355), .Z(n1284) );
  XOR U1739 ( .A(n1352), .B(n1366), .Z(n1355) );
  NAND U1740 ( .A(b[1]), .B(a[45]), .Z(n1366) );
  XOR U1741 ( .A(n1360), .B(n1367), .Z(n1354) );
  XOR U1742 ( .A(n1352), .B(n1359), .Z(n1367) );
  XNOR U1743 ( .A(n1368), .B(n1358), .Z(n1359) );
  AND U1744 ( .A(b[2]), .B(a[44]), .Z(n1368) );
  NANDN U1745 ( .A(n1369), .B(n1370), .Z(n1352) );
  XOR U1746 ( .A(n1358), .B(n1350), .Z(n1371) );
  XNOR U1747 ( .A(n1349), .B(n1345), .Z(n1372) );
  XNOR U1748 ( .A(n1344), .B(n1340), .Z(n1373) );
  XNOR U1749 ( .A(n1339), .B(n1335), .Z(n1374) );
  XNOR U1750 ( .A(n1334), .B(n1330), .Z(n1375) );
  XNOR U1751 ( .A(n1329), .B(n1325), .Z(n1376) );
  XNOR U1752 ( .A(n1324), .B(n1320), .Z(n1377) );
  XNOR U1753 ( .A(n1319), .B(n1315), .Z(n1378) );
  XNOR U1754 ( .A(n1314), .B(n1310), .Z(n1379) );
  XOR U1755 ( .A(n1309), .B(n1306), .Z(n1380) );
  XOR U1756 ( .A(n1381), .B(n1382), .Z(n1306) );
  XOR U1757 ( .A(n1304), .B(n1383), .Z(n1382) );
  XOR U1758 ( .A(n1384), .B(n1385), .Z(n1383) );
  XOR U1759 ( .A(n1386), .B(n1387), .Z(n1385) );
  NAND U1760 ( .A(b[14]), .B(a[32]), .Z(n1387) );
  AND U1761 ( .A(b[15]), .B(a[31]), .Z(n1386) );
  XOR U1762 ( .A(n1388), .B(n1384), .Z(n1381) );
  XOR U1763 ( .A(n1389), .B(n1390), .Z(n1384) );
  NOR U1764 ( .A(n1391), .B(n1392), .Z(n1389) );
  AND U1765 ( .A(b[13]), .B(a[33]), .Z(n1388) );
  XNOR U1766 ( .A(n1393), .B(n1304), .Z(n1305) );
  XOR U1767 ( .A(n1394), .B(n1395), .Z(n1304) );
  ANDN U1768 ( .B(n1396), .A(n1397), .Z(n1394) );
  AND U1769 ( .A(b[12]), .B(a[34]), .Z(n1393) );
  XNOR U1770 ( .A(n1398), .B(n1309), .Z(n1311) );
  XOR U1771 ( .A(n1399), .B(n1400), .Z(n1309) );
  ANDN U1772 ( .B(n1401), .A(n1402), .Z(n1399) );
  AND U1773 ( .A(b[11]), .B(a[35]), .Z(n1398) );
  XNOR U1774 ( .A(n1403), .B(n1314), .Z(n1316) );
  XOR U1775 ( .A(n1404), .B(n1405), .Z(n1314) );
  ANDN U1776 ( .B(n1406), .A(n1407), .Z(n1404) );
  AND U1777 ( .A(b[10]), .B(a[36]), .Z(n1403) );
  XNOR U1778 ( .A(n1408), .B(n1319), .Z(n1321) );
  XOR U1779 ( .A(n1409), .B(n1410), .Z(n1319) );
  ANDN U1780 ( .B(n1411), .A(n1412), .Z(n1409) );
  AND U1781 ( .A(b[9]), .B(a[37]), .Z(n1408) );
  XNOR U1782 ( .A(n1413), .B(n1324), .Z(n1326) );
  XOR U1783 ( .A(n1414), .B(n1415), .Z(n1324) );
  ANDN U1784 ( .B(n1416), .A(n1417), .Z(n1414) );
  AND U1785 ( .A(b[8]), .B(a[38]), .Z(n1413) );
  XNOR U1786 ( .A(n1418), .B(n1329), .Z(n1331) );
  XOR U1787 ( .A(n1419), .B(n1420), .Z(n1329) );
  ANDN U1788 ( .B(n1421), .A(n1422), .Z(n1419) );
  AND U1789 ( .A(b[7]), .B(a[39]), .Z(n1418) );
  XNOR U1790 ( .A(n1423), .B(n1334), .Z(n1336) );
  XOR U1791 ( .A(n1424), .B(n1425), .Z(n1334) );
  ANDN U1792 ( .B(n1426), .A(n1427), .Z(n1424) );
  AND U1793 ( .A(b[6]), .B(a[40]), .Z(n1423) );
  XNOR U1794 ( .A(n1428), .B(n1339), .Z(n1341) );
  XOR U1795 ( .A(n1429), .B(n1430), .Z(n1339) );
  ANDN U1796 ( .B(n1431), .A(n1432), .Z(n1429) );
  AND U1797 ( .A(b[5]), .B(a[41]), .Z(n1428) );
  XNOR U1798 ( .A(n1433), .B(n1344), .Z(n1346) );
  XOR U1799 ( .A(n1434), .B(n1435), .Z(n1344) );
  ANDN U1800 ( .B(n1436), .A(n1437), .Z(n1434) );
  AND U1801 ( .A(b[4]), .B(a[42]), .Z(n1433) );
  XNOR U1802 ( .A(n1438), .B(n1439), .Z(n1358) );
  NANDN U1803 ( .A(n1440), .B(n1441), .Z(n1439) );
  XNOR U1804 ( .A(n1442), .B(n1349), .Z(n1351) );
  XNOR U1805 ( .A(n1443), .B(n1444), .Z(n1349) );
  AND U1806 ( .A(n1445), .B(n1446), .Z(n1443) );
  AND U1807 ( .A(b[3]), .B(a[43]), .Z(n1442) );
  XOR U1808 ( .A(n1365), .B(n1364), .Z(swire[45]) );
  XOR U1809 ( .A(sreg[109]), .B(n1363), .Z(n1364) );
  XOR U1810 ( .A(n1370), .B(n1447), .Z(n1365) );
  XNOR U1811 ( .A(n1369), .B(n1363), .Z(n1447) );
  XOR U1812 ( .A(n1448), .B(n1449), .Z(n1363) );
  NOR U1813 ( .A(n1450), .B(n1451), .Z(n1448) );
  NAND U1814 ( .A(a[45]), .B(b[0]), .Z(n1369) );
  XNOR U1815 ( .A(n1440), .B(n1441), .Z(n1370) );
  XOR U1816 ( .A(n1438), .B(n1452), .Z(n1441) );
  NAND U1817 ( .A(b[1]), .B(a[44]), .Z(n1452) );
  XOR U1818 ( .A(n1446), .B(n1453), .Z(n1440) );
  XOR U1819 ( .A(n1438), .B(n1445), .Z(n1453) );
  XNOR U1820 ( .A(n1454), .B(n1444), .Z(n1445) );
  AND U1821 ( .A(b[2]), .B(a[43]), .Z(n1454) );
  NANDN U1822 ( .A(n1455), .B(n1456), .Z(n1438) );
  XOR U1823 ( .A(n1444), .B(n1436), .Z(n1457) );
  XNOR U1824 ( .A(n1435), .B(n1431), .Z(n1458) );
  XNOR U1825 ( .A(n1430), .B(n1426), .Z(n1459) );
  XNOR U1826 ( .A(n1425), .B(n1421), .Z(n1460) );
  XNOR U1827 ( .A(n1420), .B(n1416), .Z(n1461) );
  XNOR U1828 ( .A(n1415), .B(n1411), .Z(n1462) );
  XNOR U1829 ( .A(n1410), .B(n1406), .Z(n1463) );
  XNOR U1830 ( .A(n1405), .B(n1401), .Z(n1464) );
  XNOR U1831 ( .A(n1400), .B(n1396), .Z(n1465) );
  XOR U1832 ( .A(n1395), .B(n1392), .Z(n1466) );
  XOR U1833 ( .A(n1467), .B(n1468), .Z(n1392) );
  XOR U1834 ( .A(n1390), .B(n1469), .Z(n1468) );
  XOR U1835 ( .A(n1470), .B(n1471), .Z(n1469) );
  XOR U1836 ( .A(n1472), .B(n1473), .Z(n1471) );
  NAND U1837 ( .A(b[14]), .B(a[31]), .Z(n1473) );
  AND U1838 ( .A(b[15]), .B(a[30]), .Z(n1472) );
  XOR U1839 ( .A(n1474), .B(n1470), .Z(n1467) );
  XOR U1840 ( .A(n1475), .B(n1476), .Z(n1470) );
  NOR U1841 ( .A(n1477), .B(n1478), .Z(n1475) );
  AND U1842 ( .A(b[13]), .B(a[32]), .Z(n1474) );
  XNOR U1843 ( .A(n1479), .B(n1390), .Z(n1391) );
  XOR U1844 ( .A(n1480), .B(n1481), .Z(n1390) );
  ANDN U1845 ( .B(n1482), .A(n1483), .Z(n1480) );
  AND U1846 ( .A(b[12]), .B(a[33]), .Z(n1479) );
  XNOR U1847 ( .A(n1484), .B(n1395), .Z(n1397) );
  XOR U1848 ( .A(n1485), .B(n1486), .Z(n1395) );
  ANDN U1849 ( .B(n1487), .A(n1488), .Z(n1485) );
  AND U1850 ( .A(b[11]), .B(a[34]), .Z(n1484) );
  XNOR U1851 ( .A(n1489), .B(n1400), .Z(n1402) );
  XOR U1852 ( .A(n1490), .B(n1491), .Z(n1400) );
  ANDN U1853 ( .B(n1492), .A(n1493), .Z(n1490) );
  AND U1854 ( .A(b[10]), .B(a[35]), .Z(n1489) );
  XNOR U1855 ( .A(n1494), .B(n1405), .Z(n1407) );
  XOR U1856 ( .A(n1495), .B(n1496), .Z(n1405) );
  ANDN U1857 ( .B(n1497), .A(n1498), .Z(n1495) );
  AND U1858 ( .A(b[9]), .B(a[36]), .Z(n1494) );
  XNOR U1859 ( .A(n1499), .B(n1410), .Z(n1412) );
  XOR U1860 ( .A(n1500), .B(n1501), .Z(n1410) );
  ANDN U1861 ( .B(n1502), .A(n1503), .Z(n1500) );
  AND U1862 ( .A(b[8]), .B(a[37]), .Z(n1499) );
  XNOR U1863 ( .A(n1504), .B(n1415), .Z(n1417) );
  XOR U1864 ( .A(n1505), .B(n1506), .Z(n1415) );
  ANDN U1865 ( .B(n1507), .A(n1508), .Z(n1505) );
  AND U1866 ( .A(b[7]), .B(a[38]), .Z(n1504) );
  XNOR U1867 ( .A(n1509), .B(n1420), .Z(n1422) );
  XOR U1868 ( .A(n1510), .B(n1511), .Z(n1420) );
  ANDN U1869 ( .B(n1512), .A(n1513), .Z(n1510) );
  AND U1870 ( .A(b[6]), .B(a[39]), .Z(n1509) );
  XNOR U1871 ( .A(n1514), .B(n1425), .Z(n1427) );
  XOR U1872 ( .A(n1515), .B(n1516), .Z(n1425) );
  ANDN U1873 ( .B(n1517), .A(n1518), .Z(n1515) );
  AND U1874 ( .A(b[5]), .B(a[40]), .Z(n1514) );
  XNOR U1875 ( .A(n1519), .B(n1430), .Z(n1432) );
  XOR U1876 ( .A(n1520), .B(n1521), .Z(n1430) );
  ANDN U1877 ( .B(n1522), .A(n1523), .Z(n1520) );
  AND U1878 ( .A(b[4]), .B(a[41]), .Z(n1519) );
  XNOR U1879 ( .A(n1524), .B(n1525), .Z(n1444) );
  NANDN U1880 ( .A(n1526), .B(n1527), .Z(n1525) );
  XNOR U1881 ( .A(n1528), .B(n1435), .Z(n1437) );
  XNOR U1882 ( .A(n1529), .B(n1530), .Z(n1435) );
  AND U1883 ( .A(n1531), .B(n1532), .Z(n1529) );
  AND U1884 ( .A(b[3]), .B(a[42]), .Z(n1528) );
  XOR U1885 ( .A(n1451), .B(n1450), .Z(swire[44]) );
  XOR U1886 ( .A(sreg[108]), .B(n1449), .Z(n1450) );
  XOR U1887 ( .A(n1456), .B(n1533), .Z(n1451) );
  XNOR U1888 ( .A(n1455), .B(n1449), .Z(n1533) );
  XOR U1889 ( .A(n1534), .B(n1535), .Z(n1449) );
  NOR U1890 ( .A(n1536), .B(n1537), .Z(n1534) );
  NAND U1891 ( .A(a[44]), .B(b[0]), .Z(n1455) );
  XNOR U1892 ( .A(n1526), .B(n1527), .Z(n1456) );
  XOR U1893 ( .A(n1524), .B(n1538), .Z(n1527) );
  NAND U1894 ( .A(b[1]), .B(a[43]), .Z(n1538) );
  XOR U1895 ( .A(n1532), .B(n1539), .Z(n1526) );
  XOR U1896 ( .A(n1524), .B(n1531), .Z(n1539) );
  XNOR U1897 ( .A(n1540), .B(n1530), .Z(n1531) );
  AND U1898 ( .A(b[2]), .B(a[42]), .Z(n1540) );
  NANDN U1899 ( .A(n1541), .B(n1542), .Z(n1524) );
  XOR U1900 ( .A(n1530), .B(n1522), .Z(n1543) );
  XNOR U1901 ( .A(n1521), .B(n1517), .Z(n1544) );
  XNOR U1902 ( .A(n1516), .B(n1512), .Z(n1545) );
  XNOR U1903 ( .A(n1511), .B(n1507), .Z(n1546) );
  XNOR U1904 ( .A(n1506), .B(n1502), .Z(n1547) );
  XNOR U1905 ( .A(n1501), .B(n1497), .Z(n1548) );
  XNOR U1906 ( .A(n1496), .B(n1492), .Z(n1549) );
  XNOR U1907 ( .A(n1491), .B(n1487), .Z(n1550) );
  XNOR U1908 ( .A(n1486), .B(n1482), .Z(n1551) );
  XOR U1909 ( .A(n1481), .B(n1478), .Z(n1552) );
  XOR U1910 ( .A(n1553), .B(n1554), .Z(n1478) );
  XOR U1911 ( .A(n1476), .B(n1555), .Z(n1554) );
  XOR U1912 ( .A(n1556), .B(n1557), .Z(n1555) );
  XOR U1913 ( .A(n1558), .B(n1559), .Z(n1557) );
  NAND U1914 ( .A(b[14]), .B(a[30]), .Z(n1559) );
  AND U1915 ( .A(b[15]), .B(a[29]), .Z(n1558) );
  XOR U1916 ( .A(n1560), .B(n1556), .Z(n1553) );
  XOR U1917 ( .A(n1561), .B(n1562), .Z(n1556) );
  NOR U1918 ( .A(n1563), .B(n1564), .Z(n1561) );
  AND U1919 ( .A(b[13]), .B(a[31]), .Z(n1560) );
  XNOR U1920 ( .A(n1565), .B(n1476), .Z(n1477) );
  XOR U1921 ( .A(n1566), .B(n1567), .Z(n1476) );
  ANDN U1922 ( .B(n1568), .A(n1569), .Z(n1566) );
  AND U1923 ( .A(b[12]), .B(a[32]), .Z(n1565) );
  XNOR U1924 ( .A(n1570), .B(n1481), .Z(n1483) );
  XOR U1925 ( .A(n1571), .B(n1572), .Z(n1481) );
  ANDN U1926 ( .B(n1573), .A(n1574), .Z(n1571) );
  AND U1927 ( .A(b[11]), .B(a[33]), .Z(n1570) );
  XNOR U1928 ( .A(n1575), .B(n1486), .Z(n1488) );
  XOR U1929 ( .A(n1576), .B(n1577), .Z(n1486) );
  ANDN U1930 ( .B(n1578), .A(n1579), .Z(n1576) );
  AND U1931 ( .A(b[10]), .B(a[34]), .Z(n1575) );
  XNOR U1932 ( .A(n1580), .B(n1491), .Z(n1493) );
  XOR U1933 ( .A(n1581), .B(n1582), .Z(n1491) );
  ANDN U1934 ( .B(n1583), .A(n1584), .Z(n1581) );
  AND U1935 ( .A(b[9]), .B(a[35]), .Z(n1580) );
  XNOR U1936 ( .A(n1585), .B(n1496), .Z(n1498) );
  XOR U1937 ( .A(n1586), .B(n1587), .Z(n1496) );
  ANDN U1938 ( .B(n1588), .A(n1589), .Z(n1586) );
  AND U1939 ( .A(b[8]), .B(a[36]), .Z(n1585) );
  XNOR U1940 ( .A(n1590), .B(n1501), .Z(n1503) );
  XOR U1941 ( .A(n1591), .B(n1592), .Z(n1501) );
  ANDN U1942 ( .B(n1593), .A(n1594), .Z(n1591) );
  AND U1943 ( .A(b[7]), .B(a[37]), .Z(n1590) );
  XNOR U1944 ( .A(n1595), .B(n1506), .Z(n1508) );
  XOR U1945 ( .A(n1596), .B(n1597), .Z(n1506) );
  ANDN U1946 ( .B(n1598), .A(n1599), .Z(n1596) );
  AND U1947 ( .A(b[6]), .B(a[38]), .Z(n1595) );
  XNOR U1948 ( .A(n1600), .B(n1511), .Z(n1513) );
  XOR U1949 ( .A(n1601), .B(n1602), .Z(n1511) );
  ANDN U1950 ( .B(n1603), .A(n1604), .Z(n1601) );
  AND U1951 ( .A(b[5]), .B(a[39]), .Z(n1600) );
  XNOR U1952 ( .A(n1605), .B(n1516), .Z(n1518) );
  XOR U1953 ( .A(n1606), .B(n1607), .Z(n1516) );
  ANDN U1954 ( .B(n1608), .A(n1609), .Z(n1606) );
  AND U1955 ( .A(b[4]), .B(a[40]), .Z(n1605) );
  XNOR U1956 ( .A(n1610), .B(n1611), .Z(n1530) );
  NANDN U1957 ( .A(n1612), .B(n1613), .Z(n1611) );
  XNOR U1958 ( .A(n1614), .B(n1521), .Z(n1523) );
  XNOR U1959 ( .A(n1615), .B(n1616), .Z(n1521) );
  AND U1960 ( .A(n1617), .B(n1618), .Z(n1615) );
  AND U1961 ( .A(b[3]), .B(a[41]), .Z(n1614) );
  XOR U1962 ( .A(n1537), .B(n1536), .Z(swire[43]) );
  XOR U1963 ( .A(sreg[107]), .B(n1535), .Z(n1536) );
  XOR U1964 ( .A(n1542), .B(n1619), .Z(n1537) );
  XNOR U1965 ( .A(n1541), .B(n1535), .Z(n1619) );
  XOR U1966 ( .A(n1620), .B(n1621), .Z(n1535) );
  NOR U1967 ( .A(n1622), .B(n1623), .Z(n1620) );
  NAND U1968 ( .A(a[43]), .B(b[0]), .Z(n1541) );
  XNOR U1969 ( .A(n1612), .B(n1613), .Z(n1542) );
  XOR U1970 ( .A(n1610), .B(n1624), .Z(n1613) );
  NAND U1971 ( .A(b[1]), .B(a[42]), .Z(n1624) );
  XOR U1972 ( .A(n1618), .B(n1625), .Z(n1612) );
  XOR U1973 ( .A(n1610), .B(n1617), .Z(n1625) );
  XNOR U1974 ( .A(n1626), .B(n1616), .Z(n1617) );
  AND U1975 ( .A(b[2]), .B(a[41]), .Z(n1626) );
  NANDN U1976 ( .A(n1627), .B(n1628), .Z(n1610) );
  XOR U1977 ( .A(n1616), .B(n1608), .Z(n1629) );
  XNOR U1978 ( .A(n1607), .B(n1603), .Z(n1630) );
  XNOR U1979 ( .A(n1602), .B(n1598), .Z(n1631) );
  XNOR U1980 ( .A(n1597), .B(n1593), .Z(n1632) );
  XNOR U1981 ( .A(n1592), .B(n1588), .Z(n1633) );
  XNOR U1982 ( .A(n1587), .B(n1583), .Z(n1634) );
  XNOR U1983 ( .A(n1582), .B(n1578), .Z(n1635) );
  XNOR U1984 ( .A(n1577), .B(n1573), .Z(n1636) );
  XNOR U1985 ( .A(n1572), .B(n1568), .Z(n1637) );
  XOR U1986 ( .A(n1567), .B(n1564), .Z(n1638) );
  XOR U1987 ( .A(n1639), .B(n1640), .Z(n1564) );
  XOR U1988 ( .A(n1562), .B(n1641), .Z(n1640) );
  XOR U1989 ( .A(n1642), .B(n1643), .Z(n1641) );
  XOR U1990 ( .A(n1644), .B(n1645), .Z(n1643) );
  NAND U1991 ( .A(b[14]), .B(a[29]), .Z(n1645) );
  AND U1992 ( .A(b[15]), .B(a[28]), .Z(n1644) );
  XOR U1993 ( .A(n1646), .B(n1642), .Z(n1639) );
  XOR U1994 ( .A(n1647), .B(n1648), .Z(n1642) );
  NOR U1995 ( .A(n1649), .B(n1650), .Z(n1647) );
  AND U1996 ( .A(b[13]), .B(a[30]), .Z(n1646) );
  XNOR U1997 ( .A(n1651), .B(n1562), .Z(n1563) );
  XOR U1998 ( .A(n1652), .B(n1653), .Z(n1562) );
  ANDN U1999 ( .B(n1654), .A(n1655), .Z(n1652) );
  AND U2000 ( .A(b[12]), .B(a[31]), .Z(n1651) );
  XNOR U2001 ( .A(n1656), .B(n1567), .Z(n1569) );
  XOR U2002 ( .A(n1657), .B(n1658), .Z(n1567) );
  ANDN U2003 ( .B(n1659), .A(n1660), .Z(n1657) );
  AND U2004 ( .A(b[11]), .B(a[32]), .Z(n1656) );
  XNOR U2005 ( .A(n1661), .B(n1572), .Z(n1574) );
  XOR U2006 ( .A(n1662), .B(n1663), .Z(n1572) );
  ANDN U2007 ( .B(n1664), .A(n1665), .Z(n1662) );
  AND U2008 ( .A(b[10]), .B(a[33]), .Z(n1661) );
  XNOR U2009 ( .A(n1666), .B(n1577), .Z(n1579) );
  XOR U2010 ( .A(n1667), .B(n1668), .Z(n1577) );
  ANDN U2011 ( .B(n1669), .A(n1670), .Z(n1667) );
  AND U2012 ( .A(b[9]), .B(a[34]), .Z(n1666) );
  XNOR U2013 ( .A(n1671), .B(n1582), .Z(n1584) );
  XOR U2014 ( .A(n1672), .B(n1673), .Z(n1582) );
  ANDN U2015 ( .B(n1674), .A(n1675), .Z(n1672) );
  AND U2016 ( .A(b[8]), .B(a[35]), .Z(n1671) );
  XNOR U2017 ( .A(n1676), .B(n1587), .Z(n1589) );
  XOR U2018 ( .A(n1677), .B(n1678), .Z(n1587) );
  ANDN U2019 ( .B(n1679), .A(n1680), .Z(n1677) );
  AND U2020 ( .A(b[7]), .B(a[36]), .Z(n1676) );
  XNOR U2021 ( .A(n1681), .B(n1592), .Z(n1594) );
  XOR U2022 ( .A(n1682), .B(n1683), .Z(n1592) );
  ANDN U2023 ( .B(n1684), .A(n1685), .Z(n1682) );
  AND U2024 ( .A(b[6]), .B(a[37]), .Z(n1681) );
  XNOR U2025 ( .A(n1686), .B(n1597), .Z(n1599) );
  XOR U2026 ( .A(n1687), .B(n1688), .Z(n1597) );
  ANDN U2027 ( .B(n1689), .A(n1690), .Z(n1687) );
  AND U2028 ( .A(b[5]), .B(a[38]), .Z(n1686) );
  XNOR U2029 ( .A(n1691), .B(n1602), .Z(n1604) );
  XOR U2030 ( .A(n1692), .B(n1693), .Z(n1602) );
  ANDN U2031 ( .B(n1694), .A(n1695), .Z(n1692) );
  AND U2032 ( .A(b[4]), .B(a[39]), .Z(n1691) );
  XNOR U2033 ( .A(n1696), .B(n1697), .Z(n1616) );
  NANDN U2034 ( .A(n1698), .B(n1699), .Z(n1697) );
  XNOR U2035 ( .A(n1700), .B(n1607), .Z(n1609) );
  XNOR U2036 ( .A(n1701), .B(n1702), .Z(n1607) );
  AND U2037 ( .A(n1703), .B(n1704), .Z(n1701) );
  AND U2038 ( .A(b[3]), .B(a[40]), .Z(n1700) );
  XOR U2039 ( .A(n1623), .B(n1622), .Z(swire[42]) );
  XOR U2040 ( .A(sreg[106]), .B(n1621), .Z(n1622) );
  XOR U2041 ( .A(n1628), .B(n1705), .Z(n1623) );
  XNOR U2042 ( .A(n1627), .B(n1621), .Z(n1705) );
  XOR U2043 ( .A(n1706), .B(n1707), .Z(n1621) );
  NOR U2044 ( .A(n1708), .B(n1709), .Z(n1706) );
  NAND U2045 ( .A(a[42]), .B(b[0]), .Z(n1627) );
  XNOR U2046 ( .A(n1698), .B(n1699), .Z(n1628) );
  XOR U2047 ( .A(n1696), .B(n1710), .Z(n1699) );
  NAND U2048 ( .A(b[1]), .B(a[41]), .Z(n1710) );
  XOR U2049 ( .A(n1704), .B(n1711), .Z(n1698) );
  XOR U2050 ( .A(n1696), .B(n1703), .Z(n1711) );
  XNOR U2051 ( .A(n1712), .B(n1702), .Z(n1703) );
  AND U2052 ( .A(b[2]), .B(a[40]), .Z(n1712) );
  NANDN U2053 ( .A(n1713), .B(n1714), .Z(n1696) );
  XOR U2054 ( .A(n1702), .B(n1694), .Z(n1715) );
  XNOR U2055 ( .A(n1693), .B(n1689), .Z(n1716) );
  XNOR U2056 ( .A(n1688), .B(n1684), .Z(n1717) );
  XNOR U2057 ( .A(n1683), .B(n1679), .Z(n1718) );
  XNOR U2058 ( .A(n1678), .B(n1674), .Z(n1719) );
  XNOR U2059 ( .A(n1673), .B(n1669), .Z(n1720) );
  XNOR U2060 ( .A(n1668), .B(n1664), .Z(n1721) );
  XNOR U2061 ( .A(n1663), .B(n1659), .Z(n1722) );
  XNOR U2062 ( .A(n1658), .B(n1654), .Z(n1723) );
  XOR U2063 ( .A(n1653), .B(n1650), .Z(n1724) );
  XOR U2064 ( .A(n1725), .B(n1726), .Z(n1650) );
  XOR U2065 ( .A(n1648), .B(n1727), .Z(n1726) );
  XOR U2066 ( .A(n1728), .B(n1729), .Z(n1727) );
  XOR U2067 ( .A(n1730), .B(n1731), .Z(n1729) );
  NAND U2068 ( .A(b[14]), .B(a[28]), .Z(n1731) );
  AND U2069 ( .A(b[15]), .B(a[27]), .Z(n1730) );
  XOR U2070 ( .A(n1732), .B(n1728), .Z(n1725) );
  XOR U2071 ( .A(n1733), .B(n1734), .Z(n1728) );
  NOR U2072 ( .A(n1735), .B(n1736), .Z(n1733) );
  AND U2073 ( .A(b[13]), .B(a[29]), .Z(n1732) );
  XNOR U2074 ( .A(n1737), .B(n1648), .Z(n1649) );
  XOR U2075 ( .A(n1738), .B(n1739), .Z(n1648) );
  ANDN U2076 ( .B(n1740), .A(n1741), .Z(n1738) );
  AND U2077 ( .A(b[12]), .B(a[30]), .Z(n1737) );
  XNOR U2078 ( .A(n1742), .B(n1653), .Z(n1655) );
  XOR U2079 ( .A(n1743), .B(n1744), .Z(n1653) );
  ANDN U2080 ( .B(n1745), .A(n1746), .Z(n1743) );
  AND U2081 ( .A(b[11]), .B(a[31]), .Z(n1742) );
  XNOR U2082 ( .A(n1747), .B(n1658), .Z(n1660) );
  XOR U2083 ( .A(n1748), .B(n1749), .Z(n1658) );
  ANDN U2084 ( .B(n1750), .A(n1751), .Z(n1748) );
  AND U2085 ( .A(b[10]), .B(a[32]), .Z(n1747) );
  XNOR U2086 ( .A(n1752), .B(n1663), .Z(n1665) );
  XOR U2087 ( .A(n1753), .B(n1754), .Z(n1663) );
  ANDN U2088 ( .B(n1755), .A(n1756), .Z(n1753) );
  AND U2089 ( .A(b[9]), .B(a[33]), .Z(n1752) );
  XNOR U2090 ( .A(n1757), .B(n1668), .Z(n1670) );
  XOR U2091 ( .A(n1758), .B(n1759), .Z(n1668) );
  ANDN U2092 ( .B(n1760), .A(n1761), .Z(n1758) );
  AND U2093 ( .A(b[8]), .B(a[34]), .Z(n1757) );
  XNOR U2094 ( .A(n1762), .B(n1673), .Z(n1675) );
  XOR U2095 ( .A(n1763), .B(n1764), .Z(n1673) );
  ANDN U2096 ( .B(n1765), .A(n1766), .Z(n1763) );
  AND U2097 ( .A(b[7]), .B(a[35]), .Z(n1762) );
  XNOR U2098 ( .A(n1767), .B(n1678), .Z(n1680) );
  XOR U2099 ( .A(n1768), .B(n1769), .Z(n1678) );
  ANDN U2100 ( .B(n1770), .A(n1771), .Z(n1768) );
  AND U2101 ( .A(b[6]), .B(a[36]), .Z(n1767) );
  XNOR U2102 ( .A(n1772), .B(n1683), .Z(n1685) );
  XOR U2103 ( .A(n1773), .B(n1774), .Z(n1683) );
  ANDN U2104 ( .B(n1775), .A(n1776), .Z(n1773) );
  AND U2105 ( .A(b[5]), .B(a[37]), .Z(n1772) );
  XNOR U2106 ( .A(n1777), .B(n1688), .Z(n1690) );
  XOR U2107 ( .A(n1778), .B(n1779), .Z(n1688) );
  ANDN U2108 ( .B(n1780), .A(n1781), .Z(n1778) );
  AND U2109 ( .A(b[4]), .B(a[38]), .Z(n1777) );
  XNOR U2110 ( .A(n1782), .B(n1783), .Z(n1702) );
  NANDN U2111 ( .A(n1784), .B(n1785), .Z(n1783) );
  XNOR U2112 ( .A(n1786), .B(n1693), .Z(n1695) );
  XNOR U2113 ( .A(n1787), .B(n1788), .Z(n1693) );
  AND U2114 ( .A(n1789), .B(n1790), .Z(n1787) );
  AND U2115 ( .A(b[3]), .B(a[39]), .Z(n1786) );
  XOR U2116 ( .A(n1709), .B(n1708), .Z(swire[41]) );
  XOR U2117 ( .A(sreg[105]), .B(n1707), .Z(n1708) );
  XOR U2118 ( .A(n1714), .B(n1791), .Z(n1709) );
  XNOR U2119 ( .A(n1713), .B(n1707), .Z(n1791) );
  XOR U2120 ( .A(n1792), .B(n1793), .Z(n1707) );
  NOR U2121 ( .A(n1794), .B(n1795), .Z(n1792) );
  NAND U2122 ( .A(a[41]), .B(b[0]), .Z(n1713) );
  XNOR U2123 ( .A(n1784), .B(n1785), .Z(n1714) );
  XOR U2124 ( .A(n1782), .B(n1796), .Z(n1785) );
  NAND U2125 ( .A(b[1]), .B(a[40]), .Z(n1796) );
  XOR U2126 ( .A(n1790), .B(n1797), .Z(n1784) );
  XOR U2127 ( .A(n1782), .B(n1789), .Z(n1797) );
  XNOR U2128 ( .A(n1798), .B(n1788), .Z(n1789) );
  AND U2129 ( .A(b[2]), .B(a[39]), .Z(n1798) );
  NANDN U2130 ( .A(n1799), .B(n1800), .Z(n1782) );
  XOR U2131 ( .A(n1788), .B(n1780), .Z(n1801) );
  XNOR U2132 ( .A(n1779), .B(n1775), .Z(n1802) );
  XNOR U2133 ( .A(n1774), .B(n1770), .Z(n1803) );
  XNOR U2134 ( .A(n1769), .B(n1765), .Z(n1804) );
  XNOR U2135 ( .A(n1764), .B(n1760), .Z(n1805) );
  XNOR U2136 ( .A(n1759), .B(n1755), .Z(n1806) );
  XNOR U2137 ( .A(n1754), .B(n1750), .Z(n1807) );
  XNOR U2138 ( .A(n1749), .B(n1745), .Z(n1808) );
  XNOR U2139 ( .A(n1744), .B(n1740), .Z(n1809) );
  XOR U2140 ( .A(n1739), .B(n1736), .Z(n1810) );
  XOR U2141 ( .A(n1811), .B(n1812), .Z(n1736) );
  XOR U2142 ( .A(n1734), .B(n1813), .Z(n1812) );
  XOR U2143 ( .A(n1814), .B(n1815), .Z(n1813) );
  XOR U2144 ( .A(n1816), .B(n1817), .Z(n1815) );
  NAND U2145 ( .A(b[14]), .B(a[27]), .Z(n1817) );
  AND U2146 ( .A(b[15]), .B(a[26]), .Z(n1816) );
  XOR U2147 ( .A(n1818), .B(n1814), .Z(n1811) );
  XOR U2148 ( .A(n1819), .B(n1820), .Z(n1814) );
  NOR U2149 ( .A(n1821), .B(n1822), .Z(n1819) );
  AND U2150 ( .A(b[13]), .B(a[28]), .Z(n1818) );
  XNOR U2151 ( .A(n1823), .B(n1734), .Z(n1735) );
  XOR U2152 ( .A(n1824), .B(n1825), .Z(n1734) );
  ANDN U2153 ( .B(n1826), .A(n1827), .Z(n1824) );
  AND U2154 ( .A(b[12]), .B(a[29]), .Z(n1823) );
  XNOR U2155 ( .A(n1828), .B(n1739), .Z(n1741) );
  XOR U2156 ( .A(n1829), .B(n1830), .Z(n1739) );
  ANDN U2157 ( .B(n1831), .A(n1832), .Z(n1829) );
  AND U2158 ( .A(b[11]), .B(a[30]), .Z(n1828) );
  XNOR U2159 ( .A(n1833), .B(n1744), .Z(n1746) );
  XOR U2160 ( .A(n1834), .B(n1835), .Z(n1744) );
  ANDN U2161 ( .B(n1836), .A(n1837), .Z(n1834) );
  AND U2162 ( .A(b[10]), .B(a[31]), .Z(n1833) );
  XNOR U2163 ( .A(n1838), .B(n1749), .Z(n1751) );
  XOR U2164 ( .A(n1839), .B(n1840), .Z(n1749) );
  ANDN U2165 ( .B(n1841), .A(n1842), .Z(n1839) );
  AND U2166 ( .A(b[9]), .B(a[32]), .Z(n1838) );
  XNOR U2167 ( .A(n1843), .B(n1754), .Z(n1756) );
  XOR U2168 ( .A(n1844), .B(n1845), .Z(n1754) );
  ANDN U2169 ( .B(n1846), .A(n1847), .Z(n1844) );
  AND U2170 ( .A(b[8]), .B(a[33]), .Z(n1843) );
  XNOR U2171 ( .A(n1848), .B(n1759), .Z(n1761) );
  XOR U2172 ( .A(n1849), .B(n1850), .Z(n1759) );
  ANDN U2173 ( .B(n1851), .A(n1852), .Z(n1849) );
  AND U2174 ( .A(b[7]), .B(a[34]), .Z(n1848) );
  XNOR U2175 ( .A(n1853), .B(n1764), .Z(n1766) );
  XOR U2176 ( .A(n1854), .B(n1855), .Z(n1764) );
  ANDN U2177 ( .B(n1856), .A(n1857), .Z(n1854) );
  AND U2178 ( .A(b[6]), .B(a[35]), .Z(n1853) );
  XNOR U2179 ( .A(n1858), .B(n1769), .Z(n1771) );
  XOR U2180 ( .A(n1859), .B(n1860), .Z(n1769) );
  ANDN U2181 ( .B(n1861), .A(n1862), .Z(n1859) );
  AND U2182 ( .A(b[5]), .B(a[36]), .Z(n1858) );
  XNOR U2183 ( .A(n1863), .B(n1774), .Z(n1776) );
  XOR U2184 ( .A(n1864), .B(n1865), .Z(n1774) );
  ANDN U2185 ( .B(n1866), .A(n1867), .Z(n1864) );
  AND U2186 ( .A(b[4]), .B(a[37]), .Z(n1863) );
  XNOR U2187 ( .A(n1868), .B(n1869), .Z(n1788) );
  NANDN U2188 ( .A(n1870), .B(n1871), .Z(n1869) );
  XNOR U2189 ( .A(n1872), .B(n1779), .Z(n1781) );
  XNOR U2190 ( .A(n1873), .B(n1874), .Z(n1779) );
  AND U2191 ( .A(n1875), .B(n1876), .Z(n1873) );
  AND U2192 ( .A(b[3]), .B(a[38]), .Z(n1872) );
  XOR U2193 ( .A(n1795), .B(n1794), .Z(swire[40]) );
  XOR U2194 ( .A(sreg[104]), .B(n1793), .Z(n1794) );
  XOR U2195 ( .A(n1800), .B(n1877), .Z(n1795) );
  XNOR U2196 ( .A(n1799), .B(n1793), .Z(n1877) );
  XOR U2197 ( .A(n1878), .B(n1879), .Z(n1793) );
  NOR U2198 ( .A(n1880), .B(n1881), .Z(n1878) );
  NAND U2199 ( .A(a[40]), .B(b[0]), .Z(n1799) );
  XNOR U2200 ( .A(n1870), .B(n1871), .Z(n1800) );
  XOR U2201 ( .A(n1868), .B(n1882), .Z(n1871) );
  NAND U2202 ( .A(b[1]), .B(a[39]), .Z(n1882) );
  XOR U2203 ( .A(n1876), .B(n1883), .Z(n1870) );
  XOR U2204 ( .A(n1868), .B(n1875), .Z(n1883) );
  XNOR U2205 ( .A(n1884), .B(n1874), .Z(n1875) );
  AND U2206 ( .A(b[2]), .B(a[38]), .Z(n1884) );
  NANDN U2207 ( .A(n1885), .B(n1886), .Z(n1868) );
  XOR U2208 ( .A(n1874), .B(n1866), .Z(n1887) );
  XNOR U2209 ( .A(n1865), .B(n1861), .Z(n1888) );
  XNOR U2210 ( .A(n1860), .B(n1856), .Z(n1889) );
  XNOR U2211 ( .A(n1855), .B(n1851), .Z(n1890) );
  XNOR U2212 ( .A(n1850), .B(n1846), .Z(n1891) );
  XNOR U2213 ( .A(n1845), .B(n1841), .Z(n1892) );
  XNOR U2214 ( .A(n1840), .B(n1836), .Z(n1893) );
  XNOR U2215 ( .A(n1835), .B(n1831), .Z(n1894) );
  XNOR U2216 ( .A(n1830), .B(n1826), .Z(n1895) );
  XOR U2217 ( .A(n1825), .B(n1822), .Z(n1896) );
  XOR U2218 ( .A(n1897), .B(n1898), .Z(n1822) );
  XOR U2219 ( .A(n1820), .B(n1899), .Z(n1898) );
  XOR U2220 ( .A(n1900), .B(n1901), .Z(n1899) );
  XOR U2221 ( .A(n1902), .B(n1903), .Z(n1901) );
  NAND U2222 ( .A(b[14]), .B(a[26]), .Z(n1903) );
  AND U2223 ( .A(b[15]), .B(a[25]), .Z(n1902) );
  XOR U2224 ( .A(n1904), .B(n1900), .Z(n1897) );
  XOR U2225 ( .A(n1905), .B(n1906), .Z(n1900) );
  NOR U2226 ( .A(n1907), .B(n1908), .Z(n1905) );
  AND U2227 ( .A(b[13]), .B(a[27]), .Z(n1904) );
  XNOR U2228 ( .A(n1909), .B(n1820), .Z(n1821) );
  XOR U2229 ( .A(n1910), .B(n1911), .Z(n1820) );
  ANDN U2230 ( .B(n1912), .A(n1913), .Z(n1910) );
  AND U2231 ( .A(b[12]), .B(a[28]), .Z(n1909) );
  XNOR U2232 ( .A(n1914), .B(n1825), .Z(n1827) );
  XOR U2233 ( .A(n1915), .B(n1916), .Z(n1825) );
  ANDN U2234 ( .B(n1917), .A(n1918), .Z(n1915) );
  AND U2235 ( .A(b[11]), .B(a[29]), .Z(n1914) );
  XNOR U2236 ( .A(n1919), .B(n1830), .Z(n1832) );
  XOR U2237 ( .A(n1920), .B(n1921), .Z(n1830) );
  ANDN U2238 ( .B(n1922), .A(n1923), .Z(n1920) );
  AND U2239 ( .A(b[10]), .B(a[30]), .Z(n1919) );
  XNOR U2240 ( .A(n1924), .B(n1835), .Z(n1837) );
  XOR U2241 ( .A(n1925), .B(n1926), .Z(n1835) );
  ANDN U2242 ( .B(n1927), .A(n1928), .Z(n1925) );
  AND U2243 ( .A(b[9]), .B(a[31]), .Z(n1924) );
  XNOR U2244 ( .A(n1929), .B(n1840), .Z(n1842) );
  XOR U2245 ( .A(n1930), .B(n1931), .Z(n1840) );
  ANDN U2246 ( .B(n1932), .A(n1933), .Z(n1930) );
  AND U2247 ( .A(b[8]), .B(a[32]), .Z(n1929) );
  XNOR U2248 ( .A(n1934), .B(n1845), .Z(n1847) );
  XOR U2249 ( .A(n1935), .B(n1936), .Z(n1845) );
  ANDN U2250 ( .B(n1937), .A(n1938), .Z(n1935) );
  AND U2251 ( .A(b[7]), .B(a[33]), .Z(n1934) );
  XNOR U2252 ( .A(n1939), .B(n1850), .Z(n1852) );
  XOR U2253 ( .A(n1940), .B(n1941), .Z(n1850) );
  ANDN U2254 ( .B(n1942), .A(n1943), .Z(n1940) );
  AND U2255 ( .A(b[6]), .B(a[34]), .Z(n1939) );
  XNOR U2256 ( .A(n1944), .B(n1855), .Z(n1857) );
  XOR U2257 ( .A(n1945), .B(n1946), .Z(n1855) );
  ANDN U2258 ( .B(n1947), .A(n1948), .Z(n1945) );
  AND U2259 ( .A(b[5]), .B(a[35]), .Z(n1944) );
  XNOR U2260 ( .A(n1949), .B(n1860), .Z(n1862) );
  XOR U2261 ( .A(n1950), .B(n1951), .Z(n1860) );
  ANDN U2262 ( .B(n1952), .A(n1953), .Z(n1950) );
  AND U2263 ( .A(b[4]), .B(a[36]), .Z(n1949) );
  XNOR U2264 ( .A(n1954), .B(n1955), .Z(n1874) );
  NANDN U2265 ( .A(n1956), .B(n1957), .Z(n1955) );
  XNOR U2266 ( .A(n1958), .B(n1865), .Z(n1867) );
  XNOR U2267 ( .A(n1959), .B(n1960), .Z(n1865) );
  AND U2268 ( .A(n1961), .B(n1962), .Z(n1959) );
  AND U2269 ( .A(b[3]), .B(a[37]), .Z(n1958) );
  XOR U2270 ( .A(n1881), .B(n1880), .Z(swire[39]) );
  XOR U2271 ( .A(sreg[103]), .B(n1879), .Z(n1880) );
  XOR U2272 ( .A(n1886), .B(n1963), .Z(n1881) );
  XNOR U2273 ( .A(n1885), .B(n1879), .Z(n1963) );
  XOR U2274 ( .A(n1964), .B(n1965), .Z(n1879) );
  NOR U2275 ( .A(n1966), .B(n1967), .Z(n1964) );
  NAND U2276 ( .A(a[39]), .B(b[0]), .Z(n1885) );
  XNOR U2277 ( .A(n1956), .B(n1957), .Z(n1886) );
  XOR U2278 ( .A(n1954), .B(n1968), .Z(n1957) );
  NAND U2279 ( .A(b[1]), .B(a[38]), .Z(n1968) );
  XOR U2280 ( .A(n1962), .B(n1969), .Z(n1956) );
  XOR U2281 ( .A(n1954), .B(n1961), .Z(n1969) );
  XNOR U2282 ( .A(n1970), .B(n1960), .Z(n1961) );
  AND U2283 ( .A(b[2]), .B(a[37]), .Z(n1970) );
  NANDN U2284 ( .A(n1971), .B(n1972), .Z(n1954) );
  XOR U2285 ( .A(n1960), .B(n1952), .Z(n1973) );
  XNOR U2286 ( .A(n1951), .B(n1947), .Z(n1974) );
  XNOR U2287 ( .A(n1946), .B(n1942), .Z(n1975) );
  XNOR U2288 ( .A(n1941), .B(n1937), .Z(n1976) );
  XNOR U2289 ( .A(n1936), .B(n1932), .Z(n1977) );
  XNOR U2290 ( .A(n1931), .B(n1927), .Z(n1978) );
  XNOR U2291 ( .A(n1926), .B(n1922), .Z(n1979) );
  XNOR U2292 ( .A(n1921), .B(n1917), .Z(n1980) );
  XNOR U2293 ( .A(n1916), .B(n1912), .Z(n1981) );
  XOR U2294 ( .A(n1911), .B(n1908), .Z(n1982) );
  XOR U2295 ( .A(n1983), .B(n1984), .Z(n1908) );
  XOR U2296 ( .A(n1906), .B(n1985), .Z(n1984) );
  XOR U2297 ( .A(n1986), .B(n1987), .Z(n1985) );
  XOR U2298 ( .A(n1988), .B(n1989), .Z(n1987) );
  NAND U2299 ( .A(b[14]), .B(a[25]), .Z(n1989) );
  AND U2300 ( .A(b[15]), .B(a[24]), .Z(n1988) );
  XOR U2301 ( .A(n1990), .B(n1986), .Z(n1983) );
  XOR U2302 ( .A(n1991), .B(n1992), .Z(n1986) );
  NOR U2303 ( .A(n1993), .B(n1994), .Z(n1991) );
  AND U2304 ( .A(b[13]), .B(a[26]), .Z(n1990) );
  XNOR U2305 ( .A(n1995), .B(n1906), .Z(n1907) );
  XOR U2306 ( .A(n1996), .B(n1997), .Z(n1906) );
  ANDN U2307 ( .B(n1998), .A(n1999), .Z(n1996) );
  AND U2308 ( .A(b[12]), .B(a[27]), .Z(n1995) );
  XNOR U2309 ( .A(n2000), .B(n1911), .Z(n1913) );
  XOR U2310 ( .A(n2001), .B(n2002), .Z(n1911) );
  ANDN U2311 ( .B(n2003), .A(n2004), .Z(n2001) );
  AND U2312 ( .A(b[11]), .B(a[28]), .Z(n2000) );
  XNOR U2313 ( .A(n2005), .B(n1916), .Z(n1918) );
  XOR U2314 ( .A(n2006), .B(n2007), .Z(n1916) );
  ANDN U2315 ( .B(n2008), .A(n2009), .Z(n2006) );
  AND U2316 ( .A(b[10]), .B(a[29]), .Z(n2005) );
  XNOR U2317 ( .A(n2010), .B(n1921), .Z(n1923) );
  XOR U2318 ( .A(n2011), .B(n2012), .Z(n1921) );
  ANDN U2319 ( .B(n2013), .A(n2014), .Z(n2011) );
  AND U2320 ( .A(b[9]), .B(a[30]), .Z(n2010) );
  XNOR U2321 ( .A(n2015), .B(n1926), .Z(n1928) );
  XOR U2322 ( .A(n2016), .B(n2017), .Z(n1926) );
  ANDN U2323 ( .B(n2018), .A(n2019), .Z(n2016) );
  AND U2324 ( .A(b[8]), .B(a[31]), .Z(n2015) );
  XNOR U2325 ( .A(n2020), .B(n1931), .Z(n1933) );
  XOR U2326 ( .A(n2021), .B(n2022), .Z(n1931) );
  ANDN U2327 ( .B(n2023), .A(n2024), .Z(n2021) );
  AND U2328 ( .A(b[7]), .B(a[32]), .Z(n2020) );
  XNOR U2329 ( .A(n2025), .B(n1936), .Z(n1938) );
  XOR U2330 ( .A(n2026), .B(n2027), .Z(n1936) );
  ANDN U2331 ( .B(n2028), .A(n2029), .Z(n2026) );
  AND U2332 ( .A(b[6]), .B(a[33]), .Z(n2025) );
  XNOR U2333 ( .A(n2030), .B(n1941), .Z(n1943) );
  XOR U2334 ( .A(n2031), .B(n2032), .Z(n1941) );
  ANDN U2335 ( .B(n2033), .A(n2034), .Z(n2031) );
  AND U2336 ( .A(b[5]), .B(a[34]), .Z(n2030) );
  XNOR U2337 ( .A(n2035), .B(n1946), .Z(n1948) );
  XOR U2338 ( .A(n2036), .B(n2037), .Z(n1946) );
  ANDN U2339 ( .B(n2038), .A(n2039), .Z(n2036) );
  AND U2340 ( .A(b[4]), .B(a[35]), .Z(n2035) );
  XNOR U2341 ( .A(n2040), .B(n2041), .Z(n1960) );
  NANDN U2342 ( .A(n2042), .B(n2043), .Z(n2041) );
  XNOR U2343 ( .A(n2044), .B(n1951), .Z(n1953) );
  XNOR U2344 ( .A(n2045), .B(n2046), .Z(n1951) );
  AND U2345 ( .A(n2047), .B(n2048), .Z(n2045) );
  AND U2346 ( .A(b[3]), .B(a[36]), .Z(n2044) );
  XOR U2347 ( .A(n1967), .B(n1966), .Z(swire[38]) );
  XOR U2348 ( .A(sreg[102]), .B(n1965), .Z(n1966) );
  XOR U2349 ( .A(n1972), .B(n2049), .Z(n1967) );
  XNOR U2350 ( .A(n1971), .B(n1965), .Z(n2049) );
  XOR U2351 ( .A(n2050), .B(n2051), .Z(n1965) );
  NOR U2352 ( .A(n2052), .B(n2053), .Z(n2050) );
  NAND U2353 ( .A(a[38]), .B(b[0]), .Z(n1971) );
  XNOR U2354 ( .A(n2042), .B(n2043), .Z(n1972) );
  XOR U2355 ( .A(n2040), .B(n2054), .Z(n2043) );
  NAND U2356 ( .A(b[1]), .B(a[37]), .Z(n2054) );
  XOR U2357 ( .A(n2048), .B(n2055), .Z(n2042) );
  XOR U2358 ( .A(n2040), .B(n2047), .Z(n2055) );
  XNOR U2359 ( .A(n2056), .B(n2046), .Z(n2047) );
  AND U2360 ( .A(b[2]), .B(a[36]), .Z(n2056) );
  NANDN U2361 ( .A(n2057), .B(n2058), .Z(n2040) );
  XOR U2362 ( .A(n2046), .B(n2038), .Z(n2059) );
  XNOR U2363 ( .A(n2037), .B(n2033), .Z(n2060) );
  XNOR U2364 ( .A(n2032), .B(n2028), .Z(n2061) );
  XNOR U2365 ( .A(n2027), .B(n2023), .Z(n2062) );
  XNOR U2366 ( .A(n2022), .B(n2018), .Z(n2063) );
  XNOR U2367 ( .A(n2017), .B(n2013), .Z(n2064) );
  XNOR U2368 ( .A(n2012), .B(n2008), .Z(n2065) );
  XNOR U2369 ( .A(n2007), .B(n2003), .Z(n2066) );
  XNOR U2370 ( .A(n2002), .B(n1998), .Z(n2067) );
  XOR U2371 ( .A(n1997), .B(n1994), .Z(n2068) );
  XOR U2372 ( .A(n2069), .B(n2070), .Z(n1994) );
  XOR U2373 ( .A(n1992), .B(n2071), .Z(n2070) );
  XOR U2374 ( .A(n2072), .B(n2073), .Z(n2071) );
  XOR U2375 ( .A(n2074), .B(n2075), .Z(n2073) );
  NAND U2376 ( .A(b[14]), .B(a[24]), .Z(n2075) );
  AND U2377 ( .A(b[15]), .B(a[23]), .Z(n2074) );
  XOR U2378 ( .A(n2076), .B(n2072), .Z(n2069) );
  XOR U2379 ( .A(n2077), .B(n2078), .Z(n2072) );
  NOR U2380 ( .A(n2079), .B(n2080), .Z(n2077) );
  AND U2381 ( .A(b[13]), .B(a[25]), .Z(n2076) );
  XNOR U2382 ( .A(n2081), .B(n1992), .Z(n1993) );
  XOR U2383 ( .A(n2082), .B(n2083), .Z(n1992) );
  ANDN U2384 ( .B(n2084), .A(n2085), .Z(n2082) );
  AND U2385 ( .A(b[12]), .B(a[26]), .Z(n2081) );
  XNOR U2386 ( .A(n2086), .B(n1997), .Z(n1999) );
  XOR U2387 ( .A(n2087), .B(n2088), .Z(n1997) );
  ANDN U2388 ( .B(n2089), .A(n2090), .Z(n2087) );
  AND U2389 ( .A(b[11]), .B(a[27]), .Z(n2086) );
  XNOR U2390 ( .A(n2091), .B(n2002), .Z(n2004) );
  XOR U2391 ( .A(n2092), .B(n2093), .Z(n2002) );
  ANDN U2392 ( .B(n2094), .A(n2095), .Z(n2092) );
  AND U2393 ( .A(b[10]), .B(a[28]), .Z(n2091) );
  XNOR U2394 ( .A(n2096), .B(n2007), .Z(n2009) );
  XOR U2395 ( .A(n2097), .B(n2098), .Z(n2007) );
  ANDN U2396 ( .B(n2099), .A(n2100), .Z(n2097) );
  AND U2397 ( .A(b[9]), .B(a[29]), .Z(n2096) );
  XNOR U2398 ( .A(n2101), .B(n2012), .Z(n2014) );
  XOR U2399 ( .A(n2102), .B(n2103), .Z(n2012) );
  ANDN U2400 ( .B(n2104), .A(n2105), .Z(n2102) );
  AND U2401 ( .A(b[8]), .B(a[30]), .Z(n2101) );
  XNOR U2402 ( .A(n2106), .B(n2017), .Z(n2019) );
  XOR U2403 ( .A(n2107), .B(n2108), .Z(n2017) );
  ANDN U2404 ( .B(n2109), .A(n2110), .Z(n2107) );
  AND U2405 ( .A(b[7]), .B(a[31]), .Z(n2106) );
  XNOR U2406 ( .A(n2111), .B(n2022), .Z(n2024) );
  XOR U2407 ( .A(n2112), .B(n2113), .Z(n2022) );
  ANDN U2408 ( .B(n2114), .A(n2115), .Z(n2112) );
  AND U2409 ( .A(b[6]), .B(a[32]), .Z(n2111) );
  XNOR U2410 ( .A(n2116), .B(n2027), .Z(n2029) );
  XOR U2411 ( .A(n2117), .B(n2118), .Z(n2027) );
  ANDN U2412 ( .B(n2119), .A(n2120), .Z(n2117) );
  AND U2413 ( .A(b[5]), .B(a[33]), .Z(n2116) );
  XNOR U2414 ( .A(n2121), .B(n2032), .Z(n2034) );
  XOR U2415 ( .A(n2122), .B(n2123), .Z(n2032) );
  ANDN U2416 ( .B(n2124), .A(n2125), .Z(n2122) );
  AND U2417 ( .A(b[4]), .B(a[34]), .Z(n2121) );
  XNOR U2418 ( .A(n2126), .B(n2127), .Z(n2046) );
  NANDN U2419 ( .A(n2128), .B(n2129), .Z(n2127) );
  XNOR U2420 ( .A(n2130), .B(n2037), .Z(n2039) );
  XNOR U2421 ( .A(n2131), .B(n2132), .Z(n2037) );
  AND U2422 ( .A(n2133), .B(n2134), .Z(n2131) );
  AND U2423 ( .A(b[3]), .B(a[35]), .Z(n2130) );
  XOR U2424 ( .A(n2053), .B(n2052), .Z(swire[37]) );
  XOR U2425 ( .A(sreg[101]), .B(n2051), .Z(n2052) );
  XOR U2426 ( .A(n2058), .B(n2135), .Z(n2053) );
  XNOR U2427 ( .A(n2057), .B(n2051), .Z(n2135) );
  XOR U2428 ( .A(n2136), .B(n2137), .Z(n2051) );
  NOR U2429 ( .A(n2138), .B(n2139), .Z(n2136) );
  NAND U2430 ( .A(a[37]), .B(b[0]), .Z(n2057) );
  XNOR U2431 ( .A(n2128), .B(n2129), .Z(n2058) );
  XOR U2432 ( .A(n2126), .B(n2140), .Z(n2129) );
  NAND U2433 ( .A(b[1]), .B(a[36]), .Z(n2140) );
  XOR U2434 ( .A(n2134), .B(n2141), .Z(n2128) );
  XOR U2435 ( .A(n2126), .B(n2133), .Z(n2141) );
  XNOR U2436 ( .A(n2142), .B(n2132), .Z(n2133) );
  AND U2437 ( .A(b[2]), .B(a[35]), .Z(n2142) );
  NANDN U2438 ( .A(n2143), .B(n2144), .Z(n2126) );
  XOR U2439 ( .A(n2132), .B(n2124), .Z(n2145) );
  XNOR U2440 ( .A(n2123), .B(n2119), .Z(n2146) );
  XNOR U2441 ( .A(n2118), .B(n2114), .Z(n2147) );
  XNOR U2442 ( .A(n2113), .B(n2109), .Z(n2148) );
  XNOR U2443 ( .A(n2108), .B(n2104), .Z(n2149) );
  XNOR U2444 ( .A(n2103), .B(n2099), .Z(n2150) );
  XNOR U2445 ( .A(n2098), .B(n2094), .Z(n2151) );
  XNOR U2446 ( .A(n2093), .B(n2089), .Z(n2152) );
  XNOR U2447 ( .A(n2088), .B(n2084), .Z(n2153) );
  XOR U2448 ( .A(n2083), .B(n2080), .Z(n2154) );
  XOR U2449 ( .A(n2155), .B(n2156), .Z(n2080) );
  XOR U2450 ( .A(n2078), .B(n2157), .Z(n2156) );
  XOR U2451 ( .A(n2158), .B(n2159), .Z(n2157) );
  XOR U2452 ( .A(n2160), .B(n2161), .Z(n2159) );
  NAND U2453 ( .A(b[14]), .B(a[23]), .Z(n2161) );
  AND U2454 ( .A(b[15]), .B(a[22]), .Z(n2160) );
  XOR U2455 ( .A(n2162), .B(n2158), .Z(n2155) );
  XOR U2456 ( .A(n2163), .B(n2164), .Z(n2158) );
  NOR U2457 ( .A(n2165), .B(n2166), .Z(n2163) );
  AND U2458 ( .A(b[13]), .B(a[24]), .Z(n2162) );
  XNOR U2459 ( .A(n2167), .B(n2078), .Z(n2079) );
  XOR U2460 ( .A(n2168), .B(n2169), .Z(n2078) );
  ANDN U2461 ( .B(n2170), .A(n2171), .Z(n2168) );
  AND U2462 ( .A(b[12]), .B(a[25]), .Z(n2167) );
  XNOR U2463 ( .A(n2172), .B(n2083), .Z(n2085) );
  XOR U2464 ( .A(n2173), .B(n2174), .Z(n2083) );
  ANDN U2465 ( .B(n2175), .A(n2176), .Z(n2173) );
  AND U2466 ( .A(b[11]), .B(a[26]), .Z(n2172) );
  XNOR U2467 ( .A(n2177), .B(n2088), .Z(n2090) );
  XOR U2468 ( .A(n2178), .B(n2179), .Z(n2088) );
  ANDN U2469 ( .B(n2180), .A(n2181), .Z(n2178) );
  AND U2470 ( .A(b[10]), .B(a[27]), .Z(n2177) );
  XNOR U2471 ( .A(n2182), .B(n2093), .Z(n2095) );
  XOR U2472 ( .A(n2183), .B(n2184), .Z(n2093) );
  ANDN U2473 ( .B(n2185), .A(n2186), .Z(n2183) );
  AND U2474 ( .A(b[9]), .B(a[28]), .Z(n2182) );
  XNOR U2475 ( .A(n2187), .B(n2098), .Z(n2100) );
  XOR U2476 ( .A(n2188), .B(n2189), .Z(n2098) );
  ANDN U2477 ( .B(n2190), .A(n2191), .Z(n2188) );
  AND U2478 ( .A(b[8]), .B(a[29]), .Z(n2187) );
  XNOR U2479 ( .A(n2192), .B(n2103), .Z(n2105) );
  XOR U2480 ( .A(n2193), .B(n2194), .Z(n2103) );
  ANDN U2481 ( .B(n2195), .A(n2196), .Z(n2193) );
  AND U2482 ( .A(b[7]), .B(a[30]), .Z(n2192) );
  XNOR U2483 ( .A(n2197), .B(n2108), .Z(n2110) );
  XOR U2484 ( .A(n2198), .B(n2199), .Z(n2108) );
  ANDN U2485 ( .B(n2200), .A(n2201), .Z(n2198) );
  AND U2486 ( .A(b[6]), .B(a[31]), .Z(n2197) );
  XNOR U2487 ( .A(n2202), .B(n2113), .Z(n2115) );
  XOR U2488 ( .A(n2203), .B(n2204), .Z(n2113) );
  ANDN U2489 ( .B(n2205), .A(n2206), .Z(n2203) );
  AND U2490 ( .A(b[5]), .B(a[32]), .Z(n2202) );
  XNOR U2491 ( .A(n2207), .B(n2118), .Z(n2120) );
  XOR U2492 ( .A(n2208), .B(n2209), .Z(n2118) );
  ANDN U2493 ( .B(n2210), .A(n2211), .Z(n2208) );
  AND U2494 ( .A(b[4]), .B(a[33]), .Z(n2207) );
  XNOR U2495 ( .A(n2212), .B(n2213), .Z(n2132) );
  NANDN U2496 ( .A(n2214), .B(n2215), .Z(n2213) );
  XNOR U2497 ( .A(n2216), .B(n2123), .Z(n2125) );
  XNOR U2498 ( .A(n2217), .B(n2218), .Z(n2123) );
  AND U2499 ( .A(n2219), .B(n2220), .Z(n2217) );
  AND U2500 ( .A(b[3]), .B(a[34]), .Z(n2216) );
  XOR U2501 ( .A(n2139), .B(n2138), .Z(swire[36]) );
  XOR U2502 ( .A(sreg[100]), .B(n2137), .Z(n2138) );
  XOR U2503 ( .A(n2144), .B(n2221), .Z(n2139) );
  XNOR U2504 ( .A(n2143), .B(n2137), .Z(n2221) );
  XOR U2505 ( .A(n2222), .B(n2223), .Z(n2137) );
  NOR U2506 ( .A(n2224), .B(n2225), .Z(n2222) );
  NAND U2507 ( .A(a[36]), .B(b[0]), .Z(n2143) );
  XNOR U2508 ( .A(n2214), .B(n2215), .Z(n2144) );
  XOR U2509 ( .A(n2212), .B(n2226), .Z(n2215) );
  NAND U2510 ( .A(b[1]), .B(a[35]), .Z(n2226) );
  XOR U2511 ( .A(n2220), .B(n2227), .Z(n2214) );
  XOR U2512 ( .A(n2212), .B(n2219), .Z(n2227) );
  XNOR U2513 ( .A(n2228), .B(n2218), .Z(n2219) );
  AND U2514 ( .A(b[2]), .B(a[34]), .Z(n2228) );
  NANDN U2515 ( .A(n2229), .B(n2230), .Z(n2212) );
  XOR U2516 ( .A(n2218), .B(n2210), .Z(n2231) );
  XNOR U2517 ( .A(n2209), .B(n2205), .Z(n2232) );
  XNOR U2518 ( .A(n2204), .B(n2200), .Z(n2233) );
  XNOR U2519 ( .A(n2199), .B(n2195), .Z(n2234) );
  XNOR U2520 ( .A(n2194), .B(n2190), .Z(n2235) );
  XNOR U2521 ( .A(n2189), .B(n2185), .Z(n2236) );
  XNOR U2522 ( .A(n2184), .B(n2180), .Z(n2237) );
  XNOR U2523 ( .A(n2179), .B(n2175), .Z(n2238) );
  XNOR U2524 ( .A(n2174), .B(n2170), .Z(n2239) );
  XOR U2525 ( .A(n2169), .B(n2166), .Z(n2240) );
  XOR U2526 ( .A(n2241), .B(n2242), .Z(n2166) );
  XOR U2527 ( .A(n2164), .B(n2243), .Z(n2242) );
  XOR U2528 ( .A(n2244), .B(n2245), .Z(n2243) );
  XOR U2529 ( .A(n2246), .B(n2247), .Z(n2245) );
  NAND U2530 ( .A(b[14]), .B(a[22]), .Z(n2247) );
  AND U2531 ( .A(b[15]), .B(a[21]), .Z(n2246) );
  XOR U2532 ( .A(n2248), .B(n2244), .Z(n2241) );
  XOR U2533 ( .A(n2249), .B(n2250), .Z(n2244) );
  NOR U2534 ( .A(n2251), .B(n2252), .Z(n2249) );
  AND U2535 ( .A(b[13]), .B(a[23]), .Z(n2248) );
  XNOR U2536 ( .A(n2253), .B(n2164), .Z(n2165) );
  XOR U2537 ( .A(n2254), .B(n2255), .Z(n2164) );
  ANDN U2538 ( .B(n2256), .A(n2257), .Z(n2254) );
  AND U2539 ( .A(b[12]), .B(a[24]), .Z(n2253) );
  XNOR U2540 ( .A(n2258), .B(n2169), .Z(n2171) );
  XOR U2541 ( .A(n2259), .B(n2260), .Z(n2169) );
  ANDN U2542 ( .B(n2261), .A(n2262), .Z(n2259) );
  AND U2543 ( .A(b[11]), .B(a[25]), .Z(n2258) );
  XNOR U2544 ( .A(n2263), .B(n2174), .Z(n2176) );
  XOR U2545 ( .A(n2264), .B(n2265), .Z(n2174) );
  ANDN U2546 ( .B(n2266), .A(n2267), .Z(n2264) );
  AND U2547 ( .A(b[10]), .B(a[26]), .Z(n2263) );
  XNOR U2548 ( .A(n2268), .B(n2179), .Z(n2181) );
  XOR U2549 ( .A(n2269), .B(n2270), .Z(n2179) );
  ANDN U2550 ( .B(n2271), .A(n2272), .Z(n2269) );
  AND U2551 ( .A(b[9]), .B(a[27]), .Z(n2268) );
  XNOR U2552 ( .A(n2273), .B(n2184), .Z(n2186) );
  XOR U2553 ( .A(n2274), .B(n2275), .Z(n2184) );
  ANDN U2554 ( .B(n2276), .A(n2277), .Z(n2274) );
  AND U2555 ( .A(b[8]), .B(a[28]), .Z(n2273) );
  XNOR U2556 ( .A(n2278), .B(n2189), .Z(n2191) );
  XOR U2557 ( .A(n2279), .B(n2280), .Z(n2189) );
  ANDN U2558 ( .B(n2281), .A(n2282), .Z(n2279) );
  AND U2559 ( .A(b[7]), .B(a[29]), .Z(n2278) );
  XNOR U2560 ( .A(n2283), .B(n2194), .Z(n2196) );
  XOR U2561 ( .A(n2284), .B(n2285), .Z(n2194) );
  ANDN U2562 ( .B(n2286), .A(n2287), .Z(n2284) );
  AND U2563 ( .A(b[6]), .B(a[30]), .Z(n2283) );
  XNOR U2564 ( .A(n2288), .B(n2199), .Z(n2201) );
  XOR U2565 ( .A(n2289), .B(n2290), .Z(n2199) );
  ANDN U2566 ( .B(n2291), .A(n2292), .Z(n2289) );
  AND U2567 ( .A(b[5]), .B(a[31]), .Z(n2288) );
  XNOR U2568 ( .A(n2293), .B(n2204), .Z(n2206) );
  XOR U2569 ( .A(n2294), .B(n2295), .Z(n2204) );
  ANDN U2570 ( .B(n2296), .A(n2297), .Z(n2294) );
  AND U2571 ( .A(b[4]), .B(a[32]), .Z(n2293) );
  XNOR U2572 ( .A(n2298), .B(n2299), .Z(n2218) );
  NANDN U2573 ( .A(n2300), .B(n2301), .Z(n2299) );
  XNOR U2574 ( .A(n2302), .B(n2209), .Z(n2211) );
  XNOR U2575 ( .A(n2303), .B(n2304), .Z(n2209) );
  AND U2576 ( .A(n2305), .B(n2306), .Z(n2303) );
  AND U2577 ( .A(b[3]), .B(a[33]), .Z(n2302) );
  XOR U2578 ( .A(n2225), .B(n2224), .Z(swire[35]) );
  XOR U2579 ( .A(sreg[99]), .B(n2223), .Z(n2224) );
  XOR U2580 ( .A(n2230), .B(n2307), .Z(n2225) );
  XNOR U2581 ( .A(n2229), .B(n2223), .Z(n2307) );
  XOR U2582 ( .A(n2308), .B(n2309), .Z(n2223) );
  NOR U2583 ( .A(n2310), .B(n2311), .Z(n2308) );
  NAND U2584 ( .A(a[35]), .B(b[0]), .Z(n2229) );
  XNOR U2585 ( .A(n2300), .B(n2301), .Z(n2230) );
  XOR U2586 ( .A(n2298), .B(n2312), .Z(n2301) );
  NAND U2587 ( .A(b[1]), .B(a[34]), .Z(n2312) );
  XOR U2588 ( .A(n2306), .B(n2313), .Z(n2300) );
  XOR U2589 ( .A(n2298), .B(n2305), .Z(n2313) );
  XNOR U2590 ( .A(n2314), .B(n2304), .Z(n2305) );
  AND U2591 ( .A(b[2]), .B(a[33]), .Z(n2314) );
  NANDN U2592 ( .A(n2315), .B(n2316), .Z(n2298) );
  XOR U2593 ( .A(n2304), .B(n2296), .Z(n2317) );
  XNOR U2594 ( .A(n2295), .B(n2291), .Z(n2318) );
  XNOR U2595 ( .A(n2290), .B(n2286), .Z(n2319) );
  XNOR U2596 ( .A(n2285), .B(n2281), .Z(n2320) );
  XNOR U2597 ( .A(n2280), .B(n2276), .Z(n2321) );
  XNOR U2598 ( .A(n2275), .B(n2271), .Z(n2322) );
  XNOR U2599 ( .A(n2270), .B(n2266), .Z(n2323) );
  XNOR U2600 ( .A(n2265), .B(n2261), .Z(n2324) );
  XNOR U2601 ( .A(n2260), .B(n2256), .Z(n2325) );
  XOR U2602 ( .A(n2255), .B(n2252), .Z(n2326) );
  XOR U2603 ( .A(n2327), .B(n2328), .Z(n2252) );
  XOR U2604 ( .A(n2250), .B(n2329), .Z(n2328) );
  XOR U2605 ( .A(n2330), .B(n2331), .Z(n2329) );
  XOR U2606 ( .A(n2332), .B(n2333), .Z(n2331) );
  NAND U2607 ( .A(b[14]), .B(a[21]), .Z(n2333) );
  AND U2608 ( .A(b[15]), .B(a[20]), .Z(n2332) );
  XOR U2609 ( .A(n2334), .B(n2330), .Z(n2327) );
  XOR U2610 ( .A(n2335), .B(n2336), .Z(n2330) );
  NOR U2611 ( .A(n2337), .B(n2338), .Z(n2335) );
  AND U2612 ( .A(b[13]), .B(a[22]), .Z(n2334) );
  XNOR U2613 ( .A(n2339), .B(n2250), .Z(n2251) );
  XOR U2614 ( .A(n2340), .B(n2341), .Z(n2250) );
  ANDN U2615 ( .B(n2342), .A(n2343), .Z(n2340) );
  AND U2616 ( .A(b[12]), .B(a[23]), .Z(n2339) );
  XNOR U2617 ( .A(n2344), .B(n2255), .Z(n2257) );
  XOR U2618 ( .A(n2345), .B(n2346), .Z(n2255) );
  ANDN U2619 ( .B(n2347), .A(n2348), .Z(n2345) );
  AND U2620 ( .A(b[11]), .B(a[24]), .Z(n2344) );
  XNOR U2621 ( .A(n2349), .B(n2260), .Z(n2262) );
  XOR U2622 ( .A(n2350), .B(n2351), .Z(n2260) );
  ANDN U2623 ( .B(n2352), .A(n2353), .Z(n2350) );
  AND U2624 ( .A(b[10]), .B(a[25]), .Z(n2349) );
  XNOR U2625 ( .A(n2354), .B(n2265), .Z(n2267) );
  XOR U2626 ( .A(n2355), .B(n2356), .Z(n2265) );
  ANDN U2627 ( .B(n2357), .A(n2358), .Z(n2355) );
  AND U2628 ( .A(b[9]), .B(a[26]), .Z(n2354) );
  XNOR U2629 ( .A(n2359), .B(n2270), .Z(n2272) );
  XOR U2630 ( .A(n2360), .B(n2361), .Z(n2270) );
  ANDN U2631 ( .B(n2362), .A(n2363), .Z(n2360) );
  AND U2632 ( .A(b[8]), .B(a[27]), .Z(n2359) );
  XNOR U2633 ( .A(n2364), .B(n2275), .Z(n2277) );
  XOR U2634 ( .A(n2365), .B(n2366), .Z(n2275) );
  ANDN U2635 ( .B(n2367), .A(n2368), .Z(n2365) );
  AND U2636 ( .A(b[7]), .B(a[28]), .Z(n2364) );
  XNOR U2637 ( .A(n2369), .B(n2280), .Z(n2282) );
  XOR U2638 ( .A(n2370), .B(n2371), .Z(n2280) );
  ANDN U2639 ( .B(n2372), .A(n2373), .Z(n2370) );
  AND U2640 ( .A(b[6]), .B(a[29]), .Z(n2369) );
  XNOR U2641 ( .A(n2374), .B(n2285), .Z(n2287) );
  XOR U2642 ( .A(n2375), .B(n2376), .Z(n2285) );
  ANDN U2643 ( .B(n2377), .A(n2378), .Z(n2375) );
  AND U2644 ( .A(b[5]), .B(a[30]), .Z(n2374) );
  XNOR U2645 ( .A(n2379), .B(n2290), .Z(n2292) );
  XOR U2646 ( .A(n2380), .B(n2381), .Z(n2290) );
  ANDN U2647 ( .B(n2382), .A(n2383), .Z(n2380) );
  AND U2648 ( .A(b[4]), .B(a[31]), .Z(n2379) );
  XNOR U2649 ( .A(n2384), .B(n2385), .Z(n2304) );
  NANDN U2650 ( .A(n2386), .B(n2387), .Z(n2385) );
  XNOR U2651 ( .A(n2388), .B(n2295), .Z(n2297) );
  XNOR U2652 ( .A(n2389), .B(n2390), .Z(n2295) );
  AND U2653 ( .A(n2391), .B(n2392), .Z(n2389) );
  AND U2654 ( .A(b[3]), .B(a[32]), .Z(n2388) );
  XOR U2655 ( .A(n2311), .B(n2310), .Z(swire[34]) );
  XOR U2656 ( .A(sreg[98]), .B(n2309), .Z(n2310) );
  XOR U2657 ( .A(n2316), .B(n2393), .Z(n2311) );
  XNOR U2658 ( .A(n2315), .B(n2309), .Z(n2393) );
  XOR U2659 ( .A(n2394), .B(n2395), .Z(n2309) );
  NOR U2660 ( .A(n2396), .B(n2397), .Z(n2394) );
  NAND U2661 ( .A(a[34]), .B(b[0]), .Z(n2315) );
  XNOR U2662 ( .A(n2386), .B(n2387), .Z(n2316) );
  XOR U2663 ( .A(n2384), .B(n2398), .Z(n2387) );
  NAND U2664 ( .A(b[1]), .B(a[33]), .Z(n2398) );
  XOR U2665 ( .A(n2392), .B(n2399), .Z(n2386) );
  XOR U2666 ( .A(n2384), .B(n2391), .Z(n2399) );
  XNOR U2667 ( .A(n2400), .B(n2390), .Z(n2391) );
  AND U2668 ( .A(b[2]), .B(a[32]), .Z(n2400) );
  NANDN U2669 ( .A(n2401), .B(n2402), .Z(n2384) );
  XOR U2670 ( .A(n2390), .B(n2382), .Z(n2403) );
  XNOR U2671 ( .A(n2381), .B(n2377), .Z(n2404) );
  XNOR U2672 ( .A(n2376), .B(n2372), .Z(n2405) );
  XNOR U2673 ( .A(n2371), .B(n2367), .Z(n2406) );
  XNOR U2674 ( .A(n2366), .B(n2362), .Z(n2407) );
  XNOR U2675 ( .A(n2361), .B(n2357), .Z(n2408) );
  XNOR U2676 ( .A(n2356), .B(n2352), .Z(n2409) );
  XNOR U2677 ( .A(n2351), .B(n2347), .Z(n2410) );
  XNOR U2678 ( .A(n2346), .B(n2342), .Z(n2411) );
  XOR U2679 ( .A(n2341), .B(n2338), .Z(n2412) );
  XOR U2680 ( .A(n2413), .B(n2414), .Z(n2338) );
  XOR U2681 ( .A(n2336), .B(n2415), .Z(n2414) );
  XOR U2682 ( .A(n2416), .B(n2417), .Z(n2415) );
  XOR U2683 ( .A(n2418), .B(n2419), .Z(n2417) );
  NAND U2684 ( .A(b[14]), .B(a[20]), .Z(n2419) );
  AND U2685 ( .A(b[15]), .B(a[19]), .Z(n2418) );
  XOR U2686 ( .A(n2420), .B(n2416), .Z(n2413) );
  XOR U2687 ( .A(n2421), .B(n2422), .Z(n2416) );
  NOR U2688 ( .A(n2423), .B(n2424), .Z(n2421) );
  AND U2689 ( .A(b[13]), .B(a[21]), .Z(n2420) );
  XNOR U2690 ( .A(n2425), .B(n2336), .Z(n2337) );
  XOR U2691 ( .A(n2426), .B(n2427), .Z(n2336) );
  ANDN U2692 ( .B(n2428), .A(n2429), .Z(n2426) );
  AND U2693 ( .A(b[12]), .B(a[22]), .Z(n2425) );
  XNOR U2694 ( .A(n2430), .B(n2341), .Z(n2343) );
  XOR U2695 ( .A(n2431), .B(n2432), .Z(n2341) );
  ANDN U2696 ( .B(n2433), .A(n2434), .Z(n2431) );
  AND U2697 ( .A(b[11]), .B(a[23]), .Z(n2430) );
  XNOR U2698 ( .A(n2435), .B(n2346), .Z(n2348) );
  XOR U2699 ( .A(n2436), .B(n2437), .Z(n2346) );
  ANDN U2700 ( .B(n2438), .A(n2439), .Z(n2436) );
  AND U2701 ( .A(b[10]), .B(a[24]), .Z(n2435) );
  XNOR U2702 ( .A(n2440), .B(n2351), .Z(n2353) );
  XOR U2703 ( .A(n2441), .B(n2442), .Z(n2351) );
  ANDN U2704 ( .B(n2443), .A(n2444), .Z(n2441) );
  AND U2705 ( .A(b[9]), .B(a[25]), .Z(n2440) );
  XNOR U2706 ( .A(n2445), .B(n2356), .Z(n2358) );
  XOR U2707 ( .A(n2446), .B(n2447), .Z(n2356) );
  ANDN U2708 ( .B(n2448), .A(n2449), .Z(n2446) );
  AND U2709 ( .A(b[8]), .B(a[26]), .Z(n2445) );
  XNOR U2710 ( .A(n2450), .B(n2361), .Z(n2363) );
  XOR U2711 ( .A(n2451), .B(n2452), .Z(n2361) );
  ANDN U2712 ( .B(n2453), .A(n2454), .Z(n2451) );
  AND U2713 ( .A(b[7]), .B(a[27]), .Z(n2450) );
  XNOR U2714 ( .A(n2455), .B(n2366), .Z(n2368) );
  XOR U2715 ( .A(n2456), .B(n2457), .Z(n2366) );
  ANDN U2716 ( .B(n2458), .A(n2459), .Z(n2456) );
  AND U2717 ( .A(b[6]), .B(a[28]), .Z(n2455) );
  XNOR U2718 ( .A(n2460), .B(n2371), .Z(n2373) );
  XOR U2719 ( .A(n2461), .B(n2462), .Z(n2371) );
  ANDN U2720 ( .B(n2463), .A(n2464), .Z(n2461) );
  AND U2721 ( .A(b[5]), .B(a[29]), .Z(n2460) );
  XNOR U2722 ( .A(n2465), .B(n2376), .Z(n2378) );
  XOR U2723 ( .A(n2466), .B(n2467), .Z(n2376) );
  ANDN U2724 ( .B(n2468), .A(n2469), .Z(n2466) );
  AND U2725 ( .A(b[4]), .B(a[30]), .Z(n2465) );
  XNOR U2726 ( .A(n2470), .B(n2471), .Z(n2390) );
  NANDN U2727 ( .A(n2472), .B(n2473), .Z(n2471) );
  XNOR U2728 ( .A(n2474), .B(n2381), .Z(n2383) );
  XNOR U2729 ( .A(n2475), .B(n2476), .Z(n2381) );
  AND U2730 ( .A(n2477), .B(n2478), .Z(n2475) );
  AND U2731 ( .A(b[3]), .B(a[31]), .Z(n2474) );
  XOR U2732 ( .A(n2397), .B(n2396), .Z(swire[33]) );
  XOR U2733 ( .A(sreg[97]), .B(n2395), .Z(n2396) );
  XOR U2734 ( .A(n2402), .B(n2479), .Z(n2397) );
  XNOR U2735 ( .A(n2401), .B(n2395), .Z(n2479) );
  XOR U2736 ( .A(n2480), .B(n2481), .Z(n2395) );
  NOR U2737 ( .A(n2482), .B(n2483), .Z(n2480) );
  NAND U2738 ( .A(a[33]), .B(b[0]), .Z(n2401) );
  XNOR U2739 ( .A(n2472), .B(n2473), .Z(n2402) );
  XOR U2740 ( .A(n2470), .B(n2484), .Z(n2473) );
  NAND U2741 ( .A(b[1]), .B(a[32]), .Z(n2484) );
  XOR U2742 ( .A(n2478), .B(n2485), .Z(n2472) );
  XOR U2743 ( .A(n2470), .B(n2477), .Z(n2485) );
  XNOR U2744 ( .A(n2486), .B(n2476), .Z(n2477) );
  AND U2745 ( .A(b[2]), .B(a[31]), .Z(n2486) );
  NANDN U2746 ( .A(n2487), .B(n2488), .Z(n2470) );
  XOR U2747 ( .A(n2476), .B(n2468), .Z(n2489) );
  XNOR U2748 ( .A(n2467), .B(n2463), .Z(n2490) );
  XNOR U2749 ( .A(n2462), .B(n2458), .Z(n2491) );
  XNOR U2750 ( .A(n2457), .B(n2453), .Z(n2492) );
  XNOR U2751 ( .A(n2452), .B(n2448), .Z(n2493) );
  XNOR U2752 ( .A(n2447), .B(n2443), .Z(n2494) );
  XNOR U2753 ( .A(n2442), .B(n2438), .Z(n2495) );
  XNOR U2754 ( .A(n2437), .B(n2433), .Z(n2496) );
  XNOR U2755 ( .A(n2432), .B(n2428), .Z(n2497) );
  XOR U2756 ( .A(n2427), .B(n2424), .Z(n2498) );
  XOR U2757 ( .A(n2499), .B(n2500), .Z(n2424) );
  XOR U2758 ( .A(n2422), .B(n2501), .Z(n2500) );
  XOR U2759 ( .A(n2502), .B(n2503), .Z(n2501) );
  XOR U2760 ( .A(n2504), .B(n2505), .Z(n2503) );
  NAND U2761 ( .A(b[14]), .B(a[19]), .Z(n2505) );
  AND U2762 ( .A(b[15]), .B(a[18]), .Z(n2504) );
  XOR U2763 ( .A(n2506), .B(n2502), .Z(n2499) );
  XOR U2764 ( .A(n2507), .B(n2508), .Z(n2502) );
  NOR U2765 ( .A(n2509), .B(n2510), .Z(n2507) );
  AND U2766 ( .A(b[13]), .B(a[20]), .Z(n2506) );
  XNOR U2767 ( .A(n2511), .B(n2422), .Z(n2423) );
  XOR U2768 ( .A(n2512), .B(n2513), .Z(n2422) );
  ANDN U2769 ( .B(n2514), .A(n2515), .Z(n2512) );
  AND U2770 ( .A(b[12]), .B(a[21]), .Z(n2511) );
  XNOR U2771 ( .A(n2516), .B(n2427), .Z(n2429) );
  XOR U2772 ( .A(n2517), .B(n2518), .Z(n2427) );
  ANDN U2773 ( .B(n2519), .A(n2520), .Z(n2517) );
  AND U2774 ( .A(b[11]), .B(a[22]), .Z(n2516) );
  XNOR U2775 ( .A(n2521), .B(n2432), .Z(n2434) );
  XOR U2776 ( .A(n2522), .B(n2523), .Z(n2432) );
  ANDN U2777 ( .B(n2524), .A(n2525), .Z(n2522) );
  AND U2778 ( .A(b[10]), .B(a[23]), .Z(n2521) );
  XNOR U2779 ( .A(n2526), .B(n2437), .Z(n2439) );
  XOR U2780 ( .A(n2527), .B(n2528), .Z(n2437) );
  ANDN U2781 ( .B(n2529), .A(n2530), .Z(n2527) );
  AND U2782 ( .A(b[9]), .B(a[24]), .Z(n2526) );
  XNOR U2783 ( .A(n2531), .B(n2442), .Z(n2444) );
  XOR U2784 ( .A(n2532), .B(n2533), .Z(n2442) );
  ANDN U2785 ( .B(n2534), .A(n2535), .Z(n2532) );
  AND U2786 ( .A(b[8]), .B(a[25]), .Z(n2531) );
  XNOR U2787 ( .A(n2536), .B(n2447), .Z(n2449) );
  XOR U2788 ( .A(n2537), .B(n2538), .Z(n2447) );
  ANDN U2789 ( .B(n2539), .A(n2540), .Z(n2537) );
  AND U2790 ( .A(b[7]), .B(a[26]), .Z(n2536) );
  XNOR U2791 ( .A(n2541), .B(n2452), .Z(n2454) );
  XOR U2792 ( .A(n2542), .B(n2543), .Z(n2452) );
  ANDN U2793 ( .B(n2544), .A(n2545), .Z(n2542) );
  AND U2794 ( .A(b[6]), .B(a[27]), .Z(n2541) );
  XNOR U2795 ( .A(n2546), .B(n2457), .Z(n2459) );
  XOR U2796 ( .A(n2547), .B(n2548), .Z(n2457) );
  ANDN U2797 ( .B(n2549), .A(n2550), .Z(n2547) );
  AND U2798 ( .A(b[5]), .B(a[28]), .Z(n2546) );
  XNOR U2799 ( .A(n2551), .B(n2462), .Z(n2464) );
  XOR U2800 ( .A(n2552), .B(n2553), .Z(n2462) );
  ANDN U2801 ( .B(n2554), .A(n2555), .Z(n2552) );
  AND U2802 ( .A(b[4]), .B(a[29]), .Z(n2551) );
  XNOR U2803 ( .A(n2556), .B(n2557), .Z(n2476) );
  NANDN U2804 ( .A(n2558), .B(n2559), .Z(n2557) );
  XNOR U2805 ( .A(n2560), .B(n2467), .Z(n2469) );
  XNOR U2806 ( .A(n2561), .B(n2562), .Z(n2467) );
  AND U2807 ( .A(n2563), .B(n2564), .Z(n2561) );
  AND U2808 ( .A(b[3]), .B(a[30]), .Z(n2560) );
  XOR U2809 ( .A(n2483), .B(n2482), .Z(swire[32]) );
  XOR U2810 ( .A(sreg[96]), .B(n2481), .Z(n2482) );
  XOR U2811 ( .A(n2488), .B(n2565), .Z(n2483) );
  XNOR U2812 ( .A(n2487), .B(n2481), .Z(n2565) );
  XOR U2813 ( .A(n2566), .B(n2567), .Z(n2481) );
  NOR U2814 ( .A(n2568), .B(n2569), .Z(n2566) );
  NAND U2815 ( .A(a[32]), .B(b[0]), .Z(n2487) );
  XNOR U2816 ( .A(n2558), .B(n2559), .Z(n2488) );
  XOR U2817 ( .A(n2556), .B(n2570), .Z(n2559) );
  NAND U2818 ( .A(b[1]), .B(a[31]), .Z(n2570) );
  XOR U2819 ( .A(n2564), .B(n2571), .Z(n2558) );
  XOR U2820 ( .A(n2556), .B(n2563), .Z(n2571) );
  XNOR U2821 ( .A(n2572), .B(n2562), .Z(n2563) );
  AND U2822 ( .A(b[2]), .B(a[30]), .Z(n2572) );
  NANDN U2823 ( .A(n2573), .B(n2574), .Z(n2556) );
  XOR U2824 ( .A(n2562), .B(n2554), .Z(n2575) );
  XNOR U2825 ( .A(n2553), .B(n2549), .Z(n2576) );
  XNOR U2826 ( .A(n2548), .B(n2544), .Z(n2577) );
  XNOR U2827 ( .A(n2543), .B(n2539), .Z(n2578) );
  XNOR U2828 ( .A(n2538), .B(n2534), .Z(n2579) );
  XNOR U2829 ( .A(n2533), .B(n2529), .Z(n2580) );
  XNOR U2830 ( .A(n2528), .B(n2524), .Z(n2581) );
  XNOR U2831 ( .A(n2523), .B(n2519), .Z(n2582) );
  XNOR U2832 ( .A(n2518), .B(n2514), .Z(n2583) );
  XOR U2833 ( .A(n2513), .B(n2510), .Z(n2584) );
  XOR U2834 ( .A(n2585), .B(n2586), .Z(n2510) );
  XOR U2835 ( .A(n2508), .B(n2587), .Z(n2586) );
  XOR U2836 ( .A(n2588), .B(n2589), .Z(n2587) );
  XOR U2837 ( .A(n2590), .B(n2591), .Z(n2589) );
  NAND U2838 ( .A(b[14]), .B(a[18]), .Z(n2591) );
  AND U2839 ( .A(b[15]), .B(a[17]), .Z(n2590) );
  XOR U2840 ( .A(n2592), .B(n2588), .Z(n2585) );
  XOR U2841 ( .A(n2593), .B(n2594), .Z(n2588) );
  NOR U2842 ( .A(n2595), .B(n2596), .Z(n2593) );
  AND U2843 ( .A(b[13]), .B(a[19]), .Z(n2592) );
  XNOR U2844 ( .A(n2597), .B(n2508), .Z(n2509) );
  XOR U2845 ( .A(n2598), .B(n2599), .Z(n2508) );
  ANDN U2846 ( .B(n2600), .A(n2601), .Z(n2598) );
  AND U2847 ( .A(b[12]), .B(a[20]), .Z(n2597) );
  XNOR U2848 ( .A(n2602), .B(n2513), .Z(n2515) );
  XOR U2849 ( .A(n2603), .B(n2604), .Z(n2513) );
  ANDN U2850 ( .B(n2605), .A(n2606), .Z(n2603) );
  AND U2851 ( .A(b[11]), .B(a[21]), .Z(n2602) );
  XNOR U2852 ( .A(n2607), .B(n2518), .Z(n2520) );
  XOR U2853 ( .A(n2608), .B(n2609), .Z(n2518) );
  ANDN U2854 ( .B(n2610), .A(n2611), .Z(n2608) );
  AND U2855 ( .A(b[10]), .B(a[22]), .Z(n2607) );
  XNOR U2856 ( .A(n2612), .B(n2523), .Z(n2525) );
  XOR U2857 ( .A(n2613), .B(n2614), .Z(n2523) );
  ANDN U2858 ( .B(n2615), .A(n2616), .Z(n2613) );
  AND U2859 ( .A(b[9]), .B(a[23]), .Z(n2612) );
  XNOR U2860 ( .A(n2617), .B(n2528), .Z(n2530) );
  XOR U2861 ( .A(n2618), .B(n2619), .Z(n2528) );
  ANDN U2862 ( .B(n2620), .A(n2621), .Z(n2618) );
  AND U2863 ( .A(b[8]), .B(a[24]), .Z(n2617) );
  XNOR U2864 ( .A(n2622), .B(n2533), .Z(n2535) );
  XOR U2865 ( .A(n2623), .B(n2624), .Z(n2533) );
  ANDN U2866 ( .B(n2625), .A(n2626), .Z(n2623) );
  AND U2867 ( .A(b[7]), .B(a[25]), .Z(n2622) );
  XNOR U2868 ( .A(n2627), .B(n2538), .Z(n2540) );
  XOR U2869 ( .A(n2628), .B(n2629), .Z(n2538) );
  ANDN U2870 ( .B(n2630), .A(n2631), .Z(n2628) );
  AND U2871 ( .A(b[6]), .B(a[26]), .Z(n2627) );
  XNOR U2872 ( .A(n2632), .B(n2543), .Z(n2545) );
  XOR U2873 ( .A(n2633), .B(n2634), .Z(n2543) );
  ANDN U2874 ( .B(n2635), .A(n2636), .Z(n2633) );
  AND U2875 ( .A(b[5]), .B(a[27]), .Z(n2632) );
  XNOR U2876 ( .A(n2637), .B(n2548), .Z(n2550) );
  XOR U2877 ( .A(n2638), .B(n2639), .Z(n2548) );
  ANDN U2878 ( .B(n2640), .A(n2641), .Z(n2638) );
  AND U2879 ( .A(b[4]), .B(a[28]), .Z(n2637) );
  XNOR U2880 ( .A(n2642), .B(n2643), .Z(n2562) );
  NANDN U2881 ( .A(n2644), .B(n2645), .Z(n2643) );
  XNOR U2882 ( .A(n2646), .B(n2553), .Z(n2555) );
  XNOR U2883 ( .A(n2647), .B(n2648), .Z(n2553) );
  AND U2884 ( .A(n2649), .B(n2650), .Z(n2647) );
  AND U2885 ( .A(b[3]), .B(a[29]), .Z(n2646) );
  XOR U2886 ( .A(n2569), .B(n2568), .Z(swire[31]) );
  XOR U2887 ( .A(sreg[95]), .B(n2567), .Z(n2568) );
  XOR U2888 ( .A(n2574), .B(n2651), .Z(n2569) );
  XNOR U2889 ( .A(n2573), .B(n2567), .Z(n2651) );
  XOR U2890 ( .A(n2652), .B(n2653), .Z(n2567) );
  NOR U2891 ( .A(n2654), .B(n2655), .Z(n2652) );
  NAND U2892 ( .A(a[31]), .B(b[0]), .Z(n2573) );
  XNOR U2893 ( .A(n2644), .B(n2645), .Z(n2574) );
  XOR U2894 ( .A(n2642), .B(n2656), .Z(n2645) );
  NAND U2895 ( .A(b[1]), .B(a[30]), .Z(n2656) );
  XOR U2896 ( .A(n2650), .B(n2657), .Z(n2644) );
  XOR U2897 ( .A(n2642), .B(n2649), .Z(n2657) );
  XNOR U2898 ( .A(n2658), .B(n2648), .Z(n2649) );
  AND U2899 ( .A(b[2]), .B(a[29]), .Z(n2658) );
  NANDN U2900 ( .A(n2659), .B(n2660), .Z(n2642) );
  XOR U2901 ( .A(n2648), .B(n2640), .Z(n2661) );
  XNOR U2902 ( .A(n2639), .B(n2635), .Z(n2662) );
  XNOR U2903 ( .A(n2634), .B(n2630), .Z(n2663) );
  XNOR U2904 ( .A(n2629), .B(n2625), .Z(n2664) );
  XNOR U2905 ( .A(n2624), .B(n2620), .Z(n2665) );
  XNOR U2906 ( .A(n2619), .B(n2615), .Z(n2666) );
  XNOR U2907 ( .A(n2614), .B(n2610), .Z(n2667) );
  XNOR U2908 ( .A(n2609), .B(n2605), .Z(n2668) );
  XNOR U2909 ( .A(n2604), .B(n2600), .Z(n2669) );
  XOR U2910 ( .A(n2599), .B(n2596), .Z(n2670) );
  XOR U2911 ( .A(n2671), .B(n2672), .Z(n2596) );
  XOR U2912 ( .A(n2594), .B(n2673), .Z(n2672) );
  XOR U2913 ( .A(n2674), .B(n2675), .Z(n2673) );
  XOR U2914 ( .A(n2676), .B(n2677), .Z(n2675) );
  NAND U2915 ( .A(b[14]), .B(a[17]), .Z(n2677) );
  AND U2916 ( .A(b[15]), .B(a[16]), .Z(n2676) );
  XOR U2917 ( .A(n2678), .B(n2674), .Z(n2671) );
  XOR U2918 ( .A(n2679), .B(n2680), .Z(n2674) );
  NOR U2919 ( .A(n2681), .B(n2682), .Z(n2679) );
  AND U2920 ( .A(b[13]), .B(a[18]), .Z(n2678) );
  XNOR U2921 ( .A(n2683), .B(n2594), .Z(n2595) );
  XOR U2922 ( .A(n2684), .B(n2685), .Z(n2594) );
  ANDN U2923 ( .B(n2686), .A(n2687), .Z(n2684) );
  AND U2924 ( .A(b[12]), .B(a[19]), .Z(n2683) );
  XNOR U2925 ( .A(n2688), .B(n2599), .Z(n2601) );
  XOR U2926 ( .A(n2689), .B(n2690), .Z(n2599) );
  ANDN U2927 ( .B(n2691), .A(n2692), .Z(n2689) );
  AND U2928 ( .A(b[11]), .B(a[20]), .Z(n2688) );
  XNOR U2929 ( .A(n2693), .B(n2604), .Z(n2606) );
  XOR U2930 ( .A(n2694), .B(n2695), .Z(n2604) );
  ANDN U2931 ( .B(n2696), .A(n2697), .Z(n2694) );
  AND U2932 ( .A(b[10]), .B(a[21]), .Z(n2693) );
  XNOR U2933 ( .A(n2698), .B(n2609), .Z(n2611) );
  XOR U2934 ( .A(n2699), .B(n2700), .Z(n2609) );
  ANDN U2935 ( .B(n2701), .A(n2702), .Z(n2699) );
  AND U2936 ( .A(b[9]), .B(a[22]), .Z(n2698) );
  XNOR U2937 ( .A(n2703), .B(n2614), .Z(n2616) );
  XOR U2938 ( .A(n2704), .B(n2705), .Z(n2614) );
  ANDN U2939 ( .B(n2706), .A(n2707), .Z(n2704) );
  AND U2940 ( .A(b[8]), .B(a[23]), .Z(n2703) );
  XNOR U2941 ( .A(n2708), .B(n2619), .Z(n2621) );
  XOR U2942 ( .A(n2709), .B(n2710), .Z(n2619) );
  ANDN U2943 ( .B(n2711), .A(n2712), .Z(n2709) );
  AND U2944 ( .A(b[7]), .B(a[24]), .Z(n2708) );
  XNOR U2945 ( .A(n2713), .B(n2624), .Z(n2626) );
  XOR U2946 ( .A(n2714), .B(n2715), .Z(n2624) );
  ANDN U2947 ( .B(n2716), .A(n2717), .Z(n2714) );
  AND U2948 ( .A(b[6]), .B(a[25]), .Z(n2713) );
  XNOR U2949 ( .A(n2718), .B(n2629), .Z(n2631) );
  XOR U2950 ( .A(n2719), .B(n2720), .Z(n2629) );
  ANDN U2951 ( .B(n2721), .A(n2722), .Z(n2719) );
  AND U2952 ( .A(b[5]), .B(a[26]), .Z(n2718) );
  XNOR U2953 ( .A(n2723), .B(n2634), .Z(n2636) );
  XOR U2954 ( .A(n2724), .B(n2725), .Z(n2634) );
  ANDN U2955 ( .B(n2726), .A(n2727), .Z(n2724) );
  AND U2956 ( .A(b[4]), .B(a[27]), .Z(n2723) );
  XNOR U2957 ( .A(n2728), .B(n2729), .Z(n2648) );
  NANDN U2958 ( .A(n2730), .B(n2731), .Z(n2729) );
  XNOR U2959 ( .A(n2732), .B(n2639), .Z(n2641) );
  XNOR U2960 ( .A(n2733), .B(n2734), .Z(n2639) );
  AND U2961 ( .A(n2735), .B(n2736), .Z(n2733) );
  AND U2962 ( .A(b[3]), .B(a[28]), .Z(n2732) );
  XOR U2963 ( .A(n2655), .B(n2654), .Z(swire[30]) );
  XOR U2964 ( .A(sreg[94]), .B(n2653), .Z(n2654) );
  XOR U2965 ( .A(n2660), .B(n2737), .Z(n2655) );
  XNOR U2966 ( .A(n2659), .B(n2653), .Z(n2737) );
  XOR U2967 ( .A(n2738), .B(n2739), .Z(n2653) );
  NOR U2968 ( .A(n2740), .B(n2741), .Z(n2738) );
  NAND U2969 ( .A(a[30]), .B(b[0]), .Z(n2659) );
  XNOR U2970 ( .A(n2730), .B(n2731), .Z(n2660) );
  XOR U2971 ( .A(n2728), .B(n2742), .Z(n2731) );
  NAND U2972 ( .A(b[1]), .B(a[29]), .Z(n2742) );
  XOR U2973 ( .A(n2736), .B(n2743), .Z(n2730) );
  XOR U2974 ( .A(n2728), .B(n2735), .Z(n2743) );
  XNOR U2975 ( .A(n2744), .B(n2734), .Z(n2735) );
  AND U2976 ( .A(b[2]), .B(a[28]), .Z(n2744) );
  NANDN U2977 ( .A(n2745), .B(n2746), .Z(n2728) );
  XOR U2978 ( .A(n2734), .B(n2726), .Z(n2747) );
  XNOR U2979 ( .A(n2725), .B(n2721), .Z(n2748) );
  XNOR U2980 ( .A(n2720), .B(n2716), .Z(n2749) );
  XNOR U2981 ( .A(n2715), .B(n2711), .Z(n2750) );
  XNOR U2982 ( .A(n2710), .B(n2706), .Z(n2751) );
  XNOR U2983 ( .A(n2705), .B(n2701), .Z(n2752) );
  XNOR U2984 ( .A(n2700), .B(n2696), .Z(n2753) );
  XNOR U2985 ( .A(n2695), .B(n2691), .Z(n2754) );
  XNOR U2986 ( .A(n2690), .B(n2686), .Z(n2755) );
  XOR U2987 ( .A(n2685), .B(n2682), .Z(n2756) );
  XOR U2988 ( .A(n2757), .B(n2758), .Z(n2682) );
  XOR U2989 ( .A(n2680), .B(n2759), .Z(n2758) );
  XOR U2990 ( .A(n2760), .B(n2761), .Z(n2759) );
  XOR U2991 ( .A(n2762), .B(n2763), .Z(n2761) );
  NAND U2992 ( .A(b[14]), .B(a[16]), .Z(n2763) );
  AND U2993 ( .A(b[15]), .B(a[15]), .Z(n2762) );
  XOR U2994 ( .A(n2764), .B(n2760), .Z(n2757) );
  XOR U2995 ( .A(n2765), .B(n2766), .Z(n2760) );
  NOR U2996 ( .A(n2767), .B(n2768), .Z(n2765) );
  AND U2997 ( .A(b[13]), .B(a[17]), .Z(n2764) );
  XNOR U2998 ( .A(n2769), .B(n2680), .Z(n2681) );
  XOR U2999 ( .A(n2770), .B(n2771), .Z(n2680) );
  ANDN U3000 ( .B(n2772), .A(n2773), .Z(n2770) );
  AND U3001 ( .A(b[12]), .B(a[18]), .Z(n2769) );
  XNOR U3002 ( .A(n2774), .B(n2685), .Z(n2687) );
  XOR U3003 ( .A(n2775), .B(n2776), .Z(n2685) );
  ANDN U3004 ( .B(n2777), .A(n2778), .Z(n2775) );
  AND U3005 ( .A(b[11]), .B(a[19]), .Z(n2774) );
  XNOR U3006 ( .A(n2779), .B(n2690), .Z(n2692) );
  XOR U3007 ( .A(n2780), .B(n2781), .Z(n2690) );
  ANDN U3008 ( .B(n2782), .A(n2783), .Z(n2780) );
  AND U3009 ( .A(b[10]), .B(a[20]), .Z(n2779) );
  XNOR U3010 ( .A(n2784), .B(n2695), .Z(n2697) );
  XOR U3011 ( .A(n2785), .B(n2786), .Z(n2695) );
  ANDN U3012 ( .B(n2787), .A(n2788), .Z(n2785) );
  AND U3013 ( .A(b[9]), .B(a[21]), .Z(n2784) );
  XNOR U3014 ( .A(n2789), .B(n2700), .Z(n2702) );
  XOR U3015 ( .A(n2790), .B(n2791), .Z(n2700) );
  ANDN U3016 ( .B(n2792), .A(n2793), .Z(n2790) );
  AND U3017 ( .A(b[8]), .B(a[22]), .Z(n2789) );
  XNOR U3018 ( .A(n2794), .B(n2705), .Z(n2707) );
  XOR U3019 ( .A(n2795), .B(n2796), .Z(n2705) );
  ANDN U3020 ( .B(n2797), .A(n2798), .Z(n2795) );
  AND U3021 ( .A(b[7]), .B(a[23]), .Z(n2794) );
  XNOR U3022 ( .A(n2799), .B(n2710), .Z(n2712) );
  XOR U3023 ( .A(n2800), .B(n2801), .Z(n2710) );
  ANDN U3024 ( .B(n2802), .A(n2803), .Z(n2800) );
  AND U3025 ( .A(b[6]), .B(a[24]), .Z(n2799) );
  XNOR U3026 ( .A(n2804), .B(n2715), .Z(n2717) );
  XOR U3027 ( .A(n2805), .B(n2806), .Z(n2715) );
  ANDN U3028 ( .B(n2807), .A(n2808), .Z(n2805) );
  AND U3029 ( .A(b[5]), .B(a[25]), .Z(n2804) );
  XNOR U3030 ( .A(n2809), .B(n2720), .Z(n2722) );
  XOR U3031 ( .A(n2810), .B(n2811), .Z(n2720) );
  ANDN U3032 ( .B(n2812), .A(n2813), .Z(n2810) );
  AND U3033 ( .A(b[4]), .B(a[26]), .Z(n2809) );
  XNOR U3034 ( .A(n2814), .B(n2815), .Z(n2734) );
  NANDN U3035 ( .A(n2816), .B(n2817), .Z(n2815) );
  XNOR U3036 ( .A(n2818), .B(n2725), .Z(n2727) );
  XNOR U3037 ( .A(n2819), .B(n2820), .Z(n2725) );
  AND U3038 ( .A(n2821), .B(n2822), .Z(n2819) );
  AND U3039 ( .A(b[3]), .B(a[27]), .Z(n2818) );
  XOR U3040 ( .A(n2741), .B(n2740), .Z(swire[29]) );
  XOR U3041 ( .A(sreg[93]), .B(n2739), .Z(n2740) );
  XOR U3042 ( .A(n2746), .B(n2823), .Z(n2741) );
  XNOR U3043 ( .A(n2745), .B(n2739), .Z(n2823) );
  XOR U3044 ( .A(n2824), .B(n2825), .Z(n2739) );
  NOR U3045 ( .A(n2826), .B(n2827), .Z(n2824) );
  NAND U3046 ( .A(a[29]), .B(b[0]), .Z(n2745) );
  XNOR U3047 ( .A(n2816), .B(n2817), .Z(n2746) );
  XOR U3048 ( .A(n2814), .B(n2828), .Z(n2817) );
  NAND U3049 ( .A(b[1]), .B(a[28]), .Z(n2828) );
  XOR U3050 ( .A(n2822), .B(n2829), .Z(n2816) );
  XOR U3051 ( .A(n2814), .B(n2821), .Z(n2829) );
  XNOR U3052 ( .A(n2830), .B(n2820), .Z(n2821) );
  AND U3053 ( .A(b[2]), .B(a[27]), .Z(n2830) );
  NANDN U3054 ( .A(n2831), .B(n2832), .Z(n2814) );
  XOR U3055 ( .A(n2820), .B(n2812), .Z(n2833) );
  XNOR U3056 ( .A(n2811), .B(n2807), .Z(n2834) );
  XNOR U3057 ( .A(n2806), .B(n2802), .Z(n2835) );
  XNOR U3058 ( .A(n2801), .B(n2797), .Z(n2836) );
  XNOR U3059 ( .A(n2796), .B(n2792), .Z(n2837) );
  XNOR U3060 ( .A(n2791), .B(n2787), .Z(n2838) );
  XNOR U3061 ( .A(n2786), .B(n2782), .Z(n2839) );
  XNOR U3062 ( .A(n2781), .B(n2777), .Z(n2840) );
  XNOR U3063 ( .A(n2776), .B(n2772), .Z(n2841) );
  XOR U3064 ( .A(n2771), .B(n2768), .Z(n2842) );
  XOR U3065 ( .A(n2843), .B(n2844), .Z(n2768) );
  XOR U3066 ( .A(n2766), .B(n2845), .Z(n2844) );
  XOR U3067 ( .A(n2846), .B(n2847), .Z(n2845) );
  XOR U3068 ( .A(n2848), .B(n2849), .Z(n2847) );
  NAND U3069 ( .A(b[14]), .B(a[15]), .Z(n2849) );
  AND U3070 ( .A(b[15]), .B(a[14]), .Z(n2848) );
  XOR U3071 ( .A(n2850), .B(n2846), .Z(n2843) );
  XOR U3072 ( .A(n2851), .B(n2852), .Z(n2846) );
  NOR U3073 ( .A(n2853), .B(n2854), .Z(n2851) );
  AND U3074 ( .A(b[13]), .B(a[16]), .Z(n2850) );
  XNOR U3075 ( .A(n2855), .B(n2766), .Z(n2767) );
  XOR U3076 ( .A(n2856), .B(n2857), .Z(n2766) );
  ANDN U3077 ( .B(n2858), .A(n2859), .Z(n2856) );
  AND U3078 ( .A(b[12]), .B(a[17]), .Z(n2855) );
  XNOR U3079 ( .A(n2860), .B(n2771), .Z(n2773) );
  XOR U3080 ( .A(n2861), .B(n2862), .Z(n2771) );
  ANDN U3081 ( .B(n2863), .A(n2864), .Z(n2861) );
  AND U3082 ( .A(b[11]), .B(a[18]), .Z(n2860) );
  XNOR U3083 ( .A(n2865), .B(n2776), .Z(n2778) );
  XOR U3084 ( .A(n2866), .B(n2867), .Z(n2776) );
  ANDN U3085 ( .B(n2868), .A(n2869), .Z(n2866) );
  AND U3086 ( .A(b[10]), .B(a[19]), .Z(n2865) );
  XNOR U3087 ( .A(n2870), .B(n2781), .Z(n2783) );
  XOR U3088 ( .A(n2871), .B(n2872), .Z(n2781) );
  ANDN U3089 ( .B(n2873), .A(n2874), .Z(n2871) );
  AND U3090 ( .A(b[9]), .B(a[20]), .Z(n2870) );
  XNOR U3091 ( .A(n2875), .B(n2786), .Z(n2788) );
  XOR U3092 ( .A(n2876), .B(n2877), .Z(n2786) );
  ANDN U3093 ( .B(n2878), .A(n2879), .Z(n2876) );
  AND U3094 ( .A(b[8]), .B(a[21]), .Z(n2875) );
  XNOR U3095 ( .A(n2880), .B(n2791), .Z(n2793) );
  XOR U3096 ( .A(n2881), .B(n2882), .Z(n2791) );
  ANDN U3097 ( .B(n2883), .A(n2884), .Z(n2881) );
  AND U3098 ( .A(b[7]), .B(a[22]), .Z(n2880) );
  XNOR U3099 ( .A(n2885), .B(n2796), .Z(n2798) );
  XOR U3100 ( .A(n2886), .B(n2887), .Z(n2796) );
  ANDN U3101 ( .B(n2888), .A(n2889), .Z(n2886) );
  AND U3102 ( .A(b[6]), .B(a[23]), .Z(n2885) );
  XNOR U3103 ( .A(n2890), .B(n2801), .Z(n2803) );
  XOR U3104 ( .A(n2891), .B(n2892), .Z(n2801) );
  ANDN U3105 ( .B(n2893), .A(n2894), .Z(n2891) );
  AND U3106 ( .A(b[5]), .B(a[24]), .Z(n2890) );
  XNOR U3107 ( .A(n2895), .B(n2806), .Z(n2808) );
  XOR U3108 ( .A(n2896), .B(n2897), .Z(n2806) );
  ANDN U3109 ( .B(n2898), .A(n2899), .Z(n2896) );
  AND U3110 ( .A(b[4]), .B(a[25]), .Z(n2895) );
  XNOR U3111 ( .A(n2900), .B(n2901), .Z(n2820) );
  NANDN U3112 ( .A(n2902), .B(n2903), .Z(n2901) );
  XNOR U3113 ( .A(n2904), .B(n2811), .Z(n2813) );
  XNOR U3114 ( .A(n2905), .B(n2906), .Z(n2811) );
  AND U3115 ( .A(n2907), .B(n2908), .Z(n2905) );
  AND U3116 ( .A(b[3]), .B(a[26]), .Z(n2904) );
  XOR U3117 ( .A(n2827), .B(n2826), .Z(swire[28]) );
  XOR U3118 ( .A(sreg[92]), .B(n2825), .Z(n2826) );
  XOR U3119 ( .A(n2832), .B(n2909), .Z(n2827) );
  XNOR U3120 ( .A(n2831), .B(n2825), .Z(n2909) );
  XOR U3121 ( .A(n2910), .B(n2911), .Z(n2825) );
  NOR U3122 ( .A(n2912), .B(n2913), .Z(n2910) );
  NAND U3123 ( .A(a[28]), .B(b[0]), .Z(n2831) );
  XNOR U3124 ( .A(n2902), .B(n2903), .Z(n2832) );
  XOR U3125 ( .A(n2900), .B(n2914), .Z(n2903) );
  NAND U3126 ( .A(b[1]), .B(a[27]), .Z(n2914) );
  XOR U3127 ( .A(n2908), .B(n2915), .Z(n2902) );
  XOR U3128 ( .A(n2900), .B(n2907), .Z(n2915) );
  XNOR U3129 ( .A(n2916), .B(n2906), .Z(n2907) );
  AND U3130 ( .A(b[2]), .B(a[26]), .Z(n2916) );
  NANDN U3131 ( .A(n2917), .B(n2918), .Z(n2900) );
  XOR U3132 ( .A(n2906), .B(n2898), .Z(n2919) );
  XNOR U3133 ( .A(n2897), .B(n2893), .Z(n2920) );
  XNOR U3134 ( .A(n2892), .B(n2888), .Z(n2921) );
  XNOR U3135 ( .A(n2887), .B(n2883), .Z(n2922) );
  XNOR U3136 ( .A(n2882), .B(n2878), .Z(n2923) );
  XNOR U3137 ( .A(n2877), .B(n2873), .Z(n2924) );
  XNOR U3138 ( .A(n2872), .B(n2868), .Z(n2925) );
  XNOR U3139 ( .A(n2867), .B(n2863), .Z(n2926) );
  XNOR U3140 ( .A(n2862), .B(n2858), .Z(n2927) );
  XOR U3141 ( .A(n2857), .B(n2854), .Z(n2928) );
  XOR U3142 ( .A(n2929), .B(n2930), .Z(n2854) );
  XOR U3143 ( .A(n2852), .B(n2931), .Z(n2930) );
  XOR U3144 ( .A(n2932), .B(n2933), .Z(n2931) );
  XOR U3145 ( .A(n2934), .B(n2935), .Z(n2933) );
  NAND U3146 ( .A(b[14]), .B(a[14]), .Z(n2935) );
  AND U3147 ( .A(b[15]), .B(a[13]), .Z(n2934) );
  XOR U3148 ( .A(n2936), .B(n2932), .Z(n2929) );
  XOR U3149 ( .A(n2937), .B(n2938), .Z(n2932) );
  NOR U3150 ( .A(n2939), .B(n2940), .Z(n2937) );
  AND U3151 ( .A(b[13]), .B(a[15]), .Z(n2936) );
  XNOR U3152 ( .A(n2941), .B(n2852), .Z(n2853) );
  XOR U3153 ( .A(n2942), .B(n2943), .Z(n2852) );
  ANDN U3154 ( .B(n2944), .A(n2945), .Z(n2942) );
  AND U3155 ( .A(b[12]), .B(a[16]), .Z(n2941) );
  XNOR U3156 ( .A(n2946), .B(n2857), .Z(n2859) );
  XOR U3157 ( .A(n2947), .B(n2948), .Z(n2857) );
  ANDN U3158 ( .B(n2949), .A(n2950), .Z(n2947) );
  AND U3159 ( .A(b[11]), .B(a[17]), .Z(n2946) );
  XNOR U3160 ( .A(n2951), .B(n2862), .Z(n2864) );
  XOR U3161 ( .A(n2952), .B(n2953), .Z(n2862) );
  ANDN U3162 ( .B(n2954), .A(n2955), .Z(n2952) );
  AND U3163 ( .A(b[10]), .B(a[18]), .Z(n2951) );
  XNOR U3164 ( .A(n2956), .B(n2867), .Z(n2869) );
  XOR U3165 ( .A(n2957), .B(n2958), .Z(n2867) );
  ANDN U3166 ( .B(n2959), .A(n2960), .Z(n2957) );
  AND U3167 ( .A(b[9]), .B(a[19]), .Z(n2956) );
  XNOR U3168 ( .A(n2961), .B(n2872), .Z(n2874) );
  XOR U3169 ( .A(n2962), .B(n2963), .Z(n2872) );
  ANDN U3170 ( .B(n2964), .A(n2965), .Z(n2962) );
  AND U3171 ( .A(b[8]), .B(a[20]), .Z(n2961) );
  XNOR U3172 ( .A(n2966), .B(n2877), .Z(n2879) );
  XOR U3173 ( .A(n2967), .B(n2968), .Z(n2877) );
  ANDN U3174 ( .B(n2969), .A(n2970), .Z(n2967) );
  AND U3175 ( .A(b[7]), .B(a[21]), .Z(n2966) );
  XNOR U3176 ( .A(n2971), .B(n2882), .Z(n2884) );
  XOR U3177 ( .A(n2972), .B(n2973), .Z(n2882) );
  ANDN U3178 ( .B(n2974), .A(n2975), .Z(n2972) );
  AND U3179 ( .A(b[6]), .B(a[22]), .Z(n2971) );
  XNOR U3180 ( .A(n2976), .B(n2887), .Z(n2889) );
  XOR U3181 ( .A(n2977), .B(n2978), .Z(n2887) );
  ANDN U3182 ( .B(n2979), .A(n2980), .Z(n2977) );
  AND U3183 ( .A(b[5]), .B(a[23]), .Z(n2976) );
  XNOR U3184 ( .A(n2981), .B(n2892), .Z(n2894) );
  XOR U3185 ( .A(n2982), .B(n2983), .Z(n2892) );
  ANDN U3186 ( .B(n2984), .A(n2985), .Z(n2982) );
  AND U3187 ( .A(b[4]), .B(a[24]), .Z(n2981) );
  XNOR U3188 ( .A(n2986), .B(n2987), .Z(n2906) );
  NANDN U3189 ( .A(n2988), .B(n2989), .Z(n2987) );
  XNOR U3190 ( .A(n2990), .B(n2897), .Z(n2899) );
  XNOR U3191 ( .A(n2991), .B(n2992), .Z(n2897) );
  AND U3192 ( .A(n2993), .B(n2994), .Z(n2991) );
  AND U3193 ( .A(b[3]), .B(a[25]), .Z(n2990) );
  XOR U3194 ( .A(n2913), .B(n2912), .Z(swire[27]) );
  XOR U3195 ( .A(sreg[91]), .B(n2911), .Z(n2912) );
  XOR U3196 ( .A(n2918), .B(n2995), .Z(n2913) );
  XNOR U3197 ( .A(n2917), .B(n2911), .Z(n2995) );
  XOR U3198 ( .A(n2996), .B(n2997), .Z(n2911) );
  NOR U3199 ( .A(n2998), .B(n2999), .Z(n2996) );
  NAND U3200 ( .A(a[27]), .B(b[0]), .Z(n2917) );
  XNOR U3201 ( .A(n2988), .B(n2989), .Z(n2918) );
  XOR U3202 ( .A(n2986), .B(n3000), .Z(n2989) );
  NAND U3203 ( .A(b[1]), .B(a[26]), .Z(n3000) );
  XOR U3204 ( .A(n2994), .B(n3001), .Z(n2988) );
  XOR U3205 ( .A(n2986), .B(n2993), .Z(n3001) );
  XNOR U3206 ( .A(n3002), .B(n2992), .Z(n2993) );
  AND U3207 ( .A(b[2]), .B(a[25]), .Z(n3002) );
  NANDN U3208 ( .A(n3003), .B(n3004), .Z(n2986) );
  XOR U3209 ( .A(n2992), .B(n2984), .Z(n3005) );
  XNOR U3210 ( .A(n2983), .B(n2979), .Z(n3006) );
  XNOR U3211 ( .A(n2978), .B(n2974), .Z(n3007) );
  XNOR U3212 ( .A(n2973), .B(n2969), .Z(n3008) );
  XNOR U3213 ( .A(n2968), .B(n2964), .Z(n3009) );
  XNOR U3214 ( .A(n2963), .B(n2959), .Z(n3010) );
  XNOR U3215 ( .A(n2958), .B(n2954), .Z(n3011) );
  XNOR U3216 ( .A(n2953), .B(n2949), .Z(n3012) );
  XNOR U3217 ( .A(n2948), .B(n2944), .Z(n3013) );
  XOR U3218 ( .A(n2943), .B(n2940), .Z(n3014) );
  XOR U3219 ( .A(n3015), .B(n3016), .Z(n2940) );
  XOR U3220 ( .A(n2938), .B(n3017), .Z(n3016) );
  XOR U3221 ( .A(n3018), .B(n3019), .Z(n3017) );
  XOR U3222 ( .A(n3020), .B(n3021), .Z(n3019) );
  NAND U3223 ( .A(b[14]), .B(a[13]), .Z(n3021) );
  AND U3224 ( .A(b[15]), .B(a[12]), .Z(n3020) );
  XOR U3225 ( .A(n3022), .B(n3018), .Z(n3015) );
  XOR U3226 ( .A(n3023), .B(n3024), .Z(n3018) );
  NOR U3227 ( .A(n3025), .B(n3026), .Z(n3023) );
  AND U3228 ( .A(b[13]), .B(a[14]), .Z(n3022) );
  XNOR U3229 ( .A(n3027), .B(n2938), .Z(n2939) );
  XOR U3230 ( .A(n3028), .B(n3029), .Z(n2938) );
  ANDN U3231 ( .B(n3030), .A(n3031), .Z(n3028) );
  AND U3232 ( .A(b[12]), .B(a[15]), .Z(n3027) );
  XNOR U3233 ( .A(n3032), .B(n2943), .Z(n2945) );
  XOR U3234 ( .A(n3033), .B(n3034), .Z(n2943) );
  ANDN U3235 ( .B(n3035), .A(n3036), .Z(n3033) );
  AND U3236 ( .A(b[11]), .B(a[16]), .Z(n3032) );
  XNOR U3237 ( .A(n3037), .B(n2948), .Z(n2950) );
  XOR U3238 ( .A(n3038), .B(n3039), .Z(n2948) );
  ANDN U3239 ( .B(n3040), .A(n3041), .Z(n3038) );
  AND U3240 ( .A(b[10]), .B(a[17]), .Z(n3037) );
  XNOR U3241 ( .A(n3042), .B(n2953), .Z(n2955) );
  XOR U3242 ( .A(n3043), .B(n3044), .Z(n2953) );
  ANDN U3243 ( .B(n3045), .A(n3046), .Z(n3043) );
  AND U3244 ( .A(b[9]), .B(a[18]), .Z(n3042) );
  XNOR U3245 ( .A(n3047), .B(n2958), .Z(n2960) );
  XOR U3246 ( .A(n3048), .B(n3049), .Z(n2958) );
  ANDN U3247 ( .B(n3050), .A(n3051), .Z(n3048) );
  AND U3248 ( .A(b[8]), .B(a[19]), .Z(n3047) );
  XNOR U3249 ( .A(n3052), .B(n2963), .Z(n2965) );
  XOR U3250 ( .A(n3053), .B(n3054), .Z(n2963) );
  ANDN U3251 ( .B(n3055), .A(n3056), .Z(n3053) );
  AND U3252 ( .A(b[7]), .B(a[20]), .Z(n3052) );
  XNOR U3253 ( .A(n3057), .B(n2968), .Z(n2970) );
  XOR U3254 ( .A(n3058), .B(n3059), .Z(n2968) );
  ANDN U3255 ( .B(n3060), .A(n3061), .Z(n3058) );
  AND U3256 ( .A(b[6]), .B(a[21]), .Z(n3057) );
  XNOR U3257 ( .A(n3062), .B(n2973), .Z(n2975) );
  XOR U3258 ( .A(n3063), .B(n3064), .Z(n2973) );
  ANDN U3259 ( .B(n3065), .A(n3066), .Z(n3063) );
  AND U3260 ( .A(b[5]), .B(a[22]), .Z(n3062) );
  XNOR U3261 ( .A(n3067), .B(n2978), .Z(n2980) );
  XOR U3262 ( .A(n3068), .B(n3069), .Z(n2978) );
  ANDN U3263 ( .B(n3070), .A(n3071), .Z(n3068) );
  AND U3264 ( .A(b[4]), .B(a[23]), .Z(n3067) );
  XNOR U3265 ( .A(n3072), .B(n3073), .Z(n2992) );
  NANDN U3266 ( .A(n3074), .B(n3075), .Z(n3073) );
  XNOR U3267 ( .A(n3076), .B(n2983), .Z(n2985) );
  XNOR U3268 ( .A(n3077), .B(n3078), .Z(n2983) );
  AND U3269 ( .A(n3079), .B(n3080), .Z(n3077) );
  AND U3270 ( .A(b[3]), .B(a[24]), .Z(n3076) );
  XOR U3271 ( .A(n2999), .B(n2998), .Z(swire[26]) );
  XOR U3272 ( .A(sreg[90]), .B(n2997), .Z(n2998) );
  XOR U3273 ( .A(n3004), .B(n3081), .Z(n2999) );
  XNOR U3274 ( .A(n3003), .B(n2997), .Z(n3081) );
  XOR U3275 ( .A(n3082), .B(n3083), .Z(n2997) );
  NOR U3276 ( .A(n3084), .B(n3085), .Z(n3082) );
  NAND U3277 ( .A(a[26]), .B(b[0]), .Z(n3003) );
  XNOR U3278 ( .A(n3074), .B(n3075), .Z(n3004) );
  XOR U3279 ( .A(n3072), .B(n3086), .Z(n3075) );
  NAND U3280 ( .A(b[1]), .B(a[25]), .Z(n3086) );
  XOR U3281 ( .A(n3080), .B(n3087), .Z(n3074) );
  XOR U3282 ( .A(n3072), .B(n3079), .Z(n3087) );
  XNOR U3283 ( .A(n3088), .B(n3078), .Z(n3079) );
  AND U3284 ( .A(b[2]), .B(a[24]), .Z(n3088) );
  NANDN U3285 ( .A(n3089), .B(n3090), .Z(n3072) );
  XOR U3286 ( .A(n3078), .B(n3070), .Z(n3091) );
  XNOR U3287 ( .A(n3069), .B(n3065), .Z(n3092) );
  XNOR U3288 ( .A(n3064), .B(n3060), .Z(n3093) );
  XNOR U3289 ( .A(n3059), .B(n3055), .Z(n3094) );
  XNOR U3290 ( .A(n3054), .B(n3050), .Z(n3095) );
  XNOR U3291 ( .A(n3049), .B(n3045), .Z(n3096) );
  XNOR U3292 ( .A(n3044), .B(n3040), .Z(n3097) );
  XNOR U3293 ( .A(n3039), .B(n3035), .Z(n3098) );
  XNOR U3294 ( .A(n3034), .B(n3030), .Z(n3099) );
  XOR U3295 ( .A(n3029), .B(n3026), .Z(n3100) );
  XOR U3296 ( .A(n3101), .B(n3102), .Z(n3026) );
  XOR U3297 ( .A(n3024), .B(n3103), .Z(n3102) );
  XOR U3298 ( .A(n3104), .B(n3105), .Z(n3103) );
  XOR U3299 ( .A(n3106), .B(n3107), .Z(n3105) );
  NAND U3300 ( .A(b[14]), .B(a[12]), .Z(n3107) );
  AND U3301 ( .A(b[15]), .B(a[11]), .Z(n3106) );
  XOR U3302 ( .A(n3108), .B(n3104), .Z(n3101) );
  XOR U3303 ( .A(n3109), .B(n3110), .Z(n3104) );
  NOR U3304 ( .A(n3111), .B(n3112), .Z(n3109) );
  AND U3305 ( .A(b[13]), .B(a[13]), .Z(n3108) );
  XNOR U3306 ( .A(n3113), .B(n3024), .Z(n3025) );
  XOR U3307 ( .A(n3114), .B(n3115), .Z(n3024) );
  ANDN U3308 ( .B(n3116), .A(n3117), .Z(n3114) );
  AND U3309 ( .A(b[12]), .B(a[14]), .Z(n3113) );
  XNOR U3310 ( .A(n3118), .B(n3029), .Z(n3031) );
  XOR U3311 ( .A(n3119), .B(n3120), .Z(n3029) );
  ANDN U3312 ( .B(n3121), .A(n3122), .Z(n3119) );
  AND U3313 ( .A(b[11]), .B(a[15]), .Z(n3118) );
  XNOR U3314 ( .A(n3123), .B(n3034), .Z(n3036) );
  XOR U3315 ( .A(n3124), .B(n3125), .Z(n3034) );
  ANDN U3316 ( .B(n3126), .A(n3127), .Z(n3124) );
  AND U3317 ( .A(b[10]), .B(a[16]), .Z(n3123) );
  XNOR U3318 ( .A(n3128), .B(n3039), .Z(n3041) );
  XOR U3319 ( .A(n3129), .B(n3130), .Z(n3039) );
  ANDN U3320 ( .B(n3131), .A(n3132), .Z(n3129) );
  AND U3321 ( .A(b[9]), .B(a[17]), .Z(n3128) );
  XNOR U3322 ( .A(n3133), .B(n3044), .Z(n3046) );
  XOR U3323 ( .A(n3134), .B(n3135), .Z(n3044) );
  ANDN U3324 ( .B(n3136), .A(n3137), .Z(n3134) );
  AND U3325 ( .A(b[8]), .B(a[18]), .Z(n3133) );
  XNOR U3326 ( .A(n3138), .B(n3049), .Z(n3051) );
  XOR U3327 ( .A(n3139), .B(n3140), .Z(n3049) );
  ANDN U3328 ( .B(n3141), .A(n3142), .Z(n3139) );
  AND U3329 ( .A(b[7]), .B(a[19]), .Z(n3138) );
  XNOR U3330 ( .A(n3143), .B(n3054), .Z(n3056) );
  XOR U3331 ( .A(n3144), .B(n3145), .Z(n3054) );
  ANDN U3332 ( .B(n3146), .A(n3147), .Z(n3144) );
  AND U3333 ( .A(b[6]), .B(a[20]), .Z(n3143) );
  XNOR U3334 ( .A(n3148), .B(n3059), .Z(n3061) );
  XOR U3335 ( .A(n3149), .B(n3150), .Z(n3059) );
  ANDN U3336 ( .B(n3151), .A(n3152), .Z(n3149) );
  AND U3337 ( .A(b[5]), .B(a[21]), .Z(n3148) );
  XNOR U3338 ( .A(n3153), .B(n3064), .Z(n3066) );
  XOR U3339 ( .A(n3154), .B(n3155), .Z(n3064) );
  ANDN U3340 ( .B(n3156), .A(n3157), .Z(n3154) );
  AND U3341 ( .A(b[4]), .B(a[22]), .Z(n3153) );
  XNOR U3342 ( .A(n3158), .B(n3159), .Z(n3078) );
  NANDN U3343 ( .A(n3160), .B(n3161), .Z(n3159) );
  XNOR U3344 ( .A(n3162), .B(n3069), .Z(n3071) );
  XNOR U3345 ( .A(n3163), .B(n3164), .Z(n3069) );
  AND U3346 ( .A(n3165), .B(n3166), .Z(n3163) );
  AND U3347 ( .A(b[3]), .B(a[23]), .Z(n3162) );
  XOR U3348 ( .A(n3085), .B(n3084), .Z(swire[25]) );
  XOR U3349 ( .A(sreg[89]), .B(n3083), .Z(n3084) );
  XOR U3350 ( .A(n3090), .B(n3167), .Z(n3085) );
  XNOR U3351 ( .A(n3089), .B(n3083), .Z(n3167) );
  XOR U3352 ( .A(n3168), .B(n3169), .Z(n3083) );
  NOR U3353 ( .A(n3170), .B(n3171), .Z(n3168) );
  NAND U3354 ( .A(a[25]), .B(b[0]), .Z(n3089) );
  XNOR U3355 ( .A(n3160), .B(n3161), .Z(n3090) );
  XOR U3356 ( .A(n3158), .B(n3172), .Z(n3161) );
  NAND U3357 ( .A(b[1]), .B(a[24]), .Z(n3172) );
  XOR U3358 ( .A(n3166), .B(n3173), .Z(n3160) );
  XOR U3359 ( .A(n3158), .B(n3165), .Z(n3173) );
  XNOR U3360 ( .A(n3174), .B(n3164), .Z(n3165) );
  AND U3361 ( .A(b[2]), .B(a[23]), .Z(n3174) );
  NANDN U3362 ( .A(n3175), .B(n3176), .Z(n3158) );
  XOR U3363 ( .A(n3164), .B(n3156), .Z(n3177) );
  XNOR U3364 ( .A(n3155), .B(n3151), .Z(n3178) );
  XNOR U3365 ( .A(n3150), .B(n3146), .Z(n3179) );
  XNOR U3366 ( .A(n3145), .B(n3141), .Z(n3180) );
  XNOR U3367 ( .A(n3140), .B(n3136), .Z(n3181) );
  XNOR U3368 ( .A(n3135), .B(n3131), .Z(n3182) );
  XNOR U3369 ( .A(n3130), .B(n3126), .Z(n3183) );
  XNOR U3370 ( .A(n3125), .B(n3121), .Z(n3184) );
  XNOR U3371 ( .A(n3120), .B(n3116), .Z(n3185) );
  XOR U3372 ( .A(n3115), .B(n3112), .Z(n3186) );
  XOR U3373 ( .A(n3187), .B(n3188), .Z(n3112) );
  XOR U3374 ( .A(n3110), .B(n3189), .Z(n3188) );
  XOR U3375 ( .A(n3190), .B(n3191), .Z(n3189) );
  XOR U3376 ( .A(n3192), .B(n3193), .Z(n3191) );
  NAND U3377 ( .A(b[14]), .B(a[11]), .Z(n3193) );
  AND U3378 ( .A(b[15]), .B(a[10]), .Z(n3192) );
  XOR U3379 ( .A(n3194), .B(n3190), .Z(n3187) );
  XOR U3380 ( .A(n3195), .B(n3196), .Z(n3190) );
  NOR U3381 ( .A(n3197), .B(n3198), .Z(n3195) );
  AND U3382 ( .A(b[13]), .B(a[12]), .Z(n3194) );
  XNOR U3383 ( .A(n3199), .B(n3110), .Z(n3111) );
  XOR U3384 ( .A(n3200), .B(n3201), .Z(n3110) );
  ANDN U3385 ( .B(n3202), .A(n3203), .Z(n3200) );
  AND U3386 ( .A(b[12]), .B(a[13]), .Z(n3199) );
  XNOR U3387 ( .A(n3204), .B(n3115), .Z(n3117) );
  XOR U3388 ( .A(n3205), .B(n3206), .Z(n3115) );
  ANDN U3389 ( .B(n3207), .A(n3208), .Z(n3205) );
  AND U3390 ( .A(b[11]), .B(a[14]), .Z(n3204) );
  XNOR U3391 ( .A(n3209), .B(n3120), .Z(n3122) );
  XOR U3392 ( .A(n3210), .B(n3211), .Z(n3120) );
  ANDN U3393 ( .B(n3212), .A(n3213), .Z(n3210) );
  AND U3394 ( .A(b[10]), .B(a[15]), .Z(n3209) );
  XNOR U3395 ( .A(n3214), .B(n3125), .Z(n3127) );
  XOR U3396 ( .A(n3215), .B(n3216), .Z(n3125) );
  ANDN U3397 ( .B(n3217), .A(n3218), .Z(n3215) );
  AND U3398 ( .A(b[9]), .B(a[16]), .Z(n3214) );
  XNOR U3399 ( .A(n3219), .B(n3130), .Z(n3132) );
  XOR U3400 ( .A(n3220), .B(n3221), .Z(n3130) );
  ANDN U3401 ( .B(n3222), .A(n3223), .Z(n3220) );
  AND U3402 ( .A(b[8]), .B(a[17]), .Z(n3219) );
  XNOR U3403 ( .A(n3224), .B(n3135), .Z(n3137) );
  XOR U3404 ( .A(n3225), .B(n3226), .Z(n3135) );
  ANDN U3405 ( .B(n3227), .A(n3228), .Z(n3225) );
  AND U3406 ( .A(b[7]), .B(a[18]), .Z(n3224) );
  XNOR U3407 ( .A(n3229), .B(n3140), .Z(n3142) );
  XOR U3408 ( .A(n3230), .B(n3231), .Z(n3140) );
  ANDN U3409 ( .B(n3232), .A(n3233), .Z(n3230) );
  AND U3410 ( .A(b[6]), .B(a[19]), .Z(n3229) );
  XNOR U3411 ( .A(n3234), .B(n3145), .Z(n3147) );
  XOR U3412 ( .A(n3235), .B(n3236), .Z(n3145) );
  ANDN U3413 ( .B(n3237), .A(n3238), .Z(n3235) );
  AND U3414 ( .A(b[5]), .B(a[20]), .Z(n3234) );
  XNOR U3415 ( .A(n3239), .B(n3150), .Z(n3152) );
  XOR U3416 ( .A(n3240), .B(n3241), .Z(n3150) );
  ANDN U3417 ( .B(n3242), .A(n3243), .Z(n3240) );
  AND U3418 ( .A(b[4]), .B(a[21]), .Z(n3239) );
  XNOR U3419 ( .A(n3244), .B(n3245), .Z(n3164) );
  NANDN U3420 ( .A(n3246), .B(n3247), .Z(n3245) );
  XNOR U3421 ( .A(n3248), .B(n3155), .Z(n3157) );
  XNOR U3422 ( .A(n3249), .B(n3250), .Z(n3155) );
  AND U3423 ( .A(n3251), .B(n3252), .Z(n3249) );
  AND U3424 ( .A(b[3]), .B(a[22]), .Z(n3248) );
  XOR U3425 ( .A(n3171), .B(n3170), .Z(swire[24]) );
  XOR U3426 ( .A(sreg[88]), .B(n3169), .Z(n3170) );
  XOR U3427 ( .A(n3176), .B(n3253), .Z(n3171) );
  XNOR U3428 ( .A(n3175), .B(n3169), .Z(n3253) );
  XOR U3429 ( .A(n3254), .B(n3255), .Z(n3169) );
  NOR U3430 ( .A(n3256), .B(n3257), .Z(n3254) );
  NAND U3431 ( .A(a[24]), .B(b[0]), .Z(n3175) );
  XNOR U3432 ( .A(n3246), .B(n3247), .Z(n3176) );
  XOR U3433 ( .A(n3244), .B(n3258), .Z(n3247) );
  NAND U3434 ( .A(b[1]), .B(a[23]), .Z(n3258) );
  XOR U3435 ( .A(n3252), .B(n3259), .Z(n3246) );
  XOR U3436 ( .A(n3244), .B(n3251), .Z(n3259) );
  XNOR U3437 ( .A(n3260), .B(n3250), .Z(n3251) );
  AND U3438 ( .A(b[2]), .B(a[22]), .Z(n3260) );
  NANDN U3439 ( .A(n3261), .B(n3262), .Z(n3244) );
  XOR U3440 ( .A(n3250), .B(n3242), .Z(n3263) );
  XNOR U3441 ( .A(n3241), .B(n3237), .Z(n3264) );
  XNOR U3442 ( .A(n3236), .B(n3232), .Z(n3265) );
  XNOR U3443 ( .A(n3231), .B(n3227), .Z(n3266) );
  XNOR U3444 ( .A(n3226), .B(n3222), .Z(n3267) );
  XNOR U3445 ( .A(n3221), .B(n3217), .Z(n3268) );
  XNOR U3446 ( .A(n3216), .B(n3212), .Z(n3269) );
  XNOR U3447 ( .A(n3211), .B(n3207), .Z(n3270) );
  XNOR U3448 ( .A(n3206), .B(n3202), .Z(n3271) );
  XOR U3449 ( .A(n3201), .B(n3198), .Z(n3272) );
  XOR U3450 ( .A(n3273), .B(n3274), .Z(n3198) );
  XOR U3451 ( .A(n3196), .B(n3275), .Z(n3274) );
  XOR U3452 ( .A(n3276), .B(n3277), .Z(n3275) );
  XOR U3453 ( .A(n3278), .B(n3279), .Z(n3277) );
  NAND U3454 ( .A(b[14]), .B(a[10]), .Z(n3279) );
  AND U3455 ( .A(b[15]), .B(a[9]), .Z(n3278) );
  XOR U3456 ( .A(n3280), .B(n3276), .Z(n3273) );
  XOR U3457 ( .A(n3281), .B(n3282), .Z(n3276) );
  NOR U3458 ( .A(n3283), .B(n3284), .Z(n3281) );
  AND U3459 ( .A(b[13]), .B(a[11]), .Z(n3280) );
  XNOR U3460 ( .A(n3285), .B(n3196), .Z(n3197) );
  XOR U3461 ( .A(n3286), .B(n3287), .Z(n3196) );
  ANDN U3462 ( .B(n3288), .A(n3289), .Z(n3286) );
  AND U3463 ( .A(b[12]), .B(a[12]), .Z(n3285) );
  XNOR U3464 ( .A(n3290), .B(n3201), .Z(n3203) );
  XOR U3465 ( .A(n3291), .B(n3292), .Z(n3201) );
  ANDN U3466 ( .B(n3293), .A(n3294), .Z(n3291) );
  AND U3467 ( .A(b[11]), .B(a[13]), .Z(n3290) );
  XNOR U3468 ( .A(n3295), .B(n3206), .Z(n3208) );
  XOR U3469 ( .A(n3296), .B(n3297), .Z(n3206) );
  ANDN U3470 ( .B(n3298), .A(n3299), .Z(n3296) );
  AND U3471 ( .A(b[10]), .B(a[14]), .Z(n3295) );
  XNOR U3472 ( .A(n3300), .B(n3211), .Z(n3213) );
  XOR U3473 ( .A(n3301), .B(n3302), .Z(n3211) );
  ANDN U3474 ( .B(n3303), .A(n3304), .Z(n3301) );
  AND U3475 ( .A(b[9]), .B(a[15]), .Z(n3300) );
  XNOR U3476 ( .A(n3305), .B(n3216), .Z(n3218) );
  XOR U3477 ( .A(n3306), .B(n3307), .Z(n3216) );
  ANDN U3478 ( .B(n3308), .A(n3309), .Z(n3306) );
  AND U3479 ( .A(b[8]), .B(a[16]), .Z(n3305) );
  XNOR U3480 ( .A(n3310), .B(n3221), .Z(n3223) );
  XOR U3481 ( .A(n3311), .B(n3312), .Z(n3221) );
  ANDN U3482 ( .B(n3313), .A(n3314), .Z(n3311) );
  AND U3483 ( .A(b[7]), .B(a[17]), .Z(n3310) );
  XNOR U3484 ( .A(n3315), .B(n3226), .Z(n3228) );
  XOR U3485 ( .A(n3316), .B(n3317), .Z(n3226) );
  ANDN U3486 ( .B(n3318), .A(n3319), .Z(n3316) );
  AND U3487 ( .A(b[6]), .B(a[18]), .Z(n3315) );
  XNOR U3488 ( .A(n3320), .B(n3231), .Z(n3233) );
  XOR U3489 ( .A(n3321), .B(n3322), .Z(n3231) );
  ANDN U3490 ( .B(n3323), .A(n3324), .Z(n3321) );
  AND U3491 ( .A(b[5]), .B(a[19]), .Z(n3320) );
  XNOR U3492 ( .A(n3325), .B(n3236), .Z(n3238) );
  XOR U3493 ( .A(n3326), .B(n3327), .Z(n3236) );
  ANDN U3494 ( .B(n3328), .A(n3329), .Z(n3326) );
  AND U3495 ( .A(b[4]), .B(a[20]), .Z(n3325) );
  XNOR U3496 ( .A(n3330), .B(n3331), .Z(n3250) );
  NANDN U3497 ( .A(n3332), .B(n3333), .Z(n3331) );
  XNOR U3498 ( .A(n3334), .B(n3241), .Z(n3243) );
  XNOR U3499 ( .A(n3335), .B(n3336), .Z(n3241) );
  AND U3500 ( .A(n3337), .B(n3338), .Z(n3335) );
  AND U3501 ( .A(b[3]), .B(a[21]), .Z(n3334) );
  XOR U3502 ( .A(n3257), .B(n3256), .Z(swire[23]) );
  XOR U3503 ( .A(sreg[87]), .B(n3255), .Z(n3256) );
  XOR U3504 ( .A(n3262), .B(n3339), .Z(n3257) );
  XNOR U3505 ( .A(n3261), .B(n3255), .Z(n3339) );
  XOR U3506 ( .A(n3340), .B(n3341), .Z(n3255) );
  NOR U3507 ( .A(n3342), .B(n3343), .Z(n3340) );
  NAND U3508 ( .A(a[23]), .B(b[0]), .Z(n3261) );
  XNOR U3509 ( .A(n3332), .B(n3333), .Z(n3262) );
  XOR U3510 ( .A(n3330), .B(n3344), .Z(n3333) );
  NAND U3511 ( .A(b[1]), .B(a[22]), .Z(n3344) );
  XOR U3512 ( .A(n3338), .B(n3345), .Z(n3332) );
  XOR U3513 ( .A(n3330), .B(n3337), .Z(n3345) );
  XNOR U3514 ( .A(n3346), .B(n3336), .Z(n3337) );
  AND U3515 ( .A(b[2]), .B(a[21]), .Z(n3346) );
  NANDN U3516 ( .A(n3347), .B(n3348), .Z(n3330) );
  XOR U3517 ( .A(n3336), .B(n3328), .Z(n3349) );
  XNOR U3518 ( .A(n3327), .B(n3323), .Z(n3350) );
  XNOR U3519 ( .A(n3322), .B(n3318), .Z(n3351) );
  XNOR U3520 ( .A(n3317), .B(n3313), .Z(n3352) );
  XNOR U3521 ( .A(n3312), .B(n3308), .Z(n3353) );
  XNOR U3522 ( .A(n3307), .B(n3303), .Z(n3354) );
  XNOR U3523 ( .A(n3302), .B(n3298), .Z(n3355) );
  XNOR U3524 ( .A(n3297), .B(n3293), .Z(n3356) );
  XNOR U3525 ( .A(n3292), .B(n3288), .Z(n3357) );
  XOR U3526 ( .A(n3287), .B(n3284), .Z(n3358) );
  XOR U3527 ( .A(n3359), .B(n3360), .Z(n3284) );
  XOR U3528 ( .A(n3282), .B(n3361), .Z(n3360) );
  XOR U3529 ( .A(n3362), .B(n3363), .Z(n3361) );
  XOR U3530 ( .A(n3364), .B(n3365), .Z(n3363) );
  NAND U3531 ( .A(b[14]), .B(a[9]), .Z(n3365) );
  AND U3532 ( .A(b[15]), .B(a[8]), .Z(n3364) );
  XOR U3533 ( .A(n3366), .B(n3362), .Z(n3359) );
  XOR U3534 ( .A(n3367), .B(n3368), .Z(n3362) );
  NOR U3535 ( .A(n3369), .B(n3370), .Z(n3367) );
  AND U3536 ( .A(b[13]), .B(a[10]), .Z(n3366) );
  XNOR U3537 ( .A(n3371), .B(n3282), .Z(n3283) );
  XOR U3538 ( .A(n3372), .B(n3373), .Z(n3282) );
  ANDN U3539 ( .B(n3374), .A(n3375), .Z(n3372) );
  AND U3540 ( .A(b[12]), .B(a[11]), .Z(n3371) );
  XNOR U3541 ( .A(n3376), .B(n3287), .Z(n3289) );
  XOR U3542 ( .A(n3377), .B(n3378), .Z(n3287) );
  ANDN U3543 ( .B(n3379), .A(n3380), .Z(n3377) );
  AND U3544 ( .A(b[11]), .B(a[12]), .Z(n3376) );
  XNOR U3545 ( .A(n3381), .B(n3292), .Z(n3294) );
  XOR U3546 ( .A(n3382), .B(n3383), .Z(n3292) );
  ANDN U3547 ( .B(n3384), .A(n3385), .Z(n3382) );
  AND U3548 ( .A(b[10]), .B(a[13]), .Z(n3381) );
  XNOR U3549 ( .A(n3386), .B(n3297), .Z(n3299) );
  XOR U3550 ( .A(n3387), .B(n3388), .Z(n3297) );
  ANDN U3551 ( .B(n3389), .A(n3390), .Z(n3387) );
  AND U3552 ( .A(b[9]), .B(a[14]), .Z(n3386) );
  XNOR U3553 ( .A(n3391), .B(n3302), .Z(n3304) );
  XOR U3554 ( .A(n3392), .B(n3393), .Z(n3302) );
  ANDN U3555 ( .B(n3394), .A(n3395), .Z(n3392) );
  AND U3556 ( .A(b[8]), .B(a[15]), .Z(n3391) );
  XNOR U3557 ( .A(n3396), .B(n3307), .Z(n3309) );
  XOR U3558 ( .A(n3397), .B(n3398), .Z(n3307) );
  ANDN U3559 ( .B(n3399), .A(n3400), .Z(n3397) );
  AND U3560 ( .A(b[7]), .B(a[16]), .Z(n3396) );
  XNOR U3561 ( .A(n3401), .B(n3312), .Z(n3314) );
  XOR U3562 ( .A(n3402), .B(n3403), .Z(n3312) );
  ANDN U3563 ( .B(n3404), .A(n3405), .Z(n3402) );
  AND U3564 ( .A(b[6]), .B(a[17]), .Z(n3401) );
  XNOR U3565 ( .A(n3406), .B(n3317), .Z(n3319) );
  XOR U3566 ( .A(n3407), .B(n3408), .Z(n3317) );
  ANDN U3567 ( .B(n3409), .A(n3410), .Z(n3407) );
  AND U3568 ( .A(b[5]), .B(a[18]), .Z(n3406) );
  XNOR U3569 ( .A(n3411), .B(n3322), .Z(n3324) );
  XOR U3570 ( .A(n3412), .B(n3413), .Z(n3322) );
  ANDN U3571 ( .B(n3414), .A(n3415), .Z(n3412) );
  AND U3572 ( .A(b[4]), .B(a[19]), .Z(n3411) );
  XNOR U3573 ( .A(n3416), .B(n3417), .Z(n3336) );
  NANDN U3574 ( .A(n3418), .B(n3419), .Z(n3417) );
  XNOR U3575 ( .A(n3420), .B(n3327), .Z(n3329) );
  XNOR U3576 ( .A(n3421), .B(n3422), .Z(n3327) );
  AND U3577 ( .A(n3423), .B(n3424), .Z(n3421) );
  AND U3578 ( .A(b[3]), .B(a[20]), .Z(n3420) );
  XOR U3579 ( .A(n3343), .B(n3342), .Z(swire[22]) );
  XOR U3580 ( .A(sreg[86]), .B(n3341), .Z(n3342) );
  XOR U3581 ( .A(n3348), .B(n3425), .Z(n3343) );
  XNOR U3582 ( .A(n3347), .B(n3341), .Z(n3425) );
  XOR U3583 ( .A(n3426), .B(n3427), .Z(n3341) );
  NOR U3584 ( .A(n3428), .B(n3429), .Z(n3426) );
  NAND U3585 ( .A(a[22]), .B(b[0]), .Z(n3347) );
  XNOR U3586 ( .A(n3418), .B(n3419), .Z(n3348) );
  XOR U3587 ( .A(n3416), .B(n3430), .Z(n3419) );
  NAND U3588 ( .A(b[1]), .B(a[21]), .Z(n3430) );
  XOR U3589 ( .A(n3424), .B(n3431), .Z(n3418) );
  XOR U3590 ( .A(n3416), .B(n3423), .Z(n3431) );
  XNOR U3591 ( .A(n3432), .B(n3422), .Z(n3423) );
  AND U3592 ( .A(b[2]), .B(a[20]), .Z(n3432) );
  NANDN U3593 ( .A(n3433), .B(n3434), .Z(n3416) );
  XOR U3594 ( .A(n3422), .B(n3414), .Z(n3435) );
  XNOR U3595 ( .A(n3413), .B(n3409), .Z(n3436) );
  XNOR U3596 ( .A(n3408), .B(n3404), .Z(n3437) );
  XNOR U3597 ( .A(n3403), .B(n3399), .Z(n3438) );
  XNOR U3598 ( .A(n3398), .B(n3394), .Z(n3439) );
  XNOR U3599 ( .A(n3393), .B(n3389), .Z(n3440) );
  XNOR U3600 ( .A(n3388), .B(n3384), .Z(n3441) );
  XNOR U3601 ( .A(n3383), .B(n3379), .Z(n3442) );
  XNOR U3602 ( .A(n3378), .B(n3374), .Z(n3443) );
  XOR U3603 ( .A(n3373), .B(n3370), .Z(n3444) );
  XOR U3604 ( .A(n3445), .B(n3446), .Z(n3370) );
  XOR U3605 ( .A(n3368), .B(n3447), .Z(n3446) );
  XOR U3606 ( .A(n3448), .B(n3449), .Z(n3447) );
  XOR U3607 ( .A(n3450), .B(n3451), .Z(n3449) );
  NAND U3608 ( .A(b[14]), .B(a[8]), .Z(n3451) );
  AND U3609 ( .A(b[15]), .B(a[7]), .Z(n3450) );
  XOR U3610 ( .A(n3452), .B(n3448), .Z(n3445) );
  XOR U3611 ( .A(n3453), .B(n3454), .Z(n3448) );
  NOR U3612 ( .A(n3455), .B(n3456), .Z(n3453) );
  AND U3613 ( .A(b[13]), .B(a[9]), .Z(n3452) );
  XNOR U3614 ( .A(n3457), .B(n3368), .Z(n3369) );
  XOR U3615 ( .A(n3458), .B(n3459), .Z(n3368) );
  ANDN U3616 ( .B(n3460), .A(n3461), .Z(n3458) );
  AND U3617 ( .A(b[12]), .B(a[10]), .Z(n3457) );
  XNOR U3618 ( .A(n3462), .B(n3373), .Z(n3375) );
  XOR U3619 ( .A(n3463), .B(n3464), .Z(n3373) );
  ANDN U3620 ( .B(n3465), .A(n3466), .Z(n3463) );
  AND U3621 ( .A(b[11]), .B(a[11]), .Z(n3462) );
  XNOR U3622 ( .A(n3467), .B(n3378), .Z(n3380) );
  XOR U3623 ( .A(n3468), .B(n3469), .Z(n3378) );
  ANDN U3624 ( .B(n3470), .A(n3471), .Z(n3468) );
  AND U3625 ( .A(b[10]), .B(a[12]), .Z(n3467) );
  XNOR U3626 ( .A(n3472), .B(n3383), .Z(n3385) );
  XOR U3627 ( .A(n3473), .B(n3474), .Z(n3383) );
  ANDN U3628 ( .B(n3475), .A(n3476), .Z(n3473) );
  AND U3629 ( .A(b[9]), .B(a[13]), .Z(n3472) );
  XNOR U3630 ( .A(n3477), .B(n3388), .Z(n3390) );
  XOR U3631 ( .A(n3478), .B(n3479), .Z(n3388) );
  ANDN U3632 ( .B(n3480), .A(n3481), .Z(n3478) );
  AND U3633 ( .A(b[8]), .B(a[14]), .Z(n3477) );
  XNOR U3634 ( .A(n3482), .B(n3393), .Z(n3395) );
  XOR U3635 ( .A(n3483), .B(n3484), .Z(n3393) );
  ANDN U3636 ( .B(n3485), .A(n3486), .Z(n3483) );
  AND U3637 ( .A(b[7]), .B(a[15]), .Z(n3482) );
  XNOR U3638 ( .A(n3487), .B(n3398), .Z(n3400) );
  XOR U3639 ( .A(n3488), .B(n3489), .Z(n3398) );
  ANDN U3640 ( .B(n3490), .A(n3491), .Z(n3488) );
  AND U3641 ( .A(b[6]), .B(a[16]), .Z(n3487) );
  XNOR U3642 ( .A(n3492), .B(n3403), .Z(n3405) );
  XOR U3643 ( .A(n3493), .B(n3494), .Z(n3403) );
  ANDN U3644 ( .B(n3495), .A(n3496), .Z(n3493) );
  AND U3645 ( .A(b[5]), .B(a[17]), .Z(n3492) );
  XNOR U3646 ( .A(n3497), .B(n3408), .Z(n3410) );
  XOR U3647 ( .A(n3498), .B(n3499), .Z(n3408) );
  ANDN U3648 ( .B(n3500), .A(n3501), .Z(n3498) );
  AND U3649 ( .A(b[4]), .B(a[18]), .Z(n3497) );
  XNOR U3650 ( .A(n3502), .B(n3503), .Z(n3422) );
  NANDN U3651 ( .A(n3504), .B(n3505), .Z(n3503) );
  XNOR U3652 ( .A(n3506), .B(n3413), .Z(n3415) );
  XNOR U3653 ( .A(n3507), .B(n3508), .Z(n3413) );
  AND U3654 ( .A(n3509), .B(n3510), .Z(n3507) );
  AND U3655 ( .A(b[3]), .B(a[19]), .Z(n3506) );
  XOR U3656 ( .A(n3429), .B(n3428), .Z(swire[21]) );
  XOR U3657 ( .A(sreg[85]), .B(n3427), .Z(n3428) );
  XOR U3658 ( .A(n3434), .B(n3511), .Z(n3429) );
  XNOR U3659 ( .A(n3433), .B(n3427), .Z(n3511) );
  XOR U3660 ( .A(n3512), .B(n3513), .Z(n3427) );
  NOR U3661 ( .A(n3514), .B(n3515), .Z(n3512) );
  NAND U3662 ( .A(a[21]), .B(b[0]), .Z(n3433) );
  XNOR U3663 ( .A(n3504), .B(n3505), .Z(n3434) );
  XOR U3664 ( .A(n3502), .B(n3516), .Z(n3505) );
  NAND U3665 ( .A(b[1]), .B(a[20]), .Z(n3516) );
  XOR U3666 ( .A(n3510), .B(n3517), .Z(n3504) );
  XOR U3667 ( .A(n3502), .B(n3509), .Z(n3517) );
  XNOR U3668 ( .A(n3518), .B(n3508), .Z(n3509) );
  AND U3669 ( .A(b[2]), .B(a[19]), .Z(n3518) );
  NANDN U3670 ( .A(n3519), .B(n3520), .Z(n3502) );
  XOR U3671 ( .A(n3508), .B(n3500), .Z(n3521) );
  XNOR U3672 ( .A(n3499), .B(n3495), .Z(n3522) );
  XNOR U3673 ( .A(n3494), .B(n3490), .Z(n3523) );
  XNOR U3674 ( .A(n3489), .B(n3485), .Z(n3524) );
  XNOR U3675 ( .A(n3484), .B(n3480), .Z(n3525) );
  XNOR U3676 ( .A(n3479), .B(n3475), .Z(n3526) );
  XNOR U3677 ( .A(n3474), .B(n3470), .Z(n3527) );
  XNOR U3678 ( .A(n3469), .B(n3465), .Z(n3528) );
  XNOR U3679 ( .A(n3464), .B(n3460), .Z(n3529) );
  XOR U3680 ( .A(n3459), .B(n3456), .Z(n3530) );
  XOR U3681 ( .A(n3531), .B(n3532), .Z(n3456) );
  XOR U3682 ( .A(n3454), .B(n3533), .Z(n3532) );
  XOR U3683 ( .A(n3534), .B(n3535), .Z(n3533) );
  XOR U3684 ( .A(n3536), .B(n3537), .Z(n3535) );
  NAND U3685 ( .A(b[14]), .B(a[7]), .Z(n3537) );
  AND U3686 ( .A(b[15]), .B(a[6]), .Z(n3536) );
  XOR U3687 ( .A(n3538), .B(n3534), .Z(n3531) );
  XOR U3688 ( .A(n3539), .B(n3540), .Z(n3534) );
  NOR U3689 ( .A(n3541), .B(n3542), .Z(n3539) );
  AND U3690 ( .A(b[13]), .B(a[8]), .Z(n3538) );
  XNOR U3691 ( .A(n3543), .B(n3454), .Z(n3455) );
  XOR U3692 ( .A(n3544), .B(n3545), .Z(n3454) );
  ANDN U3693 ( .B(n3546), .A(n3547), .Z(n3544) );
  AND U3694 ( .A(b[12]), .B(a[9]), .Z(n3543) );
  XNOR U3695 ( .A(n3548), .B(n3459), .Z(n3461) );
  XOR U3696 ( .A(n3549), .B(n3550), .Z(n3459) );
  ANDN U3697 ( .B(n3551), .A(n3552), .Z(n3549) );
  AND U3698 ( .A(b[11]), .B(a[10]), .Z(n3548) );
  XNOR U3699 ( .A(n3553), .B(n3464), .Z(n3466) );
  XOR U3700 ( .A(n3554), .B(n3555), .Z(n3464) );
  ANDN U3701 ( .B(n3556), .A(n3557), .Z(n3554) );
  AND U3702 ( .A(b[10]), .B(a[11]), .Z(n3553) );
  XNOR U3703 ( .A(n3558), .B(n3469), .Z(n3471) );
  XOR U3704 ( .A(n3559), .B(n3560), .Z(n3469) );
  ANDN U3705 ( .B(n3561), .A(n3562), .Z(n3559) );
  AND U3706 ( .A(b[9]), .B(a[12]), .Z(n3558) );
  XNOR U3707 ( .A(n3563), .B(n3474), .Z(n3476) );
  XOR U3708 ( .A(n3564), .B(n3565), .Z(n3474) );
  ANDN U3709 ( .B(n3566), .A(n3567), .Z(n3564) );
  AND U3710 ( .A(b[8]), .B(a[13]), .Z(n3563) );
  XNOR U3711 ( .A(n3568), .B(n3479), .Z(n3481) );
  XOR U3712 ( .A(n3569), .B(n3570), .Z(n3479) );
  ANDN U3713 ( .B(n3571), .A(n3572), .Z(n3569) );
  AND U3714 ( .A(b[7]), .B(a[14]), .Z(n3568) );
  XNOR U3715 ( .A(n3573), .B(n3484), .Z(n3486) );
  XOR U3716 ( .A(n3574), .B(n3575), .Z(n3484) );
  ANDN U3717 ( .B(n3576), .A(n3577), .Z(n3574) );
  AND U3718 ( .A(b[6]), .B(a[15]), .Z(n3573) );
  XNOR U3719 ( .A(n3578), .B(n3489), .Z(n3491) );
  XOR U3720 ( .A(n3579), .B(n3580), .Z(n3489) );
  ANDN U3721 ( .B(n3581), .A(n3582), .Z(n3579) );
  AND U3722 ( .A(b[5]), .B(a[16]), .Z(n3578) );
  XNOR U3723 ( .A(n3583), .B(n3494), .Z(n3496) );
  XOR U3724 ( .A(n3584), .B(n3585), .Z(n3494) );
  ANDN U3725 ( .B(n3586), .A(n3587), .Z(n3584) );
  AND U3726 ( .A(b[4]), .B(a[17]), .Z(n3583) );
  XNOR U3727 ( .A(n3588), .B(n3589), .Z(n3508) );
  NANDN U3728 ( .A(n3590), .B(n3591), .Z(n3589) );
  XNOR U3729 ( .A(n3592), .B(n3499), .Z(n3501) );
  XNOR U3730 ( .A(n3593), .B(n3594), .Z(n3499) );
  AND U3731 ( .A(n3595), .B(n3596), .Z(n3593) );
  AND U3732 ( .A(b[3]), .B(a[18]), .Z(n3592) );
  XOR U3733 ( .A(n3515), .B(n3514), .Z(swire[20]) );
  XOR U3734 ( .A(sreg[84]), .B(n3513), .Z(n3514) );
  XOR U3735 ( .A(n3520), .B(n3597), .Z(n3515) );
  XNOR U3736 ( .A(n3519), .B(n3513), .Z(n3597) );
  XOR U3737 ( .A(n3598), .B(n3599), .Z(n3513) );
  NOR U3738 ( .A(n3600), .B(n3601), .Z(n3598) );
  NAND U3739 ( .A(a[20]), .B(b[0]), .Z(n3519) );
  XNOR U3740 ( .A(n3590), .B(n3591), .Z(n3520) );
  XOR U3741 ( .A(n3588), .B(n3602), .Z(n3591) );
  NAND U3742 ( .A(b[1]), .B(a[19]), .Z(n3602) );
  XOR U3743 ( .A(n3596), .B(n3603), .Z(n3590) );
  XOR U3744 ( .A(n3588), .B(n3595), .Z(n3603) );
  XNOR U3745 ( .A(n3604), .B(n3594), .Z(n3595) );
  AND U3746 ( .A(b[2]), .B(a[18]), .Z(n3604) );
  NANDN U3747 ( .A(n3605), .B(n3606), .Z(n3588) );
  XOR U3748 ( .A(n3594), .B(n3586), .Z(n3607) );
  XNOR U3749 ( .A(n3585), .B(n3581), .Z(n3608) );
  XNOR U3750 ( .A(n3580), .B(n3576), .Z(n3609) );
  XNOR U3751 ( .A(n3575), .B(n3571), .Z(n3610) );
  XNOR U3752 ( .A(n3570), .B(n3566), .Z(n3611) );
  XNOR U3753 ( .A(n3565), .B(n3561), .Z(n3612) );
  XNOR U3754 ( .A(n3560), .B(n3556), .Z(n3613) );
  XNOR U3755 ( .A(n3555), .B(n3551), .Z(n3614) );
  XNOR U3756 ( .A(n3550), .B(n3546), .Z(n3615) );
  XOR U3757 ( .A(n3545), .B(n3542), .Z(n3616) );
  XOR U3758 ( .A(n3617), .B(n3618), .Z(n3542) );
  XOR U3759 ( .A(n3540), .B(n3619), .Z(n3618) );
  XOR U3760 ( .A(n3620), .B(n3621), .Z(n3619) );
  XOR U3761 ( .A(n3622), .B(n3623), .Z(n3621) );
  NAND U3762 ( .A(b[14]), .B(a[6]), .Z(n3623) );
  AND U3763 ( .A(b[15]), .B(a[5]), .Z(n3622) );
  XOR U3764 ( .A(n3624), .B(n3620), .Z(n3617) );
  XOR U3765 ( .A(n3625), .B(n3626), .Z(n3620) );
  NOR U3766 ( .A(n3627), .B(n3628), .Z(n3625) );
  AND U3767 ( .A(b[13]), .B(a[7]), .Z(n3624) );
  XNOR U3768 ( .A(n3629), .B(n3540), .Z(n3541) );
  XOR U3769 ( .A(n3630), .B(n3631), .Z(n3540) );
  ANDN U3770 ( .B(n3632), .A(n3633), .Z(n3630) );
  AND U3771 ( .A(b[12]), .B(a[8]), .Z(n3629) );
  XNOR U3772 ( .A(n3634), .B(n3545), .Z(n3547) );
  XOR U3773 ( .A(n3635), .B(n3636), .Z(n3545) );
  ANDN U3774 ( .B(n3637), .A(n3638), .Z(n3635) );
  AND U3775 ( .A(b[11]), .B(a[9]), .Z(n3634) );
  XNOR U3776 ( .A(n3639), .B(n3550), .Z(n3552) );
  XOR U3777 ( .A(n3640), .B(n3641), .Z(n3550) );
  ANDN U3778 ( .B(n3642), .A(n3643), .Z(n3640) );
  AND U3779 ( .A(b[10]), .B(a[10]), .Z(n3639) );
  XNOR U3780 ( .A(n3644), .B(n3555), .Z(n3557) );
  XOR U3781 ( .A(n3645), .B(n3646), .Z(n3555) );
  ANDN U3782 ( .B(n3647), .A(n3648), .Z(n3645) );
  AND U3783 ( .A(b[9]), .B(a[11]), .Z(n3644) );
  XNOR U3784 ( .A(n3649), .B(n3560), .Z(n3562) );
  XOR U3785 ( .A(n3650), .B(n3651), .Z(n3560) );
  ANDN U3786 ( .B(n3652), .A(n3653), .Z(n3650) );
  AND U3787 ( .A(b[8]), .B(a[12]), .Z(n3649) );
  XNOR U3788 ( .A(n3654), .B(n3565), .Z(n3567) );
  XOR U3789 ( .A(n3655), .B(n3656), .Z(n3565) );
  ANDN U3790 ( .B(n3657), .A(n3658), .Z(n3655) );
  AND U3791 ( .A(b[7]), .B(a[13]), .Z(n3654) );
  XNOR U3792 ( .A(n3659), .B(n3570), .Z(n3572) );
  XOR U3793 ( .A(n3660), .B(n3661), .Z(n3570) );
  ANDN U3794 ( .B(n3662), .A(n3663), .Z(n3660) );
  AND U3795 ( .A(b[6]), .B(a[14]), .Z(n3659) );
  XNOR U3796 ( .A(n3664), .B(n3575), .Z(n3577) );
  XOR U3797 ( .A(n3665), .B(n3666), .Z(n3575) );
  ANDN U3798 ( .B(n3667), .A(n3668), .Z(n3665) );
  AND U3799 ( .A(b[5]), .B(a[15]), .Z(n3664) );
  XNOR U3800 ( .A(n3669), .B(n3580), .Z(n3582) );
  XOR U3801 ( .A(n3670), .B(n3671), .Z(n3580) );
  ANDN U3802 ( .B(n3672), .A(n3673), .Z(n3670) );
  AND U3803 ( .A(b[4]), .B(a[16]), .Z(n3669) );
  XNOR U3804 ( .A(n3674), .B(n3675), .Z(n3594) );
  NANDN U3805 ( .A(n3676), .B(n3677), .Z(n3675) );
  XNOR U3806 ( .A(n3678), .B(n3585), .Z(n3587) );
  XNOR U3807 ( .A(n3679), .B(n3680), .Z(n3585) );
  AND U3808 ( .A(n3681), .B(n3682), .Z(n3679) );
  AND U3809 ( .A(b[3]), .B(a[17]), .Z(n3678) );
  XOR U3810 ( .A(n3601), .B(n3600), .Z(swire[19]) );
  XOR U3811 ( .A(sreg[83]), .B(n3599), .Z(n3600) );
  XOR U3812 ( .A(n3606), .B(n3683), .Z(n3601) );
  XNOR U3813 ( .A(n3605), .B(n3599), .Z(n3683) );
  XOR U3814 ( .A(n3684), .B(n3685), .Z(n3599) );
  NOR U3815 ( .A(n3686), .B(n3687), .Z(n3684) );
  NAND U3816 ( .A(a[19]), .B(b[0]), .Z(n3605) );
  XNOR U3817 ( .A(n3676), .B(n3677), .Z(n3606) );
  XOR U3818 ( .A(n3674), .B(n3688), .Z(n3677) );
  NAND U3819 ( .A(b[1]), .B(a[18]), .Z(n3688) );
  XOR U3820 ( .A(n3682), .B(n3689), .Z(n3676) );
  XOR U3821 ( .A(n3674), .B(n3681), .Z(n3689) );
  XNOR U3822 ( .A(n3690), .B(n3680), .Z(n3681) );
  AND U3823 ( .A(b[2]), .B(a[17]), .Z(n3690) );
  NANDN U3824 ( .A(n3691), .B(n3692), .Z(n3674) );
  XOR U3825 ( .A(n3680), .B(n3672), .Z(n3693) );
  XNOR U3826 ( .A(n3671), .B(n3667), .Z(n3694) );
  XNOR U3827 ( .A(n3666), .B(n3662), .Z(n3695) );
  XNOR U3828 ( .A(n3661), .B(n3657), .Z(n3696) );
  XNOR U3829 ( .A(n3656), .B(n3652), .Z(n3697) );
  XNOR U3830 ( .A(n3651), .B(n3647), .Z(n3698) );
  XNOR U3831 ( .A(n3646), .B(n3642), .Z(n3699) );
  XNOR U3832 ( .A(n3641), .B(n3637), .Z(n3700) );
  XNOR U3833 ( .A(n3636), .B(n3632), .Z(n3701) );
  XOR U3834 ( .A(n3631), .B(n3628), .Z(n3702) );
  XOR U3835 ( .A(n3703), .B(n3704), .Z(n3628) );
  XOR U3836 ( .A(n3626), .B(n3705), .Z(n3704) );
  XOR U3837 ( .A(n3706), .B(n3707), .Z(n3705) );
  XOR U3838 ( .A(n3708), .B(n3709), .Z(n3707) );
  NAND U3839 ( .A(b[14]), .B(a[5]), .Z(n3709) );
  AND U3840 ( .A(b[15]), .B(a[4]), .Z(n3708) );
  XOR U3841 ( .A(n3710), .B(n3706), .Z(n3703) );
  XOR U3842 ( .A(n3711), .B(n3712), .Z(n3706) );
  NOR U3843 ( .A(n3713), .B(n3714), .Z(n3711) );
  AND U3844 ( .A(b[13]), .B(a[6]), .Z(n3710) );
  XNOR U3845 ( .A(n3715), .B(n3626), .Z(n3627) );
  XOR U3846 ( .A(n3716), .B(n3717), .Z(n3626) );
  ANDN U3847 ( .B(n3718), .A(n3719), .Z(n3716) );
  AND U3848 ( .A(b[12]), .B(a[7]), .Z(n3715) );
  XNOR U3849 ( .A(n3720), .B(n3631), .Z(n3633) );
  XOR U3850 ( .A(n3721), .B(n3722), .Z(n3631) );
  ANDN U3851 ( .B(n3723), .A(n3724), .Z(n3721) );
  AND U3852 ( .A(b[11]), .B(a[8]), .Z(n3720) );
  XNOR U3853 ( .A(n3725), .B(n3636), .Z(n3638) );
  XOR U3854 ( .A(n3726), .B(n3727), .Z(n3636) );
  ANDN U3855 ( .B(n3728), .A(n3729), .Z(n3726) );
  AND U3856 ( .A(b[10]), .B(a[9]), .Z(n3725) );
  XNOR U3857 ( .A(n3730), .B(n3641), .Z(n3643) );
  XOR U3858 ( .A(n3731), .B(n3732), .Z(n3641) );
  ANDN U3859 ( .B(n3733), .A(n3734), .Z(n3731) );
  AND U3860 ( .A(b[9]), .B(a[10]), .Z(n3730) );
  XNOR U3861 ( .A(n3735), .B(n3646), .Z(n3648) );
  XOR U3862 ( .A(n3736), .B(n3737), .Z(n3646) );
  ANDN U3863 ( .B(n3738), .A(n3739), .Z(n3736) );
  AND U3864 ( .A(b[8]), .B(a[11]), .Z(n3735) );
  XNOR U3865 ( .A(n3740), .B(n3651), .Z(n3653) );
  XOR U3866 ( .A(n3741), .B(n3742), .Z(n3651) );
  ANDN U3867 ( .B(n3743), .A(n3744), .Z(n3741) );
  AND U3868 ( .A(b[7]), .B(a[12]), .Z(n3740) );
  XNOR U3869 ( .A(n3745), .B(n3656), .Z(n3658) );
  XOR U3870 ( .A(n3746), .B(n3747), .Z(n3656) );
  ANDN U3871 ( .B(n3748), .A(n3749), .Z(n3746) );
  AND U3872 ( .A(b[6]), .B(a[13]), .Z(n3745) );
  XNOR U3873 ( .A(n3750), .B(n3661), .Z(n3663) );
  XOR U3874 ( .A(n3751), .B(n3752), .Z(n3661) );
  ANDN U3875 ( .B(n3753), .A(n3754), .Z(n3751) );
  AND U3876 ( .A(b[5]), .B(a[14]), .Z(n3750) );
  XNOR U3877 ( .A(n3755), .B(n3666), .Z(n3668) );
  XOR U3878 ( .A(n3756), .B(n3757), .Z(n3666) );
  ANDN U3879 ( .B(n3758), .A(n3759), .Z(n3756) );
  AND U3880 ( .A(b[4]), .B(a[15]), .Z(n3755) );
  XNOR U3881 ( .A(n3760), .B(n3761), .Z(n3680) );
  NANDN U3882 ( .A(n3762), .B(n3763), .Z(n3761) );
  XNOR U3883 ( .A(n3764), .B(n3671), .Z(n3673) );
  XNOR U3884 ( .A(n3765), .B(n3766), .Z(n3671) );
  AND U3885 ( .A(n3767), .B(n3768), .Z(n3765) );
  AND U3886 ( .A(b[3]), .B(a[16]), .Z(n3764) );
  XOR U3887 ( .A(n3687), .B(n3686), .Z(swire[18]) );
  XOR U3888 ( .A(sreg[82]), .B(n3685), .Z(n3686) );
  XOR U3889 ( .A(n3692), .B(n3769), .Z(n3687) );
  XNOR U3890 ( .A(n3691), .B(n3685), .Z(n3769) );
  XOR U3891 ( .A(n3770), .B(n3771), .Z(n3685) );
  NOR U3892 ( .A(n3772), .B(n3773), .Z(n3770) );
  NAND U3893 ( .A(a[18]), .B(b[0]), .Z(n3691) );
  XNOR U3894 ( .A(n3762), .B(n3763), .Z(n3692) );
  XOR U3895 ( .A(n3760), .B(n3774), .Z(n3763) );
  NAND U3896 ( .A(b[1]), .B(a[17]), .Z(n3774) );
  XOR U3897 ( .A(n3768), .B(n3775), .Z(n3762) );
  XOR U3898 ( .A(n3760), .B(n3767), .Z(n3775) );
  XNOR U3899 ( .A(n3776), .B(n3766), .Z(n3767) );
  AND U3900 ( .A(b[2]), .B(a[16]), .Z(n3776) );
  NANDN U3901 ( .A(n3777), .B(n3778), .Z(n3760) );
  XOR U3902 ( .A(n3766), .B(n3758), .Z(n3779) );
  XNOR U3903 ( .A(n3757), .B(n3753), .Z(n3780) );
  XNOR U3904 ( .A(n3752), .B(n3748), .Z(n3781) );
  XNOR U3905 ( .A(n3747), .B(n3743), .Z(n3782) );
  XNOR U3906 ( .A(n3742), .B(n3738), .Z(n3783) );
  XNOR U3907 ( .A(n3737), .B(n3733), .Z(n3784) );
  XNOR U3908 ( .A(n3732), .B(n3728), .Z(n3785) );
  XNOR U3909 ( .A(n3727), .B(n3723), .Z(n3786) );
  XNOR U3910 ( .A(n3722), .B(n3718), .Z(n3787) );
  XOR U3911 ( .A(n3717), .B(n3714), .Z(n3788) );
  XOR U3912 ( .A(n3789), .B(n3790), .Z(n3714) );
  XOR U3913 ( .A(n3712), .B(n3791), .Z(n3790) );
  XOR U3914 ( .A(n3792), .B(n3793), .Z(n3791) );
  XOR U3915 ( .A(n3794), .B(n3795), .Z(n3793) );
  NAND U3916 ( .A(b[14]), .B(a[4]), .Z(n3795) );
  AND U3917 ( .A(b[15]), .B(a[3]), .Z(n3794) );
  XOR U3918 ( .A(n3796), .B(n3792), .Z(n3789) );
  XOR U3919 ( .A(n3797), .B(n3798), .Z(n3792) );
  NOR U3920 ( .A(n3799), .B(n3800), .Z(n3797) );
  AND U3921 ( .A(b[13]), .B(a[5]), .Z(n3796) );
  XNOR U3922 ( .A(n3801), .B(n3712), .Z(n3713) );
  XOR U3923 ( .A(n3802), .B(n3803), .Z(n3712) );
  ANDN U3924 ( .B(n3804), .A(n3805), .Z(n3802) );
  AND U3925 ( .A(b[12]), .B(a[6]), .Z(n3801) );
  XNOR U3926 ( .A(n3806), .B(n3717), .Z(n3719) );
  XOR U3927 ( .A(n3807), .B(n3808), .Z(n3717) );
  ANDN U3928 ( .B(n3809), .A(n3810), .Z(n3807) );
  AND U3929 ( .A(b[11]), .B(a[7]), .Z(n3806) );
  XNOR U3930 ( .A(n3811), .B(n3722), .Z(n3724) );
  XOR U3931 ( .A(n3812), .B(n3813), .Z(n3722) );
  ANDN U3932 ( .B(n3814), .A(n3815), .Z(n3812) );
  AND U3933 ( .A(b[10]), .B(a[8]), .Z(n3811) );
  XNOR U3934 ( .A(n3816), .B(n3727), .Z(n3729) );
  XOR U3935 ( .A(n3817), .B(n3818), .Z(n3727) );
  ANDN U3936 ( .B(n3819), .A(n3820), .Z(n3817) );
  AND U3937 ( .A(b[9]), .B(a[9]), .Z(n3816) );
  XNOR U3938 ( .A(n3821), .B(n3732), .Z(n3734) );
  XOR U3939 ( .A(n3822), .B(n3823), .Z(n3732) );
  ANDN U3940 ( .B(n3824), .A(n3825), .Z(n3822) );
  AND U3941 ( .A(b[8]), .B(a[10]), .Z(n3821) );
  XNOR U3942 ( .A(n3826), .B(n3737), .Z(n3739) );
  XOR U3943 ( .A(n3827), .B(n3828), .Z(n3737) );
  ANDN U3944 ( .B(n3829), .A(n3830), .Z(n3827) );
  AND U3945 ( .A(b[7]), .B(a[11]), .Z(n3826) );
  XNOR U3946 ( .A(n3831), .B(n3742), .Z(n3744) );
  XOR U3947 ( .A(n3832), .B(n3833), .Z(n3742) );
  ANDN U3948 ( .B(n3834), .A(n3835), .Z(n3832) );
  AND U3949 ( .A(b[6]), .B(a[12]), .Z(n3831) );
  XNOR U3950 ( .A(n3836), .B(n3747), .Z(n3749) );
  XOR U3951 ( .A(n3837), .B(n3838), .Z(n3747) );
  ANDN U3952 ( .B(n3839), .A(n3840), .Z(n3837) );
  AND U3953 ( .A(b[5]), .B(a[13]), .Z(n3836) );
  XNOR U3954 ( .A(n3841), .B(n3752), .Z(n3754) );
  XOR U3955 ( .A(n3842), .B(n3843), .Z(n3752) );
  ANDN U3956 ( .B(n3844), .A(n3845), .Z(n3842) );
  AND U3957 ( .A(b[4]), .B(a[14]), .Z(n3841) );
  XNOR U3958 ( .A(n3846), .B(n3847), .Z(n3766) );
  NANDN U3959 ( .A(n3848), .B(n3849), .Z(n3847) );
  XNOR U3960 ( .A(n3850), .B(n3757), .Z(n3759) );
  XNOR U3961 ( .A(n3851), .B(n3852), .Z(n3757) );
  AND U3962 ( .A(n3853), .B(n3854), .Z(n3851) );
  AND U3963 ( .A(b[3]), .B(a[15]), .Z(n3850) );
  XOR U3964 ( .A(n3773), .B(n3772), .Z(swire[17]) );
  XOR U3965 ( .A(sreg[81]), .B(n3771), .Z(n3772) );
  XOR U3966 ( .A(n3778), .B(n3855), .Z(n3773) );
  XNOR U3967 ( .A(n3777), .B(n3771), .Z(n3855) );
  XOR U3968 ( .A(n3856), .B(n3857), .Z(n3771) );
  NOR U3969 ( .A(n3858), .B(n3859), .Z(n3856) );
  NAND U3970 ( .A(a[17]), .B(b[0]), .Z(n3777) );
  XNOR U3971 ( .A(n3848), .B(n3849), .Z(n3778) );
  XOR U3972 ( .A(n3846), .B(n3860), .Z(n3849) );
  NAND U3973 ( .A(b[1]), .B(a[16]), .Z(n3860) );
  XOR U3974 ( .A(n3854), .B(n3861), .Z(n3848) );
  XOR U3975 ( .A(n3846), .B(n3853), .Z(n3861) );
  XNOR U3976 ( .A(n3862), .B(n3852), .Z(n3853) );
  AND U3977 ( .A(b[2]), .B(a[15]), .Z(n3862) );
  NANDN U3978 ( .A(n3863), .B(n3864), .Z(n3846) );
  XOR U3979 ( .A(n3852), .B(n3844), .Z(n3865) );
  XNOR U3980 ( .A(n3843), .B(n3839), .Z(n3866) );
  XNOR U3981 ( .A(n3838), .B(n3834), .Z(n3867) );
  XNOR U3982 ( .A(n3833), .B(n3829), .Z(n3868) );
  XNOR U3983 ( .A(n3828), .B(n3824), .Z(n3869) );
  XNOR U3984 ( .A(n3823), .B(n3819), .Z(n3870) );
  XNOR U3985 ( .A(n3818), .B(n3814), .Z(n3871) );
  XNOR U3986 ( .A(n3813), .B(n3809), .Z(n3872) );
  XNOR U3987 ( .A(n3808), .B(n3804), .Z(n3873) );
  XOR U3988 ( .A(n3803), .B(n3800), .Z(n3874) );
  XOR U3989 ( .A(n3875), .B(n3876), .Z(n3800) );
  XOR U3990 ( .A(n3798), .B(n3877), .Z(n3876) );
  XOR U3991 ( .A(n3878), .B(n3879), .Z(n3877) );
  XOR U3992 ( .A(n3880), .B(n3881), .Z(n3879) );
  NAND U3993 ( .A(b[14]), .B(a[3]), .Z(n3881) );
  AND U3994 ( .A(b[15]), .B(a[2]), .Z(n3880) );
  XOR U3995 ( .A(n3882), .B(n3878), .Z(n3875) );
  XOR U3996 ( .A(n3883), .B(n3884), .Z(n3878) );
  NOR U3997 ( .A(n3885), .B(n3886), .Z(n3883) );
  AND U3998 ( .A(b[13]), .B(a[4]), .Z(n3882) );
  XNOR U3999 ( .A(n3887), .B(n3798), .Z(n3799) );
  XOR U4000 ( .A(n3888), .B(n3889), .Z(n3798) );
  ANDN U4001 ( .B(n3890), .A(n3891), .Z(n3888) );
  AND U4002 ( .A(b[12]), .B(a[5]), .Z(n3887) );
  XNOR U4003 ( .A(n3892), .B(n3803), .Z(n3805) );
  XOR U4004 ( .A(n3893), .B(n3894), .Z(n3803) );
  ANDN U4005 ( .B(n3895), .A(n3896), .Z(n3893) );
  AND U4006 ( .A(b[11]), .B(a[6]), .Z(n3892) );
  XNOR U4007 ( .A(n3897), .B(n3808), .Z(n3810) );
  XOR U4008 ( .A(n3898), .B(n3899), .Z(n3808) );
  ANDN U4009 ( .B(n3900), .A(n3901), .Z(n3898) );
  AND U4010 ( .A(b[10]), .B(a[7]), .Z(n3897) );
  XNOR U4011 ( .A(n3902), .B(n3813), .Z(n3815) );
  XOR U4012 ( .A(n3903), .B(n3904), .Z(n3813) );
  ANDN U4013 ( .B(n3905), .A(n3906), .Z(n3903) );
  AND U4014 ( .A(b[9]), .B(a[8]), .Z(n3902) );
  XNOR U4015 ( .A(n3907), .B(n3818), .Z(n3820) );
  XOR U4016 ( .A(n3908), .B(n3909), .Z(n3818) );
  ANDN U4017 ( .B(n3910), .A(n3911), .Z(n3908) );
  AND U4018 ( .A(b[8]), .B(a[9]), .Z(n3907) );
  XNOR U4019 ( .A(n3912), .B(n3823), .Z(n3825) );
  XOR U4020 ( .A(n3913), .B(n3914), .Z(n3823) );
  ANDN U4021 ( .B(n3915), .A(n3916), .Z(n3913) );
  AND U4022 ( .A(b[7]), .B(a[10]), .Z(n3912) );
  XNOR U4023 ( .A(n3917), .B(n3828), .Z(n3830) );
  XOR U4024 ( .A(n3918), .B(n3919), .Z(n3828) );
  ANDN U4025 ( .B(n3920), .A(n3921), .Z(n3918) );
  AND U4026 ( .A(b[6]), .B(a[11]), .Z(n3917) );
  XNOR U4027 ( .A(n3922), .B(n3833), .Z(n3835) );
  XOR U4028 ( .A(n3923), .B(n3924), .Z(n3833) );
  ANDN U4029 ( .B(n3925), .A(n3926), .Z(n3923) );
  AND U4030 ( .A(b[5]), .B(a[12]), .Z(n3922) );
  XNOR U4031 ( .A(n3927), .B(n3838), .Z(n3840) );
  XOR U4032 ( .A(n3928), .B(n3929), .Z(n3838) );
  ANDN U4033 ( .B(n3930), .A(n3931), .Z(n3928) );
  AND U4034 ( .A(b[4]), .B(a[13]), .Z(n3927) );
  XNOR U4035 ( .A(n3932), .B(n3933), .Z(n3852) );
  NANDN U4036 ( .A(n3934), .B(n3935), .Z(n3933) );
  XNOR U4037 ( .A(n3936), .B(n3843), .Z(n3845) );
  XNOR U4038 ( .A(n3937), .B(n3938), .Z(n3843) );
  AND U4039 ( .A(n3939), .B(n3940), .Z(n3937) );
  AND U4040 ( .A(b[3]), .B(a[14]), .Z(n3936) );
  XOR U4041 ( .A(n3859), .B(n3858), .Z(swire[16]) );
  XOR U4042 ( .A(sreg[80]), .B(n3857), .Z(n3858) );
  XOR U4043 ( .A(n3864), .B(n3941), .Z(n3859) );
  XNOR U4044 ( .A(n3863), .B(n3857), .Z(n3941) );
  XOR U4045 ( .A(n3942), .B(n3943), .Z(n3857) );
  NOR U4046 ( .A(n3944), .B(n3945), .Z(n3942) );
  NAND U4047 ( .A(a[16]), .B(b[0]), .Z(n3863) );
  XNOR U4048 ( .A(n3934), .B(n3935), .Z(n3864) );
  XOR U4049 ( .A(n3932), .B(n3946), .Z(n3935) );
  NAND U4050 ( .A(b[1]), .B(a[15]), .Z(n3946) );
  XOR U4051 ( .A(n3940), .B(n3947), .Z(n3934) );
  XOR U4052 ( .A(n3932), .B(n3939), .Z(n3947) );
  XNOR U4053 ( .A(n3948), .B(n3938), .Z(n3939) );
  AND U4054 ( .A(b[2]), .B(a[14]), .Z(n3948) );
  NANDN U4055 ( .A(n3949), .B(n3950), .Z(n3932) );
  XOR U4056 ( .A(n3938), .B(n3930), .Z(n3951) );
  XNOR U4057 ( .A(n3929), .B(n3925), .Z(n3952) );
  XNOR U4058 ( .A(n3924), .B(n3920), .Z(n3953) );
  XNOR U4059 ( .A(n3919), .B(n3915), .Z(n3954) );
  XNOR U4060 ( .A(n3914), .B(n3910), .Z(n3955) );
  XNOR U4061 ( .A(n3909), .B(n3905), .Z(n3956) );
  XNOR U4062 ( .A(n3904), .B(n3900), .Z(n3957) );
  XNOR U4063 ( .A(n3899), .B(n3895), .Z(n3958) );
  XNOR U4064 ( .A(n3894), .B(n3890), .Z(n3959) );
  XOR U4065 ( .A(n3889), .B(n3886), .Z(n3960) );
  XOR U4066 ( .A(n3961), .B(n3962), .Z(n3886) );
  XOR U4067 ( .A(n3884), .B(n3963), .Z(n3962) );
  XOR U4068 ( .A(n3964), .B(n3965), .Z(n3963) );
  XOR U4069 ( .A(n3966), .B(n3967), .Z(n3965) );
  NAND U4070 ( .A(b[14]), .B(a[2]), .Z(n3967) );
  AND U4071 ( .A(b[15]), .B(a[1]), .Z(n3966) );
  XOR U4072 ( .A(n3968), .B(n3964), .Z(n3961) );
  XOR U4073 ( .A(n3969), .B(n3970), .Z(n3964) );
  NOR U4074 ( .A(n3971), .B(n3972), .Z(n3969) );
  AND U4075 ( .A(b[13]), .B(a[3]), .Z(n3968) );
  XNOR U4076 ( .A(n3973), .B(n3884), .Z(n3885) );
  XOR U4077 ( .A(n3974), .B(n3975), .Z(n3884) );
  ANDN U4078 ( .B(n3976), .A(n3977), .Z(n3974) );
  AND U4079 ( .A(b[12]), .B(a[4]), .Z(n3973) );
  XNOR U4080 ( .A(n3978), .B(n3889), .Z(n3891) );
  XOR U4081 ( .A(n3979), .B(n3980), .Z(n3889) );
  ANDN U4082 ( .B(n3981), .A(n3982), .Z(n3979) );
  AND U4083 ( .A(b[11]), .B(a[5]), .Z(n3978) );
  XNOR U4084 ( .A(n3983), .B(n3894), .Z(n3896) );
  XOR U4085 ( .A(n3984), .B(n3985), .Z(n3894) );
  ANDN U4086 ( .B(n3986), .A(n3987), .Z(n3984) );
  AND U4087 ( .A(b[10]), .B(a[6]), .Z(n3983) );
  XNOR U4088 ( .A(n3988), .B(n3899), .Z(n3901) );
  XOR U4089 ( .A(n3989), .B(n3990), .Z(n3899) );
  ANDN U4090 ( .B(n3991), .A(n3992), .Z(n3989) );
  AND U4091 ( .A(b[9]), .B(a[7]), .Z(n3988) );
  XNOR U4092 ( .A(n3993), .B(n3904), .Z(n3906) );
  XOR U4093 ( .A(n3994), .B(n3995), .Z(n3904) );
  ANDN U4094 ( .B(n3996), .A(n3997), .Z(n3994) );
  AND U4095 ( .A(b[8]), .B(a[8]), .Z(n3993) );
  XNOR U4096 ( .A(n3998), .B(n3909), .Z(n3911) );
  XOR U4097 ( .A(n3999), .B(n4000), .Z(n3909) );
  ANDN U4098 ( .B(n4001), .A(n4002), .Z(n3999) );
  AND U4099 ( .A(b[7]), .B(a[9]), .Z(n3998) );
  XNOR U4100 ( .A(n4003), .B(n3914), .Z(n3916) );
  XOR U4101 ( .A(n4004), .B(n4005), .Z(n3914) );
  ANDN U4102 ( .B(n4006), .A(n4007), .Z(n4004) );
  AND U4103 ( .A(b[6]), .B(a[10]), .Z(n4003) );
  XNOR U4104 ( .A(n4008), .B(n3919), .Z(n3921) );
  XOR U4105 ( .A(n4009), .B(n4010), .Z(n3919) );
  ANDN U4106 ( .B(n4011), .A(n4012), .Z(n4009) );
  AND U4107 ( .A(b[5]), .B(a[11]), .Z(n4008) );
  XNOR U4108 ( .A(n4013), .B(n3924), .Z(n3926) );
  XOR U4109 ( .A(n4014), .B(n4015), .Z(n3924) );
  ANDN U4110 ( .B(n4016), .A(n4017), .Z(n4014) );
  AND U4111 ( .A(b[4]), .B(a[12]), .Z(n4013) );
  XNOR U4112 ( .A(n4018), .B(n4019), .Z(n3938) );
  NANDN U4113 ( .A(n4020), .B(n4021), .Z(n4019) );
  XNOR U4114 ( .A(n4022), .B(n3929), .Z(n3931) );
  XNOR U4115 ( .A(n4023), .B(n4024), .Z(n3929) );
  AND U4116 ( .A(n4025), .B(n4026), .Z(n4023) );
  AND U4117 ( .A(b[3]), .B(a[13]), .Z(n4022) );
  XOR U4118 ( .A(n3945), .B(n3944), .Z(c[63]) );
  XOR U4119 ( .A(sreg[79]), .B(n3943), .Z(n3944) );
  XOR U4120 ( .A(n3950), .B(n4027), .Z(n3945) );
  XNOR U4121 ( .A(n3949), .B(n3943), .Z(n4027) );
  XOR U4122 ( .A(n4028), .B(n4029), .Z(n3943) );
  NOR U4123 ( .A(n4030), .B(n4031), .Z(n4028) );
  NAND U4124 ( .A(a[15]), .B(b[0]), .Z(n3949) );
  XNOR U4125 ( .A(n4020), .B(n4021), .Z(n3950) );
  XOR U4126 ( .A(n4018), .B(n4032), .Z(n4021) );
  NAND U4127 ( .A(b[1]), .B(a[14]), .Z(n4032) );
  XOR U4128 ( .A(n4026), .B(n4033), .Z(n4020) );
  XOR U4129 ( .A(n4018), .B(n4025), .Z(n4033) );
  XNOR U4130 ( .A(n4034), .B(n4024), .Z(n4025) );
  AND U4131 ( .A(b[2]), .B(a[13]), .Z(n4034) );
  NANDN U4132 ( .A(n4035), .B(n4036), .Z(n4018) );
  XOR U4133 ( .A(n4024), .B(n4016), .Z(n4037) );
  XNOR U4134 ( .A(n4015), .B(n4011), .Z(n4038) );
  XNOR U4135 ( .A(n4010), .B(n4006), .Z(n4039) );
  XNOR U4136 ( .A(n4005), .B(n4001), .Z(n4040) );
  XNOR U4137 ( .A(n4000), .B(n3996), .Z(n4041) );
  XNOR U4138 ( .A(n3995), .B(n3991), .Z(n4042) );
  XNOR U4139 ( .A(n3990), .B(n3986), .Z(n4043) );
  XNOR U4140 ( .A(n3985), .B(n3981), .Z(n4044) );
  XNOR U4141 ( .A(n3980), .B(n3976), .Z(n4045) );
  XOR U4142 ( .A(n3975), .B(n3972), .Z(n4046) );
  XOR U4143 ( .A(n4047), .B(n4048), .Z(n3972) );
  XOR U4144 ( .A(n3970), .B(n4049), .Z(n4048) );
  XOR U4145 ( .A(n4050), .B(n4051), .Z(n4049) );
  XOR U4146 ( .A(n4052), .B(n4053), .Z(n4051) );
  NAND U4147 ( .A(b[14]), .B(a[1]), .Z(n4053) );
  AND U4148 ( .A(b[15]), .B(a[0]), .Z(n4052) );
  XOR U4149 ( .A(n4054), .B(n4050), .Z(n4047) );
  XOR U4150 ( .A(n4055), .B(n4056), .Z(n4050) );
  NOR U4151 ( .A(n4057), .B(n4058), .Z(n4055) );
  AND U4152 ( .A(b[13]), .B(a[2]), .Z(n4054) );
  XNOR U4153 ( .A(n4059), .B(n3970), .Z(n3971) );
  XOR U4154 ( .A(n4060), .B(n4061), .Z(n3970) );
  ANDN U4155 ( .B(n4062), .A(n4063), .Z(n4060) );
  AND U4156 ( .A(b[12]), .B(a[3]), .Z(n4059) );
  XNOR U4157 ( .A(n4064), .B(n3975), .Z(n3977) );
  XOR U4158 ( .A(n4065), .B(n4066), .Z(n3975) );
  ANDN U4159 ( .B(n4067), .A(n4068), .Z(n4065) );
  AND U4160 ( .A(b[11]), .B(a[4]), .Z(n4064) );
  XNOR U4161 ( .A(n4069), .B(n3980), .Z(n3982) );
  XOR U4162 ( .A(n4070), .B(n4071), .Z(n3980) );
  ANDN U4163 ( .B(n4072), .A(n4073), .Z(n4070) );
  AND U4164 ( .A(b[10]), .B(a[5]), .Z(n4069) );
  XNOR U4165 ( .A(n4074), .B(n3985), .Z(n3987) );
  XOR U4166 ( .A(n4075), .B(n4076), .Z(n3985) );
  ANDN U4167 ( .B(n4077), .A(n4078), .Z(n4075) );
  AND U4168 ( .A(b[9]), .B(a[6]), .Z(n4074) );
  XNOR U4169 ( .A(n4079), .B(n3990), .Z(n3992) );
  XOR U4170 ( .A(n4080), .B(n4081), .Z(n3990) );
  ANDN U4171 ( .B(n4082), .A(n4083), .Z(n4080) );
  AND U4172 ( .A(b[8]), .B(a[7]), .Z(n4079) );
  XNOR U4173 ( .A(n4084), .B(n3995), .Z(n3997) );
  XOR U4174 ( .A(n4085), .B(n4086), .Z(n3995) );
  ANDN U4175 ( .B(n4087), .A(n4088), .Z(n4085) );
  AND U4176 ( .A(b[7]), .B(a[8]), .Z(n4084) );
  XNOR U4177 ( .A(n4089), .B(n4000), .Z(n4002) );
  XOR U4178 ( .A(n4090), .B(n4091), .Z(n4000) );
  ANDN U4179 ( .B(n4092), .A(n4093), .Z(n4090) );
  AND U4180 ( .A(b[6]), .B(a[9]), .Z(n4089) );
  XNOR U4181 ( .A(n4094), .B(n4005), .Z(n4007) );
  XOR U4182 ( .A(n4095), .B(n4096), .Z(n4005) );
  ANDN U4183 ( .B(n4097), .A(n4098), .Z(n4095) );
  AND U4184 ( .A(b[5]), .B(a[10]), .Z(n4094) );
  XNOR U4185 ( .A(n4099), .B(n4010), .Z(n4012) );
  XOR U4186 ( .A(n4100), .B(n4101), .Z(n4010) );
  ANDN U4187 ( .B(n4102), .A(n4103), .Z(n4100) );
  AND U4188 ( .A(b[4]), .B(a[11]), .Z(n4099) );
  XNOR U4189 ( .A(n4104), .B(n4105), .Z(n4024) );
  NANDN U4190 ( .A(n4106), .B(n4107), .Z(n4105) );
  XNOR U4191 ( .A(n4108), .B(n4015), .Z(n4017) );
  XNOR U4192 ( .A(n4109), .B(n4110), .Z(n4015) );
  AND U4193 ( .A(n4111), .B(n4112), .Z(n4109) );
  AND U4194 ( .A(b[3]), .B(a[12]), .Z(n4108) );
  XOR U4195 ( .A(n4031), .B(n4030), .Z(c[62]) );
  XOR U4196 ( .A(sreg[78]), .B(n4029), .Z(n4030) );
  XOR U4197 ( .A(n4036), .B(n4113), .Z(n4031) );
  XNOR U4198 ( .A(n4035), .B(n4029), .Z(n4113) );
  XOR U4199 ( .A(n4114), .B(n4115), .Z(n4029) );
  NOR U4200 ( .A(n4116), .B(n4117), .Z(n4114) );
  NAND U4201 ( .A(a[14]), .B(b[0]), .Z(n4035) );
  XNOR U4202 ( .A(n4106), .B(n4107), .Z(n4036) );
  XOR U4203 ( .A(n4104), .B(n4118), .Z(n4107) );
  NAND U4204 ( .A(b[1]), .B(a[13]), .Z(n4118) );
  XOR U4205 ( .A(n4112), .B(n4119), .Z(n4106) );
  XOR U4206 ( .A(n4104), .B(n4111), .Z(n4119) );
  XNOR U4207 ( .A(n4120), .B(n4110), .Z(n4111) );
  AND U4208 ( .A(b[2]), .B(a[12]), .Z(n4120) );
  NANDN U4209 ( .A(n4121), .B(n4122), .Z(n4104) );
  XOR U4210 ( .A(n4110), .B(n4102), .Z(n4123) );
  XNOR U4211 ( .A(n4101), .B(n4097), .Z(n4124) );
  XNOR U4212 ( .A(n4096), .B(n4092), .Z(n4125) );
  XNOR U4213 ( .A(n4091), .B(n4087), .Z(n4126) );
  XNOR U4214 ( .A(n4086), .B(n4082), .Z(n4127) );
  XNOR U4215 ( .A(n4081), .B(n4077), .Z(n4128) );
  XNOR U4216 ( .A(n4076), .B(n4072), .Z(n4129) );
  XNOR U4217 ( .A(n4071), .B(n4067), .Z(n4130) );
  XNOR U4218 ( .A(n4066), .B(n4062), .Z(n4131) );
  XOR U4219 ( .A(n4061), .B(n4058), .Z(n4132) );
  XOR U4220 ( .A(n4133), .B(n4134), .Z(n4058) );
  XOR U4221 ( .A(n4056), .B(n4135), .Z(n4134) );
  XOR U4222 ( .A(n4136), .B(n4137), .Z(n4135) );
  AND U4223 ( .A(b[14]), .B(a[0]), .Z(n4136) );
  XNOR U4224 ( .A(n4138), .B(n4137), .Z(n4133) );
  XOR U4225 ( .A(n4139), .B(n4140), .Z(n4137) );
  NOR U4226 ( .A(n4141), .B(n4142), .Z(n4139) );
  AND U4227 ( .A(b[13]), .B(a[1]), .Z(n4138) );
  XNOR U4228 ( .A(n4143), .B(n4056), .Z(n4057) );
  XOR U4229 ( .A(n4144), .B(n4145), .Z(n4056) );
  NOR U4230 ( .A(n4146), .B(n4147), .Z(n4144) );
  AND U4231 ( .A(b[12]), .B(a[2]), .Z(n4143) );
  XNOR U4232 ( .A(n4148), .B(n4061), .Z(n4063) );
  XOR U4233 ( .A(n4149), .B(n4150), .Z(n4061) );
  ANDN U4234 ( .B(n4151), .A(n4152), .Z(n4149) );
  AND U4235 ( .A(b[11]), .B(a[3]), .Z(n4148) );
  XNOR U4236 ( .A(n4153), .B(n4066), .Z(n4068) );
  XOR U4237 ( .A(n4154), .B(n4155), .Z(n4066) );
  ANDN U4238 ( .B(n4156), .A(n4157), .Z(n4154) );
  AND U4239 ( .A(b[10]), .B(a[4]), .Z(n4153) );
  XNOR U4240 ( .A(n4158), .B(n4071), .Z(n4073) );
  XOR U4241 ( .A(n4159), .B(n4160), .Z(n4071) );
  ANDN U4242 ( .B(n4161), .A(n4162), .Z(n4159) );
  AND U4243 ( .A(b[9]), .B(a[5]), .Z(n4158) );
  XNOR U4244 ( .A(n4163), .B(n4076), .Z(n4078) );
  XOR U4245 ( .A(n4164), .B(n4165), .Z(n4076) );
  ANDN U4246 ( .B(n4166), .A(n4167), .Z(n4164) );
  AND U4247 ( .A(b[8]), .B(a[6]), .Z(n4163) );
  XNOR U4248 ( .A(n4168), .B(n4081), .Z(n4083) );
  XOR U4249 ( .A(n4169), .B(n4170), .Z(n4081) );
  ANDN U4250 ( .B(n4171), .A(n4172), .Z(n4169) );
  AND U4251 ( .A(b[7]), .B(a[7]), .Z(n4168) );
  XNOR U4252 ( .A(n4173), .B(n4086), .Z(n4088) );
  XOR U4253 ( .A(n4174), .B(n4175), .Z(n4086) );
  ANDN U4254 ( .B(n4176), .A(n4177), .Z(n4174) );
  AND U4255 ( .A(b[6]), .B(a[8]), .Z(n4173) );
  XNOR U4256 ( .A(n4178), .B(n4091), .Z(n4093) );
  XOR U4257 ( .A(n4179), .B(n4180), .Z(n4091) );
  ANDN U4258 ( .B(n4181), .A(n4182), .Z(n4179) );
  AND U4259 ( .A(b[5]), .B(a[9]), .Z(n4178) );
  XNOR U4260 ( .A(n4183), .B(n4096), .Z(n4098) );
  XOR U4261 ( .A(n4184), .B(n4185), .Z(n4096) );
  ANDN U4262 ( .B(n4186), .A(n4187), .Z(n4184) );
  AND U4263 ( .A(b[4]), .B(a[10]), .Z(n4183) );
  XNOR U4264 ( .A(n4188), .B(n4189), .Z(n4110) );
  NANDN U4265 ( .A(n4190), .B(n4191), .Z(n4189) );
  XNOR U4266 ( .A(n4192), .B(n4101), .Z(n4103) );
  XNOR U4267 ( .A(n4193), .B(n4194), .Z(n4101) );
  AND U4268 ( .A(n4195), .B(n4196), .Z(n4193) );
  AND U4269 ( .A(b[3]), .B(a[11]), .Z(n4192) );
  XOR U4270 ( .A(n4117), .B(n4116), .Z(c[61]) );
  XOR U4271 ( .A(sreg[77]), .B(n4115), .Z(n4116) );
  XOR U4272 ( .A(n4122), .B(n4197), .Z(n4117) );
  XNOR U4273 ( .A(n4121), .B(n4115), .Z(n4197) );
  XOR U4274 ( .A(n4198), .B(n4199), .Z(n4115) );
  NOR U4275 ( .A(n4200), .B(n4201), .Z(n4198) );
  NAND U4276 ( .A(a[13]), .B(b[0]), .Z(n4121) );
  XNOR U4277 ( .A(n4190), .B(n4191), .Z(n4122) );
  XOR U4278 ( .A(n4188), .B(n4202), .Z(n4191) );
  NAND U4279 ( .A(b[1]), .B(a[12]), .Z(n4202) );
  XOR U4280 ( .A(n4196), .B(n4203), .Z(n4190) );
  XOR U4281 ( .A(n4188), .B(n4195), .Z(n4203) );
  XNOR U4282 ( .A(n4204), .B(n4194), .Z(n4195) );
  AND U4283 ( .A(b[2]), .B(a[11]), .Z(n4204) );
  NANDN U4284 ( .A(n4205), .B(n4206), .Z(n4188) );
  XOR U4285 ( .A(n4194), .B(n4186), .Z(n4207) );
  XNOR U4286 ( .A(n4185), .B(n4181), .Z(n4208) );
  XNOR U4287 ( .A(n4180), .B(n4176), .Z(n4209) );
  XNOR U4288 ( .A(n4175), .B(n4171), .Z(n4210) );
  XNOR U4289 ( .A(n4170), .B(n4166), .Z(n4211) );
  XNOR U4290 ( .A(n4165), .B(n4161), .Z(n4212) );
  XNOR U4291 ( .A(n4160), .B(n4156), .Z(n4213) );
  XNOR U4292 ( .A(n4155), .B(n4151), .Z(n4214) );
  XOR U4293 ( .A(n4150), .B(n4147), .Z(n4215) );
  XOR U4294 ( .A(n4141), .B(n4216), .Z(n4147) );
  XNOR U4295 ( .A(n4145), .B(n4142), .Z(n4216) );
  XNOR U4296 ( .A(n4217), .B(n4140), .Z(n4142) );
  AND U4297 ( .A(b[13]), .B(a[0]), .Z(n4217) );
  XNOR U4298 ( .A(n4218), .B(n4140), .Z(n4141) );
  XOR U4299 ( .A(n4219), .B(n4220), .Z(n4140) );
  NOR U4300 ( .A(n4221), .B(n4222), .Z(n4219) );
  AND U4301 ( .A(b[12]), .B(a[1]), .Z(n4218) );
  XNOR U4302 ( .A(n4223), .B(n4145), .Z(n4146) );
  XOR U4303 ( .A(n4224), .B(n4225), .Z(n4145) );
  NOR U4304 ( .A(n4226), .B(n4227), .Z(n4224) );
  AND U4305 ( .A(b[11]), .B(a[2]), .Z(n4223) );
  XNOR U4306 ( .A(n4228), .B(n4150), .Z(n4152) );
  XOR U4307 ( .A(n4229), .B(n4230), .Z(n4150) );
  ANDN U4308 ( .B(n4231), .A(n4232), .Z(n4229) );
  AND U4309 ( .A(b[10]), .B(a[3]), .Z(n4228) );
  XNOR U4310 ( .A(n4233), .B(n4155), .Z(n4157) );
  XOR U4311 ( .A(n4234), .B(n4235), .Z(n4155) );
  ANDN U4312 ( .B(n4236), .A(n4237), .Z(n4234) );
  AND U4313 ( .A(b[9]), .B(a[4]), .Z(n4233) );
  XNOR U4314 ( .A(n4238), .B(n4160), .Z(n4162) );
  XOR U4315 ( .A(n4239), .B(n4240), .Z(n4160) );
  ANDN U4316 ( .B(n4241), .A(n4242), .Z(n4239) );
  AND U4317 ( .A(b[8]), .B(a[5]), .Z(n4238) );
  XNOR U4318 ( .A(n4243), .B(n4165), .Z(n4167) );
  XOR U4319 ( .A(n4244), .B(n4245), .Z(n4165) );
  ANDN U4320 ( .B(n4246), .A(n4247), .Z(n4244) );
  AND U4321 ( .A(b[7]), .B(a[6]), .Z(n4243) );
  XNOR U4322 ( .A(n4248), .B(n4170), .Z(n4172) );
  XOR U4323 ( .A(n4249), .B(n4250), .Z(n4170) );
  ANDN U4324 ( .B(n4251), .A(n4252), .Z(n4249) );
  AND U4325 ( .A(b[6]), .B(a[7]), .Z(n4248) );
  XNOR U4326 ( .A(n4253), .B(n4175), .Z(n4177) );
  XOR U4327 ( .A(n4254), .B(n4255), .Z(n4175) );
  ANDN U4328 ( .B(n4256), .A(n4257), .Z(n4254) );
  AND U4329 ( .A(b[5]), .B(a[8]), .Z(n4253) );
  XNOR U4330 ( .A(n4258), .B(n4180), .Z(n4182) );
  XOR U4331 ( .A(n4259), .B(n4260), .Z(n4180) );
  ANDN U4332 ( .B(n4261), .A(n4262), .Z(n4259) );
  AND U4333 ( .A(b[4]), .B(a[9]), .Z(n4258) );
  XNOR U4334 ( .A(n4263), .B(n4264), .Z(n4194) );
  NANDN U4335 ( .A(n4265), .B(n4266), .Z(n4264) );
  XNOR U4336 ( .A(n4267), .B(n4185), .Z(n4187) );
  XNOR U4337 ( .A(n4268), .B(n4269), .Z(n4185) );
  AND U4338 ( .A(n4270), .B(n4271), .Z(n4268) );
  AND U4339 ( .A(b[3]), .B(a[10]), .Z(n4267) );
  XOR U4340 ( .A(n4201), .B(n4200), .Z(c[60]) );
  XOR U4341 ( .A(sreg[76]), .B(n4199), .Z(n4200) );
  XOR U4342 ( .A(n4206), .B(n4272), .Z(n4201) );
  XNOR U4343 ( .A(n4205), .B(n4199), .Z(n4272) );
  XOR U4344 ( .A(n4273), .B(n4274), .Z(n4199) );
  NOR U4345 ( .A(n4275), .B(n4276), .Z(n4273) );
  NAND U4346 ( .A(a[12]), .B(b[0]), .Z(n4205) );
  XNOR U4347 ( .A(n4265), .B(n4266), .Z(n4206) );
  XOR U4348 ( .A(n4263), .B(n4277), .Z(n4266) );
  NAND U4349 ( .A(b[1]), .B(a[11]), .Z(n4277) );
  XOR U4350 ( .A(n4271), .B(n4278), .Z(n4265) );
  XOR U4351 ( .A(n4263), .B(n4270), .Z(n4278) );
  XNOR U4352 ( .A(n4279), .B(n4269), .Z(n4270) );
  AND U4353 ( .A(b[2]), .B(a[10]), .Z(n4279) );
  NANDN U4354 ( .A(n4280), .B(n4281), .Z(n4263) );
  XOR U4355 ( .A(n4269), .B(n4261), .Z(n4282) );
  XNOR U4356 ( .A(n4260), .B(n4256), .Z(n4283) );
  XNOR U4357 ( .A(n4255), .B(n4251), .Z(n4284) );
  XNOR U4358 ( .A(n4250), .B(n4246), .Z(n4285) );
  XNOR U4359 ( .A(n4245), .B(n4241), .Z(n4286) );
  XNOR U4360 ( .A(n4240), .B(n4236), .Z(n4287) );
  XNOR U4361 ( .A(n4235), .B(n4231), .Z(n4288) );
  XOR U4362 ( .A(n4230), .B(n4227), .Z(n4289) );
  XOR U4363 ( .A(n4221), .B(n4290), .Z(n4227) );
  XNOR U4364 ( .A(n4225), .B(n4222), .Z(n4290) );
  XNOR U4365 ( .A(n4291), .B(n4220), .Z(n4222) );
  AND U4366 ( .A(b[12]), .B(a[0]), .Z(n4291) );
  XNOR U4367 ( .A(n4292), .B(n4220), .Z(n4221) );
  XOR U4368 ( .A(n4293), .B(n4294), .Z(n4220) );
  NOR U4369 ( .A(n4295), .B(n4296), .Z(n4293) );
  AND U4370 ( .A(b[11]), .B(a[1]), .Z(n4292) );
  XNOR U4371 ( .A(n4297), .B(n4225), .Z(n4226) );
  XOR U4372 ( .A(n4298), .B(n4299), .Z(n4225) );
  NOR U4373 ( .A(n4300), .B(n4301), .Z(n4298) );
  AND U4374 ( .A(b[10]), .B(a[2]), .Z(n4297) );
  XNOR U4375 ( .A(n4302), .B(n4230), .Z(n4232) );
  XOR U4376 ( .A(n4303), .B(n4304), .Z(n4230) );
  ANDN U4377 ( .B(n4305), .A(n4306), .Z(n4303) );
  AND U4378 ( .A(b[9]), .B(a[3]), .Z(n4302) );
  XNOR U4379 ( .A(n4307), .B(n4235), .Z(n4237) );
  XOR U4380 ( .A(n4308), .B(n4309), .Z(n4235) );
  ANDN U4381 ( .B(n4310), .A(n4311), .Z(n4308) );
  AND U4382 ( .A(b[8]), .B(a[4]), .Z(n4307) );
  XNOR U4383 ( .A(n4312), .B(n4240), .Z(n4242) );
  XOR U4384 ( .A(n4313), .B(n4314), .Z(n4240) );
  ANDN U4385 ( .B(n4315), .A(n4316), .Z(n4313) );
  AND U4386 ( .A(b[7]), .B(a[5]), .Z(n4312) );
  XNOR U4387 ( .A(n4317), .B(n4245), .Z(n4247) );
  XOR U4388 ( .A(n4318), .B(n4319), .Z(n4245) );
  ANDN U4389 ( .B(n4320), .A(n4321), .Z(n4318) );
  AND U4390 ( .A(b[6]), .B(a[6]), .Z(n4317) );
  XNOR U4391 ( .A(n4322), .B(n4250), .Z(n4252) );
  XOR U4392 ( .A(n4323), .B(n4324), .Z(n4250) );
  ANDN U4393 ( .B(n4325), .A(n4326), .Z(n4323) );
  AND U4394 ( .A(b[5]), .B(a[7]), .Z(n4322) );
  XNOR U4395 ( .A(n4327), .B(n4255), .Z(n4257) );
  XOR U4396 ( .A(n4328), .B(n4329), .Z(n4255) );
  ANDN U4397 ( .B(n4330), .A(n4331), .Z(n4328) );
  AND U4398 ( .A(b[4]), .B(a[8]), .Z(n4327) );
  XNOR U4399 ( .A(n4332), .B(n4333), .Z(n4269) );
  NANDN U4400 ( .A(n4334), .B(n4335), .Z(n4333) );
  XNOR U4401 ( .A(n4336), .B(n4260), .Z(n4262) );
  XNOR U4402 ( .A(n4337), .B(n4338), .Z(n4260) );
  AND U4403 ( .A(n4339), .B(n4340), .Z(n4337) );
  AND U4404 ( .A(b[3]), .B(a[9]), .Z(n4336) );
  XOR U4405 ( .A(n4276), .B(n4275), .Z(c[59]) );
  XOR U4406 ( .A(sreg[75]), .B(n4274), .Z(n4275) );
  XOR U4407 ( .A(n4281), .B(n4341), .Z(n4276) );
  XNOR U4408 ( .A(n4280), .B(n4274), .Z(n4341) );
  XOR U4409 ( .A(n4342), .B(n4343), .Z(n4274) );
  NOR U4410 ( .A(n4344), .B(n4345), .Z(n4342) );
  NAND U4411 ( .A(a[11]), .B(b[0]), .Z(n4280) );
  XNOR U4412 ( .A(n4334), .B(n4335), .Z(n4281) );
  XOR U4413 ( .A(n4332), .B(n4346), .Z(n4335) );
  NAND U4414 ( .A(b[1]), .B(a[10]), .Z(n4346) );
  XOR U4415 ( .A(n4340), .B(n4347), .Z(n4334) );
  XOR U4416 ( .A(n4332), .B(n4339), .Z(n4347) );
  XNOR U4417 ( .A(n4348), .B(n4338), .Z(n4339) );
  AND U4418 ( .A(b[2]), .B(a[9]), .Z(n4348) );
  NANDN U4419 ( .A(n4349), .B(n4350), .Z(n4332) );
  XOR U4420 ( .A(n4338), .B(n4330), .Z(n4351) );
  XNOR U4421 ( .A(n4329), .B(n4325), .Z(n4352) );
  XNOR U4422 ( .A(n4324), .B(n4320), .Z(n4353) );
  XNOR U4423 ( .A(n4319), .B(n4315), .Z(n4354) );
  XNOR U4424 ( .A(n4314), .B(n4310), .Z(n4355) );
  XNOR U4425 ( .A(n4309), .B(n4305), .Z(n4356) );
  XOR U4426 ( .A(n4304), .B(n4301), .Z(n4357) );
  XOR U4427 ( .A(n4295), .B(n4358), .Z(n4301) );
  XNOR U4428 ( .A(n4299), .B(n4296), .Z(n4358) );
  XNOR U4429 ( .A(n4359), .B(n4294), .Z(n4296) );
  AND U4430 ( .A(b[11]), .B(a[0]), .Z(n4359) );
  XNOR U4431 ( .A(n4360), .B(n4294), .Z(n4295) );
  XOR U4432 ( .A(n4361), .B(n4362), .Z(n4294) );
  NOR U4433 ( .A(n4363), .B(n4364), .Z(n4361) );
  AND U4434 ( .A(b[10]), .B(a[1]), .Z(n4360) );
  XNOR U4435 ( .A(n4365), .B(n4299), .Z(n4300) );
  XOR U4436 ( .A(n4366), .B(n4367), .Z(n4299) );
  NOR U4437 ( .A(n4368), .B(n4369), .Z(n4366) );
  AND U4438 ( .A(b[9]), .B(a[2]), .Z(n4365) );
  XNOR U4439 ( .A(n4370), .B(n4304), .Z(n4306) );
  XOR U4440 ( .A(n4371), .B(n4372), .Z(n4304) );
  ANDN U4441 ( .B(n4373), .A(n4374), .Z(n4371) );
  AND U4442 ( .A(b[8]), .B(a[3]), .Z(n4370) );
  XNOR U4443 ( .A(n4375), .B(n4309), .Z(n4311) );
  XOR U4444 ( .A(n4376), .B(n4377), .Z(n4309) );
  ANDN U4445 ( .B(n4378), .A(n4379), .Z(n4376) );
  AND U4446 ( .A(b[7]), .B(a[4]), .Z(n4375) );
  XNOR U4447 ( .A(n4380), .B(n4314), .Z(n4316) );
  XOR U4448 ( .A(n4381), .B(n4382), .Z(n4314) );
  ANDN U4449 ( .B(n4383), .A(n4384), .Z(n4381) );
  AND U4450 ( .A(b[6]), .B(a[5]), .Z(n4380) );
  XNOR U4451 ( .A(n4385), .B(n4319), .Z(n4321) );
  XOR U4452 ( .A(n4386), .B(n4387), .Z(n4319) );
  ANDN U4453 ( .B(n4388), .A(n4389), .Z(n4386) );
  AND U4454 ( .A(b[5]), .B(a[6]), .Z(n4385) );
  XNOR U4455 ( .A(n4390), .B(n4324), .Z(n4326) );
  XOR U4456 ( .A(n4391), .B(n4392), .Z(n4324) );
  ANDN U4457 ( .B(n4393), .A(n4394), .Z(n4391) );
  AND U4458 ( .A(b[4]), .B(a[7]), .Z(n4390) );
  XNOR U4459 ( .A(n4395), .B(n4396), .Z(n4338) );
  NANDN U4460 ( .A(n4397), .B(n4398), .Z(n4396) );
  XNOR U4461 ( .A(n4399), .B(n4329), .Z(n4331) );
  XNOR U4462 ( .A(n4400), .B(n4401), .Z(n4329) );
  AND U4463 ( .A(n4402), .B(n4403), .Z(n4400) );
  AND U4464 ( .A(b[3]), .B(a[8]), .Z(n4399) );
  XOR U4465 ( .A(n4345), .B(n4344), .Z(c[58]) );
  XOR U4466 ( .A(sreg[74]), .B(n4343), .Z(n4344) );
  XOR U4467 ( .A(n4350), .B(n4404), .Z(n4345) );
  XNOR U4468 ( .A(n4349), .B(n4343), .Z(n4404) );
  XOR U4469 ( .A(n4405), .B(n4406), .Z(n4343) );
  NOR U4470 ( .A(n4407), .B(n4408), .Z(n4405) );
  NAND U4471 ( .A(a[10]), .B(b[0]), .Z(n4349) );
  XNOR U4472 ( .A(n4397), .B(n4398), .Z(n4350) );
  XOR U4473 ( .A(n4395), .B(n4409), .Z(n4398) );
  NAND U4474 ( .A(b[1]), .B(a[9]), .Z(n4409) );
  XOR U4475 ( .A(n4403), .B(n4410), .Z(n4397) );
  XOR U4476 ( .A(n4395), .B(n4402), .Z(n4410) );
  XNOR U4477 ( .A(n4411), .B(n4401), .Z(n4402) );
  AND U4478 ( .A(b[2]), .B(a[8]), .Z(n4411) );
  NANDN U4479 ( .A(n4412), .B(n4413), .Z(n4395) );
  XOR U4480 ( .A(n4401), .B(n4393), .Z(n4414) );
  XNOR U4481 ( .A(n4392), .B(n4388), .Z(n4415) );
  XNOR U4482 ( .A(n4387), .B(n4383), .Z(n4416) );
  XNOR U4483 ( .A(n4382), .B(n4378), .Z(n4417) );
  XNOR U4484 ( .A(n4377), .B(n4373), .Z(n4418) );
  XOR U4485 ( .A(n4372), .B(n4369), .Z(n4419) );
  XOR U4486 ( .A(n4363), .B(n4420), .Z(n4369) );
  XNOR U4487 ( .A(n4367), .B(n4364), .Z(n4420) );
  XNOR U4488 ( .A(n4421), .B(n4362), .Z(n4364) );
  AND U4489 ( .A(b[10]), .B(a[0]), .Z(n4421) );
  XNOR U4490 ( .A(n4422), .B(n4362), .Z(n4363) );
  XOR U4491 ( .A(n4423), .B(n4424), .Z(n4362) );
  NOR U4492 ( .A(n4425), .B(n4426), .Z(n4423) );
  AND U4493 ( .A(b[9]), .B(a[1]), .Z(n4422) );
  XNOR U4494 ( .A(n4427), .B(n4367), .Z(n4368) );
  XOR U4495 ( .A(n4428), .B(n4429), .Z(n4367) );
  NOR U4496 ( .A(n4430), .B(n4431), .Z(n4428) );
  AND U4497 ( .A(b[8]), .B(a[2]), .Z(n4427) );
  XNOR U4498 ( .A(n4432), .B(n4372), .Z(n4374) );
  XOR U4499 ( .A(n4433), .B(n4434), .Z(n4372) );
  ANDN U4500 ( .B(n4435), .A(n4436), .Z(n4433) );
  AND U4501 ( .A(b[7]), .B(a[3]), .Z(n4432) );
  XNOR U4502 ( .A(n4437), .B(n4377), .Z(n4379) );
  XOR U4503 ( .A(n4438), .B(n4439), .Z(n4377) );
  ANDN U4504 ( .B(n4440), .A(n4441), .Z(n4438) );
  AND U4505 ( .A(b[6]), .B(a[4]), .Z(n4437) );
  XNOR U4506 ( .A(n4442), .B(n4382), .Z(n4384) );
  XOR U4507 ( .A(n4443), .B(n4444), .Z(n4382) );
  ANDN U4508 ( .B(n4445), .A(n4446), .Z(n4443) );
  AND U4509 ( .A(b[5]), .B(a[5]), .Z(n4442) );
  XNOR U4510 ( .A(n4447), .B(n4387), .Z(n4389) );
  XOR U4511 ( .A(n4448), .B(n4449), .Z(n4387) );
  ANDN U4512 ( .B(n4450), .A(n4451), .Z(n4448) );
  AND U4513 ( .A(b[4]), .B(a[6]), .Z(n4447) );
  XNOR U4514 ( .A(n4452), .B(n4453), .Z(n4401) );
  NANDN U4515 ( .A(n4454), .B(n4455), .Z(n4453) );
  XNOR U4516 ( .A(n4456), .B(n4392), .Z(n4394) );
  XNOR U4517 ( .A(n4457), .B(n4458), .Z(n4392) );
  AND U4518 ( .A(n4459), .B(n4460), .Z(n4457) );
  AND U4519 ( .A(b[3]), .B(a[7]), .Z(n4456) );
  XOR U4520 ( .A(n4408), .B(n4407), .Z(c[57]) );
  XOR U4521 ( .A(sreg[73]), .B(n4406), .Z(n4407) );
  XOR U4522 ( .A(n4413), .B(n4461), .Z(n4408) );
  XNOR U4523 ( .A(n4412), .B(n4406), .Z(n4461) );
  XOR U4524 ( .A(n4462), .B(n4463), .Z(n4406) );
  NOR U4525 ( .A(n4464), .B(n4465), .Z(n4462) );
  NAND U4526 ( .A(a[9]), .B(b[0]), .Z(n4412) );
  XNOR U4527 ( .A(n4454), .B(n4455), .Z(n4413) );
  XOR U4528 ( .A(n4452), .B(n4466), .Z(n4455) );
  NAND U4529 ( .A(b[1]), .B(a[8]), .Z(n4466) );
  XOR U4530 ( .A(n4460), .B(n4467), .Z(n4454) );
  XOR U4531 ( .A(n4452), .B(n4459), .Z(n4467) );
  XNOR U4532 ( .A(n4468), .B(n4458), .Z(n4459) );
  AND U4533 ( .A(b[2]), .B(a[7]), .Z(n4468) );
  NANDN U4534 ( .A(n4469), .B(n4470), .Z(n4452) );
  XOR U4535 ( .A(n4458), .B(n4450), .Z(n4471) );
  XNOR U4536 ( .A(n4449), .B(n4445), .Z(n4472) );
  XNOR U4537 ( .A(n4444), .B(n4440), .Z(n4473) );
  XNOR U4538 ( .A(n4439), .B(n4435), .Z(n4474) );
  XOR U4539 ( .A(n4434), .B(n4431), .Z(n4475) );
  XOR U4540 ( .A(n4425), .B(n4476), .Z(n4431) );
  XNOR U4541 ( .A(n4429), .B(n4426), .Z(n4476) );
  XNOR U4542 ( .A(n4477), .B(n4424), .Z(n4426) );
  AND U4543 ( .A(b[9]), .B(a[0]), .Z(n4477) );
  XNOR U4544 ( .A(n4478), .B(n4424), .Z(n4425) );
  XOR U4545 ( .A(n4479), .B(n4480), .Z(n4424) );
  NOR U4546 ( .A(n4481), .B(n4482), .Z(n4479) );
  AND U4547 ( .A(b[8]), .B(a[1]), .Z(n4478) );
  XNOR U4548 ( .A(n4483), .B(n4429), .Z(n4430) );
  XOR U4549 ( .A(n4484), .B(n4485), .Z(n4429) );
  NOR U4550 ( .A(n4486), .B(n4487), .Z(n4484) );
  AND U4551 ( .A(b[7]), .B(a[2]), .Z(n4483) );
  XNOR U4552 ( .A(n4488), .B(n4434), .Z(n4436) );
  XOR U4553 ( .A(n4489), .B(n4490), .Z(n4434) );
  ANDN U4554 ( .B(n4491), .A(n4492), .Z(n4489) );
  AND U4555 ( .A(b[6]), .B(a[3]), .Z(n4488) );
  XNOR U4556 ( .A(n4493), .B(n4439), .Z(n4441) );
  XOR U4557 ( .A(n4494), .B(n4495), .Z(n4439) );
  ANDN U4558 ( .B(n4496), .A(n4497), .Z(n4494) );
  AND U4559 ( .A(b[5]), .B(a[4]), .Z(n4493) );
  XNOR U4560 ( .A(n4498), .B(n4444), .Z(n4446) );
  XOR U4561 ( .A(n4499), .B(n4500), .Z(n4444) );
  ANDN U4562 ( .B(n4501), .A(n4502), .Z(n4499) );
  AND U4563 ( .A(b[4]), .B(a[5]), .Z(n4498) );
  XNOR U4564 ( .A(n4503), .B(n4504), .Z(n4458) );
  NANDN U4565 ( .A(n4505), .B(n4506), .Z(n4504) );
  XNOR U4566 ( .A(n4507), .B(n4449), .Z(n4451) );
  XNOR U4567 ( .A(n4508), .B(n4509), .Z(n4449) );
  AND U4568 ( .A(n4510), .B(n4511), .Z(n4508) );
  AND U4569 ( .A(b[3]), .B(a[6]), .Z(n4507) );
  XOR U4570 ( .A(n4465), .B(n4464), .Z(c[56]) );
  XOR U4571 ( .A(sreg[72]), .B(n4463), .Z(n4464) );
  XOR U4572 ( .A(n4470), .B(n4512), .Z(n4465) );
  XNOR U4573 ( .A(n4469), .B(n4463), .Z(n4512) );
  XOR U4574 ( .A(n4513), .B(n4514), .Z(n4463) );
  NOR U4575 ( .A(n4515), .B(n4516), .Z(n4513) );
  NAND U4576 ( .A(a[8]), .B(b[0]), .Z(n4469) );
  XNOR U4577 ( .A(n4505), .B(n4506), .Z(n4470) );
  XOR U4578 ( .A(n4503), .B(n4517), .Z(n4506) );
  NAND U4579 ( .A(b[1]), .B(a[7]), .Z(n4517) );
  XOR U4580 ( .A(n4511), .B(n4518), .Z(n4505) );
  XOR U4581 ( .A(n4503), .B(n4510), .Z(n4518) );
  XNOR U4582 ( .A(n4519), .B(n4509), .Z(n4510) );
  AND U4583 ( .A(b[2]), .B(a[6]), .Z(n4519) );
  NANDN U4584 ( .A(n4520), .B(n4521), .Z(n4503) );
  XOR U4585 ( .A(n4509), .B(n4501), .Z(n4522) );
  XNOR U4586 ( .A(n4500), .B(n4496), .Z(n4523) );
  XNOR U4587 ( .A(n4495), .B(n4491), .Z(n4524) );
  XOR U4588 ( .A(n4490), .B(n4487), .Z(n4525) );
  XOR U4589 ( .A(n4481), .B(n4526), .Z(n4487) );
  XNOR U4590 ( .A(n4485), .B(n4482), .Z(n4526) );
  XNOR U4591 ( .A(n4527), .B(n4480), .Z(n4482) );
  AND U4592 ( .A(b[8]), .B(a[0]), .Z(n4527) );
  XNOR U4593 ( .A(n4528), .B(n4480), .Z(n4481) );
  XOR U4594 ( .A(n4529), .B(n4530), .Z(n4480) );
  NOR U4595 ( .A(n4531), .B(n4532), .Z(n4529) );
  AND U4596 ( .A(b[7]), .B(a[1]), .Z(n4528) );
  XNOR U4597 ( .A(n4533), .B(n4485), .Z(n4486) );
  XOR U4598 ( .A(n4534), .B(n4535), .Z(n4485) );
  NOR U4599 ( .A(n4536), .B(n4537), .Z(n4534) );
  AND U4600 ( .A(b[6]), .B(a[2]), .Z(n4533) );
  XNOR U4601 ( .A(n4538), .B(n4490), .Z(n4492) );
  XOR U4602 ( .A(n4539), .B(n4540), .Z(n4490) );
  ANDN U4603 ( .B(n4541), .A(n4542), .Z(n4539) );
  AND U4604 ( .A(b[5]), .B(a[3]), .Z(n4538) );
  XNOR U4605 ( .A(n4543), .B(n4495), .Z(n4497) );
  XOR U4606 ( .A(n4544), .B(n4545), .Z(n4495) );
  ANDN U4607 ( .B(n4546), .A(n4547), .Z(n4544) );
  AND U4608 ( .A(b[4]), .B(a[4]), .Z(n4543) );
  XNOR U4609 ( .A(n4548), .B(n4549), .Z(n4509) );
  NANDN U4610 ( .A(n4550), .B(n4551), .Z(n4549) );
  XNOR U4611 ( .A(n4552), .B(n4500), .Z(n4502) );
  XNOR U4612 ( .A(n4553), .B(n4554), .Z(n4500) );
  AND U4613 ( .A(n4555), .B(n4556), .Z(n4553) );
  AND U4614 ( .A(b[3]), .B(a[5]), .Z(n4552) );
  XOR U4615 ( .A(n4516), .B(n4515), .Z(c[55]) );
  XOR U4616 ( .A(sreg[71]), .B(n4514), .Z(n4515) );
  XOR U4617 ( .A(n4521), .B(n4557), .Z(n4516) );
  XNOR U4618 ( .A(n4520), .B(n4514), .Z(n4557) );
  XOR U4619 ( .A(n4558), .B(n4559), .Z(n4514) );
  NOR U4620 ( .A(n4560), .B(n4561), .Z(n4558) );
  NAND U4621 ( .A(a[7]), .B(b[0]), .Z(n4520) );
  XNOR U4622 ( .A(n4550), .B(n4551), .Z(n4521) );
  XOR U4623 ( .A(n4548), .B(n4562), .Z(n4551) );
  NAND U4624 ( .A(b[1]), .B(a[6]), .Z(n4562) );
  XOR U4625 ( .A(n4556), .B(n4563), .Z(n4550) );
  XOR U4626 ( .A(n4548), .B(n4555), .Z(n4563) );
  XNOR U4627 ( .A(n4564), .B(n4554), .Z(n4555) );
  AND U4628 ( .A(b[2]), .B(a[5]), .Z(n4564) );
  NANDN U4629 ( .A(n4565), .B(n4566), .Z(n4548) );
  XOR U4630 ( .A(n4554), .B(n4546), .Z(n4567) );
  XNOR U4631 ( .A(n4545), .B(n4541), .Z(n4568) );
  XOR U4632 ( .A(n4540), .B(n4537), .Z(n4569) );
  XOR U4633 ( .A(n4531), .B(n4570), .Z(n4537) );
  XNOR U4634 ( .A(n4535), .B(n4532), .Z(n4570) );
  XNOR U4635 ( .A(n4571), .B(n4530), .Z(n4532) );
  AND U4636 ( .A(b[7]), .B(a[0]), .Z(n4571) );
  XNOR U4637 ( .A(n4572), .B(n4530), .Z(n4531) );
  XOR U4638 ( .A(n4573), .B(n4574), .Z(n4530) );
  NOR U4639 ( .A(n4575), .B(n4576), .Z(n4573) );
  AND U4640 ( .A(b[6]), .B(a[1]), .Z(n4572) );
  XNOR U4641 ( .A(n4577), .B(n4535), .Z(n4536) );
  XOR U4642 ( .A(n4578), .B(n4579), .Z(n4535) );
  NOR U4643 ( .A(n4580), .B(n4581), .Z(n4578) );
  AND U4644 ( .A(b[5]), .B(a[2]), .Z(n4577) );
  XNOR U4645 ( .A(n4582), .B(n4540), .Z(n4542) );
  XOR U4646 ( .A(n4583), .B(n4584), .Z(n4540) );
  ANDN U4647 ( .B(n4585), .A(n4586), .Z(n4583) );
  AND U4648 ( .A(b[4]), .B(a[3]), .Z(n4582) );
  XNOR U4649 ( .A(n4587), .B(n4588), .Z(n4554) );
  NANDN U4650 ( .A(n4589), .B(n4590), .Z(n4588) );
  XNOR U4651 ( .A(n4591), .B(n4545), .Z(n4547) );
  XNOR U4652 ( .A(n4592), .B(n4593), .Z(n4545) );
  AND U4653 ( .A(n4594), .B(n4595), .Z(n4592) );
  AND U4654 ( .A(b[3]), .B(a[4]), .Z(n4591) );
  XOR U4655 ( .A(n4561), .B(n4560), .Z(c[54]) );
  XOR U4656 ( .A(sreg[70]), .B(n4559), .Z(n4560) );
  XOR U4657 ( .A(n4566), .B(n4596), .Z(n4561) );
  XNOR U4658 ( .A(n4565), .B(n4559), .Z(n4596) );
  XOR U4659 ( .A(n4597), .B(n4598), .Z(n4559) );
  NOR U4660 ( .A(n4599), .B(n4600), .Z(n4597) );
  NAND U4661 ( .A(a[6]), .B(b[0]), .Z(n4565) );
  XNOR U4662 ( .A(n4589), .B(n4590), .Z(n4566) );
  XOR U4663 ( .A(n4587), .B(n4601), .Z(n4590) );
  NAND U4664 ( .A(b[1]), .B(a[5]), .Z(n4601) );
  XOR U4665 ( .A(n4595), .B(n4602), .Z(n4589) );
  XOR U4666 ( .A(n4587), .B(n4594), .Z(n4602) );
  XNOR U4667 ( .A(n4603), .B(n4593), .Z(n4594) );
  AND U4668 ( .A(b[2]), .B(a[4]), .Z(n4603) );
  NANDN U4669 ( .A(n4604), .B(n4605), .Z(n4587) );
  XOR U4670 ( .A(n4593), .B(n4585), .Z(n4606) );
  XOR U4671 ( .A(n4584), .B(n4581), .Z(n4607) );
  XOR U4672 ( .A(n4575), .B(n4608), .Z(n4581) );
  XNOR U4673 ( .A(n4579), .B(n4576), .Z(n4608) );
  XNOR U4674 ( .A(n4609), .B(n4574), .Z(n4576) );
  AND U4675 ( .A(b[6]), .B(a[0]), .Z(n4609) );
  XNOR U4676 ( .A(n4610), .B(n4574), .Z(n4575) );
  XOR U4677 ( .A(n4611), .B(n4612), .Z(n4574) );
  NOR U4678 ( .A(n4613), .B(n4614), .Z(n4611) );
  AND U4679 ( .A(b[5]), .B(a[1]), .Z(n4610) );
  XNOR U4680 ( .A(n4615), .B(n4579), .Z(n4580) );
  XOR U4681 ( .A(n4616), .B(n4617), .Z(n4579) );
  NOR U4682 ( .A(n4618), .B(n4619), .Z(n4616) );
  AND U4683 ( .A(b[4]), .B(a[2]), .Z(n4615) );
  XNOR U4684 ( .A(n4620), .B(n4621), .Z(n4593) );
  NANDN U4685 ( .A(n4622), .B(n4623), .Z(n4621) );
  XNOR U4686 ( .A(n4624), .B(n4584), .Z(n4586) );
  XNOR U4687 ( .A(n4625), .B(n4626), .Z(n4584) );
  AND U4688 ( .A(n4627), .B(n4628), .Z(n4625) );
  AND U4689 ( .A(b[3]), .B(a[3]), .Z(n4624) );
  XOR U4690 ( .A(n4600), .B(n4599), .Z(c[53]) );
  XOR U4691 ( .A(sreg[69]), .B(n4598), .Z(n4599) );
  XOR U4692 ( .A(n4605), .B(n4629), .Z(n4600) );
  XNOR U4693 ( .A(n4604), .B(n4598), .Z(n4629) );
  XOR U4694 ( .A(n4630), .B(n4631), .Z(n4598) );
  NOR U4695 ( .A(n4632), .B(n4633), .Z(n4630) );
  NAND U4696 ( .A(a[5]), .B(b[0]), .Z(n4604) );
  XNOR U4697 ( .A(n4622), .B(n4623), .Z(n4605) );
  XOR U4698 ( .A(n4620), .B(n4634), .Z(n4623) );
  NAND U4699 ( .A(b[1]), .B(a[4]), .Z(n4634) );
  XOR U4700 ( .A(n4628), .B(n4635), .Z(n4622) );
  XOR U4701 ( .A(n4620), .B(n4627), .Z(n4635) );
  XNOR U4702 ( .A(n4636), .B(n4626), .Z(n4627) );
  AND U4703 ( .A(b[2]), .B(a[3]), .Z(n4636) );
  NANDN U4704 ( .A(n4637), .B(n4638), .Z(n4620) );
  XNOR U4705 ( .A(n4626), .B(n4619), .Z(n4639) );
  XOR U4706 ( .A(n4613), .B(n4640), .Z(n4619) );
  XNOR U4707 ( .A(n4617), .B(n4614), .Z(n4640) );
  XNOR U4708 ( .A(n4641), .B(n4612), .Z(n4614) );
  AND U4709 ( .A(b[5]), .B(a[0]), .Z(n4641) );
  XNOR U4710 ( .A(n4642), .B(n4612), .Z(n4613) );
  XOR U4711 ( .A(n4643), .B(n4644), .Z(n4612) );
  NOR U4712 ( .A(n4645), .B(n4646), .Z(n4643) );
  AND U4713 ( .A(b[4]), .B(a[1]), .Z(n4642) );
  XNOR U4714 ( .A(n4647), .B(n4648), .Z(n4626) );
  NANDN U4715 ( .A(n4649), .B(n4650), .Z(n4648) );
  XNOR U4716 ( .A(n4651), .B(n4617), .Z(n4618) );
  XNOR U4717 ( .A(n4652), .B(n4653), .Z(n4617) );
  AND U4718 ( .A(n4654), .B(n4655), .Z(n4652) );
  AND U4719 ( .A(b[3]), .B(a[2]), .Z(n4651) );
  XOR U4720 ( .A(n4633), .B(n4632), .Z(c[52]) );
  XOR U4721 ( .A(sreg[68]), .B(n4631), .Z(n4632) );
  XOR U4722 ( .A(n4638), .B(n4656), .Z(n4633) );
  XNOR U4723 ( .A(n4637), .B(n4631), .Z(n4656) );
  XOR U4724 ( .A(n4657), .B(n4658), .Z(n4631) );
  NOR U4725 ( .A(n4659), .B(n4660), .Z(n4657) );
  NAND U4726 ( .A(a[4]), .B(b[0]), .Z(n4637) );
  XNOR U4727 ( .A(n4649), .B(n4650), .Z(n4638) );
  XOR U4728 ( .A(n4647), .B(n4661), .Z(n4650) );
  NAND U4729 ( .A(b[1]), .B(a[3]), .Z(n4661) );
  XOR U4730 ( .A(n4655), .B(n4662), .Z(n4649) );
  XOR U4731 ( .A(n4647), .B(n4654), .Z(n4662) );
  XNOR U4732 ( .A(n4663), .B(n4653), .Z(n4654) );
  AND U4733 ( .A(b[2]), .B(a[2]), .Z(n4663) );
  NANDN U4734 ( .A(n4664), .B(n4665), .Z(n4647) );
  XNOR U4735 ( .A(n4645), .B(n4666), .Z(n4655) );
  XOR U4736 ( .A(n4653), .B(n4646), .Z(n4666) );
  XNOR U4737 ( .A(n4667), .B(n4644), .Z(n4646) );
  AND U4738 ( .A(b[4]), .B(a[0]), .Z(n4667) );
  XNOR U4739 ( .A(n4668), .B(n4669), .Z(n4653) );
  NANDN U4740 ( .A(n4670), .B(n4671), .Z(n4669) );
  XNOR U4741 ( .A(n4672), .B(n4644), .Z(n4645) );
  XNOR U4742 ( .A(n4673), .B(n4674), .Z(n4644) );
  ANDN U4743 ( .B(n4675), .A(n4676), .Z(n4673) );
  AND U4744 ( .A(b[3]), .B(a[1]), .Z(n4672) );
  XOR U4745 ( .A(n4660), .B(n4659), .Z(c[51]) );
  XOR U4746 ( .A(sreg[67]), .B(n4658), .Z(n4659) );
  XOR U4747 ( .A(n4665), .B(n4677), .Z(n4660) );
  XNOR U4748 ( .A(n4664), .B(n4658), .Z(n4677) );
  XNOR U4749 ( .A(n4678), .B(n4679), .Z(n4658) );
  NOR U4750 ( .A(n4680), .B(n4681), .Z(n4678) );
  NAND U4751 ( .A(a[3]), .B(b[0]), .Z(n4664) );
  XNOR U4752 ( .A(n4670), .B(n4671), .Z(n4665) );
  XOR U4753 ( .A(n4668), .B(n4682), .Z(n4671) );
  NAND U4754 ( .A(b[1]), .B(a[2]), .Z(n4682) );
  XNOR U4755 ( .A(n4675), .B(n4683), .Z(n4670) );
  XOR U4756 ( .A(n4668), .B(n4676), .Z(n4683) );
  XOR U4757 ( .A(n4684), .B(n4674), .Z(n4676) );
  AND U4758 ( .A(b[2]), .B(a[1]), .Z(n4684) );
  NANDN U4759 ( .A(n4685), .B(n4686), .Z(n4668) );
  XNOR U4760 ( .A(n4687), .B(n4674), .Z(n4675) );
  ANDN U4761 ( .B(n4688), .A(n4689), .Z(n4674) );
  NANDN U4762 ( .A(n4690), .B(n4691), .Z(n4688) );
  AND U4763 ( .A(b[3]), .B(a[0]), .Z(n4687) );
  XOR U4764 ( .A(n4681), .B(n4680), .Z(c[50]) );
  XNOR U4765 ( .A(sreg[66]), .B(n4679), .Z(n4680) );
  XOR U4766 ( .A(n4686), .B(n4692), .Z(n4681) );
  XNOR U4767 ( .A(n4693), .B(n4694), .Z(n4679) );
  NAND U4768 ( .A(n4695), .B(n4696), .Z(n4694) );
  NAND U4769 ( .A(a[2]), .B(b[0]), .Z(n4685) );
  XNOR U4770 ( .A(n4690), .B(n4691), .Z(n4686) );
  XOR U4771 ( .A(n4697), .B(n4689), .Z(n4691) );
  AND U4772 ( .A(b[2]), .B(a[0]), .Z(n4697) );
  NAND U4773 ( .A(n4698), .B(a[1]), .Z(n4690) );
  ANDN U4774 ( .B(b[1]), .A(n4689), .Z(n4698) );
  NOR U4775 ( .A(n4699), .B(n4700), .Z(n4689) );
  XOR U4776 ( .A(n4695), .B(n4696), .Z(c[49]) );
  XOR U4777 ( .A(sreg[65]), .B(n4693), .Z(n4696) );
  XNOR U4778 ( .A(n4693), .B(n4701), .Z(n4695) );
  XNOR U4779 ( .A(n4700), .B(n4699), .Z(n4701) );
  NAND U4780 ( .A(b[0]), .B(a[1]), .Z(n4699) );
  NAND U4781 ( .A(a[0]), .B(b[1]), .Z(n4700) );
  ANDN U4782 ( .B(sreg[64]), .A(n4702), .Z(n4693) );
  XNOR U4783 ( .A(sreg[64]), .B(n4702), .Z(c[48]) );
  NAND U4784 ( .A(a[0]), .B(b[0]), .Z(n4702) );
endmodule

