
module compare_N16384_CC32 ( clk, rst, x, y, g, e );
  input [511:0] x;
  input [511:0] y;
  input clk, rst;
  output g, e;
  wire   ebreg, n4, n5, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611;

  DFF ebreg_reg ( .D(n5), .CLK(clk), .RST(rst), .Q(ebreg) );
  DFF greg_reg ( .D(n4), .CLK(clk), .RST(rst), .Q(g) );
  NANDN U10 ( .A(n2158), .B(n2177), .Z(n8) );
  NAND U11 ( .A(n2178), .B(n8), .Z(n9) );
  ANDN U12 ( .B(n9), .A(n2179), .Z(n10) );
  NANDN U13 ( .A(n10), .B(n2180), .Z(n11) );
  NANDN U14 ( .A(n2157), .B(n11), .Z(n12) );
  NAND U15 ( .A(n2181), .B(n12), .Z(n13) );
  NANDN U16 ( .A(n2156), .B(n13), .Z(n14) );
  NAND U17 ( .A(n2182), .B(n14), .Z(n15) );
  ANDN U18 ( .B(n15), .A(n2183), .Z(n16) );
  NANDN U19 ( .A(n16), .B(n2184), .Z(n17) );
  NANDN U20 ( .A(n2155), .B(n17), .Z(n18) );
  NAND U21 ( .A(n2185), .B(n18), .Z(n19) );
  NANDN U22 ( .A(n2154), .B(n19), .Z(n2186) );
  NANDN U23 ( .A(n2145), .B(n2210), .Z(n20) );
  NAND U24 ( .A(n2211), .B(n20), .Z(n21) );
  NANDN U25 ( .A(n2212), .B(n21), .Z(n22) );
  AND U26 ( .A(n2144), .B(n2143), .Z(n23) );
  NAND U27 ( .A(n22), .B(n23), .Z(n24) );
  NANDN U28 ( .A(n2213), .B(n24), .Z(n25) );
  NAND U29 ( .A(n2214), .B(n25), .Z(n26) );
  NANDN U30 ( .A(n2142), .B(n26), .Z(n27) );
  AND U31 ( .A(n2215), .B(n27), .Z(n28) );
  OR U32 ( .A(n2141), .B(n28), .Z(n29) );
  NAND U33 ( .A(n2216), .B(n29), .Z(n30) );
  NAND U34 ( .A(n2217), .B(n30), .Z(n31) );
  AND U35 ( .A(n2140), .B(n2139), .Z(n32) );
  NAND U36 ( .A(n31), .B(n32), .Z(n33) );
  NAND U37 ( .A(n2218), .B(n33), .Z(n2219) );
  NAND U38 ( .A(n2242), .B(n2241), .Z(n34) );
  NANDN U39 ( .A(n2243), .B(n34), .Z(n35) );
  AND U40 ( .A(n2244), .B(n35), .Z(n36) );
  OR U41 ( .A(n2130), .B(n36), .Z(n37) );
  NAND U42 ( .A(n2245), .B(n37), .Z(n38) );
  NANDN U43 ( .A(n2129), .B(n38), .Z(n39) );
  NAND U44 ( .A(n2246), .B(n39), .Z(n40) );
  NANDN U45 ( .A(n2247), .B(n40), .Z(n41) );
  AND U46 ( .A(n2248), .B(n41), .Z(n42) );
  NANDN U47 ( .A(n42), .B(n2249), .Z(n43) );
  AND U48 ( .A(n2250), .B(n43), .Z(n44) );
  OR U49 ( .A(n2128), .B(n44), .Z(n45) );
  NAND U50 ( .A(n2251), .B(n45), .Z(n46) );
  NANDN U51 ( .A(n2252), .B(n46), .Z(n2253) );
  NAND U52 ( .A(n2276), .B(n2275), .Z(n47) );
  NAND U53 ( .A(n2277), .B(n47), .Z(n48) );
  NANDN U54 ( .A(n2119), .B(n48), .Z(n49) );
  NAND U55 ( .A(n2278), .B(n49), .Z(n50) );
  NANDN U56 ( .A(n2279), .B(n50), .Z(n51) );
  AND U57 ( .A(n2280), .B(n51), .Z(n52) );
  NANDN U58 ( .A(n52), .B(n2281), .Z(n53) );
  NAND U59 ( .A(n2282), .B(n53), .Z(n54) );
  NANDN U60 ( .A(n2118), .B(n54), .Z(n55) );
  NAND U61 ( .A(n2283), .B(n55), .Z(n56) );
  NANDN U62 ( .A(n2284), .B(n56), .Z(n57) );
  AND U63 ( .A(n2285), .B(n57), .Z(n58) );
  OR U64 ( .A(n2117), .B(n58), .Z(n59) );
  NAND U65 ( .A(n2286), .B(n59), .Z(n60) );
  NAND U66 ( .A(n2287), .B(n60), .Z(n2288) );
  NAND U67 ( .A(n2314), .B(n2315), .Z(n61) );
  NAND U68 ( .A(n2317), .B(n61), .Z(n62) );
  AND U69 ( .A(n2318), .B(n62), .Z(n63) );
  OR U70 ( .A(n2109), .B(n63), .Z(n64) );
  NAND U71 ( .A(n2319), .B(n64), .Z(n65) );
  NANDN U72 ( .A(n2108), .B(n65), .Z(n66) );
  NAND U73 ( .A(n2320), .B(n66), .Z(n67) );
  NANDN U74 ( .A(n2321), .B(n67), .Z(n68) );
  AND U75 ( .A(n2322), .B(n68), .Z(n69) );
  AND U76 ( .A(n2324), .B(n2325), .Z(n70) );
  NANDN U77 ( .A(n69), .B(n2323), .Z(n71) );
  AND U78 ( .A(n70), .B(n71), .Z(n72) );
  OR U79 ( .A(n2107), .B(n72), .Z(n73) );
  NAND U80 ( .A(n2326), .B(n73), .Z(n74) );
  NANDN U81 ( .A(n2106), .B(n74), .Z(n2327) );
  NANDN U82 ( .A(n2098), .B(n2352), .Z(n75) );
  NAND U83 ( .A(n2353), .B(n75), .Z(n76) );
  NANDN U84 ( .A(n2097), .B(n76), .Z(n77) );
  NAND U85 ( .A(n2354), .B(n77), .Z(n78) );
  NAND U86 ( .A(n2355), .B(n78), .Z(n79) );
  AND U87 ( .A(n2356), .B(n79), .Z(n80) );
  NANDN U88 ( .A(n80), .B(n2357), .Z(n81) );
  NAND U89 ( .A(n2358), .B(n81), .Z(n82) );
  NANDN U90 ( .A(n2096), .B(n82), .Z(n83) );
  NAND U91 ( .A(n2359), .B(n83), .Z(n84) );
  NANDN U92 ( .A(n2360), .B(n84), .Z(n85) );
  AND U93 ( .A(n2361), .B(n85), .Z(n86) );
  NANDN U94 ( .A(n86), .B(n2362), .Z(n87) );
  NAND U95 ( .A(n2363), .B(n87), .Z(n88) );
  NANDN U96 ( .A(n2095), .B(n88), .Z(n2364) );
  NAND U97 ( .A(n2393), .B(n2392), .Z(n89) );
  NAND U98 ( .A(n2394), .B(n89), .Z(n90) );
  NAND U99 ( .A(n2395), .B(n90), .Z(n91) );
  NAND U100 ( .A(n2396), .B(n91), .Z(n92) );
  NAND U101 ( .A(n2397), .B(n92), .Z(n93) );
  AND U102 ( .A(n2398), .B(n93), .Z(n94) );
  OR U103 ( .A(n2088), .B(n94), .Z(n95) );
  NAND U104 ( .A(n2399), .B(n95), .Z(n96) );
  NANDN U105 ( .A(n2087), .B(n96), .Z(n97) );
  NAND U106 ( .A(n2400), .B(n97), .Z(n98) );
  NANDN U107 ( .A(n2401), .B(n98), .Z(n99) );
  AND U108 ( .A(n2402), .B(n99), .Z(n100) );
  OR U109 ( .A(n2086), .B(n100), .Z(n101) );
  NAND U110 ( .A(n2403), .B(n101), .Z(n102) );
  NANDN U111 ( .A(n2085), .B(n102), .Z(n2404) );
  NAND U112 ( .A(n2428), .B(n2427), .Z(n103) );
  AND U113 ( .A(n2429), .B(n103), .Z(n104) );
  NAND U114 ( .A(n104), .B(n2430), .Z(n105) );
  NAND U115 ( .A(n2431), .B(n105), .Z(n106) );
  NAND U116 ( .A(n2432), .B(n106), .Z(n107) );
  ANDN U117 ( .B(n107), .A(n2433), .Z(n108) );
  ANDN U118 ( .B(n2075), .A(n108), .Z(n109) );
  NAND U119 ( .A(n2074), .B(n109), .Z(n110) );
  AND U120 ( .A(n2434), .B(n110), .Z(n111) );
  NANDN U121 ( .A(n111), .B(n2435), .Z(n112) );
  NANDN U122 ( .A(n2073), .B(n112), .Z(n113) );
  NAND U123 ( .A(n2436), .B(n113), .Z(n114) );
  NANDN U124 ( .A(n2072), .B(n114), .Z(n115) );
  NAND U125 ( .A(n2437), .B(n115), .Z(n116) );
  AND U126 ( .A(n2439), .B(n116), .Z(n117) );
  NANDN U127 ( .A(n2438), .B(n117), .Z(n2440) );
  NAND U128 ( .A(n2466), .B(n2465), .Z(n118) );
  NANDN U129 ( .A(n2467), .B(n118), .Z(n119) );
  NAND U130 ( .A(n2468), .B(n119), .Z(n120) );
  NANDN U131 ( .A(n2064), .B(n120), .Z(n121) );
  NAND U132 ( .A(n2469), .B(n121), .Z(n122) );
  ANDN U133 ( .B(n122), .A(n2063), .Z(n123) );
  NANDN U134 ( .A(n123), .B(n2470), .Z(n124) );
  NAND U135 ( .A(n2471), .B(n124), .Z(n125) );
  NAND U136 ( .A(n2472), .B(n125), .Z(n126) );
  NANDN U137 ( .A(n2062), .B(n126), .Z(n127) );
  NAND U138 ( .A(n2473), .B(n127), .Z(n128) );
  ANDN U139 ( .B(n128), .A(n2061), .Z(n129) );
  NANDN U140 ( .A(n129), .B(n2474), .Z(n130) );
  NAND U141 ( .A(n2475), .B(n130), .Z(n131) );
  NAND U142 ( .A(n2476), .B(n131), .Z(n2477) );
  NAND U143 ( .A(n2503), .B(n2504), .Z(n132) );
  NAND U144 ( .A(n2505), .B(n132), .Z(n133) );
  ANDN U145 ( .B(n133), .A(n2052), .Z(n134) );
  NANDN U146 ( .A(n134), .B(n2506), .Z(n135) );
  NANDN U147 ( .A(n2507), .B(n135), .Z(n136) );
  NAND U148 ( .A(n2508), .B(n136), .Z(n137) );
  NANDN U149 ( .A(n2051), .B(n137), .Z(n138) );
  NAND U150 ( .A(n2509), .B(n138), .Z(n139) );
  ANDN U151 ( .B(n139), .A(n2050), .Z(n140) );
  NANDN U152 ( .A(n140), .B(n2510), .Z(n141) );
  ANDN U153 ( .B(n141), .A(n2511), .Z(n142) );
  NANDN U154 ( .A(n142), .B(n2512), .Z(n143) );
  NANDN U155 ( .A(n2049), .B(n143), .Z(n144) );
  NAND U156 ( .A(n2513), .B(n144), .Z(n2514) );
  NANDN U157 ( .A(n2040), .B(n2538), .Z(n145) );
  NAND U158 ( .A(n2539), .B(n145), .Z(n146) );
  NANDN U159 ( .A(n2540), .B(n146), .Z(n147) );
  NAND U160 ( .A(n2541), .B(n147), .Z(n148) );
  NAND U161 ( .A(n2542), .B(n148), .Z(n149) );
  AND U162 ( .A(n2543), .B(n149), .Z(n150) );
  OR U163 ( .A(n2039), .B(n150), .Z(n151) );
  NAND U164 ( .A(n2544), .B(n151), .Z(n152) );
  NANDN U165 ( .A(n2545), .B(n152), .Z(n153) );
  NAND U166 ( .A(n2546), .B(n153), .Z(n154) );
  NANDN U167 ( .A(n2038), .B(n154), .Z(n155) );
  AND U168 ( .A(n2547), .B(n155), .Z(n156) );
  OR U169 ( .A(n2037), .B(n156), .Z(n157) );
  AND U170 ( .A(n2548), .B(n157), .Z(n2551) );
  NANDN U171 ( .A(n2030), .B(n2575), .Z(n158) );
  NAND U172 ( .A(n2576), .B(n158), .Z(n159) );
  NAND U173 ( .A(n2577), .B(n159), .Z(n160) );
  NAND U174 ( .A(n2578), .B(n160), .Z(n161) );
  NAND U175 ( .A(n2579), .B(n161), .Z(n162) );
  AND U176 ( .A(n2580), .B(n162), .Z(n163) );
  NANDN U177 ( .A(n163), .B(n2581), .Z(n164) );
  NAND U178 ( .A(n2582), .B(n164), .Z(n165) );
  NANDN U179 ( .A(n2029), .B(n165), .Z(n166) );
  NAND U180 ( .A(n2583), .B(n166), .Z(n167) );
  NANDN U181 ( .A(n2584), .B(n167), .Z(n168) );
  AND U182 ( .A(n2585), .B(n168), .Z(n169) );
  OR U183 ( .A(n2028), .B(n169), .Z(n170) );
  NAND U184 ( .A(n2586), .B(n170), .Z(n171) );
  NANDN U185 ( .A(n2027), .B(n171), .Z(n2587) );
  NAND U186 ( .A(n2162), .B(n2163), .Z(n2164) );
  NAND U187 ( .A(n2186), .B(n2187), .Z(n172) );
  NAND U188 ( .A(n2189), .B(n172), .Z(n173) );
  AND U189 ( .A(n2190), .B(n173), .Z(n174) );
  OR U190 ( .A(n2153), .B(n174), .Z(n175) );
  NAND U191 ( .A(n2191), .B(n175), .Z(n176) );
  NANDN U192 ( .A(n2152), .B(n176), .Z(n177) );
  NAND U193 ( .A(n2192), .B(n177), .Z(n178) );
  NANDN U194 ( .A(n2193), .B(n178), .Z(n179) );
  AND U195 ( .A(n2194), .B(n179), .Z(n180) );
  OR U196 ( .A(n2151), .B(n180), .Z(n181) );
  AND U197 ( .A(n2195), .B(n181), .Z(n182) );
  OR U198 ( .A(n2150), .B(n182), .Z(n183) );
  NAND U199 ( .A(n2196), .B(n183), .Z(n184) );
  NANDN U200 ( .A(n2197), .B(n184), .Z(n2198) );
  NAND U201 ( .A(n2219), .B(n2220), .Z(n185) );
  NANDN U202 ( .A(n2138), .B(n185), .Z(n186) );
  AND U203 ( .A(n2221), .B(n186), .Z(n187) );
  NANDN U204 ( .A(n187), .B(n2222), .Z(n188) );
  NAND U205 ( .A(n2223), .B(n188), .Z(n189) );
  NANDN U206 ( .A(n2224), .B(n189), .Z(n190) );
  NAND U207 ( .A(n2225), .B(n190), .Z(n191) );
  NANDN U208 ( .A(n2137), .B(n191), .Z(n192) );
  AND U209 ( .A(n2226), .B(n192), .Z(n193) );
  OR U210 ( .A(n2136), .B(n193), .Z(n194) );
  AND U211 ( .A(n2227), .B(n194), .Z(n195) );
  OR U212 ( .A(n195), .B(n2228), .Z(n196) );
  NAND U213 ( .A(n2229), .B(n196), .Z(n197) );
  NANDN U214 ( .A(n2135), .B(n197), .Z(n2230) );
  NOR U215 ( .A(n2127), .B(n2255), .Z(n198) );
  NAND U216 ( .A(n2253), .B(n2254), .Z(n199) );
  AND U217 ( .A(n198), .B(n199), .Z(n200) );
  NANDN U218 ( .A(n200), .B(n2256), .Z(n201) );
  NANDN U219 ( .A(n2126), .B(n201), .Z(n202) );
  NAND U220 ( .A(n2257), .B(n202), .Z(n203) );
  NANDN U221 ( .A(n2125), .B(n203), .Z(n204) );
  NAND U222 ( .A(n2258), .B(n204), .Z(n205) );
  ANDN U223 ( .B(n205), .A(n2259), .Z(n206) );
  NANDN U224 ( .A(n206), .B(n2260), .Z(n207) );
  NANDN U225 ( .A(n2124), .B(n207), .Z(n208) );
  NAND U226 ( .A(n2261), .B(n208), .Z(n209) );
  NANDN U227 ( .A(n2123), .B(n209), .Z(n2262) );
  NAND U228 ( .A(n2288), .B(n2289), .Z(n210) );
  NAND U229 ( .A(n2291), .B(n210), .Z(n211) );
  NAND U230 ( .A(n2292), .B(n211), .Z(n212) );
  NAND U231 ( .A(n2293), .B(n212), .Z(n213) );
  NAND U232 ( .A(n2294), .B(n213), .Z(n214) );
  ANDN U233 ( .B(n214), .A(n2116), .Z(n215) );
  NANDN U234 ( .A(n215), .B(n2295), .Z(n216) );
  NANDN U235 ( .A(n2296), .B(n216), .Z(n217) );
  NAND U236 ( .A(n2297), .B(n217), .Z(n218) );
  NANDN U237 ( .A(n2115), .B(n218), .Z(n219) );
  NAND U238 ( .A(n2298), .B(n219), .Z(n220) );
  ANDN U239 ( .B(n220), .A(n2114), .Z(n221) );
  NANDN U240 ( .A(n221), .B(n2299), .Z(n222) );
  NAND U241 ( .A(n2300), .B(n222), .Z(n223) );
  NAND U242 ( .A(n2301), .B(n223), .Z(n224) );
  NAND U243 ( .A(n2302), .B(n224), .Z(n2303) );
  NAND U244 ( .A(n2327), .B(n2328), .Z(n225) );
  NAND U245 ( .A(n2329), .B(n225), .Z(n226) );
  AND U246 ( .A(n2330), .B(n226), .Z(n227) );
  OR U247 ( .A(n2105), .B(n227), .Z(n228) );
  NAND U248 ( .A(n2331), .B(n228), .Z(n229) );
  NANDN U249 ( .A(n2104), .B(n229), .Z(n230) );
  NAND U250 ( .A(n2332), .B(n230), .Z(n231) );
  AND U251 ( .A(n2334), .B(n231), .Z(n232) );
  NANDN U252 ( .A(n2333), .B(n232), .Z(n233) );
  NAND U253 ( .A(n2335), .B(n233), .Z(n234) );
  NAND U254 ( .A(n2336), .B(n234), .Z(n235) );
  AND U255 ( .A(n2337), .B(n235), .Z(n236) );
  OR U256 ( .A(n2103), .B(n236), .Z(n237) );
  NAND U257 ( .A(n2338), .B(n237), .Z(n238) );
  NANDN U258 ( .A(n2102), .B(n238), .Z(n2339) );
  NAND U259 ( .A(n2364), .B(n2365), .Z(n239) );
  NAND U260 ( .A(n2367), .B(n239), .Z(n240) );
  AND U261 ( .A(n2368), .B(n240), .Z(n241) );
  OR U262 ( .A(n2094), .B(n241), .Z(n242) );
  NAND U263 ( .A(n2369), .B(n242), .Z(n243) );
  NANDN U264 ( .A(n2093), .B(n243), .Z(n244) );
  AND U265 ( .A(n2370), .B(n2371), .Z(n245) );
  NAND U266 ( .A(n244), .B(n245), .Z(n246) );
  NANDN U267 ( .A(n2092), .B(n246), .Z(n247) );
  AND U268 ( .A(n2372), .B(n2373), .Z(n248) );
  NAND U269 ( .A(n247), .B(n248), .Z(n249) );
  NANDN U270 ( .A(n2091), .B(n249), .Z(n250) );
  NAND U271 ( .A(n2374), .B(n250), .Z(n251) );
  AND U272 ( .A(n2376), .B(n251), .Z(n252) );
  NANDN U273 ( .A(n2375), .B(n252), .Z(n2377) );
  NAND U274 ( .A(n2082), .B(n2083), .Z(n253) );
  NAND U275 ( .A(n2405), .B(n2404), .Z(n254) );
  NANDN U276 ( .A(n2406), .B(n254), .Z(n255) );
  NAND U277 ( .A(n2407), .B(n255), .Z(n256) );
  NANDN U278 ( .A(n2084), .B(n256), .Z(n257) );
  NAND U279 ( .A(n2408), .B(n257), .Z(n258) );
  AND U280 ( .A(n2409), .B(n258), .Z(n259) );
  NANDN U281 ( .A(n259), .B(n2410), .Z(n260) );
  ANDN U282 ( .B(n260), .A(n2411), .Z(n261) );
  ANDN U283 ( .B(n2413), .A(n2412), .Z(n262) );
  OR U284 ( .A(n253), .B(n261), .Z(n263) );
  AND U285 ( .A(n262), .B(n263), .Z(n264) );
  NANDN U286 ( .A(n264), .B(n2414), .Z(n265) );
  NANDN U287 ( .A(n2415), .B(n265), .Z(n266) );
  NAND U288 ( .A(n2416), .B(n266), .Z(n2417) );
  NAND U289 ( .A(n2440), .B(n2441), .Z(n267) );
  NAND U290 ( .A(n2442), .B(n267), .Z(n268) );
  NAND U291 ( .A(n2443), .B(n268), .Z(n269) );
  NAND U292 ( .A(n2444), .B(n269), .Z(n270) );
  NAND U293 ( .A(n2445), .B(n270), .Z(n271) );
  ANDN U294 ( .B(n271), .A(n2071), .Z(n272) );
  NANDN U295 ( .A(n272), .B(n2446), .Z(n273) );
  NANDN U296 ( .A(n2447), .B(n273), .Z(n274) );
  NAND U297 ( .A(n2448), .B(n274), .Z(n275) );
  NANDN U298 ( .A(n2070), .B(n275), .Z(n276) );
  NAND U299 ( .A(n2449), .B(n276), .Z(n277) );
  ANDN U300 ( .B(n277), .A(n2069), .Z(n278) );
  NANDN U301 ( .A(n278), .B(n2450), .Z(n279) );
  NAND U302 ( .A(n2451), .B(n279), .Z(n280) );
  NAND U303 ( .A(n2452), .B(n280), .Z(n281) );
  NAND U304 ( .A(n2453), .B(n281), .Z(n2454) );
  NAND U305 ( .A(n2478), .B(n2477), .Z(n282) );
  NAND U306 ( .A(n2479), .B(n282), .Z(n283) );
  ANDN U307 ( .B(n283), .A(n2059), .Z(n284) );
  NANDN U308 ( .A(n284), .B(n2480), .Z(n285) );
  NAND U309 ( .A(n2481), .B(n285), .Z(n286) );
  NAND U310 ( .A(n2482), .B(n286), .Z(n287) );
  NANDN U311 ( .A(n2058), .B(n287), .Z(n288) );
  NAND U312 ( .A(n2483), .B(n288), .Z(n289) );
  ANDN U313 ( .B(n289), .A(n2057), .Z(n290) );
  ANDN U314 ( .B(n2484), .A(n290), .Z(n291) );
  NAND U315 ( .A(n2485), .B(n291), .Z(n292) );
  ANDN U316 ( .B(n292), .A(n2056), .Z(n293) );
  NANDN U317 ( .A(n293), .B(n2486), .Z(n294) );
  NANDN U318 ( .A(n2487), .B(n294), .Z(n295) );
  NAND U319 ( .A(n2488), .B(n295), .Z(n2489) );
  NANDN U320 ( .A(n2048), .B(n2514), .Z(n296) );
  NAND U321 ( .A(n2515), .B(n296), .Z(n297) );
  NAND U322 ( .A(n2516), .B(n297), .Z(n298) );
  NAND U323 ( .A(n2517), .B(n298), .Z(n299) );
  NANDN U324 ( .A(n2047), .B(n299), .Z(n300) );
  AND U325 ( .A(n2518), .B(n300), .Z(n301) );
  OR U326 ( .A(n2046), .B(n301), .Z(n302) );
  AND U327 ( .A(n2519), .B(n302), .Z(n303) );
  NOR U328 ( .A(n2520), .B(n303), .Z(n304) );
  NAND U329 ( .A(n2521), .B(n304), .Z(n305) );
  AND U330 ( .A(n2522), .B(n305), .Z(n306) );
  NANDN U331 ( .A(n306), .B(n2523), .Z(n307) );
  NAND U332 ( .A(n2524), .B(n307), .Z(n308) );
  NANDN U333 ( .A(n2045), .B(n308), .Z(n309) );
  NAND U334 ( .A(n2525), .B(n309), .Z(n2526) );
  NANDN U335 ( .A(n2551), .B(n2550), .Z(n310) );
  NAND U336 ( .A(n2552), .B(n310), .Z(n311) );
  NAND U337 ( .A(n2553), .B(n311), .Z(n312) );
  NAND U338 ( .A(n2554), .B(n312), .Z(n313) );
  NANDN U339 ( .A(n2036), .B(n313), .Z(n314) );
  AND U340 ( .A(n2555), .B(n314), .Z(n315) );
  OR U341 ( .A(n315), .B(n2556), .Z(n316) );
  NAND U342 ( .A(n2557), .B(n316), .Z(n317) );
  NANDN U343 ( .A(n2035), .B(n317), .Z(n318) );
  NAND U344 ( .A(n2558), .B(n318), .Z(n319) );
  NANDN U345 ( .A(n2034), .B(n319), .Z(n320) );
  AND U346 ( .A(n2559), .B(n320), .Z(n321) );
  OR U347 ( .A(n321), .B(n2560), .Z(n322) );
  NAND U348 ( .A(n2561), .B(n322), .Z(n323) );
  NAND U349 ( .A(n2562), .B(n323), .Z(n2563) );
  NAND U350 ( .A(n2587), .B(n2588), .Z(n324) );
  NAND U351 ( .A(n2590), .B(n324), .Z(n325) );
  NAND U352 ( .A(n2591), .B(n325), .Z(n326) );
  NAND U353 ( .A(n2592), .B(n326), .Z(n327) );
  NAND U354 ( .A(n2593), .B(n327), .Z(n328) );
  ANDN U355 ( .B(n328), .A(n2026), .Z(n329) );
  NANDN U356 ( .A(n329), .B(n2594), .Z(n330) );
  NANDN U357 ( .A(n2595), .B(n330), .Z(n331) );
  NAND U358 ( .A(n2596), .B(n331), .Z(n332) );
  NANDN U359 ( .A(n2025), .B(n332), .Z(n333) );
  NAND U360 ( .A(n2597), .B(n333), .Z(n334) );
  ANDN U361 ( .B(n334), .A(n2024), .Z(n335) );
  NANDN U362 ( .A(n335), .B(n2598), .Z(n336) );
  NANDN U363 ( .A(n2599), .B(n336), .Z(n337) );
  NAND U364 ( .A(n2600), .B(n337), .Z(n2601) );
  AND U365 ( .A(n2165), .B(n2166), .Z(n338) );
  NANDN U366 ( .A(n2161), .B(n2164), .Z(n339) );
  NAND U367 ( .A(n338), .B(n339), .Z(n340) );
  NAND U368 ( .A(n2167), .B(n340), .Z(n341) );
  NAND U369 ( .A(n2168), .B(n341), .Z(n342) );
  ANDN U370 ( .B(n342), .A(n2169), .Z(n343) );
  NANDN U371 ( .A(n343), .B(n2170), .Z(n344) );
  NANDN U372 ( .A(n2160), .B(n344), .Z(n345) );
  NAND U373 ( .A(n2171), .B(n345), .Z(n346) );
  NANDN U374 ( .A(n2159), .B(n346), .Z(n347) );
  NAND U375 ( .A(n2172), .B(n347), .Z(n348) );
  ANDN U376 ( .B(n348), .A(n2173), .Z(n349) );
  NANDN U377 ( .A(n349), .B(n2174), .Z(n350) );
  NAND U378 ( .A(n2175), .B(n350), .Z(n351) );
  NAND U379 ( .A(n2176), .B(n351), .Z(n2177) );
  NAND U380 ( .A(n2199), .B(n2198), .Z(n352) );
  NAND U381 ( .A(n2200), .B(n352), .Z(n353) );
  NAND U382 ( .A(n2201), .B(n353), .Z(n354) );
  NANDN U383 ( .A(n2149), .B(n354), .Z(n355) );
  NAND U384 ( .A(n2202), .B(n355), .Z(n356) );
  ANDN U385 ( .B(n356), .A(n2203), .Z(n357) );
  NANDN U386 ( .A(n357), .B(n2204), .Z(n358) );
  NANDN U387 ( .A(n2148), .B(n358), .Z(n359) );
  NAND U388 ( .A(n2205), .B(n359), .Z(n360) );
  NANDN U389 ( .A(n2147), .B(n360), .Z(n361) );
  NAND U390 ( .A(n2206), .B(n361), .Z(n362) );
  AND U391 ( .A(n2207), .B(n362), .Z(n363) );
  NANDN U392 ( .A(n363), .B(n2208), .Z(n364) );
  NANDN U393 ( .A(n2146), .B(n364), .Z(n365) );
  NAND U394 ( .A(n2209), .B(n365), .Z(n2210) );
  NAND U395 ( .A(n2231), .B(n2230), .Z(n366) );
  NAND U396 ( .A(n2232), .B(n366), .Z(n367) );
  AND U397 ( .A(n2233), .B(n367), .Z(n368) );
  OR U398 ( .A(n368), .B(n2234), .Z(n369) );
  NAND U399 ( .A(n2235), .B(n369), .Z(n370) );
  NANDN U400 ( .A(n2134), .B(n370), .Z(n371) );
  NAND U401 ( .A(n2236), .B(n371), .Z(n372) );
  NANDN U402 ( .A(n2133), .B(n372), .Z(n373) );
  AND U403 ( .A(n2237), .B(n373), .Z(n374) );
  OR U404 ( .A(n374), .B(n2238), .Z(n375) );
  AND U405 ( .A(n2239), .B(n375), .Z(n376) );
  OR U406 ( .A(n2132), .B(n376), .Z(n377) );
  NAND U407 ( .A(n2240), .B(n377), .Z(n378) );
  NANDN U408 ( .A(n2131), .B(n378), .Z(n2241) );
  NAND U409 ( .A(n2263), .B(n2262), .Z(n379) );
  NANDN U410 ( .A(n2264), .B(n379), .Z(n380) );
  NAND U411 ( .A(n2265), .B(n380), .Z(n381) );
  NAND U412 ( .A(n2266), .B(n381), .Z(n382) );
  NAND U413 ( .A(n2267), .B(n382), .Z(n383) );
  ANDN U414 ( .B(n383), .A(n2122), .Z(n384) );
  NANDN U415 ( .A(n384), .B(n2268), .Z(n385) );
  NAND U416 ( .A(n2269), .B(n385), .Z(n386) );
  NAND U417 ( .A(n2270), .B(n386), .Z(n387) );
  NANDN U418 ( .A(n2121), .B(n387), .Z(n388) );
  NAND U419 ( .A(n2271), .B(n388), .Z(n389) );
  ANDN U420 ( .B(n389), .A(n2120), .Z(n390) );
  NANDN U421 ( .A(n390), .B(n2272), .Z(n391) );
  NANDN U422 ( .A(n2273), .B(n391), .Z(n392) );
  NAND U423 ( .A(n2274), .B(n392), .Z(n2275) );
  NAND U424 ( .A(n2303), .B(n2304), .Z(n393) );
  NANDN U425 ( .A(n2113), .B(n393), .Z(n394) );
  AND U426 ( .A(n2305), .B(n394), .Z(n395) );
  OR U427 ( .A(n395), .B(n2306), .Z(n396) );
  NAND U428 ( .A(n2307), .B(n396), .Z(n397) );
  NANDN U429 ( .A(n2112), .B(n397), .Z(n398) );
  NAND U430 ( .A(n2308), .B(n398), .Z(n399) );
  NAND U431 ( .A(n2309), .B(n399), .Z(n400) );
  AND U432 ( .A(n2310), .B(n400), .Z(n401) );
  OR U433 ( .A(n401), .B(n2311), .Z(n402) );
  AND U434 ( .A(n2312), .B(n402), .Z(n403) );
  OR U435 ( .A(n2111), .B(n403), .Z(n404) );
  NAND U436 ( .A(n2313), .B(n404), .Z(n405) );
  NANDN U437 ( .A(n2110), .B(n405), .Z(n2314) );
  NAND U438 ( .A(n2340), .B(n2339), .Z(n406) );
  NANDN U439 ( .A(n2341), .B(n406), .Z(n407) );
  NAND U440 ( .A(n2342), .B(n407), .Z(n408) );
  NANDN U441 ( .A(n2101), .B(n408), .Z(n409) );
  NAND U442 ( .A(n2343), .B(n409), .Z(n410) );
  ANDN U443 ( .B(n410), .A(n2100), .Z(n411) );
  NANDN U444 ( .A(n411), .B(n2344), .Z(n412) );
  NAND U445 ( .A(n2345), .B(n412), .Z(n413) );
  NAND U446 ( .A(n2346), .B(n413), .Z(n414) );
  NAND U447 ( .A(n2347), .B(n414), .Z(n415) );
  NAND U448 ( .A(n2348), .B(n415), .Z(n416) );
  ANDN U449 ( .B(n416), .A(n2099), .Z(n417) );
  NANDN U450 ( .A(n417), .B(n2349), .Z(n418) );
  NANDN U451 ( .A(n2350), .B(n418), .Z(n419) );
  NAND U452 ( .A(n2351), .B(n419), .Z(n2352) );
  ANDN U453 ( .B(n2381), .A(n2380), .Z(n420) );
  NAND U454 ( .A(n2377), .B(n2378), .Z(n421) );
  AND U455 ( .A(n420), .B(n421), .Z(n422) );
  NANDN U456 ( .A(x[255]), .B(y[255]), .Z(n423) );
  NANDN U457 ( .A(n422), .B(n423), .Z(n424) );
  ANDN U458 ( .B(n424), .A(n2382), .Z(n425) );
  NANDN U459 ( .A(n425), .B(n2383), .Z(n426) );
  NAND U460 ( .A(n2384), .B(n426), .Z(n427) );
  NAND U461 ( .A(n2385), .B(n427), .Z(n428) );
  NAND U462 ( .A(n2386), .B(n428), .Z(n429) );
  NAND U463 ( .A(n2387), .B(n429), .Z(n430) );
  ANDN U464 ( .B(n430), .A(n2388), .Z(n431) );
  NANDN U465 ( .A(n431), .B(n2389), .Z(n432) );
  NANDN U466 ( .A(n2090), .B(n432), .Z(n433) );
  NAND U467 ( .A(n2390), .B(n433), .Z(n434) );
  ANDN U468 ( .B(n434), .A(n2391), .Z(n2392) );
  ANDN U469 ( .B(n2417), .A(n2081), .Z(n435) );
  NAND U470 ( .A(n2418), .B(n435), .Z(n436) );
  NAND U471 ( .A(n2419), .B(n436), .Z(n437) );
  AND U472 ( .A(n2421), .B(n2420), .Z(n438) );
  NANDN U473 ( .A(n2080), .B(n437), .Z(n439) );
  NAND U474 ( .A(n438), .B(n439), .Z(n440) );
  NANDN U475 ( .A(n2079), .B(n440), .Z(n441) );
  NAND U476 ( .A(n2422), .B(n441), .Z(n442) );
  ANDN U477 ( .B(n442), .A(n2078), .Z(n443) );
  NANDN U478 ( .A(n443), .B(n2423), .Z(n444) );
  ANDN U479 ( .B(n444), .A(n2424), .Z(n445) );
  NANDN U480 ( .A(n445), .B(n2425), .Z(n446) );
  NANDN U481 ( .A(n2077), .B(n446), .Z(n447) );
  NAND U482 ( .A(n2426), .B(n447), .Z(n2427) );
  NAND U483 ( .A(n2454), .B(n2455), .Z(n448) );
  NANDN U484 ( .A(n2068), .B(n448), .Z(n449) );
  AND U485 ( .A(n2456), .B(n449), .Z(n450) );
  OR U486 ( .A(n450), .B(n2457), .Z(n451) );
  NAND U487 ( .A(n2458), .B(n451), .Z(n452) );
  NAND U488 ( .A(n2459), .B(n452), .Z(n453) );
  NAND U489 ( .A(n2460), .B(n453), .Z(n454) );
  NANDN U490 ( .A(n2067), .B(n454), .Z(n455) );
  AND U491 ( .A(n2461), .B(n455), .Z(n456) );
  OR U492 ( .A(n456), .B(n2462), .Z(n457) );
  AND U493 ( .A(n2463), .B(n457), .Z(n458) );
  OR U494 ( .A(n2066), .B(n458), .Z(n459) );
  NAND U495 ( .A(n2464), .B(n459), .Z(n460) );
  NANDN U496 ( .A(n2065), .B(n460), .Z(n2465) );
  NAND U497 ( .A(n2490), .B(n2489), .Z(n461) );
  NAND U498 ( .A(n2491), .B(n461), .Z(n462) );
  ANDN U499 ( .B(n462), .A(n2054), .Z(n463) );
  NANDN U500 ( .A(n463), .B(n2492), .Z(n464) );
  NANDN U501 ( .A(n2493), .B(n464), .Z(n465) );
  NAND U502 ( .A(n2494), .B(n465), .Z(n466) );
  NAND U503 ( .A(n2495), .B(n466), .Z(n467) );
  NAND U504 ( .A(n2496), .B(n467), .Z(n468) );
  ANDN U505 ( .B(n468), .A(n2497), .Z(n469) );
  NANDN U506 ( .A(n2053), .B(n469), .Z(n470) );
  NAND U507 ( .A(n2498), .B(n470), .Z(n471) );
  AND U508 ( .A(n2499), .B(n471), .Z(n472) );
  NANDN U509 ( .A(n472), .B(n2500), .Z(n473) );
  NANDN U510 ( .A(n2501), .B(n473), .Z(n474) );
  NAND U511 ( .A(n2502), .B(n474), .Z(n2503) );
  NANDN U512 ( .A(n2044), .B(n2526), .Z(n475) );
  NAND U513 ( .A(n2527), .B(n475), .Z(n476) );
  ANDN U514 ( .B(n476), .A(n2528), .Z(n477) );
  ANDN U515 ( .B(n2043), .A(n477), .Z(n478) );
  NAND U516 ( .A(n2042), .B(n478), .Z(n479) );
  ANDN U517 ( .B(n479), .A(n2529), .Z(n480) );
  NANDN U518 ( .A(n480), .B(n2530), .Z(n481) );
  NAND U519 ( .A(n2531), .B(n481), .Z(n482) );
  NAND U520 ( .A(n2532), .B(n482), .Z(n483) );
  NANDN U521 ( .A(n2041), .B(n483), .Z(n484) );
  NAND U522 ( .A(n2533), .B(n484), .Z(n485) );
  ANDN U523 ( .B(n485), .A(n2534), .Z(n486) );
  NANDN U524 ( .A(n486), .B(n2535), .Z(n487) );
  NAND U525 ( .A(n2536), .B(n487), .Z(n488) );
  NAND U526 ( .A(n2537), .B(n488), .Z(n2538) );
  NAND U527 ( .A(n2563), .B(n2564), .Z(n489) );
  NANDN U528 ( .A(n2033), .B(n489), .Z(n490) );
  AND U529 ( .A(n2565), .B(n490), .Z(n491) );
  OR U530 ( .A(n491), .B(n2566), .Z(n492) );
  NAND U531 ( .A(n2567), .B(n492), .Z(n493) );
  ANDN U532 ( .B(n493), .A(n2032), .Z(n494) );
  NANDN U533 ( .A(n2568), .B(n494), .Z(n495) );
  NAND U534 ( .A(n2569), .B(n495), .Z(n496) );
  AND U535 ( .A(n2570), .B(n496), .Z(n497) );
  NANDN U536 ( .A(n497), .B(n2571), .Z(n498) );
  ANDN U537 ( .B(n498), .A(n2031), .Z(n499) );
  NANDN U538 ( .A(n499), .B(n2572), .Z(n500) );
  NANDN U539 ( .A(n2573), .B(n500), .Z(n501) );
  NAND U540 ( .A(n2574), .B(n501), .Z(n2575) );
  ANDN U541 ( .B(n2611), .A(ebreg), .Z(n502) );
  NAND U542 ( .A(n2601), .B(n2602), .Z(n503) );
  NAND U543 ( .A(n2603), .B(n503), .Z(n504) );
  NANDN U544 ( .A(n2022), .B(n504), .Z(n505) );
  NAND U545 ( .A(n2604), .B(n505), .Z(n506) );
  NAND U546 ( .A(n2605), .B(n506), .Z(n507) );
  AND U547 ( .A(n2606), .B(n507), .Z(n508) );
  OR U548 ( .A(n508), .B(n2607), .Z(n509) );
  NAND U549 ( .A(n2608), .B(n509), .Z(n510) );
  NANDN U550 ( .A(n2021), .B(n510), .Z(n511) );
  AND U551 ( .A(n2610), .B(n2609), .Z(n512) );
  NAND U552 ( .A(n511), .B(n512), .Z(n513) );
  NANDN U553 ( .A(n2020), .B(n513), .Z(n514) );
  NAND U554 ( .A(n514), .B(n502), .Z(n515) );
  NANDN U555 ( .A(n502), .B(g), .Z(n516) );
  NAND U556 ( .A(n515), .B(n516), .Z(n4) );
  IV U557 ( .A(ebreg), .Z(e) );
  NANDN U558 ( .A(x[215]), .B(y[215]), .Z(n518) );
  NANDN U559 ( .A(x[214]), .B(y[214]), .Z(n517) );
  AND U560 ( .A(n518), .B(n517), .Z(n2342) );
  NANDN U561 ( .A(x[207]), .B(y[207]), .Z(n520) );
  NANDN U562 ( .A(x[206]), .B(y[206]), .Z(n519) );
  AND U563 ( .A(n520), .B(n519), .Z(n2335) );
  AND U564 ( .A(n2342), .B(n2335), .Z(n526) );
  NANDN U565 ( .A(x[213]), .B(y[213]), .Z(n522) );
  NANDN U566 ( .A(x[212]), .B(y[212]), .Z(n521) );
  AND U567 ( .A(n522), .B(n521), .Z(n2340) );
  NANDN U568 ( .A(y[212]), .B(x[212]), .Z(n524) );
  NANDN U569 ( .A(y[211]), .B(x[211]), .Z(n523) );
  NAND U570 ( .A(n524), .B(n523), .Z(n2102) );
  ANDN U571 ( .B(n2340), .A(n2102), .Z(n525) );
  AND U572 ( .A(n526), .B(n525), .Z(n538) );
  NANDN U573 ( .A(x[205]), .B(y[205]), .Z(n528) );
  NANDN U574 ( .A(x[204]), .B(y[204]), .Z(n527) );
  AND U575 ( .A(n528), .B(n527), .Z(n2332) );
  NANDN U576 ( .A(x[197]), .B(y[197]), .Z(n530) );
  NANDN U577 ( .A(x[196]), .B(y[196]), .Z(n529) );
  AND U578 ( .A(n530), .B(n529), .Z(n2326) );
  AND U579 ( .A(n2332), .B(n2326), .Z(n536) );
  NANDN U580 ( .A(x[199]), .B(y[199]), .Z(n532) );
  NANDN U581 ( .A(x[198]), .B(y[198]), .Z(n531) );
  AND U582 ( .A(n532), .B(n531), .Z(n2328) );
  NANDN U583 ( .A(y[204]), .B(x[204]), .Z(n534) );
  NANDN U584 ( .A(y[203]), .B(x[203]), .Z(n533) );
  NAND U585 ( .A(n534), .B(n533), .Z(n2104) );
  ANDN U586 ( .B(n2328), .A(n2104), .Z(n535) );
  AND U587 ( .A(n536), .B(n535), .Z(n537) );
  AND U588 ( .A(n538), .B(n537), .Z(n562) );
  NANDN U589 ( .A(y[222]), .B(x[222]), .Z(n540) );
  NANDN U590 ( .A(y[221]), .B(x[221]), .Z(n539) );
  AND U591 ( .A(n540), .B(n539), .Z(n2347) );
  NANDN U592 ( .A(y[216]), .B(x[216]), .Z(n542) );
  NANDN U593 ( .A(y[215]), .B(x[215]), .Z(n541) );
  NAND U594 ( .A(n542), .B(n541), .Z(n2101) );
  ANDN U595 ( .B(n2347), .A(n2101), .Z(n548) );
  NANDN U596 ( .A(x[219]), .B(y[219]), .Z(n544) );
  NANDN U597 ( .A(x[218]), .B(y[218]), .Z(n543) );
  AND U598 ( .A(n544), .B(n543), .Z(n2344) );
  NANDN U599 ( .A(y[218]), .B(x[218]), .Z(n546) );
  NANDN U600 ( .A(y[217]), .B(x[217]), .Z(n545) );
  NAND U601 ( .A(n546), .B(n545), .Z(n2100) );
  ANDN U602 ( .B(n2344), .A(n2100), .Z(n547) );
  AND U603 ( .A(n548), .B(n547), .Z(n560) );
  NANDN U604 ( .A(x[189]), .B(y[189]), .Z(n550) );
  NANDN U605 ( .A(x[188]), .B(y[188]), .Z(n549) );
  AND U606 ( .A(n550), .B(n549), .Z(n2319) );
  NANDN U607 ( .A(y[196]), .B(x[196]), .Z(n552) );
  NANDN U608 ( .A(y[195]), .B(x[195]), .Z(n551) );
  NAND U609 ( .A(n552), .B(n551), .Z(n2107) );
  ANDN U610 ( .B(n2319), .A(n2107), .Z(n558) );
  NANDN U611 ( .A(y[194]), .B(x[194]), .Z(n554) );
  NANDN U612 ( .A(y[193]), .B(x[193]), .Z(n553) );
  AND U613 ( .A(n554), .B(n553), .Z(n2323) );
  NANDN U614 ( .A(y[190]), .B(x[190]), .Z(n556) );
  NANDN U615 ( .A(y[189]), .B(x[189]), .Z(n555) );
  NAND U616 ( .A(n556), .B(n555), .Z(n2108) );
  ANDN U617 ( .B(n2323), .A(n2108), .Z(n557) );
  AND U618 ( .A(n558), .B(n557), .Z(n559) );
  AND U619 ( .A(n560), .B(n559), .Z(n561) );
  AND U620 ( .A(n562), .B(n561), .Z(n610) );
  NANDN U621 ( .A(x[179]), .B(y[179]), .Z(n564) );
  NANDN U622 ( .A(x[178]), .B(y[178]), .Z(n563) );
  AND U623 ( .A(n564), .B(n563), .Z(n2310) );
  NANDN U624 ( .A(y[184]), .B(x[184]), .Z(n566) );
  NANDN U625 ( .A(y[183]), .B(x[183]), .Z(n565) );
  NAND U626 ( .A(n566), .B(n565), .Z(n2110) );
  ANDN U627 ( .B(n2310), .A(n2110), .Z(n572) );
  NANDN U628 ( .A(x[183]), .B(y[183]), .Z(n568) );
  NANDN U629 ( .A(x[182]), .B(y[182]), .Z(n567) );
  AND U630 ( .A(n568), .B(n567), .Z(n2313) );
  NANDN U631 ( .A(y[182]), .B(x[182]), .Z(n570) );
  NANDN U632 ( .A(y[181]), .B(x[181]), .Z(n569) );
  NAND U633 ( .A(n570), .B(n569), .Z(n2111) );
  ANDN U634 ( .B(n2313), .A(n2111), .Z(n571) );
  AND U635 ( .A(n572), .B(n571), .Z(n584) );
  NANDN U636 ( .A(x[177]), .B(y[177]), .Z(n574) );
  NANDN U637 ( .A(x[176]), .B(y[176]), .Z(n573) );
  AND U638 ( .A(n574), .B(n573), .Z(n2308) );
  NANDN U639 ( .A(x[173]), .B(y[173]), .Z(n576) );
  NANDN U640 ( .A(x[172]), .B(y[172]), .Z(n575) );
  AND U641 ( .A(n576), .B(n575), .Z(n2305) );
  AND U642 ( .A(n2308), .B(n2305), .Z(n582) );
  NANDN U643 ( .A(x[175]), .B(y[175]), .Z(n578) );
  NANDN U644 ( .A(x[174]), .B(y[174]), .Z(n577) );
  AND U645 ( .A(n578), .B(n577), .Z(n2307) );
  NANDN U646 ( .A(y[174]), .B(x[174]), .Z(n580) );
  NANDN U647 ( .A(y[173]), .B(x[173]), .Z(n579) );
  NAND U648 ( .A(n580), .B(n579), .Z(n2306) );
  ANDN U649 ( .B(n2307), .A(n2306), .Z(n581) );
  AND U650 ( .A(n582), .B(n581), .Z(n583) );
  AND U651 ( .A(n584), .B(n583), .Z(n608) );
  NANDN U652 ( .A(x[185]), .B(y[185]), .Z(n586) );
  NANDN U653 ( .A(x[184]), .B(y[184]), .Z(n585) );
  AND U654 ( .A(n586), .B(n585), .Z(n2315) );
  NANDN U655 ( .A(y[188]), .B(x[188]), .Z(n588) );
  NANDN U656 ( .A(y[187]), .B(x[187]), .Z(n587) );
  NAND U657 ( .A(n588), .B(n587), .Z(n2109) );
  ANDN U658 ( .B(n2315), .A(n2109), .Z(n594) );
  NANDN U659 ( .A(x[187]), .B(y[187]), .Z(n590) );
  NANDN U660 ( .A(x[186]), .B(y[186]), .Z(n589) );
  AND U661 ( .A(n590), .B(n589), .Z(n2318) );
  NANDN U662 ( .A(y[186]), .B(x[186]), .Z(n592) );
  NANDN U663 ( .A(y[185]), .B(x[185]), .Z(n591) );
  NAND U664 ( .A(n592), .B(n591), .Z(n2316) );
  ANDN U665 ( .B(n2318), .A(n2316), .Z(n593) );
  AND U666 ( .A(n594), .B(n593), .Z(n606) );
  NANDN U667 ( .A(x[167]), .B(y[167]), .Z(n596) );
  NANDN U668 ( .A(x[166]), .B(y[166]), .Z(n595) );
  AND U669 ( .A(n596), .B(n595), .Z(n2299) );
  NANDN U670 ( .A(y[164]), .B(x[164]), .Z(n598) );
  NANDN U671 ( .A(y[163]), .B(x[163]), .Z(n597) );
  NAND U672 ( .A(n598), .B(n597), .Z(n2115) );
  ANDN U673 ( .B(n2299), .A(n2115), .Z(n604) );
  NANDN U674 ( .A(x[165]), .B(y[165]), .Z(n600) );
  NANDN U675 ( .A(x[164]), .B(y[164]), .Z(n599) );
  AND U676 ( .A(n600), .B(n599), .Z(n2298) );
  NANDN U677 ( .A(y[172]), .B(x[172]), .Z(n602) );
  NANDN U678 ( .A(y[171]), .B(x[171]), .Z(n601) );
  NAND U679 ( .A(n602), .B(n601), .Z(n2113) );
  ANDN U680 ( .B(n2298), .A(n2113), .Z(n603) );
  AND U681 ( .A(n604), .B(n603), .Z(n605) );
  AND U682 ( .A(n606), .B(n605), .Z(n607) );
  AND U683 ( .A(n608), .B(n607), .Z(n609) );
  AND U684 ( .A(n610), .B(n609), .Z(n706) );
  NANDN U685 ( .A(x[241]), .B(y[241]), .Z(n612) );
  NANDN U686 ( .A(x[240]), .B(y[240]), .Z(n611) );
  AND U687 ( .A(n612), .B(n611), .Z(n2363) );
  NANDN U688 ( .A(x[233]), .B(y[233]), .Z(n614) );
  NANDN U689 ( .A(x[232]), .B(y[232]), .Z(n613) );
  AND U690 ( .A(n614), .B(n613), .Z(n2356) );
  AND U691 ( .A(n2363), .B(n2356), .Z(n620) );
  NANDN U692 ( .A(x[237]), .B(y[237]), .Z(n616) );
  NANDN U693 ( .A(x[236]), .B(y[236]), .Z(n615) );
  AND U694 ( .A(n616), .B(n615), .Z(n2359) );
  NANDN U695 ( .A(x[235]), .B(y[235]), .Z(n618) );
  NANDN U696 ( .A(x[234]), .B(y[234]), .Z(n617) );
  AND U697 ( .A(n618), .B(n617), .Z(n2358) );
  AND U698 ( .A(n2359), .B(n2358), .Z(n619) );
  AND U699 ( .A(n620), .B(n619), .Z(n632) );
  NANDN U700 ( .A(y[232]), .B(x[232]), .Z(n622) );
  NANDN U701 ( .A(y[231]), .B(x[231]), .Z(n621) );
  AND U702 ( .A(n622), .B(n621), .Z(n2355) );
  NANDN U703 ( .A(y[226]), .B(x[226]), .Z(n624) );
  NANDN U704 ( .A(y[225]), .B(x[225]), .Z(n623) );
  NAND U705 ( .A(n624), .B(n623), .Z(n2350) );
  ANDN U706 ( .B(n2355), .A(n2350), .Z(n630) );
  NANDN U707 ( .A(x[231]), .B(y[231]), .Z(n626) );
  NANDN U708 ( .A(x[230]), .B(y[230]), .Z(n625) );
  AND U709 ( .A(n626), .B(n625), .Z(n2354) );
  NANDN U710 ( .A(y[228]), .B(x[228]), .Z(n628) );
  NANDN U711 ( .A(y[227]), .B(x[227]), .Z(n627) );
  NAND U712 ( .A(n628), .B(n627), .Z(n2098) );
  ANDN U713 ( .B(n2354), .A(n2098), .Z(n629) );
  AND U714 ( .A(n630), .B(n629), .Z(n631) );
  AND U715 ( .A(n632), .B(n631), .Z(n656) );
  NANDN U716 ( .A(x[260]), .B(y[260]), .Z(n634) );
  NANDN U717 ( .A(x[259]), .B(y[259]), .Z(n633) );
  AND U718 ( .A(n634), .B(n633), .Z(n2387) );
  NANDN U719 ( .A(y[244]), .B(x[244]), .Z(n636) );
  NANDN U720 ( .A(y[243]), .B(x[243]), .Z(n635) );
  NAND U721 ( .A(n636), .B(n635), .Z(n2366) );
  ANDN U722 ( .B(n2387), .A(n2366), .Z(n642) );
  NANDN U723 ( .A(y[259]), .B(x[259]), .Z(n638) );
  NANDN U724 ( .A(y[258]), .B(x[258]), .Z(n637) );
  AND U725 ( .A(n638), .B(n637), .Z(n2386) );
  NANDN U726 ( .A(y[246]), .B(x[246]), .Z(n640) );
  NANDN U727 ( .A(y[245]), .B(x[245]), .Z(n639) );
  NAND U728 ( .A(n640), .B(n639), .Z(n2094) );
  ANDN U729 ( .B(n2386), .A(n2094), .Z(n641) );
  AND U730 ( .A(n642), .B(n641), .Z(n654) );
  NANDN U731 ( .A(x[225]), .B(y[225]), .Z(n644) );
  NANDN U732 ( .A(x[224]), .B(y[224]), .Z(n643) );
  AND U733 ( .A(n644), .B(n643), .Z(n2349) );
  NANDN U734 ( .A(x[223]), .B(y[223]), .Z(n646) );
  NANDN U735 ( .A(x[222]), .B(y[222]), .Z(n645) );
  AND U736 ( .A(n646), .B(n645), .Z(n2348) );
  AND U737 ( .A(n2349), .B(n2348), .Z(n652) );
  NANDN U738 ( .A(x[227]), .B(y[227]), .Z(n648) );
  NANDN U739 ( .A(x[226]), .B(y[226]), .Z(n647) );
  AND U740 ( .A(n648), .B(n647), .Z(n2351) );
  NANDN U741 ( .A(y[224]), .B(x[224]), .Z(n650) );
  NANDN U742 ( .A(y[223]), .B(x[223]), .Z(n649) );
  NAND U743 ( .A(n650), .B(n649), .Z(n2099) );
  ANDN U744 ( .B(n2351), .A(n2099), .Z(n651) );
  AND U745 ( .A(n652), .B(n651), .Z(n653) );
  AND U746 ( .A(n654), .B(n653), .Z(n655) );
  AND U747 ( .A(n656), .B(n655), .Z(n704) );
  NANDN U748 ( .A(x[155]), .B(y[155]), .Z(n658) );
  NANDN U749 ( .A(x[154]), .B(y[154]), .Z(n657) );
  AND U750 ( .A(n658), .B(n657), .Z(n2289) );
  NANDN U751 ( .A(y[150]), .B(x[150]), .Z(n660) );
  NANDN U752 ( .A(y[149]), .B(x[149]), .Z(n659) );
  NAND U753 ( .A(n660), .B(n659), .Z(n2284) );
  ANDN U754 ( .B(n2289), .A(n2284), .Z(n666) );
  NANDN U755 ( .A(y[154]), .B(x[154]), .Z(n662) );
  NANDN U756 ( .A(y[153]), .B(x[153]), .Z(n661) );
  AND U757 ( .A(n662), .B(n661), .Z(n2287) );
  NANDN U758 ( .A(y[152]), .B(x[152]), .Z(n664) );
  NANDN U759 ( .A(y[151]), .B(x[151]), .Z(n663) );
  NAND U760 ( .A(n664), .B(n663), .Z(n2117) );
  ANDN U761 ( .B(n2287), .A(n2117), .Z(n665) );
  AND U762 ( .A(n666), .B(n665), .Z(n678) );
  NANDN U763 ( .A(x[149]), .B(y[149]), .Z(n668) );
  NANDN U764 ( .A(x[148]), .B(y[148]), .Z(n667) );
  AND U765 ( .A(n668), .B(n667), .Z(n2283) );
  NANDN U766 ( .A(x[141]), .B(y[141]), .Z(n670) );
  NANDN U767 ( .A(x[140]), .B(y[140]), .Z(n669) );
  AND U768 ( .A(n670), .B(n669), .Z(n2277) );
  AND U769 ( .A(n2283), .B(n2277), .Z(n676) );
  NANDN U770 ( .A(x[147]), .B(y[147]), .Z(n672) );
  NANDN U771 ( .A(x[146]), .B(y[146]), .Z(n671) );
  AND U772 ( .A(n672), .B(n671), .Z(n2282) );
  NANDN U773 ( .A(y[148]), .B(x[148]), .Z(n674) );
  NANDN U774 ( .A(y[147]), .B(x[147]), .Z(n673) );
  NAND U775 ( .A(n674), .B(n673), .Z(n2118) );
  ANDN U776 ( .B(n2282), .A(n2118), .Z(n675) );
  AND U777 ( .A(n676), .B(n675), .Z(n677) );
  AND U778 ( .A(n678), .B(n677), .Z(n702) );
  NANDN U779 ( .A(x[163]), .B(y[163]), .Z(n680) );
  NANDN U780 ( .A(x[162]), .B(y[162]), .Z(n679) );
  AND U781 ( .A(n680), .B(n679), .Z(n2297) );
  NANDN U782 ( .A(y[156]), .B(x[156]), .Z(n682) );
  NANDN U783 ( .A(y[155]), .B(x[155]), .Z(n681) );
  NAND U784 ( .A(n682), .B(n681), .Z(n2290) );
  ANDN U785 ( .B(n2297), .A(n2290), .Z(n688) );
  NANDN U786 ( .A(x[157]), .B(y[157]), .Z(n684) );
  NANDN U787 ( .A(x[156]), .B(y[156]), .Z(n683) );
  AND U788 ( .A(n684), .B(n683), .Z(n2292) );
  NANDN U789 ( .A(y[160]), .B(x[160]), .Z(n686) );
  NANDN U790 ( .A(y[159]), .B(x[159]), .Z(n685) );
  NAND U791 ( .A(n686), .B(n685), .Z(n2116) );
  ANDN U792 ( .B(n2292), .A(n2116), .Z(n687) );
  AND U793 ( .A(n688), .B(n687), .Z(n700) );
  NANDN U794 ( .A(x[139]), .B(y[139]), .Z(n690) );
  NANDN U795 ( .A(x[138]), .B(y[138]), .Z(n689) );
  AND U796 ( .A(n690), .B(n689), .Z(n2274) );
  NANDN U797 ( .A(y[138]), .B(x[138]), .Z(n692) );
  NANDN U798 ( .A(y[137]), .B(x[137]), .Z(n691) );
  NAND U799 ( .A(n692), .B(n691), .Z(n2273) );
  ANDN U800 ( .B(n2274), .A(n2273), .Z(n698) );
  NANDN U801 ( .A(y[132]), .B(x[132]), .Z(n694) );
  NANDN U802 ( .A(y[131]), .B(x[131]), .Z(n693) );
  AND U803 ( .A(n694), .B(n693), .Z(n2269) );
  NANDN U804 ( .A(y[130]), .B(x[130]), .Z(n696) );
  NANDN U805 ( .A(y[129]), .B(x[129]), .Z(n695) );
  NAND U806 ( .A(n696), .B(n695), .Z(n2122) );
  ANDN U807 ( .B(n2269), .A(n2122), .Z(n697) );
  AND U808 ( .A(n698), .B(n697), .Z(n699) );
  AND U809 ( .A(n700), .B(n699), .Z(n701) );
  AND U810 ( .A(n702), .B(n701), .Z(n703) );
  AND U811 ( .A(n704), .B(n703), .Z(n705) );
  AND U812 ( .A(n706), .B(n705), .Z(n898) );
  NANDN U813 ( .A(x[79]), .B(y[79]), .Z(n708) );
  NANDN U814 ( .A(x[78]), .B(y[78]), .Z(n707) );
  AND U815 ( .A(n708), .B(n707), .Z(n2226) );
  NANDN U816 ( .A(x[71]), .B(y[71]), .Z(n710) );
  NANDN U817 ( .A(x[70]), .B(y[70]), .Z(n709) );
  AND U818 ( .A(n710), .B(n709), .Z(n2220) );
  AND U819 ( .A(n2226), .B(n2220), .Z(n716) );
  NANDN U820 ( .A(x[73]), .B(y[73]), .Z(n712) );
  NANDN U821 ( .A(x[72]), .B(y[72]), .Z(n711) );
  AND U822 ( .A(n712), .B(n711), .Z(n2221) );
  NANDN U823 ( .A(y[72]), .B(x[72]), .Z(n714) );
  NANDN U824 ( .A(y[71]), .B(x[71]), .Z(n713) );
  NAND U825 ( .A(n714), .B(n713), .Z(n2138) );
  ANDN U826 ( .B(n2221), .A(n2138), .Z(n715) );
  AND U827 ( .A(n716), .B(n715), .Z(n728) );
  NANDN U828 ( .A(y[70]), .B(x[70]), .Z(n718) );
  NANDN U829 ( .A(y[69]), .B(x[69]), .Z(n717) );
  AND U830 ( .A(n718), .B(n717), .Z(n2218) );
  NANDN U831 ( .A(y[60]), .B(x[60]), .Z(n720) );
  NANDN U832 ( .A(y[59]), .B(x[59]), .Z(n719) );
  NAND U833 ( .A(n720), .B(n719), .Z(n2212) );
  ANDN U834 ( .B(n2218), .A(n2212), .Z(n726) );
  NANDN U835 ( .A(y[68]), .B(x[68]), .Z(n722) );
  NANDN U836 ( .A(y[67]), .B(x[67]), .Z(n721) );
  AND U837 ( .A(n722), .B(n721), .Z(n2217) );
  NANDN U838 ( .A(y[62]), .B(x[62]), .Z(n724) );
  NANDN U839 ( .A(y[61]), .B(x[61]), .Z(n723) );
  NAND U840 ( .A(n724), .B(n723), .Z(n2213) );
  ANDN U841 ( .B(n2217), .A(n2213), .Z(n725) );
  AND U842 ( .A(n726), .B(n725), .Z(n727) );
  AND U843 ( .A(n728), .B(n727), .Z(n752) );
  NANDN U844 ( .A(x[81]), .B(y[81]), .Z(n730) );
  NANDN U845 ( .A(x[80]), .B(y[80]), .Z(n729) );
  AND U846 ( .A(n730), .B(n729), .Z(n2227) );
  NANDN U847 ( .A(y[92]), .B(x[92]), .Z(n732) );
  NANDN U848 ( .A(y[91]), .B(x[91]), .Z(n731) );
  NAND U849 ( .A(n732), .B(n731), .Z(n2133) );
  ANDN U850 ( .B(n2227), .A(n2133), .Z(n738) );
  NANDN U851 ( .A(y[86]), .B(x[86]), .Z(n734) );
  NANDN U852 ( .A(y[85]), .B(x[85]), .Z(n733) );
  AND U853 ( .A(n734), .B(n733), .Z(n2232) );
  NANDN U854 ( .A(y[82]), .B(x[82]), .Z(n736) );
  NANDN U855 ( .A(y[81]), .B(x[81]), .Z(n735) );
  NAND U856 ( .A(n736), .B(n735), .Z(n2228) );
  ANDN U857 ( .B(n2232), .A(n2228), .Z(n737) );
  AND U858 ( .A(n738), .B(n737), .Z(n750) );
  NANDN U859 ( .A(x[59]), .B(y[59]), .Z(n740) );
  NANDN U860 ( .A(x[58]), .B(y[58]), .Z(n739) );
  AND U861 ( .A(n740), .B(n739), .Z(n2211) );
  NANDN U862 ( .A(x[51]), .B(y[51]), .Z(n742) );
  NANDN U863 ( .A(x[50]), .B(y[50]), .Z(n741) );
  AND U864 ( .A(n742), .B(n741), .Z(n2205) );
  AND U865 ( .A(n2211), .B(n2205), .Z(n748) );
  NANDN U866 ( .A(x[57]), .B(y[57]), .Z(n744) );
  NANDN U867 ( .A(x[56]), .B(y[56]), .Z(n743) );
  AND U868 ( .A(n744), .B(n743), .Z(n2209) );
  NANDN U869 ( .A(y[58]), .B(x[58]), .Z(n746) );
  NANDN U870 ( .A(y[57]), .B(x[57]), .Z(n745) );
  NAND U871 ( .A(n746), .B(n745), .Z(n2145) );
  ANDN U872 ( .B(n2209), .A(n2145), .Z(n747) );
  AND U873 ( .A(n748), .B(n747), .Z(n749) );
  AND U874 ( .A(n750), .B(n749), .Z(n751) );
  AND U875 ( .A(n752), .B(n751), .Z(n800) );
  NANDN U876 ( .A(x[39]), .B(y[39]), .Z(n754) );
  NANDN U877 ( .A(x[38]), .B(y[38]), .Z(n753) );
  AND U878 ( .A(n754), .B(n753), .Z(n2195) );
  NANDN U879 ( .A(y[36]), .B(x[36]), .Z(n756) );
  NANDN U880 ( .A(y[35]), .B(x[35]), .Z(n755) );
  NAND U881 ( .A(n756), .B(n755), .Z(n2193) );
  ANDN U882 ( .B(n2195), .A(n2193), .Z(n762) );
  NANDN U883 ( .A(x[37]), .B(y[37]), .Z(n758) );
  NANDN U884 ( .A(x[36]), .B(y[36]), .Z(n757) );
  AND U885 ( .A(n758), .B(n757), .Z(n2194) );
  NANDN U886 ( .A(y[38]), .B(x[38]), .Z(n760) );
  NANDN U887 ( .A(y[37]), .B(x[37]), .Z(n759) );
  NAND U888 ( .A(n760), .B(n759), .Z(n2151) );
  ANDN U889 ( .B(n2194), .A(n2151), .Z(n761) );
  AND U890 ( .A(n762), .B(n761), .Z(n774) );
  NANDN U891 ( .A(x[35]), .B(y[35]), .Z(n764) );
  NANDN U892 ( .A(x[34]), .B(y[34]), .Z(n763) );
  AND U893 ( .A(n764), .B(n763), .Z(n2192) );
  NANDN U894 ( .A(y[30]), .B(x[30]), .Z(n766) );
  NANDN U895 ( .A(y[29]), .B(x[29]), .Z(n765) );
  NAND U896 ( .A(n766), .B(n765), .Z(n2188) );
  ANDN U897 ( .B(n2192), .A(n2188), .Z(n772) );
  NANDN U898 ( .A(x[31]), .B(y[31]), .Z(n768) );
  NANDN U899 ( .A(x[30]), .B(y[30]), .Z(n767) );
  AND U900 ( .A(n768), .B(n767), .Z(n2190) );
  NANDN U901 ( .A(y[34]), .B(x[34]), .Z(n770) );
  NANDN U902 ( .A(y[33]), .B(x[33]), .Z(n769) );
  NAND U903 ( .A(n770), .B(n769), .Z(n2152) );
  ANDN U904 ( .B(n2190), .A(n2152), .Z(n771) );
  AND U905 ( .A(n772), .B(n771), .Z(n773) );
  AND U906 ( .A(n774), .B(n773), .Z(n798) );
  NANDN U907 ( .A(x[49]), .B(y[49]), .Z(n776) );
  NANDN U908 ( .A(x[48]), .B(y[48]), .Z(n775) );
  AND U909 ( .A(n776), .B(n775), .Z(n2204) );
  NANDN U910 ( .A(y[40]), .B(x[40]), .Z(n778) );
  NANDN U911 ( .A(y[39]), .B(x[39]), .Z(n777) );
  NAND U912 ( .A(n778), .B(n777), .Z(n2150) );
  ANDN U913 ( .B(n2204), .A(n2150), .Z(n784) );
  NANDN U914 ( .A(x[43]), .B(y[43]), .Z(n780) );
  NANDN U915 ( .A(x[42]), .B(y[42]), .Z(n779) );
  AND U916 ( .A(n780), .B(n779), .Z(n2199) );
  NANDN U917 ( .A(x[41]), .B(y[41]), .Z(n782) );
  NANDN U918 ( .A(x[40]), .B(y[40]), .Z(n781) );
  AND U919 ( .A(n782), .B(n781), .Z(n2196) );
  AND U920 ( .A(n2199), .B(n2196), .Z(n783) );
  AND U921 ( .A(n784), .B(n783), .Z(n796) );
  NANDN U922 ( .A(x[27]), .B(y[27]), .Z(n786) );
  NANDN U923 ( .A(x[26]), .B(y[26]), .Z(n785) );
  AND U924 ( .A(n786), .B(n785), .Z(n2185) );
  NANDN U925 ( .A(x[23]), .B(y[23]), .Z(n788) );
  NANDN U926 ( .A(x[22]), .B(y[22]), .Z(n787) );
  AND U927 ( .A(n788), .B(n787), .Z(n2182) );
  AND U928 ( .A(n2185), .B(n2182), .Z(n794) );
  NANDN U929 ( .A(x[25]), .B(y[25]), .Z(n790) );
  NANDN U930 ( .A(x[24]), .B(y[24]), .Z(n789) );
  AND U931 ( .A(n790), .B(n789), .Z(n2184) );
  NANDN U932 ( .A(y[26]), .B(x[26]), .Z(n792) );
  NANDN U933 ( .A(y[25]), .B(x[25]), .Z(n791) );
  NAND U934 ( .A(n792), .B(n791), .Z(n2155) );
  ANDN U935 ( .B(n2184), .A(n2155), .Z(n793) );
  AND U936 ( .A(n794), .B(n793), .Z(n795) );
  AND U937 ( .A(n796), .B(n795), .Z(n797) );
  AND U938 ( .A(n798), .B(n797), .Z(n799) );
  AND U939 ( .A(n800), .B(n799), .Z(n896) );
  NANDN U940 ( .A(x[113]), .B(y[113]), .Z(n802) );
  NANDN U941 ( .A(x[112]), .B(y[112]), .Z(n801) );
  AND U942 ( .A(n802), .B(n801), .Z(n2254) );
  NANDN U943 ( .A(y[104]), .B(x[104]), .Z(n804) );
  NANDN U944 ( .A(y[103]), .B(x[103]), .Z(n803) );
  NAND U945 ( .A(n804), .B(n803), .Z(n2129) );
  ANDN U946 ( .B(n2254), .A(n2129), .Z(n810) );
  NANDN U947 ( .A(x[107]), .B(y[107]), .Z(n806) );
  NANDN U948 ( .A(x[106]), .B(y[106]), .Z(n805) );
  AND U949 ( .A(n806), .B(n805), .Z(n2248) );
  NANDN U950 ( .A(x[105]), .B(y[105]), .Z(n808) );
  NANDN U951 ( .A(x[104]), .B(y[104]), .Z(n807) );
  AND U952 ( .A(n808), .B(n807), .Z(n2246) );
  AND U953 ( .A(n2248), .B(n2246), .Z(n809) );
  AND U954 ( .A(n810), .B(n809), .Z(n822) );
  NANDN U955 ( .A(x[103]), .B(y[103]), .Z(n812) );
  NANDN U956 ( .A(x[102]), .B(y[102]), .Z(n811) );
  AND U957 ( .A(n812), .B(n811), .Z(n2245) );
  NANDN U958 ( .A(x[95]), .B(y[95]), .Z(n814) );
  NANDN U959 ( .A(x[94]), .B(y[94]), .Z(n813) );
  AND U960 ( .A(n814), .B(n813), .Z(n2239) );
  AND U961 ( .A(n2245), .B(n2239), .Z(n820) );
  NANDN U962 ( .A(x[97]), .B(y[97]), .Z(n816) );
  NANDN U963 ( .A(x[96]), .B(y[96]), .Z(n815) );
  AND U964 ( .A(n816), .B(n815), .Z(n2240) );
  NANDN U965 ( .A(y[96]), .B(x[96]), .Z(n818) );
  NANDN U966 ( .A(y[95]), .B(x[95]), .Z(n817) );
  NAND U967 ( .A(n818), .B(n817), .Z(n2132) );
  ANDN U968 ( .B(n2240), .A(n2132), .Z(n819) );
  AND U969 ( .A(n820), .B(n819), .Z(n821) );
  AND U970 ( .A(n822), .B(n821), .Z(n846) );
  NANDN U971 ( .A(x[115]), .B(y[115]), .Z(n824) );
  NANDN U972 ( .A(x[114]), .B(y[114]), .Z(n823) );
  AND U973 ( .A(n824), .B(n823), .Z(n2256) );
  NANDN U974 ( .A(y[124]), .B(x[124]), .Z(n826) );
  NANDN U975 ( .A(y[123]), .B(x[123]), .Z(n825) );
  NAND U976 ( .A(n826), .B(n825), .Z(n2123) );
  ANDN U977 ( .B(n2256), .A(n2123), .Z(n832) );
  NANDN U978 ( .A(x[121]), .B(y[121]), .Z(n828) );
  NANDN U979 ( .A(x[120]), .B(y[120]), .Z(n827) );
  AND U980 ( .A(n828), .B(n827), .Z(n2260) );
  NANDN U981 ( .A(y[122]), .B(x[122]), .Z(n830) );
  NANDN U982 ( .A(y[121]), .B(x[121]), .Z(n829) );
  NAND U983 ( .A(n830), .B(n829), .Z(n2124) );
  ANDN U984 ( .B(n2260), .A(n2124), .Z(n831) );
  AND U985 ( .A(n832), .B(n831), .Z(n844) );
  NANDN U986 ( .A(x[89]), .B(y[89]), .Z(n834) );
  NANDN U987 ( .A(x[88]), .B(y[88]), .Z(n833) );
  AND U988 ( .A(n834), .B(n833), .Z(n2235) );
  NANDN U989 ( .A(y[94]), .B(x[94]), .Z(n836) );
  NANDN U990 ( .A(y[93]), .B(x[93]), .Z(n835) );
  NAND U991 ( .A(n836), .B(n835), .Z(n2238) );
  ANDN U992 ( .B(n2235), .A(n2238), .Z(n842) );
  NANDN U993 ( .A(x[93]), .B(y[93]), .Z(n838) );
  NANDN U994 ( .A(x[92]), .B(y[92]), .Z(n837) );
  AND U995 ( .A(n838), .B(n837), .Z(n2237) );
  NANDN U996 ( .A(y[90]), .B(x[90]), .Z(n840) );
  NANDN U997 ( .A(y[89]), .B(x[89]), .Z(n839) );
  NAND U998 ( .A(n840), .B(n839), .Z(n2134) );
  ANDN U999 ( .B(n2237), .A(n2134), .Z(n841) );
  AND U1000 ( .A(n842), .B(n841), .Z(n843) );
  AND U1001 ( .A(n844), .B(n843), .Z(n845) );
  AND U1002 ( .A(n846), .B(n845), .Z(n894) );
  NANDN U1003 ( .A(x[15]), .B(y[15]), .Z(n848) );
  NANDN U1004 ( .A(x[14]), .B(y[14]), .Z(n847) );
  AND U1005 ( .A(n848), .B(n847), .Z(n2176) );
  NANDN U1006 ( .A(y[18]), .B(x[18]), .Z(n850) );
  NANDN U1007 ( .A(y[17]), .B(x[17]), .Z(n849) );
  NAND U1008 ( .A(n850), .B(n849), .Z(n2179) );
  ANDN U1009 ( .B(n2176), .A(n2179), .Z(n856) );
  NANDN U1010 ( .A(x[17]), .B(y[17]), .Z(n852) );
  NANDN U1011 ( .A(x[16]), .B(y[16]), .Z(n851) );
  AND U1012 ( .A(n852), .B(n851), .Z(n2178) );
  NANDN U1013 ( .A(y[16]), .B(x[16]), .Z(n854) );
  NANDN U1014 ( .A(y[15]), .B(x[15]), .Z(n853) );
  NAND U1015 ( .A(n854), .B(n853), .Z(n2158) );
  ANDN U1016 ( .B(n2178), .A(n2158), .Z(n855) );
  AND U1017 ( .A(n856), .B(n855), .Z(n868) );
  NANDN U1018 ( .A(y[14]), .B(x[14]), .Z(n858) );
  NANDN U1019 ( .A(y[13]), .B(x[13]), .Z(n857) );
  AND U1020 ( .A(n858), .B(n857), .Z(n2175) );
  NANDN U1021 ( .A(y[6]), .B(x[6]), .Z(n860) );
  NANDN U1022 ( .A(y[5]), .B(x[5]), .Z(n859) );
  NAND U1023 ( .A(n860), .B(n859), .Z(n2169) );
  ANDN U1024 ( .B(n2175), .A(n2169), .Z(n866) );
  NANDN U1025 ( .A(x[13]), .B(y[13]), .Z(n862) );
  NANDN U1026 ( .A(x[12]), .B(y[12]), .Z(n861) );
  AND U1027 ( .A(n862), .B(n861), .Z(n2174) );
  NANDN U1028 ( .A(x[11]), .B(y[11]), .Z(n864) );
  NANDN U1029 ( .A(x[10]), .B(y[10]), .Z(n863) );
  AND U1030 ( .A(n864), .B(n863), .Z(n2172) );
  AND U1031 ( .A(n2174), .B(n2172), .Z(n865) );
  AND U1032 ( .A(n866), .B(n865), .Z(n867) );
  AND U1033 ( .A(n868), .B(n867), .Z(n892) );
  NANDN U1034 ( .A(x[19]), .B(y[19]), .Z(n870) );
  NANDN U1035 ( .A(x[18]), .B(y[18]), .Z(n869) );
  AND U1036 ( .A(n870), .B(n869), .Z(n2180) );
  NANDN U1037 ( .A(y[22]), .B(x[22]), .Z(n872) );
  NANDN U1038 ( .A(y[21]), .B(x[21]), .Z(n871) );
  NAND U1039 ( .A(n872), .B(n871), .Z(n2156) );
  ANDN U1040 ( .B(n2180), .A(n2156), .Z(n878) );
  NANDN U1041 ( .A(x[21]), .B(y[21]), .Z(n874) );
  NANDN U1042 ( .A(x[20]), .B(y[20]), .Z(n873) );
  AND U1043 ( .A(n874), .B(n873), .Z(n2181) );
  NANDN U1044 ( .A(y[24]), .B(x[24]), .Z(n876) );
  NANDN U1045 ( .A(y[23]), .B(x[23]), .Z(n875) );
  NAND U1046 ( .A(n876), .B(n875), .Z(n2183) );
  ANDN U1047 ( .B(n2181), .A(n2183), .Z(n877) );
  AND U1048 ( .A(n878), .B(n877), .Z(n890) );
  NANDN U1049 ( .A(y[4]), .B(x[4]), .Z(n880) );
  NANDN U1050 ( .A(y[3]), .B(x[3]), .Z(n879) );
  AND U1051 ( .A(n880), .B(n879), .Z(n2167) );
  NANDN U1052 ( .A(y[314]), .B(x[314]), .Z(n882) );
  NANDN U1053 ( .A(y[313]), .B(x[313]), .Z(n881) );
  NAND U1054 ( .A(n882), .B(n881), .Z(n2072) );
  ANDN U1055 ( .B(n2167), .A(n2072), .Z(n888) );
  NANDN U1056 ( .A(x[313]), .B(y[313]), .Z(n884) );
  NANDN U1057 ( .A(x[312]), .B(y[312]), .Z(n883) );
  AND U1058 ( .A(n884), .B(n883), .Z(n2436) );
  NANDN U1059 ( .A(y[2]), .B(x[2]), .Z(n886) );
  NANDN U1060 ( .A(y[1]), .B(x[1]), .Z(n885) );
  NAND U1061 ( .A(n886), .B(n885), .Z(n2161) );
  ANDN U1062 ( .B(n2436), .A(n2161), .Z(n887) );
  AND U1063 ( .A(n888), .B(n887), .Z(n889) );
  AND U1064 ( .A(n890), .B(n889), .Z(n891) );
  AND U1065 ( .A(n892), .B(n891), .Z(n893) );
  AND U1066 ( .A(n894), .B(n893), .Z(n895) );
  AND U1067 ( .A(n896), .B(n895), .Z(n897) );
  AND U1068 ( .A(n898), .B(n897), .Z(n2019) );
  NANDN U1069 ( .A(x[87]), .B(y[87]), .Z(n900) );
  NANDN U1070 ( .A(x[86]), .B(y[86]), .Z(n899) );
  AND U1071 ( .A(n900), .B(n899), .Z(n2233) );
  NANDN U1072 ( .A(y[84]), .B(x[84]), .Z(n902) );
  NANDN U1073 ( .A(y[83]), .B(x[83]), .Z(n901) );
  NAND U1074 ( .A(n902), .B(n901), .Z(n2135) );
  ANDN U1075 ( .B(n2233), .A(n2135), .Z(n908) );
  NANDN U1076 ( .A(x[85]), .B(y[85]), .Z(n904) );
  NANDN U1077 ( .A(x[84]), .B(y[84]), .Z(n903) );
  AND U1078 ( .A(n904), .B(n903), .Z(n2231) );
  NANDN U1079 ( .A(y[98]), .B(x[98]), .Z(n906) );
  NANDN U1080 ( .A(y[97]), .B(x[97]), .Z(n905) );
  NAND U1081 ( .A(n906), .B(n905), .Z(n2131) );
  ANDN U1082 ( .B(n2231), .A(n2131), .Z(n907) );
  AND U1083 ( .A(n908), .B(n907), .Z(n920) );
  NANDN U1084 ( .A(x[83]), .B(y[83]), .Z(n910) );
  NANDN U1085 ( .A(x[82]), .B(y[82]), .Z(n909) );
  AND U1086 ( .A(n910), .B(n909), .Z(n2229) );
  NANDN U1087 ( .A(y[76]), .B(x[76]), .Z(n912) );
  NANDN U1088 ( .A(y[75]), .B(x[75]), .Z(n911) );
  NAND U1089 ( .A(n912), .B(n911), .Z(n2224) );
  ANDN U1090 ( .B(n2229), .A(n2224), .Z(n918) );
  NANDN U1091 ( .A(x[77]), .B(y[77]), .Z(n914) );
  NANDN U1092 ( .A(x[76]), .B(y[76]), .Z(n913) );
  AND U1093 ( .A(n914), .B(n913), .Z(n2225) );
  NANDN U1094 ( .A(y[78]), .B(x[78]), .Z(n916) );
  NANDN U1095 ( .A(y[77]), .B(x[77]), .Z(n915) );
  NAND U1096 ( .A(n916), .B(n915), .Z(n2137) );
  ANDN U1097 ( .B(n2225), .A(n2137), .Z(n917) );
  AND U1098 ( .A(n918), .B(n917), .Z(n919) );
  AND U1099 ( .A(n920), .B(n919), .Z(n944) );
  NANDN U1100 ( .A(y[108]), .B(x[108]), .Z(n922) );
  NANDN U1101 ( .A(y[107]), .B(x[107]), .Z(n921) );
  AND U1102 ( .A(n922), .B(n921), .Z(n2249) );
  NANDN U1103 ( .A(y[88]), .B(x[88]), .Z(n924) );
  NANDN U1104 ( .A(y[87]), .B(x[87]), .Z(n923) );
  NAND U1105 ( .A(n924), .B(n923), .Z(n2234) );
  ANDN U1106 ( .B(n2249), .A(n2234), .Z(n930) );
  NANDN U1107 ( .A(x[99]), .B(y[99]), .Z(n926) );
  NANDN U1108 ( .A(x[98]), .B(y[98]), .Z(n925) );
  AND U1109 ( .A(n926), .B(n925), .Z(n2242) );
  NANDN U1110 ( .A(y[100]), .B(x[100]), .Z(n928) );
  NANDN U1111 ( .A(y[99]), .B(x[99]), .Z(n927) );
  NAND U1112 ( .A(n928), .B(n927), .Z(n2243) );
  ANDN U1113 ( .B(n2242), .A(n2243), .Z(n929) );
  AND U1114 ( .A(n930), .B(n929), .Z(n942) );
  NANDN U1115 ( .A(y[74]), .B(x[74]), .Z(n932) );
  NANDN U1116 ( .A(y[73]), .B(x[73]), .Z(n931) );
  AND U1117 ( .A(n932), .B(n931), .Z(n2222) );
  NANDN U1118 ( .A(y[66]), .B(x[66]), .Z(n934) );
  NANDN U1119 ( .A(y[65]), .B(x[65]), .Z(n933) );
  NAND U1120 ( .A(n934), .B(n933), .Z(n2141) );
  ANDN U1121 ( .B(n2222), .A(n2141), .Z(n940) );
  NANDN U1122 ( .A(x[67]), .B(y[67]), .Z(n936) );
  NANDN U1123 ( .A(x[66]), .B(y[66]), .Z(n935) );
  AND U1124 ( .A(n936), .B(n935), .Z(n2216) );
  NANDN U1125 ( .A(x[75]), .B(y[75]), .Z(n938) );
  NANDN U1126 ( .A(x[74]), .B(y[74]), .Z(n937) );
  AND U1127 ( .A(n938), .B(n937), .Z(n2223) );
  AND U1128 ( .A(n2216), .B(n2223), .Z(n939) );
  AND U1129 ( .A(n940), .B(n939), .Z(n941) );
  AND U1130 ( .A(n942), .B(n941), .Z(n943) );
  AND U1131 ( .A(n944), .B(n943), .Z(n992) );
  NANDN U1132 ( .A(x[55]), .B(y[55]), .Z(n946) );
  NANDN U1133 ( .A(x[54]), .B(y[54]), .Z(n945) );
  AND U1134 ( .A(n946), .B(n945), .Z(n2208) );
  NANDN U1135 ( .A(y[48]), .B(x[48]), .Z(n948) );
  NANDN U1136 ( .A(y[47]), .B(x[47]), .Z(n947) );
  NAND U1137 ( .A(n948), .B(n947), .Z(n2203) );
  ANDN U1138 ( .B(n2208), .A(n2203), .Z(n954) );
  NANDN U1139 ( .A(y[54]), .B(x[54]), .Z(n950) );
  NANDN U1140 ( .A(y[53]), .B(x[53]), .Z(n949) );
  AND U1141 ( .A(n950), .B(n949), .Z(n2207) );
  NANDN U1142 ( .A(y[52]), .B(x[52]), .Z(n952) );
  NANDN U1143 ( .A(y[51]), .B(x[51]), .Z(n951) );
  NAND U1144 ( .A(n952), .B(n951), .Z(n2147) );
  ANDN U1145 ( .B(n2207), .A(n2147), .Z(n953) );
  AND U1146 ( .A(n954), .B(n953), .Z(n966) );
  NANDN U1147 ( .A(x[53]), .B(y[53]), .Z(n956) );
  NANDN U1148 ( .A(x[52]), .B(y[52]), .Z(n955) );
  AND U1149 ( .A(n956), .B(n955), .Z(n2206) );
  NANDN U1150 ( .A(x[45]), .B(y[45]), .Z(n958) );
  NANDN U1151 ( .A(x[44]), .B(y[44]), .Z(n957) );
  AND U1152 ( .A(n958), .B(n957), .Z(n2201) );
  AND U1153 ( .A(n2206), .B(n2201), .Z(n964) );
  NANDN U1154 ( .A(x[47]), .B(y[47]), .Z(n960) );
  NANDN U1155 ( .A(x[46]), .B(y[46]), .Z(n959) );
  AND U1156 ( .A(n960), .B(n959), .Z(n2202) );
  NANDN U1157 ( .A(y[46]), .B(x[46]), .Z(n962) );
  NANDN U1158 ( .A(y[45]), .B(x[45]), .Z(n961) );
  NAND U1159 ( .A(n962), .B(n961), .Z(n2149) );
  ANDN U1160 ( .B(n2202), .A(n2149), .Z(n963) );
  AND U1161 ( .A(n964), .B(n963), .Z(n965) );
  AND U1162 ( .A(n966), .B(n965), .Z(n990) );
  NANDN U1163 ( .A(x[65]), .B(y[65]), .Z(n968) );
  NANDN U1164 ( .A(x[64]), .B(y[64]), .Z(n967) );
  AND U1165 ( .A(n968), .B(n967), .Z(n2215) );
  NANDN U1166 ( .A(y[64]), .B(x[64]), .Z(n970) );
  NANDN U1167 ( .A(y[63]), .B(x[63]), .Z(n969) );
  NAND U1168 ( .A(n970), .B(n969), .Z(n2142) );
  ANDN U1169 ( .B(n2215), .A(n2142), .Z(n976) );
  NANDN U1170 ( .A(x[63]), .B(y[63]), .Z(n972) );
  NANDN U1171 ( .A(x[62]), .B(y[62]), .Z(n971) );
  AND U1172 ( .A(n972), .B(n971), .Z(n2214) );
  NANDN U1173 ( .A(y[56]), .B(x[56]), .Z(n974) );
  NANDN U1174 ( .A(y[55]), .B(x[55]), .Z(n973) );
  NAND U1175 ( .A(n974), .B(n973), .Z(n2146) );
  ANDN U1176 ( .B(n2214), .A(n2146), .Z(n975) );
  AND U1177 ( .A(n976), .B(n975), .Z(n988) );
  NANDN U1178 ( .A(y[44]), .B(x[44]), .Z(n978) );
  NANDN U1179 ( .A(y[43]), .B(x[43]), .Z(n977) );
  AND U1180 ( .A(n978), .B(n977), .Z(n2200) );
  NANDN U1181 ( .A(y[28]), .B(x[28]), .Z(n980) );
  NANDN U1182 ( .A(y[27]), .B(x[27]), .Z(n979) );
  NAND U1183 ( .A(n980), .B(n979), .Z(n2154) );
  ANDN U1184 ( .B(n2200), .A(n2154), .Z(n986) );
  NANDN U1185 ( .A(x[33]), .B(y[33]), .Z(n982) );
  NANDN U1186 ( .A(x[32]), .B(y[32]), .Z(n981) );
  AND U1187 ( .A(n982), .B(n981), .Z(n2191) );
  NANDN U1188 ( .A(y[32]), .B(x[32]), .Z(n984) );
  NANDN U1189 ( .A(y[31]), .B(x[31]), .Z(n983) );
  NAND U1190 ( .A(n984), .B(n983), .Z(n2153) );
  ANDN U1191 ( .B(n2191), .A(n2153), .Z(n985) );
  AND U1192 ( .A(n986), .B(n985), .Z(n987) );
  AND U1193 ( .A(n988), .B(n987), .Z(n989) );
  AND U1194 ( .A(n990), .B(n989), .Z(n991) );
  AND U1195 ( .A(n992), .B(n991), .Z(n1088) );
  NANDN U1196 ( .A(x[125]), .B(y[125]), .Z(n994) );
  NANDN U1197 ( .A(x[124]), .B(y[124]), .Z(n993) );
  AND U1198 ( .A(n994), .B(n993), .Z(n2263) );
  NANDN U1199 ( .A(y[118]), .B(x[118]), .Z(n996) );
  NANDN U1200 ( .A(y[117]), .B(x[117]), .Z(n995) );
  NAND U1201 ( .A(n996), .B(n995), .Z(n2125) );
  ANDN U1202 ( .B(n2263), .A(n2125), .Z(n1002) );
  NANDN U1203 ( .A(x[119]), .B(y[119]), .Z(n998) );
  NANDN U1204 ( .A(x[118]), .B(y[118]), .Z(n997) );
  AND U1205 ( .A(n998), .B(n997), .Z(n2258) );
  NANDN U1206 ( .A(y[120]), .B(x[120]), .Z(n1000) );
  NANDN U1207 ( .A(y[119]), .B(x[119]), .Z(n999) );
  NAND U1208 ( .A(n1000), .B(n999), .Z(n2259) );
  ANDN U1209 ( .B(n2258), .A(n2259), .Z(n1001) );
  AND U1210 ( .A(n1002), .B(n1001), .Z(n1014) );
  NANDN U1211 ( .A(x[117]), .B(y[117]), .Z(n1004) );
  NANDN U1212 ( .A(x[116]), .B(y[116]), .Z(n1003) );
  AND U1213 ( .A(n1004), .B(n1003), .Z(n2257) );
  NANDN U1214 ( .A(y[116]), .B(x[116]), .Z(n1006) );
  NANDN U1215 ( .A(y[115]), .B(x[115]), .Z(n1005) );
  NAND U1216 ( .A(n1006), .B(n1005), .Z(n2126) );
  ANDN U1217 ( .B(n2257), .A(n2126), .Z(n1012) );
  NANDN U1218 ( .A(x[111]), .B(y[111]), .Z(n1008) );
  NANDN U1219 ( .A(x[110]), .B(y[110]), .Z(n1007) );
  AND U1220 ( .A(n1008), .B(n1007), .Z(n2251) );
  NANDN U1221 ( .A(y[112]), .B(x[112]), .Z(n1010) );
  NANDN U1222 ( .A(y[111]), .B(x[111]), .Z(n1009) );
  NAND U1223 ( .A(n1010), .B(n1009), .Z(n2252) );
  ANDN U1224 ( .B(n2251), .A(n2252), .Z(n1011) );
  AND U1225 ( .A(n1012), .B(n1011), .Z(n1013) );
  AND U1226 ( .A(n1014), .B(n1013), .Z(n1038) );
  NANDN U1227 ( .A(y[128]), .B(x[128]), .Z(n1016) );
  NANDN U1228 ( .A(y[127]), .B(x[127]), .Z(n1015) );
  AND U1229 ( .A(n1016), .B(n1015), .Z(n2266) );
  NANDN U1230 ( .A(y[126]), .B(x[126]), .Z(n1018) );
  NANDN U1231 ( .A(y[125]), .B(x[125]), .Z(n1017) );
  NAND U1232 ( .A(n1018), .B(n1017), .Z(n2264) );
  ANDN U1233 ( .B(n2266), .A(n2264), .Z(n1024) );
  NANDN U1234 ( .A(x[127]), .B(y[127]), .Z(n1020) );
  NANDN U1235 ( .A(x[126]), .B(y[126]), .Z(n1019) );
  AND U1236 ( .A(n1020), .B(n1019), .Z(n2265) );
  NANDN U1237 ( .A(x[129]), .B(y[129]), .Z(n1022) );
  NANDN U1238 ( .A(x[128]), .B(y[128]), .Z(n1021) );
  AND U1239 ( .A(n1022), .B(n1021), .Z(n2267) );
  AND U1240 ( .A(n2265), .B(n2267), .Z(n1023) );
  AND U1241 ( .A(n1024), .B(n1023), .Z(n1036) );
  NANDN U1242 ( .A(x[101]), .B(y[101]), .Z(n1026) );
  NANDN U1243 ( .A(x[100]), .B(y[100]), .Z(n1025) );
  AND U1244 ( .A(n1026), .B(n1025), .Z(n2244) );
  NANDN U1245 ( .A(y[110]), .B(x[110]), .Z(n1028) );
  NANDN U1246 ( .A(y[109]), .B(x[109]), .Z(n1027) );
  NAND U1247 ( .A(n1028), .B(n1027), .Z(n2128) );
  ANDN U1248 ( .B(n2244), .A(n2128), .Z(n1034) );
  NANDN U1249 ( .A(x[109]), .B(y[109]), .Z(n1030) );
  NANDN U1250 ( .A(x[108]), .B(y[108]), .Z(n1029) );
  AND U1251 ( .A(n1030), .B(n1029), .Z(n2250) );
  NANDN U1252 ( .A(y[102]), .B(x[102]), .Z(n1032) );
  NANDN U1253 ( .A(y[101]), .B(x[101]), .Z(n1031) );
  NAND U1254 ( .A(n1032), .B(n1031), .Z(n2130) );
  ANDN U1255 ( .B(n2250), .A(n2130), .Z(n1033) );
  AND U1256 ( .A(n1034), .B(n1033), .Z(n1035) );
  AND U1257 ( .A(n1036), .B(n1035), .Z(n1037) );
  AND U1258 ( .A(n1038), .B(n1037), .Z(n1086) );
  NANDN U1259 ( .A(x[7]), .B(y[7]), .Z(n1040) );
  NANDN U1260 ( .A(x[6]), .B(y[6]), .Z(n1039) );
  AND U1261 ( .A(n1040), .B(n1039), .Z(n2170) );
  NANDN U1262 ( .A(y[12]), .B(x[12]), .Z(n1042) );
  NANDN U1263 ( .A(y[11]), .B(x[11]), .Z(n1041) );
  NAND U1264 ( .A(n1042), .B(n1041), .Z(n2173) );
  ANDN U1265 ( .B(n2170), .A(n2173), .Z(n1048) );
  NANDN U1266 ( .A(x[5]), .B(y[5]), .Z(n1044) );
  NANDN U1267 ( .A(x[4]), .B(y[4]), .Z(n1043) );
  AND U1268 ( .A(n1044), .B(n1043), .Z(n2168) );
  NANDN U1269 ( .A(y[8]), .B(x[8]), .Z(n1046) );
  NANDN U1270 ( .A(y[7]), .B(x[7]), .Z(n1045) );
  NAND U1271 ( .A(n1046), .B(n1045), .Z(n2160) );
  ANDN U1272 ( .B(n2168), .A(n2160), .Z(n1047) );
  AND U1273 ( .A(n1048), .B(n1047), .Z(n1060) );
  NANDN U1274 ( .A(x[131]), .B(y[131]), .Z(n1050) );
  NANDN U1275 ( .A(x[130]), .B(y[130]), .Z(n1049) );
  AND U1276 ( .A(n1050), .B(n1049), .Z(n2268) );
  NANDN U1277 ( .A(y[42]), .B(x[42]), .Z(n1052) );
  NANDN U1278 ( .A(y[41]), .B(x[41]), .Z(n1051) );
  NAND U1279 ( .A(n1052), .B(n1051), .Z(n2197) );
  ANDN U1280 ( .B(n2268), .A(n2197), .Z(n1058) );
  NANDN U1281 ( .A(x[91]), .B(y[91]), .Z(n1054) );
  NANDN U1282 ( .A(x[90]), .B(y[90]), .Z(n1053) );
  AND U1283 ( .A(n1054), .B(n1053), .Z(n2236) );
  NANDN U1284 ( .A(y[80]), .B(x[80]), .Z(n1056) );
  NANDN U1285 ( .A(y[79]), .B(x[79]), .Z(n1055) );
  NAND U1286 ( .A(n1056), .B(n1055), .Z(n2136) );
  ANDN U1287 ( .B(n2236), .A(n2136), .Z(n1057) );
  AND U1288 ( .A(n1058), .B(n1057), .Z(n1059) );
  AND U1289 ( .A(n1060), .B(n1059), .Z(n1084) );
  NANDN U1290 ( .A(x[9]), .B(y[9]), .Z(n1062) );
  NANDN U1291 ( .A(x[8]), .B(y[8]), .Z(n1061) );
  AND U1292 ( .A(n1062), .B(n1061), .Z(n2171) );
  NANDN U1293 ( .A(y[20]), .B(x[20]), .Z(n1064) );
  NANDN U1294 ( .A(y[19]), .B(x[19]), .Z(n1063) );
  NAND U1295 ( .A(n1064), .B(n1063), .Z(n2157) );
  ANDN U1296 ( .B(n2171), .A(n2157), .Z(n1070) );
  NANDN U1297 ( .A(x[29]), .B(y[29]), .Z(n1066) );
  NANDN U1298 ( .A(x[28]), .B(y[28]), .Z(n1065) );
  AND U1299 ( .A(n1066), .B(n1065), .Z(n2187) );
  NANDN U1300 ( .A(y[10]), .B(x[10]), .Z(n1068) );
  NANDN U1301 ( .A(y[9]), .B(x[9]), .Z(n1067) );
  NAND U1302 ( .A(n1068), .B(n1067), .Z(n2159) );
  ANDN U1303 ( .B(n2187), .A(n2159), .Z(n1069) );
  AND U1304 ( .A(n1070), .B(n1069), .Z(n1082) );
  NANDN U1305 ( .A(x[151]), .B(y[151]), .Z(n1072) );
  NANDN U1306 ( .A(x[150]), .B(y[150]), .Z(n1071) );
  AND U1307 ( .A(n1072), .B(n1071), .Z(n2285) );
  NANDN U1308 ( .A(x[217]), .B(y[217]), .Z(n1074) );
  NANDN U1309 ( .A(x[216]), .B(y[216]), .Z(n1073) );
  AND U1310 ( .A(n1074), .B(n1073), .Z(n2343) );
  AND U1311 ( .A(n2285), .B(n2343), .Z(n1080) );
  NANDN U1312 ( .A(y[140]), .B(x[140]), .Z(n1076) );
  NANDN U1313 ( .A(y[139]), .B(x[139]), .Z(n1075) );
  AND U1314 ( .A(n1076), .B(n1075), .Z(n2276) );
  NANDN U1315 ( .A(y[166]), .B(x[166]), .Z(n1078) );
  NANDN U1316 ( .A(y[165]), .B(x[165]), .Z(n1077) );
  NAND U1317 ( .A(n1078), .B(n1077), .Z(n2114) );
  ANDN U1318 ( .B(n2276), .A(n2114), .Z(n1079) );
  AND U1319 ( .A(n1080), .B(n1079), .Z(n1081) );
  AND U1320 ( .A(n1082), .B(n1081), .Z(n1083) );
  AND U1321 ( .A(n1084), .B(n1083), .Z(n1085) );
  AND U1322 ( .A(n1086), .B(n1085), .Z(n1087) );
  AND U1323 ( .A(n1088), .B(n1087), .Z(n1280) );
  NANDN U1324 ( .A(x[489]), .B(y[489]), .Z(n1090) );
  NANDN U1325 ( .A(x[488]), .B(y[488]), .Z(n1089) );
  AND U1326 ( .A(n1090), .B(n1089), .Z(n2591) );
  NANDN U1327 ( .A(y[484]), .B(x[484]), .Z(n1092) );
  NANDN U1328 ( .A(y[483]), .B(x[483]), .Z(n1091) );
  NAND U1329 ( .A(n1092), .B(n1091), .Z(n2028) );
  ANDN U1330 ( .B(n2591), .A(n2028), .Z(n1098) );
  NANDN U1331 ( .A(x[485]), .B(y[485]), .Z(n1094) );
  NANDN U1332 ( .A(x[484]), .B(y[484]), .Z(n1093) );
  AND U1333 ( .A(n1094), .B(n1093), .Z(n2586) );
  NANDN U1334 ( .A(y[488]), .B(x[488]), .Z(n1096) );
  NANDN U1335 ( .A(y[487]), .B(x[487]), .Z(n1095) );
  NAND U1336 ( .A(n1096), .B(n1095), .Z(n2589) );
  ANDN U1337 ( .B(n2586), .A(n2589), .Z(n1097) );
  AND U1338 ( .A(n1098), .B(n1097), .Z(n1110) );
  NANDN U1339 ( .A(x[483]), .B(y[483]), .Z(n1100) );
  NANDN U1340 ( .A(x[482]), .B(y[482]), .Z(n1099) );
  AND U1341 ( .A(n1100), .B(n1099), .Z(n2585) );
  NANDN U1342 ( .A(x[473]), .B(y[473]), .Z(n1102) );
  NANDN U1343 ( .A(x[472]), .B(y[472]), .Z(n1101) );
  AND U1344 ( .A(n1102), .B(n1101), .Z(n2576) );
  AND U1345 ( .A(n2585), .B(n2576), .Z(n1108) );
  NANDN U1346 ( .A(x[481]), .B(y[481]), .Z(n1104) );
  NANDN U1347 ( .A(x[480]), .B(y[480]), .Z(n1103) );
  AND U1348 ( .A(n1104), .B(n1103), .Z(n2583) );
  NANDN U1349 ( .A(x[475]), .B(y[475]), .Z(n1106) );
  NANDN U1350 ( .A(x[474]), .B(y[474]), .Z(n1105) );
  AND U1351 ( .A(n1106), .B(n1105), .Z(n2578) );
  AND U1352 ( .A(n2583), .B(n2578), .Z(n1107) );
  AND U1353 ( .A(n1108), .B(n1107), .Z(n1109) );
  AND U1354 ( .A(n1110), .B(n1109), .Z(n1134) );
  NANDN U1355 ( .A(x[497]), .B(y[497]), .Z(n1112) );
  NANDN U1356 ( .A(x[496]), .B(y[496]), .Z(n1111) );
  AND U1357 ( .A(n1112), .B(n1111), .Z(n2597) );
  NANDN U1358 ( .A(x[493]), .B(y[493]), .Z(n1114) );
  NANDN U1359 ( .A(x[492]), .B(y[492]), .Z(n1113) );
  AND U1360 ( .A(n1114), .B(n1113), .Z(n2594) );
  AND U1361 ( .A(n2597), .B(n2594), .Z(n1120) );
  NANDN U1362 ( .A(x[495]), .B(y[495]), .Z(n1116) );
  NANDN U1363 ( .A(x[494]), .B(y[494]), .Z(n1115) );
  AND U1364 ( .A(n1116), .B(n1115), .Z(n2596) );
  NANDN U1365 ( .A(y[496]), .B(x[496]), .Z(n1118) );
  NANDN U1366 ( .A(y[495]), .B(x[495]), .Z(n1117) );
  NAND U1367 ( .A(n1118), .B(n1117), .Z(n2025) );
  ANDN U1368 ( .B(n2596), .A(n2025), .Z(n1119) );
  AND U1369 ( .A(n1120), .B(n1119), .Z(n1132) );
  NANDN U1370 ( .A(x[471]), .B(y[471]), .Z(n1122) );
  NANDN U1371 ( .A(x[470]), .B(y[470]), .Z(n1121) );
  AND U1372 ( .A(n1122), .B(n1121), .Z(n2574) );
  NANDN U1373 ( .A(x[463]), .B(y[463]), .Z(n1124) );
  NANDN U1374 ( .A(x[462]), .B(y[462]), .Z(n1123) );
  AND U1375 ( .A(n1124), .B(n1123), .Z(n2567) );
  AND U1376 ( .A(n2574), .B(n2567), .Z(n1130) );
  NANDN U1377 ( .A(x[467]), .B(y[467]), .Z(n1126) );
  NANDN U1378 ( .A(x[466]), .B(y[466]), .Z(n1125) );
  AND U1379 ( .A(n1126), .B(n1125), .Z(n2571) );
  NANDN U1380 ( .A(x[465]), .B(y[465]), .Z(n1128) );
  NANDN U1381 ( .A(x[464]), .B(y[464]), .Z(n1127) );
  AND U1382 ( .A(n1128), .B(n1127), .Z(n2569) );
  AND U1383 ( .A(n2571), .B(n2569), .Z(n1129) );
  AND U1384 ( .A(n1130), .B(n1129), .Z(n1131) );
  AND U1385 ( .A(n1132), .B(n1131), .Z(n1133) );
  AND U1386 ( .A(n1134), .B(n1133), .Z(n1182) );
  NANDN U1387 ( .A(x[441]), .B(y[441]), .Z(n1136) );
  NANDN U1388 ( .A(x[440]), .B(y[440]), .Z(n1135) );
  AND U1389 ( .A(n1136), .B(n1135), .Z(n2547) );
  NANDN U1390 ( .A(y[452]), .B(x[452]), .Z(n1138) );
  NANDN U1391 ( .A(y[451]), .B(x[451]), .Z(n1137) );
  NAND U1392 ( .A(n1138), .B(n1137), .Z(n2035) );
  ANDN U1393 ( .B(n2547), .A(n2035), .Z(n1144) );
  NANDN U1394 ( .A(x[451]), .B(y[451]), .Z(n1140) );
  NANDN U1395 ( .A(x[450]), .B(y[450]), .Z(n1139) );
  AND U1396 ( .A(n1140), .B(n1139), .Z(n2557) );
  NANDN U1397 ( .A(x[445]), .B(y[445]), .Z(n1142) );
  NANDN U1398 ( .A(x[444]), .B(y[444]), .Z(n1141) );
  AND U1399 ( .A(n1142), .B(n1141), .Z(n2552) );
  AND U1400 ( .A(n2557), .B(n2552), .Z(n1143) );
  AND U1401 ( .A(n1144), .B(n1143), .Z(n1156) );
  NANDN U1402 ( .A(x[437]), .B(y[437]), .Z(n1146) );
  NANDN U1403 ( .A(x[436]), .B(y[436]), .Z(n1145) );
  AND U1404 ( .A(n1146), .B(n1145), .Z(n2544) );
  NANDN U1405 ( .A(y[440]), .B(x[440]), .Z(n1148) );
  NANDN U1406 ( .A(y[439]), .B(x[439]), .Z(n1147) );
  NAND U1407 ( .A(n1148), .B(n1147), .Z(n2038) );
  ANDN U1408 ( .B(n2544), .A(n2038), .Z(n1154) );
  NANDN U1409 ( .A(x[443]), .B(y[443]), .Z(n1150) );
  NANDN U1410 ( .A(x[442]), .B(y[442]), .Z(n1149) );
  AND U1411 ( .A(n1150), .B(n1149), .Z(n2548) );
  NANDN U1412 ( .A(x[439]), .B(y[439]), .Z(n1152) );
  NANDN U1413 ( .A(x[438]), .B(y[438]), .Z(n1151) );
  AND U1414 ( .A(n1152), .B(n1151), .Z(n2546) );
  AND U1415 ( .A(n2548), .B(n2546), .Z(n1153) );
  AND U1416 ( .A(n1154), .B(n1153), .Z(n1155) );
  AND U1417 ( .A(n1156), .B(n1155), .Z(n1180) );
  NANDN U1418 ( .A(x[457]), .B(y[457]), .Z(n1158) );
  NANDN U1419 ( .A(x[456]), .B(y[456]), .Z(n1157) );
  AND U1420 ( .A(n1158), .B(n1157), .Z(n2561) );
  NANDN U1421 ( .A(x[453]), .B(y[453]), .Z(n1160) );
  NANDN U1422 ( .A(x[452]), .B(y[452]), .Z(n1159) );
  AND U1423 ( .A(n1160), .B(n1159), .Z(n2558) );
  AND U1424 ( .A(n2561), .B(n2558), .Z(n1166) );
  NANDN U1425 ( .A(x[455]), .B(y[455]), .Z(n1162) );
  NANDN U1426 ( .A(x[454]), .B(y[454]), .Z(n1161) );
  AND U1427 ( .A(n1162), .B(n1161), .Z(n2559) );
  NANDN U1428 ( .A(y[454]), .B(x[454]), .Z(n1164) );
  NANDN U1429 ( .A(y[453]), .B(x[453]), .Z(n1163) );
  NAND U1430 ( .A(n1164), .B(n1163), .Z(n2034) );
  ANDN U1431 ( .B(n2559), .A(n2034), .Z(n1165) );
  AND U1432 ( .A(n1166), .B(n1165), .Z(n1178) );
  NANDN U1433 ( .A(y[434]), .B(x[434]), .Z(n1168) );
  NANDN U1434 ( .A(y[433]), .B(x[433]), .Z(n1167) );
  AND U1435 ( .A(n1168), .B(n1167), .Z(n2542) );
  NANDN U1436 ( .A(y[430]), .B(x[430]), .Z(n1170) );
  NANDN U1437 ( .A(y[429]), .B(x[429]), .Z(n1169) );
  NAND U1438 ( .A(n1170), .B(n1169), .Z(n2040) );
  ANDN U1439 ( .B(n2542), .A(n2040), .Z(n1176) );
  NANDN U1440 ( .A(x[431]), .B(y[431]), .Z(n1172) );
  NANDN U1441 ( .A(x[430]), .B(y[430]), .Z(n1171) );
  AND U1442 ( .A(n1172), .B(n1171), .Z(n2539) );
  NANDN U1443 ( .A(y[432]), .B(x[432]), .Z(n1174) );
  NANDN U1444 ( .A(y[431]), .B(x[431]), .Z(n1173) );
  NAND U1445 ( .A(n1174), .B(n1173), .Z(n2540) );
  ANDN U1446 ( .B(n2539), .A(n2540), .Z(n1175) );
  AND U1447 ( .A(n1176), .B(n1175), .Z(n1177) );
  AND U1448 ( .A(n1178), .B(n1177), .Z(n1179) );
  AND U1449 ( .A(n1180), .B(n1179), .Z(n1181) );
  AND U1450 ( .A(n1182), .B(n1181), .Z(n1278) );
  NANDN U1451 ( .A(x[387]), .B(y[387]), .Z(n1184) );
  NANDN U1452 ( .A(x[386]), .B(y[386]), .Z(n1183) );
  AND U1453 ( .A(n1184), .B(n1183), .Z(n2502) );
  NANDN U1454 ( .A(y[482]), .B(x[482]), .Z(n1186) );
  NANDN U1455 ( .A(y[481]), .B(x[481]), .Z(n1185) );
  NAND U1456 ( .A(n1186), .B(n1185), .Z(n2584) );
  ANDN U1457 ( .B(n2502), .A(n2584), .Z(n1192) );
  NANDN U1458 ( .A(x[429]), .B(y[429]), .Z(n1188) );
  NANDN U1459 ( .A(x[428]), .B(y[428]), .Z(n1187) );
  AND U1460 ( .A(n1188), .B(n1187), .Z(n2537) );
  NANDN U1461 ( .A(y[444]), .B(x[444]), .Z(n1190) );
  NANDN U1462 ( .A(y[443]), .B(x[443]), .Z(n1189) );
  NAND U1463 ( .A(n1190), .B(n1189), .Z(n2549) );
  ANDN U1464 ( .B(n2537), .A(n2549), .Z(n1191) );
  AND U1465 ( .A(n1192), .B(n1191), .Z(n1204) );
  NANDN U1466 ( .A(x[507]), .B(y[507]), .Z(n1194) );
  NANDN U1467 ( .A(x[506]), .B(y[506]), .Z(n1193) );
  AND U1468 ( .A(n1194), .B(n1193), .Z(n2606) );
  NANDN U1469 ( .A(y[494]), .B(x[494]), .Z(n1196) );
  NANDN U1470 ( .A(y[493]), .B(x[493]), .Z(n1195) );
  NAND U1471 ( .A(n1196), .B(n1195), .Z(n2595) );
  ANDN U1472 ( .B(n2606), .A(n2595), .Z(n1202) );
  NANDN U1473 ( .A(x[509]), .B(y[509]), .Z(n1198) );
  NANDN U1474 ( .A(x[508]), .B(y[508]), .Z(n1197) );
  AND U1475 ( .A(n1198), .B(n1197), .Z(n2608) );
  NANDN U1476 ( .A(y[510]), .B(x[510]), .Z(n1200) );
  NANDN U1477 ( .A(y[509]), .B(x[509]), .Z(n1199) );
  NAND U1478 ( .A(n1200), .B(n1199), .Z(n2021) );
  ANDN U1479 ( .B(n2608), .A(n2021), .Z(n1201) );
  AND U1480 ( .A(n1202), .B(n1201), .Z(n1203) );
  AND U1481 ( .A(n1204), .B(n1203), .Z(n1228) );
  NANDN U1482 ( .A(x[350]), .B(y[350]), .Z(n1206) );
  NANDN U1483 ( .A(x[349]), .B(y[349]), .Z(n1205) );
  AND U1484 ( .A(n1206), .B(n1205), .Z(n2469) );
  NANDN U1485 ( .A(y[236]), .B(x[236]), .Z(n1208) );
  NANDN U1486 ( .A(y[235]), .B(x[235]), .Z(n1207) );
  NAND U1487 ( .A(n1208), .B(n1207), .Z(n2096) );
  ANDN U1488 ( .B(n2469), .A(n2096), .Z(n1214) );
  NANDN U1489 ( .A(y[318]), .B(x[318]), .Z(n1210) );
  NANDN U1490 ( .A(y[317]), .B(x[317]), .Z(n1209) );
  AND U1491 ( .A(n1210), .B(n1209), .Z(n2442) );
  NANDN U1492 ( .A(y[339]), .B(x[339]), .Z(n1212) );
  NANDN U1493 ( .A(y[338]), .B(x[338]), .Z(n1211) );
  NAND U1494 ( .A(n1212), .B(n1211), .Z(n2067) );
  ANDN U1495 ( .B(n2442), .A(n2067), .Z(n1213) );
  AND U1496 ( .A(n1214), .B(n1213), .Z(n1226) );
  NANDN U1497 ( .A(y[506]), .B(x[506]), .Z(n1216) );
  NANDN U1498 ( .A(y[505]), .B(x[505]), .Z(n1215) );
  AND U1499 ( .A(n1216), .B(n1215), .Z(n2605) );
  NANDN U1500 ( .A(y[500]), .B(x[500]), .Z(n1218) );
  NANDN U1501 ( .A(y[499]), .B(x[499]), .Z(n1217) );
  NAND U1502 ( .A(n1218), .B(n1217), .Z(n2599) );
  ANDN U1503 ( .B(n2605), .A(n2599), .Z(n1224) );
  NANDN U1504 ( .A(x[501]), .B(y[501]), .Z(n1220) );
  NANDN U1505 ( .A(x[500]), .B(y[500]), .Z(n1219) );
  AND U1506 ( .A(n1220), .B(n1219), .Z(n2600) );
  NANDN U1507 ( .A(y[504]), .B(x[504]), .Z(n1222) );
  NANDN U1508 ( .A(y[503]), .B(x[503]), .Z(n1221) );
  NAND U1509 ( .A(n1222), .B(n1221), .Z(n2022) );
  ANDN U1510 ( .B(n2600), .A(n2022), .Z(n1223) );
  AND U1511 ( .A(n1224), .B(n1223), .Z(n1225) );
  AND U1512 ( .A(n1226), .B(n1225), .Z(n1227) );
  AND U1513 ( .A(n1228), .B(n1227), .Z(n1276) );
  NANDN U1514 ( .A(x[409]), .B(y[409]), .Z(n1230) );
  NANDN U1515 ( .A(x[408]), .B(y[408]), .Z(n1229) );
  AND U1516 ( .A(n1230), .B(n1229), .Z(n2519) );
  NANDN U1517 ( .A(y[418]), .B(x[418]), .Z(n1232) );
  NANDN U1518 ( .A(y[417]), .B(x[417]), .Z(n1231) );
  NAND U1519 ( .A(n1232), .B(n1231), .Z(n2528) );
  ANDN U1520 ( .B(n2519), .A(n2528), .Z(n1238) );
  NANDN U1521 ( .A(x[411]), .B(y[411]), .Z(n1234) );
  NANDN U1522 ( .A(x[410]), .B(y[410]), .Z(n1233) );
  AND U1523 ( .A(n1234), .B(n1233), .Z(n2522) );
  NANDN U1524 ( .A(y[414]), .B(x[414]), .Z(n1236) );
  NANDN U1525 ( .A(y[413]), .B(x[413]), .Z(n1235) );
  NAND U1526 ( .A(n1236), .B(n1235), .Z(n2045) );
  ANDN U1527 ( .B(n2522), .A(n2045), .Z(n1237) );
  AND U1528 ( .A(n1238), .B(n1237), .Z(n1250) );
  NANDN U1529 ( .A(x[401]), .B(y[401]), .Z(n1240) );
  NANDN U1530 ( .A(x[400]), .B(y[400]), .Z(n1239) );
  AND U1531 ( .A(n1240), .B(n1239), .Z(n2513) );
  NANDN U1532 ( .A(y[408]), .B(x[408]), .Z(n1242) );
  NANDN U1533 ( .A(y[407]), .B(x[407]), .Z(n1241) );
  NAND U1534 ( .A(n1242), .B(n1241), .Z(n2046) );
  ANDN U1535 ( .B(n2513), .A(n2046), .Z(n1248) );
  NANDN U1536 ( .A(x[407]), .B(y[407]), .Z(n1244) );
  NANDN U1537 ( .A(x[406]), .B(y[406]), .Z(n1243) );
  AND U1538 ( .A(n1244), .B(n1243), .Z(n2518) );
  NANDN U1539 ( .A(y[402]), .B(x[402]), .Z(n1246) );
  NANDN U1540 ( .A(y[401]), .B(x[401]), .Z(n1245) );
  NAND U1541 ( .A(n1246), .B(n1245), .Z(n2048) );
  ANDN U1542 ( .B(n2518), .A(n2048), .Z(n1247) );
  AND U1543 ( .A(n1248), .B(n1247), .Z(n1249) );
  AND U1544 ( .A(n1250), .B(n1249), .Z(n1274) );
  NANDN U1545 ( .A(y[428]), .B(x[428]), .Z(n1252) );
  NANDN U1546 ( .A(y[427]), .B(x[427]), .Z(n1251) );
  AND U1547 ( .A(n1252), .B(n1251), .Z(n2536) );
  NANDN U1548 ( .A(y[420]), .B(x[420]), .Z(n1254) );
  NANDN U1549 ( .A(y[419]), .B(x[419]), .Z(n1253) );
  NAND U1550 ( .A(n1254), .B(n1253), .Z(n2529) );
  ANDN U1551 ( .B(n2536), .A(n2529), .Z(n1260) );
  NANDN U1552 ( .A(x[423]), .B(y[423]), .Z(n1256) );
  NANDN U1553 ( .A(x[422]), .B(y[422]), .Z(n1255) );
  AND U1554 ( .A(n1256), .B(n1255), .Z(n2532) );
  NANDN U1555 ( .A(y[424]), .B(x[424]), .Z(n1258) );
  NANDN U1556 ( .A(y[423]), .B(x[423]), .Z(n1257) );
  NAND U1557 ( .A(n1258), .B(n1257), .Z(n2041) );
  ANDN U1558 ( .B(n2532), .A(n2041), .Z(n1259) );
  AND U1559 ( .A(n1260), .B(n1259), .Z(n1272) );
  NANDN U1560 ( .A(x[399]), .B(y[399]), .Z(n1262) );
  NANDN U1561 ( .A(x[398]), .B(y[398]), .Z(n1261) );
  AND U1562 ( .A(n1262), .B(n1261), .Z(n2512) );
  NANDN U1563 ( .A(y[394]), .B(x[394]), .Z(n1264) );
  NANDN U1564 ( .A(y[393]), .B(x[393]), .Z(n1263) );
  NAND U1565 ( .A(n1264), .B(n1263), .Z(n2051) );
  ANDN U1566 ( .B(n2512), .A(n2051), .Z(n1270) );
  NANDN U1567 ( .A(x[397]), .B(y[397]), .Z(n1266) );
  NANDN U1568 ( .A(x[396]), .B(y[396]), .Z(n1265) );
  AND U1569 ( .A(n1266), .B(n1265), .Z(n2510) );
  NANDN U1570 ( .A(x[395]), .B(y[395]), .Z(n1268) );
  NANDN U1571 ( .A(x[394]), .B(y[394]), .Z(n1267) );
  AND U1572 ( .A(n1268), .B(n1267), .Z(n2509) );
  AND U1573 ( .A(n2510), .B(n2509), .Z(n1269) );
  AND U1574 ( .A(n1270), .B(n1269), .Z(n1271) );
  AND U1575 ( .A(n1272), .B(n1271), .Z(n1273) );
  AND U1576 ( .A(n1274), .B(n1273), .Z(n1275) );
  AND U1577 ( .A(n1276), .B(n1275), .Z(n1277) );
  AND U1578 ( .A(n1278), .B(n1277), .Z(n1279) );
  AND U1579 ( .A(n1280), .B(n1279), .Z(n1664) );
  NANDN U1580 ( .A(y[240]), .B(x[240]), .Z(n1282) );
  NANDN U1581 ( .A(y[239]), .B(x[239]), .Z(n1281) );
  AND U1582 ( .A(n1282), .B(n1281), .Z(n2362) );
  NANDN U1583 ( .A(y[238]), .B(x[238]), .Z(n1284) );
  NANDN U1584 ( .A(y[237]), .B(x[237]), .Z(n1283) );
  NAND U1585 ( .A(n1284), .B(n1283), .Z(n2360) );
  ANDN U1586 ( .B(n2362), .A(n2360), .Z(n1290) );
  NANDN U1587 ( .A(x[239]), .B(y[239]), .Z(n1286) );
  NANDN U1588 ( .A(x[238]), .B(y[238]), .Z(n1285) );
  AND U1589 ( .A(n1286), .B(n1285), .Z(n2361) );
  NANDN U1590 ( .A(y[242]), .B(x[242]), .Z(n1288) );
  NANDN U1591 ( .A(y[241]), .B(x[241]), .Z(n1287) );
  NAND U1592 ( .A(n1288), .B(n1287), .Z(n2095) );
  ANDN U1593 ( .B(n2361), .A(n2095), .Z(n1289) );
  AND U1594 ( .A(n1290), .B(n1289), .Z(n1302) );
  NANDN U1595 ( .A(y[234]), .B(x[234]), .Z(n1292) );
  NANDN U1596 ( .A(y[233]), .B(x[233]), .Z(n1291) );
  AND U1597 ( .A(n1292), .B(n1291), .Z(n2357) );
  NANDN U1598 ( .A(y[230]), .B(x[230]), .Z(n1294) );
  NANDN U1599 ( .A(y[229]), .B(x[229]), .Z(n1293) );
  NAND U1600 ( .A(n1294), .B(n1293), .Z(n2097) );
  ANDN U1601 ( .B(n2357), .A(n2097), .Z(n1300) );
  NANDN U1602 ( .A(x[229]), .B(y[229]), .Z(n1296) );
  NANDN U1603 ( .A(x[228]), .B(y[228]), .Z(n1295) );
  AND U1604 ( .A(n1296), .B(n1295), .Z(n2353) );
  NANDN U1605 ( .A(x[221]), .B(y[221]), .Z(n1298) );
  NANDN U1606 ( .A(x[220]), .B(y[220]), .Z(n1297) );
  AND U1607 ( .A(n1298), .B(n1297), .Z(n2346) );
  AND U1608 ( .A(n2353), .B(n2346), .Z(n1299) );
  AND U1609 ( .A(n1300), .B(n1299), .Z(n1301) );
  AND U1610 ( .A(n1302), .B(n1301), .Z(n1326) );
  NANDN U1611 ( .A(x[243]), .B(y[243]), .Z(n1304) );
  NANDN U1612 ( .A(x[242]), .B(y[242]), .Z(n1303) );
  AND U1613 ( .A(n1304), .B(n1303), .Z(n2365) );
  NANDN U1614 ( .A(y[248]), .B(x[248]), .Z(n1306) );
  NANDN U1615 ( .A(y[247]), .B(x[247]), .Z(n1305) );
  NAND U1616 ( .A(n1306), .B(n1305), .Z(n2093) );
  ANDN U1617 ( .B(n2365), .A(n2093), .Z(n1312) );
  NANDN U1618 ( .A(x[254]), .B(y[254]), .Z(n1308) );
  NANDN U1619 ( .A(x[253]), .B(y[253]), .Z(n1307) );
  AND U1620 ( .A(n1308), .B(n1307), .Z(n2378) );
  NANDN U1621 ( .A(x[247]), .B(y[247]), .Z(n1310) );
  NANDN U1622 ( .A(x[246]), .B(y[246]), .Z(n1309) );
  AND U1623 ( .A(n1310), .B(n1309), .Z(n2369) );
  AND U1624 ( .A(n2378), .B(n2369), .Z(n1311) );
  AND U1625 ( .A(n1312), .B(n1311), .Z(n1324) );
  NANDN U1626 ( .A(y[220]), .B(x[220]), .Z(n1314) );
  NANDN U1627 ( .A(y[219]), .B(x[219]), .Z(n1313) );
  AND U1628 ( .A(n1314), .B(n1313), .Z(n2345) );
  NANDN U1629 ( .A(y[210]), .B(x[210]), .Z(n1316) );
  NANDN U1630 ( .A(y[209]), .B(x[209]), .Z(n1315) );
  NAND U1631 ( .A(n1316), .B(n1315), .Z(n2103) );
  ANDN U1632 ( .B(n2345), .A(n2103), .Z(n1322) );
  NANDN U1633 ( .A(x[211]), .B(y[211]), .Z(n1318) );
  NANDN U1634 ( .A(x[210]), .B(y[210]), .Z(n1317) );
  AND U1635 ( .A(n1318), .B(n1317), .Z(n2338) );
  NANDN U1636 ( .A(y[214]), .B(x[214]), .Z(n1320) );
  NANDN U1637 ( .A(y[213]), .B(x[213]), .Z(n1319) );
  NAND U1638 ( .A(n1320), .B(n1319), .Z(n2341) );
  ANDN U1639 ( .B(n2338), .A(n2341), .Z(n1321) );
  AND U1640 ( .A(n1322), .B(n1321), .Z(n1323) );
  AND U1641 ( .A(n1324), .B(n1323), .Z(n1325) );
  AND U1642 ( .A(n1326), .B(n1325), .Z(n1374) );
  NANDN U1643 ( .A(x[203]), .B(y[203]), .Z(n1328) );
  NANDN U1644 ( .A(x[202]), .B(y[202]), .Z(n1327) );
  AND U1645 ( .A(n1328), .B(n1327), .Z(n2331) );
  NANDN U1646 ( .A(y[192]), .B(x[192]), .Z(n1330) );
  NANDN U1647 ( .A(y[191]), .B(x[191]), .Z(n1329) );
  NAND U1648 ( .A(n1330), .B(n1329), .Z(n2321) );
  ANDN U1649 ( .B(n2331), .A(n2321), .Z(n1336) );
  NANDN U1650 ( .A(y[200]), .B(x[200]), .Z(n1332) );
  NANDN U1651 ( .A(y[199]), .B(x[199]), .Z(n1331) );
  AND U1652 ( .A(n1332), .B(n1331), .Z(n2329) );
  NANDN U1653 ( .A(y[198]), .B(x[198]), .Z(n1334) );
  NANDN U1654 ( .A(y[197]), .B(x[197]), .Z(n1333) );
  NAND U1655 ( .A(n1334), .B(n1333), .Z(n2106) );
  ANDN U1656 ( .B(n2329), .A(n2106), .Z(n1335) );
  AND U1657 ( .A(n1336), .B(n1335), .Z(n1348) );
  NANDN U1658 ( .A(x[191]), .B(y[191]), .Z(n1338) );
  NANDN U1659 ( .A(x[190]), .B(y[190]), .Z(n1337) );
  AND U1660 ( .A(n1338), .B(n1337), .Z(n2320) );
  NANDN U1661 ( .A(y[180]), .B(x[180]), .Z(n1340) );
  NANDN U1662 ( .A(y[179]), .B(x[179]), .Z(n1339) );
  NAND U1663 ( .A(n1340), .B(n1339), .Z(n2311) );
  ANDN U1664 ( .B(n2320), .A(n2311), .Z(n1346) );
  NANDN U1665 ( .A(x[193]), .B(y[193]), .Z(n1342) );
  NANDN U1666 ( .A(x[192]), .B(y[192]), .Z(n1341) );
  AND U1667 ( .A(n1342), .B(n1341), .Z(n2322) );
  NANDN U1668 ( .A(x[181]), .B(y[181]), .Z(n1344) );
  NANDN U1669 ( .A(x[180]), .B(y[180]), .Z(n1343) );
  AND U1670 ( .A(n1344), .B(n1343), .Z(n2312) );
  AND U1671 ( .A(n2322), .B(n2312), .Z(n1345) );
  AND U1672 ( .A(n1346), .B(n1345), .Z(n1347) );
  AND U1673 ( .A(n1348), .B(n1347), .Z(n1372) );
  NANDN U1674 ( .A(x[209]), .B(y[209]), .Z(n1350) );
  NANDN U1675 ( .A(x[208]), .B(y[208]), .Z(n1349) );
  AND U1676 ( .A(n1350), .B(n1349), .Z(n2337) );
  NANDN U1677 ( .A(x[201]), .B(y[201]), .Z(n1352) );
  NANDN U1678 ( .A(x[200]), .B(y[200]), .Z(n1351) );
  AND U1679 ( .A(n1352), .B(n1351), .Z(n2330) );
  AND U1680 ( .A(n2337), .B(n2330), .Z(n1358) );
  NANDN U1681 ( .A(y[208]), .B(x[208]), .Z(n1354) );
  NANDN U1682 ( .A(y[207]), .B(x[207]), .Z(n1353) );
  AND U1683 ( .A(n1354), .B(n1353), .Z(n2336) );
  NANDN U1684 ( .A(y[202]), .B(x[202]), .Z(n1356) );
  NANDN U1685 ( .A(y[201]), .B(x[201]), .Z(n1355) );
  NAND U1686 ( .A(n1356), .B(n1355), .Z(n2105) );
  ANDN U1687 ( .B(n2336), .A(n2105), .Z(n1357) );
  AND U1688 ( .A(n1358), .B(n1357), .Z(n1370) );
  NANDN U1689 ( .A(x[171]), .B(y[171]), .Z(n1360) );
  NANDN U1690 ( .A(x[170]), .B(y[170]), .Z(n1359) );
  AND U1691 ( .A(n1360), .B(n1359), .Z(n2304) );
  NANDN U1692 ( .A(x[169]), .B(y[169]), .Z(n1362) );
  NANDN U1693 ( .A(x[168]), .B(y[168]), .Z(n1361) );
  AND U1694 ( .A(n1362), .B(n1361), .Z(n2301) );
  AND U1695 ( .A(n2304), .B(n2301), .Z(n1368) );
  NANDN U1696 ( .A(y[170]), .B(x[170]), .Z(n1364) );
  NANDN U1697 ( .A(y[169]), .B(x[169]), .Z(n1363) );
  AND U1698 ( .A(n1364), .B(n1363), .Z(n2302) );
  NANDN U1699 ( .A(y[176]), .B(x[176]), .Z(n1366) );
  NANDN U1700 ( .A(y[175]), .B(x[175]), .Z(n1365) );
  NAND U1701 ( .A(n1366), .B(n1365), .Z(n2112) );
  ANDN U1702 ( .B(n2302), .A(n2112), .Z(n1367) );
  AND U1703 ( .A(n1368), .B(n1367), .Z(n1369) );
  AND U1704 ( .A(n1370), .B(n1369), .Z(n1371) );
  AND U1705 ( .A(n1372), .B(n1371), .Z(n1373) );
  AND U1706 ( .A(n1374), .B(n1373), .Z(n1470) );
  NANDN U1707 ( .A(x[280]), .B(y[280]), .Z(n1376) );
  NANDN U1708 ( .A(x[279]), .B(y[279]), .Z(n1375) );
  AND U1709 ( .A(n1376), .B(n1375), .Z(n2405) );
  NANDN U1710 ( .A(y[290]), .B(x[290]), .Z(n1378) );
  NANDN U1711 ( .A(y[289]), .B(x[289]), .Z(n1377) );
  NAND U1712 ( .A(n1378), .B(n1377), .Z(n2415) );
  ANDN U1713 ( .B(n2405), .A(n2415), .Z(n1384) );
  NANDN U1714 ( .A(x[289]), .B(y[289]), .Z(n1380) );
  NANDN U1715 ( .A(x[288]), .B(y[288]), .Z(n1379) );
  AND U1716 ( .A(n1380), .B(n1379), .Z(n2414) );
  NANDN U1717 ( .A(x[285]), .B(y[285]), .Z(n1382) );
  NANDN U1718 ( .A(x[284]), .B(y[284]), .Z(n1381) );
  AND U1719 ( .A(n1382), .B(n1381), .Z(n2410) );
  AND U1720 ( .A(n2414), .B(n2410), .Z(n1383) );
  AND U1721 ( .A(n1384), .B(n1383), .Z(n1396) );
  NANDN U1722 ( .A(x[270]), .B(y[270]), .Z(n1386) );
  NANDN U1723 ( .A(x[269]), .B(y[269]), .Z(n1385) );
  AND U1724 ( .A(n1386), .B(n1385), .Z(n2398) );
  NANDN U1725 ( .A(y[286]), .B(x[286]), .Z(n1388) );
  NANDN U1726 ( .A(y[285]), .B(x[285]), .Z(n1387) );
  NAND U1727 ( .A(n1388), .B(n1387), .Z(n2411) );
  ANDN U1728 ( .B(n2398), .A(n2411), .Z(n1394) );
  NANDN U1729 ( .A(x[272]), .B(y[272]), .Z(n1390) );
  NANDN U1730 ( .A(x[271]), .B(y[271]), .Z(n1389) );
  AND U1731 ( .A(n1390), .B(n1389), .Z(n2399) );
  NANDN U1732 ( .A(y[271]), .B(x[271]), .Z(n1392) );
  NANDN U1733 ( .A(y[270]), .B(x[270]), .Z(n1391) );
  NAND U1734 ( .A(n1392), .B(n1391), .Z(n2088) );
  ANDN U1735 ( .B(n2399), .A(n2088), .Z(n1393) );
  AND U1736 ( .A(n1394), .B(n1393), .Z(n1395) );
  AND U1737 ( .A(n1396), .B(n1395), .Z(n1420) );
  NANDN U1738 ( .A(x[299]), .B(y[299]), .Z(n1398) );
  NANDN U1739 ( .A(x[298]), .B(y[298]), .Z(n1397) );
  AND U1740 ( .A(n1398), .B(n1397), .Z(n2423) );
  NANDN U1741 ( .A(y[300]), .B(x[300]), .Z(n1400) );
  NANDN U1742 ( .A(y[299]), .B(x[299]), .Z(n1399) );
  NAND U1743 ( .A(n1400), .B(n1399), .Z(n2424) );
  ANDN U1744 ( .B(n2423), .A(n2424), .Z(n1406) );
  NANDN U1745 ( .A(x[297]), .B(y[297]), .Z(n1402) );
  NANDN U1746 ( .A(x[296]), .B(y[296]), .Z(n1401) );
  AND U1747 ( .A(n1402), .B(n1401), .Z(n2422) );
  NANDN U1748 ( .A(y[298]), .B(x[298]), .Z(n1404) );
  NANDN U1749 ( .A(y[297]), .B(x[297]), .Z(n1403) );
  NAND U1750 ( .A(n1404), .B(n1403), .Z(n2078) );
  ANDN U1751 ( .B(n2422), .A(n2078), .Z(n1405) );
  AND U1752 ( .A(n1406), .B(n1405), .Z(n1418) );
  NANDN U1753 ( .A(y[267]), .B(x[267]), .Z(n1408) );
  NANDN U1754 ( .A(y[266]), .B(x[266]), .Z(n1407) );
  AND U1755 ( .A(n1408), .B(n1407), .Z(n2395) );
  NANDN U1756 ( .A(y[250]), .B(x[250]), .Z(n1410) );
  NANDN U1757 ( .A(y[249]), .B(x[249]), .Z(n1409) );
  NAND U1758 ( .A(n1410), .B(n1409), .Z(n2092) );
  ANDN U1759 ( .B(n2395), .A(n2092), .Z(n1416) );
  NANDN U1760 ( .A(x[266]), .B(y[266]), .Z(n1412) );
  NANDN U1761 ( .A(x[265]), .B(y[265]), .Z(n1411) );
  AND U1762 ( .A(n1412), .B(n1411), .Z(n2394) );
  NANDN U1763 ( .A(x[256]), .B(y[256]), .Z(n1414) );
  NANDN U1764 ( .A(x[257]), .B(y[257]), .Z(n1413) );
  AND U1765 ( .A(n1414), .B(n1413), .Z(n2383) );
  AND U1766 ( .A(n2394), .B(n2383), .Z(n1415) );
  AND U1767 ( .A(n1416), .B(n1415), .Z(n1417) );
  AND U1768 ( .A(n1418), .B(n1417), .Z(n1419) );
  AND U1769 ( .A(n1420), .B(n1419), .Z(n1468) );
  NANDN U1770 ( .A(y[158]), .B(x[158]), .Z(n1422) );
  NANDN U1771 ( .A(y[157]), .B(x[157]), .Z(n1421) );
  AND U1772 ( .A(n1422), .B(n1421), .Z(n2293) );
  NANDN U1773 ( .A(y[144]), .B(x[144]), .Z(n1424) );
  NANDN U1774 ( .A(y[143]), .B(x[143]), .Z(n1423) );
  NAND U1775 ( .A(n1424), .B(n1423), .Z(n2279) );
  ANDN U1776 ( .B(n2293), .A(n2279), .Z(n1430) );
  NANDN U1777 ( .A(x[153]), .B(y[153]), .Z(n1426) );
  NANDN U1778 ( .A(x[152]), .B(y[152]), .Z(n1425) );
  AND U1779 ( .A(n1426), .B(n1425), .Z(n2286) );
  NANDN U1780 ( .A(x[145]), .B(y[145]), .Z(n1428) );
  NANDN U1781 ( .A(x[144]), .B(y[144]), .Z(n1427) );
  AND U1782 ( .A(n1428), .B(n1427), .Z(n2280) );
  AND U1783 ( .A(n2286), .B(n2280), .Z(n1429) );
  AND U1784 ( .A(n1430), .B(n1429), .Z(n1442) );
  NANDN U1785 ( .A(y[146]), .B(x[146]), .Z(n1432) );
  NANDN U1786 ( .A(y[145]), .B(x[145]), .Z(n1431) );
  AND U1787 ( .A(n1432), .B(n1431), .Z(n2281) );
  NANDN U1788 ( .A(y[136]), .B(x[136]), .Z(n1434) );
  NANDN U1789 ( .A(y[135]), .B(x[135]), .Z(n1433) );
  NAND U1790 ( .A(n1434), .B(n1433), .Z(n2120) );
  ANDN U1791 ( .B(n2281), .A(n2120), .Z(n1440) );
  NANDN U1792 ( .A(x[143]), .B(y[143]), .Z(n1436) );
  NANDN U1793 ( .A(x[142]), .B(y[142]), .Z(n1435) );
  AND U1794 ( .A(n1436), .B(n1435), .Z(n2278) );
  NANDN U1795 ( .A(y[142]), .B(x[142]), .Z(n1438) );
  NANDN U1796 ( .A(y[141]), .B(x[141]), .Z(n1437) );
  NAND U1797 ( .A(n1438), .B(n1437), .Z(n2119) );
  ANDN U1798 ( .B(n2278), .A(n2119), .Z(n1439) );
  AND U1799 ( .A(n1440), .B(n1439), .Z(n1441) );
  AND U1800 ( .A(n1442), .B(n1441), .Z(n1466) );
  NANDN U1801 ( .A(y[168]), .B(x[168]), .Z(n1444) );
  NANDN U1802 ( .A(y[167]), .B(x[167]), .Z(n1443) );
  AND U1803 ( .A(n1444), .B(n1443), .Z(n2300) );
  NANDN U1804 ( .A(y[162]), .B(x[162]), .Z(n1446) );
  NANDN U1805 ( .A(y[161]), .B(x[161]), .Z(n1445) );
  NAND U1806 ( .A(n1446), .B(n1445), .Z(n2296) );
  ANDN U1807 ( .B(n2300), .A(n2296), .Z(n1452) );
  NANDN U1808 ( .A(x[161]), .B(y[161]), .Z(n1448) );
  NANDN U1809 ( .A(x[160]), .B(y[160]), .Z(n1447) );
  AND U1810 ( .A(n1448), .B(n1447), .Z(n2295) );
  NANDN U1811 ( .A(x[159]), .B(y[159]), .Z(n1450) );
  NANDN U1812 ( .A(x[158]), .B(y[158]), .Z(n1449) );
  AND U1813 ( .A(n1450), .B(n1449), .Z(n2294) );
  AND U1814 ( .A(n2295), .B(n2294), .Z(n1451) );
  AND U1815 ( .A(n1452), .B(n1451), .Z(n1464) );
  NANDN U1816 ( .A(x[135]), .B(y[135]), .Z(n1454) );
  NANDN U1817 ( .A(x[134]), .B(y[134]), .Z(n1453) );
  AND U1818 ( .A(n1454), .B(n1453), .Z(n2271) );
  NANDN U1819 ( .A(x[133]), .B(y[133]), .Z(n1456) );
  NANDN U1820 ( .A(x[132]), .B(y[132]), .Z(n1455) );
  AND U1821 ( .A(n1456), .B(n1455), .Z(n2270) );
  AND U1822 ( .A(n2271), .B(n2270), .Z(n1462) );
  NANDN U1823 ( .A(x[137]), .B(y[137]), .Z(n1458) );
  NANDN U1824 ( .A(x[136]), .B(y[136]), .Z(n1457) );
  AND U1825 ( .A(n1458), .B(n1457), .Z(n2272) );
  NANDN U1826 ( .A(y[134]), .B(x[134]), .Z(n1460) );
  NANDN U1827 ( .A(y[133]), .B(x[133]), .Z(n1459) );
  NAND U1828 ( .A(n1460), .B(n1459), .Z(n2121) );
  ANDN U1829 ( .B(n2272), .A(n2121), .Z(n1461) );
  AND U1830 ( .A(n1462), .B(n1461), .Z(n1463) );
  AND U1831 ( .A(n1464), .B(n1463), .Z(n1465) );
  AND U1832 ( .A(n1466), .B(n1465), .Z(n1467) );
  AND U1833 ( .A(n1468), .B(n1467), .Z(n1469) );
  AND U1834 ( .A(n1470), .B(n1469), .Z(n1662) );
  NANDN U1835 ( .A(x[340]), .B(y[340]), .Z(n1472) );
  NANDN U1836 ( .A(x[339]), .B(y[339]), .Z(n1471) );
  AND U1837 ( .A(n1472), .B(n1471), .Z(n2461) );
  NANDN U1838 ( .A(y[347]), .B(x[347]), .Z(n1474) );
  NANDN U1839 ( .A(y[346]), .B(x[346]), .Z(n1473) );
  NAND U1840 ( .A(n1474), .B(n1473), .Z(n2467) );
  ANDN U1841 ( .B(n2461), .A(n2467), .Z(n1480) );
  NANDN U1842 ( .A(x[346]), .B(y[346]), .Z(n1476) );
  NANDN U1843 ( .A(x[345]), .B(y[345]), .Z(n1475) );
  AND U1844 ( .A(n1476), .B(n1475), .Z(n2466) );
  NANDN U1845 ( .A(y[345]), .B(x[345]), .Z(n1478) );
  NANDN U1846 ( .A(y[344]), .B(x[344]), .Z(n1477) );
  NAND U1847 ( .A(n1478), .B(n1477), .Z(n2065) );
  ANDN U1848 ( .B(n2466), .A(n2065), .Z(n1479) );
  AND U1849 ( .A(n1480), .B(n1479), .Z(n1492) );
  NANDN U1850 ( .A(x[338]), .B(y[338]), .Z(n1482) );
  NANDN U1851 ( .A(x[337]), .B(y[337]), .Z(n1481) );
  AND U1852 ( .A(n1482), .B(n1481), .Z(n2460) );
  NANDN U1853 ( .A(x[330]), .B(y[330]), .Z(n1484) );
  NANDN U1854 ( .A(x[329]), .B(y[329]), .Z(n1483) );
  AND U1855 ( .A(n1484), .B(n1483), .Z(n2452) );
  AND U1856 ( .A(n2460), .B(n2452), .Z(n1490) );
  NANDN U1857 ( .A(x[334]), .B(y[334]), .Z(n1486) );
  NANDN U1858 ( .A(x[333]), .B(y[333]), .Z(n1485) );
  AND U1859 ( .A(n1486), .B(n1485), .Z(n2456) );
  NANDN U1860 ( .A(y[333]), .B(x[333]), .Z(n1488) );
  NANDN U1861 ( .A(y[332]), .B(x[332]), .Z(n1487) );
  NAND U1862 ( .A(n1488), .B(n1487), .Z(n2068) );
  ANDN U1863 ( .B(n2456), .A(n2068), .Z(n1489) );
  AND U1864 ( .A(n1490), .B(n1489), .Z(n1491) );
  AND U1865 ( .A(n1492), .B(n1491), .Z(n1516) );
  NANDN U1866 ( .A(x[358]), .B(y[358]), .Z(n1494) );
  NANDN U1867 ( .A(x[357]), .B(y[357]), .Z(n1493) );
  AND U1868 ( .A(n1494), .B(n1493), .Z(n2474) );
  NANDN U1869 ( .A(y[349]), .B(x[349]), .Z(n1496) );
  NANDN U1870 ( .A(y[348]), .B(x[348]), .Z(n1495) );
  NAND U1871 ( .A(n1496), .B(n1495), .Z(n2064) );
  ANDN U1872 ( .B(n2474), .A(n2064), .Z(n1502) );
  NANDN U1873 ( .A(x[354]), .B(y[354]), .Z(n1498) );
  NANDN U1874 ( .A(x[353]), .B(y[353]), .Z(n1497) );
  AND U1875 ( .A(n1498), .B(n1497), .Z(n2472) );
  NANDN U1876 ( .A(y[351]), .B(x[351]), .Z(n1500) );
  NANDN U1877 ( .A(y[350]), .B(x[350]), .Z(n1499) );
  NAND U1878 ( .A(n1500), .B(n1499), .Z(n2063) );
  ANDN U1879 ( .B(n2472), .A(n2063), .Z(n1501) );
  AND U1880 ( .A(n1502), .B(n1501), .Z(n1514) );
  NANDN U1881 ( .A(y[329]), .B(x[329]), .Z(n1504) );
  NANDN U1882 ( .A(y[328]), .B(x[328]), .Z(n1503) );
  AND U1883 ( .A(n1504), .B(n1503), .Z(n2451) );
  NANDN U1884 ( .A(y[324]), .B(x[324]), .Z(n1506) );
  NANDN U1885 ( .A(y[323]), .B(x[323]), .Z(n1505) );
  NAND U1886 ( .A(n1506), .B(n1505), .Z(n2447) );
  ANDN U1887 ( .B(n2451), .A(n2447), .Z(n1512) );
  NANDN U1888 ( .A(x[326]), .B(y[326]), .Z(n1508) );
  NANDN U1889 ( .A(x[327]), .B(y[327]), .Z(n1507) );
  AND U1890 ( .A(n1508), .B(n1507), .Z(n2449) );
  NANDN U1891 ( .A(x[325]), .B(y[325]), .Z(n1510) );
  NANDN U1892 ( .A(x[324]), .B(y[324]), .Z(n1509) );
  AND U1893 ( .A(n1510), .B(n1509), .Z(n2448) );
  AND U1894 ( .A(n2449), .B(n2448), .Z(n1511) );
  AND U1895 ( .A(n1512), .B(n1511), .Z(n1513) );
  AND U1896 ( .A(n1514), .B(n1513), .Z(n1515) );
  AND U1897 ( .A(n1516), .B(n1515), .Z(n1564) );
  NANDN U1898 ( .A(x[311]), .B(y[311]), .Z(n1518) );
  NANDN U1899 ( .A(x[310]), .B(y[310]), .Z(n1517) );
  AND U1900 ( .A(n1518), .B(n1517), .Z(n2435) );
  NANDN U1901 ( .A(x[307]), .B(y[307]), .Z(n1520) );
  NANDN U1902 ( .A(x[306]), .B(y[306]), .Z(n1519) );
  AND U1903 ( .A(n1520), .B(n1519), .Z(n2432) );
  AND U1904 ( .A(n2435), .B(n2432), .Z(n1526) );
  NANDN U1905 ( .A(y[310]), .B(x[310]), .Z(n1522) );
  NANDN U1906 ( .A(y[309]), .B(x[309]), .Z(n1521) );
  AND U1907 ( .A(n1522), .B(n1521), .Z(n2434) );
  NANDN U1908 ( .A(y[308]), .B(x[308]), .Z(n1524) );
  NANDN U1909 ( .A(y[307]), .B(x[307]), .Z(n1523) );
  NAND U1910 ( .A(n1524), .B(n1523), .Z(n2433) );
  ANDN U1911 ( .B(n2434), .A(n2433), .Z(n1525) );
  AND U1912 ( .A(n1526), .B(n1525), .Z(n1538) );
  NANDN U1913 ( .A(y[306]), .B(x[306]), .Z(n1528) );
  NANDN U1914 ( .A(y[305]), .B(x[305]), .Z(n1527) );
  AND U1915 ( .A(n1528), .B(n1527), .Z(n2431) );
  NANDN U1916 ( .A(y[304]), .B(x[304]), .Z(n1530) );
  NANDN U1917 ( .A(y[303]), .B(x[303]), .Z(n1529) );
  NAND U1918 ( .A(n1530), .B(n1529), .Z(n2076) );
  ANDN U1919 ( .B(n2431), .A(n2076), .Z(n1536) );
  NANDN U1920 ( .A(x[301]), .B(y[301]), .Z(n1532) );
  NANDN U1921 ( .A(x[300]), .B(y[300]), .Z(n1531) );
  AND U1922 ( .A(n1532), .B(n1531), .Z(n2425) );
  NANDN U1923 ( .A(y[302]), .B(x[302]), .Z(n1534) );
  NANDN U1924 ( .A(y[301]), .B(x[301]), .Z(n1533) );
  NAND U1925 ( .A(n1534), .B(n1533), .Z(n2077) );
  ANDN U1926 ( .B(n2425), .A(n2077), .Z(n1535) );
  AND U1927 ( .A(n1536), .B(n1535), .Z(n1537) );
  AND U1928 ( .A(n1538), .B(n1537), .Z(n1562) );
  NANDN U1929 ( .A(x[319]), .B(y[319]), .Z(n1540) );
  NANDN U1930 ( .A(x[318]), .B(y[318]), .Z(n1539) );
  AND U1931 ( .A(n1540), .B(n1539), .Z(n2443) );
  NANDN U1932 ( .A(y[312]), .B(x[312]), .Z(n1542) );
  NANDN U1933 ( .A(y[311]), .B(x[311]), .Z(n1541) );
  NAND U1934 ( .A(n1542), .B(n1541), .Z(n2073) );
  ANDN U1935 ( .B(n2443), .A(n2073), .Z(n1548) );
  NANDN U1936 ( .A(x[317]), .B(y[317]), .Z(n1544) );
  NANDN U1937 ( .A(x[316]), .B(y[316]), .Z(n1543) );
  AND U1938 ( .A(n1544), .B(n1543), .Z(n2441) );
  NANDN U1939 ( .A(x[315]), .B(y[315]), .Z(n1546) );
  NANDN U1940 ( .A(x[314]), .B(y[314]), .Z(n1545) );
  AND U1941 ( .A(n1546), .B(n1545), .Z(n2437) );
  AND U1942 ( .A(n2441), .B(n2437), .Z(n1547) );
  AND U1943 ( .A(n1548), .B(n1547), .Z(n1560) );
  NANDN U1944 ( .A(x[291]), .B(y[291]), .Z(n1550) );
  NANDN U1945 ( .A(x[290]), .B(y[290]), .Z(n1549) );
  AND U1946 ( .A(n1550), .B(n1549), .Z(n2416) );
  NANDN U1947 ( .A(y[296]), .B(x[296]), .Z(n1552) );
  NANDN U1948 ( .A(y[295]), .B(x[295]), .Z(n1551) );
  NAND U1949 ( .A(n1552), .B(n1551), .Z(n2079) );
  ANDN U1950 ( .B(n2416), .A(n2079), .Z(n1558) );
  NANDN U1951 ( .A(x[293]), .B(y[293]), .Z(n1554) );
  NANDN U1952 ( .A(x[292]), .B(y[292]), .Z(n1553) );
  AND U1953 ( .A(n1554), .B(n1553), .Z(n2419) );
  NANDN U1954 ( .A(y[294]), .B(x[294]), .Z(n1556) );
  NANDN U1955 ( .A(y[293]), .B(x[293]), .Z(n1555) );
  NAND U1956 ( .A(n1556), .B(n1555), .Z(n2080) );
  ANDN U1957 ( .B(n2419), .A(n2080), .Z(n1557) );
  AND U1958 ( .A(n1558), .B(n1557), .Z(n1559) );
  AND U1959 ( .A(n1560), .B(n1559), .Z(n1561) );
  AND U1960 ( .A(n1562), .B(n1561), .Z(n1563) );
  AND U1961 ( .A(n1564), .B(n1563), .Z(n1660) );
  NANDN U1962 ( .A(x[382]), .B(y[382]), .Z(n1566) );
  NANDN U1963 ( .A(x[381]), .B(y[381]), .Z(n1565) );
  AND U1964 ( .A(n1566), .B(n1565), .Z(n2496) );
  NANDN U1965 ( .A(y[375]), .B(x[375]), .Z(n1568) );
  NANDN U1966 ( .A(y[374]), .B(x[374]), .Z(n1567) );
  NAND U1967 ( .A(n1568), .B(n1567), .Z(n2055) );
  ANDN U1968 ( .B(n2496), .A(n2055), .Z(n1574) );
  NANDN U1969 ( .A(y[381]), .B(x[381]), .Z(n1570) );
  NANDN U1970 ( .A(y[380]), .B(x[380]), .Z(n1569) );
  AND U1971 ( .A(n1570), .B(n1569), .Z(n2495) );
  NANDN U1972 ( .A(y[379]), .B(x[379]), .Z(n1572) );
  NANDN U1973 ( .A(y[378]), .B(x[378]), .Z(n1571) );
  NAND U1974 ( .A(n1572), .B(n1571), .Z(n2493) );
  ANDN U1975 ( .B(n2495), .A(n2493), .Z(n1573) );
  AND U1976 ( .A(n1574), .B(n1573), .Z(n1586) );
  NANDN U1977 ( .A(x[372]), .B(y[372]), .Z(n1576) );
  NANDN U1978 ( .A(x[371]), .B(y[371]), .Z(n1575) );
  AND U1979 ( .A(n1576), .B(n1575), .Z(n2486) );
  NANDN U1980 ( .A(y[369]), .B(x[369]), .Z(n1578) );
  NANDN U1981 ( .A(y[368]), .B(x[368]), .Z(n1577) );
  NAND U1982 ( .A(n1578), .B(n1577), .Z(n2057) );
  ANDN U1983 ( .B(n2486), .A(n2057), .Z(n1584) );
  NANDN U1984 ( .A(x[374]), .B(y[374]), .Z(n1580) );
  NANDN U1985 ( .A(x[373]), .B(y[373]), .Z(n1579) );
  AND U1986 ( .A(n1580), .B(n1579), .Z(n2488) );
  NANDN U1987 ( .A(y[371]), .B(x[371]), .Z(n1582) );
  NANDN U1988 ( .A(y[370]), .B(x[370]), .Z(n1581) );
  NAND U1989 ( .A(n1582), .B(n1581), .Z(n2056) );
  ANDN U1990 ( .B(n2488), .A(n2056), .Z(n1583) );
  AND U1991 ( .A(n1584), .B(n1583), .Z(n1585) );
  AND U1992 ( .A(n1586), .B(n1585), .Z(n1610) );
  NANDN U1993 ( .A(x[393]), .B(y[393]), .Z(n1588) );
  NANDN U1994 ( .A(x[392]), .B(y[392]), .Z(n1587) );
  AND U1995 ( .A(n1588), .B(n1587), .Z(n2508) );
  NANDN U1996 ( .A(x[384]), .B(y[384]), .Z(n1590) );
  NANDN U1997 ( .A(x[383]), .B(y[383]), .Z(n1589) );
  AND U1998 ( .A(n1590), .B(n1589), .Z(n2498) );
  AND U1999 ( .A(n2508), .B(n2498), .Z(n1596) );
  NANDN U2000 ( .A(y[388]), .B(x[388]), .Z(n1592) );
  NANDN U2001 ( .A(y[387]), .B(x[387]), .Z(n1591) );
  AND U2002 ( .A(n1592), .B(n1591), .Z(n2504) );
  NANDN U2003 ( .A(y[386]), .B(x[386]), .Z(n1594) );
  NANDN U2004 ( .A(y[385]), .B(x[385]), .Z(n1593) );
  NAND U2005 ( .A(n1594), .B(n1593), .Z(n2501) );
  ANDN U2006 ( .B(n2504), .A(n2501), .Z(n1595) );
  AND U2007 ( .A(n1596), .B(n1595), .Z(n1608) );
  NANDN U2008 ( .A(x[368]), .B(y[368]), .Z(n1598) );
  NANDN U2009 ( .A(x[367]), .B(y[367]), .Z(n1597) );
  AND U2010 ( .A(n1598), .B(n1597), .Z(n2483) );
  NANDN U2011 ( .A(x[360]), .B(y[360]), .Z(n1600) );
  NANDN U2012 ( .A(x[359]), .B(y[359]), .Z(n1599) );
  AND U2013 ( .A(n1600), .B(n1599), .Z(n2476) );
  AND U2014 ( .A(n2483), .B(n2476), .Z(n1606) );
  NANDN U2015 ( .A(y[365]), .B(x[365]), .Z(n1602) );
  NANDN U2016 ( .A(y[364]), .B(x[364]), .Z(n1601) );
  AND U2017 ( .A(n1602), .B(n1601), .Z(n2481) );
  NANDN U2018 ( .A(y[361]), .B(x[361]), .Z(n1604) );
  NANDN U2019 ( .A(y[360]), .B(x[360]), .Z(n1603) );
  NAND U2020 ( .A(n1604), .B(n1603), .Z(n2060) );
  ANDN U2021 ( .B(n2481), .A(n2060), .Z(n1605) );
  AND U2022 ( .A(n1606), .B(n1605), .Z(n1607) );
  AND U2023 ( .A(n1608), .B(n1607), .Z(n1609) );
  AND U2024 ( .A(n1610), .B(n1609), .Z(n1658) );
  NANDN U2025 ( .A(x[278]), .B(y[278]), .Z(n1612) );
  NANDN U2026 ( .A(x[277]), .B(y[277]), .Z(n1611) );
  AND U2027 ( .A(n1612), .B(n1611), .Z(n2403) );
  NANDN U2028 ( .A(y[275]), .B(x[275]), .Z(n1614) );
  NANDN U2029 ( .A(y[274]), .B(x[274]), .Z(n1613) );
  NAND U2030 ( .A(n1614), .B(n1613), .Z(n2401) );
  ANDN U2031 ( .B(n2403), .A(n2401), .Z(n1620) );
  NANDN U2032 ( .A(x[276]), .B(y[276]), .Z(n1616) );
  NANDN U2033 ( .A(x[275]), .B(y[275]), .Z(n1615) );
  AND U2034 ( .A(n1616), .B(n1615), .Z(n2402) );
  NANDN U2035 ( .A(y[277]), .B(x[277]), .Z(n1618) );
  NANDN U2036 ( .A(y[276]), .B(x[276]), .Z(n1617) );
  NAND U2037 ( .A(n1618), .B(n1617), .Z(n2086) );
  ANDN U2038 ( .B(n2402), .A(n2086), .Z(n1619) );
  AND U2039 ( .A(n1620), .B(n1619), .Z(n1632) );
  NANDN U2040 ( .A(x[274]), .B(y[274]), .Z(n1622) );
  NANDN U2041 ( .A(x[273]), .B(y[273]), .Z(n1621) );
  AND U2042 ( .A(n1622), .B(n1621), .Z(n2400) );
  NANDN U2043 ( .A(x[264]), .B(y[264]), .Z(n1624) );
  NANDN U2044 ( .A(x[263]), .B(y[263]), .Z(n1623) );
  AND U2045 ( .A(n1624), .B(n1623), .Z(n2390) );
  AND U2046 ( .A(n2400), .B(n2390), .Z(n1630) );
  NANDN U2047 ( .A(x[268]), .B(y[268]), .Z(n1626) );
  NANDN U2048 ( .A(x[267]), .B(y[267]), .Z(n1625) );
  AND U2049 ( .A(n1626), .B(n1625), .Z(n2396) );
  NANDN U2050 ( .A(y[273]), .B(x[273]), .Z(n1628) );
  NANDN U2051 ( .A(y[272]), .B(x[272]), .Z(n1627) );
  NAND U2052 ( .A(n1628), .B(n1627), .Z(n2087) );
  ANDN U2053 ( .B(n2396), .A(n2087), .Z(n1629) );
  AND U2054 ( .A(n1630), .B(n1629), .Z(n1631) );
  AND U2055 ( .A(n1632), .B(n1631), .Z(n1656) );
  NANDN U2056 ( .A(y[284]), .B(x[284]), .Z(n1634) );
  NANDN U2057 ( .A(y[283]), .B(x[283]), .Z(n1633) );
  AND U2058 ( .A(n1634), .B(n1633), .Z(n2409) );
  NANDN U2059 ( .A(y[279]), .B(x[279]), .Z(n1636) );
  NANDN U2060 ( .A(y[278]), .B(x[278]), .Z(n1635) );
  NAND U2061 ( .A(n1636), .B(n1635), .Z(n2085) );
  ANDN U2062 ( .B(n2409), .A(n2085), .Z(n1642) );
  NANDN U2063 ( .A(x[282]), .B(y[282]), .Z(n1638) );
  NANDN U2064 ( .A(x[281]), .B(y[281]), .Z(n1637) );
  AND U2065 ( .A(n1638), .B(n1637), .Z(n2407) );
  NANDN U2066 ( .A(y[281]), .B(x[281]), .Z(n1640) );
  NANDN U2067 ( .A(y[280]), .B(x[280]), .Z(n1639) );
  NAND U2068 ( .A(n1640), .B(n1639), .Z(n2406) );
  ANDN U2069 ( .B(n2407), .A(n2406), .Z(n1641) );
  AND U2070 ( .A(n1642), .B(n1641), .Z(n1654) );
  NANDN U2071 ( .A(y[269]), .B(x[269]), .Z(n1644) );
  NANDN U2072 ( .A(y[268]), .B(x[268]), .Z(n1643) );
  AND U2073 ( .A(n1644), .B(n1643), .Z(n2397) );
  NANDN U2074 ( .A(y[261]), .B(x[261]), .Z(n1646) );
  NANDN U2075 ( .A(y[260]), .B(x[260]), .Z(n1645) );
  NAND U2076 ( .A(n1646), .B(n1645), .Z(n2388) );
  ANDN U2077 ( .B(n2397), .A(n2388), .Z(n1652) );
  NANDN U2078 ( .A(x[262]), .B(y[262]), .Z(n1648) );
  NANDN U2079 ( .A(x[261]), .B(y[261]), .Z(n1647) );
  AND U2080 ( .A(n1648), .B(n1647), .Z(n2389) );
  NANDN U2081 ( .A(y[263]), .B(x[263]), .Z(n1650) );
  NANDN U2082 ( .A(y[262]), .B(x[262]), .Z(n1649) );
  NAND U2083 ( .A(n1650), .B(n1649), .Z(n2090) );
  ANDN U2084 ( .B(n2389), .A(n2090), .Z(n1651) );
  AND U2085 ( .A(n1652), .B(n1651), .Z(n1653) );
  AND U2086 ( .A(n1654), .B(n1653), .Z(n1655) );
  AND U2087 ( .A(n1656), .B(n1655), .Z(n1657) );
  AND U2088 ( .A(n1658), .B(n1657), .Z(n1659) );
  AND U2089 ( .A(n1660), .B(n1659), .Z(n1661) );
  AND U2090 ( .A(n1662), .B(n1661), .Z(n1663) );
  AND U2091 ( .A(n1664), .B(n1663), .Z(n1712) );
  NANDN U2092 ( .A(x[366]), .B(y[366]), .Z(n1666) );
  NANDN U2093 ( .A(x[365]), .B(y[365]), .Z(n1665) );
  AND U2094 ( .A(n1666), .B(n1665), .Z(n2482) );
  NANDN U2095 ( .A(y[373]), .B(x[373]), .Z(n1668) );
  NANDN U2096 ( .A(y[372]), .B(x[372]), .Z(n1667) );
  NAND U2097 ( .A(n1668), .B(n1667), .Z(n2487) );
  ANDN U2098 ( .B(n2482), .A(n2487), .Z(n1674) );
  NANDN U2099 ( .A(x[376]), .B(y[376]), .Z(n1670) );
  NANDN U2100 ( .A(x[375]), .B(y[375]), .Z(n1669) );
  AND U2101 ( .A(n1670), .B(n1669), .Z(n2491) );
  NANDN U2102 ( .A(y[367]), .B(x[367]), .Z(n1672) );
  NANDN U2103 ( .A(y[366]), .B(x[366]), .Z(n1671) );
  NAND U2104 ( .A(n1672), .B(n1671), .Z(n2058) );
  ANDN U2105 ( .B(n2491), .A(n2058), .Z(n1673) );
  AND U2106 ( .A(n1674), .B(n1673), .Z(n1686) );
  NANDN U2107 ( .A(x[364]), .B(y[364]), .Z(n1676) );
  NANDN U2108 ( .A(x[363]), .B(y[363]), .Z(n1675) );
  AND U2109 ( .A(n1676), .B(n1675), .Z(n2480) );
  NANDN U2110 ( .A(y[363]), .B(x[363]), .Z(n1678) );
  NANDN U2111 ( .A(y[362]), .B(x[362]), .Z(n1677) );
  NAND U2112 ( .A(n1678), .B(n1677), .Z(n2059) );
  ANDN U2113 ( .B(n2480), .A(n2059), .Z(n1684) );
  NANDN U2114 ( .A(x[362]), .B(y[362]), .Z(n1680) );
  NANDN U2115 ( .A(x[361]), .B(y[361]), .Z(n1679) );
  AND U2116 ( .A(n1680), .B(n1679), .Z(n2479) );
  NANDN U2117 ( .A(y[357]), .B(x[357]), .Z(n1682) );
  NANDN U2118 ( .A(y[356]), .B(x[356]), .Z(n1681) );
  NAND U2119 ( .A(n1682), .B(n1681), .Z(n2061) );
  ANDN U2120 ( .B(n2479), .A(n2061), .Z(n1683) );
  AND U2121 ( .A(n1684), .B(n1683), .Z(n1685) );
  AND U2122 ( .A(n1686), .B(n1685), .Z(n1710) );
  NANDN U2123 ( .A(x[380]), .B(y[380]), .Z(n1688) );
  NANDN U2124 ( .A(x[379]), .B(y[379]), .Z(n1687) );
  AND U2125 ( .A(n1688), .B(n1687), .Z(n2494) );
  NANDN U2126 ( .A(y[377]), .B(x[377]), .Z(n1690) );
  NANDN U2127 ( .A(y[376]), .B(x[376]), .Z(n1689) );
  NAND U2128 ( .A(n1690), .B(n1689), .Z(n2054) );
  ANDN U2129 ( .B(n2494), .A(n2054), .Z(n1696) );
  NANDN U2130 ( .A(x[378]), .B(y[378]), .Z(n1692) );
  NANDN U2131 ( .A(x[377]), .B(y[377]), .Z(n1691) );
  AND U2132 ( .A(n1692), .B(n1691), .Z(n2492) );
  NANDN U2133 ( .A(y[390]), .B(x[390]), .Z(n1694) );
  NANDN U2134 ( .A(y[389]), .B(x[389]), .Z(n1693) );
  NAND U2135 ( .A(n1694), .B(n1693), .Z(n2052) );
  ANDN U2136 ( .B(n2492), .A(n2052), .Z(n1695) );
  AND U2137 ( .A(n1696), .B(n1695), .Z(n1708) );
  NANDN U2138 ( .A(x[356]), .B(y[356]), .Z(n1698) );
  NANDN U2139 ( .A(x[355]), .B(y[355]), .Z(n1697) );
  AND U2140 ( .A(n1698), .B(n1697), .Z(n2473) );
  NANDN U2141 ( .A(x[348]), .B(y[348]), .Z(n1700) );
  NANDN U2142 ( .A(x[347]), .B(y[347]), .Z(n1699) );
  AND U2143 ( .A(n1700), .B(n1699), .Z(n2468) );
  AND U2144 ( .A(n2473), .B(n2468), .Z(n1706) );
  NANDN U2145 ( .A(x[352]), .B(y[352]), .Z(n1702) );
  NANDN U2146 ( .A(x[351]), .B(y[351]), .Z(n1701) );
  AND U2147 ( .A(n1702), .B(n1701), .Z(n2470) );
  NANDN U2148 ( .A(y[355]), .B(x[355]), .Z(n1704) );
  NANDN U2149 ( .A(y[354]), .B(x[354]), .Z(n1703) );
  NAND U2150 ( .A(n1704), .B(n1703), .Z(n2062) );
  ANDN U2151 ( .B(n2470), .A(n2062), .Z(n1705) );
  AND U2152 ( .A(n1706), .B(n1705), .Z(n1707) );
  AND U2153 ( .A(n1708), .B(n1707), .Z(n1709) );
  AND U2154 ( .A(n1710), .B(n1709), .Z(n1711) );
  AND U2155 ( .A(n1712), .B(n1711), .Z(n2017) );
  NANDN U2156 ( .A(x[2]), .B(y[2]), .Z(n2165) );
  NANDN U2157 ( .A(x[1]), .B(y[1]), .Z(n2163) );
  AND U2158 ( .A(n2165), .B(n2163), .Z(n1714) );
  NANDN U2159 ( .A(x[0]), .B(y[0]), .Z(n1713) );
  AND U2160 ( .A(n1714), .B(n1713), .Z(n1715) );
  NANDN U2161 ( .A(x[60]), .B(y[60]), .Z(n2144) );
  AND U2162 ( .A(n1715), .B(n2144), .Z(n1716) );
  NANDN U2163 ( .A(x[61]), .B(y[61]), .Z(n2143) );
  AND U2164 ( .A(n1716), .B(n2143), .Z(n1720) );
  NANDN U2165 ( .A(x[68]), .B(y[68]), .Z(n2140) );
  NANDN U2166 ( .A(y[49]), .B(x[49]), .Z(n1718) );
  NANDN U2167 ( .A(y[50]), .B(x[50]), .Z(n1717) );
  NAND U2168 ( .A(n1718), .B(n1717), .Z(n2148) );
  ANDN U2169 ( .B(n2140), .A(n2148), .Z(n1719) );
  AND U2170 ( .A(n1720), .B(n1719), .Z(n1721) );
  ANDN U2171 ( .B(x[114]), .A(y[114]), .Z(n2127) );
  ANDN U2172 ( .B(n1721), .A(n2127), .Z(n1725) );
  NANDN U2173 ( .A(x[69]), .B(y[69]), .Z(n2139) );
  NANDN U2174 ( .A(y[106]), .B(x[106]), .Z(n1723) );
  NANDN U2175 ( .A(y[105]), .B(x[105]), .Z(n1722) );
  NAND U2176 ( .A(n1723), .B(n1722), .Z(n2247) );
  ANDN U2177 ( .B(n2139), .A(n2247), .Z(n1724) );
  AND U2178 ( .A(n1725), .B(n1724), .Z(n1726) );
  NANDN U2179 ( .A(x[194]), .B(y[194]), .Z(n2324) );
  AND U2180 ( .A(n1726), .B(n2324), .Z(n1730) );
  NANDN U2181 ( .A(x[123]), .B(y[123]), .Z(n1728) );
  NANDN U2182 ( .A(x[122]), .B(y[122]), .Z(n1727) );
  AND U2183 ( .A(n1728), .B(n1727), .Z(n2261) );
  ANDN U2184 ( .B(x[113]), .A(y[113]), .Z(n2255) );
  ANDN U2185 ( .B(n2261), .A(n2255), .Z(n1729) );
  AND U2186 ( .A(n1730), .B(n1729), .Z(n1734) );
  NANDN U2187 ( .A(x[370]), .B(y[370]), .Z(n2484) );
  NANDN U2188 ( .A(y[315]), .B(x[315]), .Z(n2439) );
  AND U2189 ( .A(n2484), .B(n2439), .Z(n1732) );
  NANDN U2190 ( .A(x[328]), .B(y[328]), .Z(n2450) );
  ANDN U2191 ( .B(x[327]), .A(y[327]), .Z(n2069) );
  ANDN U2192 ( .B(n2450), .A(n2069), .Z(n1731) );
  AND U2193 ( .A(n1732), .B(n1731), .Z(n1733) );
  AND U2194 ( .A(n1734), .B(n1733), .Z(n1747) );
  NANDN U2195 ( .A(x[305]), .B(y[305]), .Z(n2429) );
  ANDN U2196 ( .B(x[265]), .A(y[265]), .Z(n2391) );
  ANDN U2197 ( .B(n2429), .A(n2391), .Z(n1736) );
  NANDN U2198 ( .A(x[286]), .B(y[286]), .Z(n2083) );
  NANDN U2199 ( .A(y[288]), .B(x[288]), .Z(n2413) );
  AND U2200 ( .A(n2083), .B(n2413), .Z(n1735) );
  AND U2201 ( .A(n1736), .B(n1735), .Z(n1737) );
  NANDN U2202 ( .A(x[369]), .B(y[369]), .Z(n2485) );
  AND U2203 ( .A(n1737), .B(n2485), .Z(n1741) );
  NANDN U2204 ( .A(y[358]), .B(x[358]), .Z(n1739) );
  NANDN U2205 ( .A(y[359]), .B(x[359]), .Z(n1738) );
  AND U2206 ( .A(n1739), .B(n1738), .Z(n2475) );
  ANDN U2207 ( .B(x[383]), .A(y[383]), .Z(n2497) );
  ANDN U2208 ( .B(n2475), .A(n2497), .Z(n1740) );
  AND U2209 ( .A(n1741), .B(n1740), .Z(n1745) );
  NANDN U2210 ( .A(x[294]), .B(y[294]), .Z(n2420) );
  NANDN U2211 ( .A(x[304]), .B(y[304]), .Z(n2430) );
  AND U2212 ( .A(n2420), .B(n2430), .Z(n1743) );
  NANDN U2213 ( .A(x[309]), .B(y[309]), .Z(n2075) );
  ANDN U2214 ( .B(x[291]), .A(y[291]), .Z(n2081) );
  ANDN U2215 ( .B(n2075), .A(n2081), .Z(n1742) );
  AND U2216 ( .A(n1743), .B(n1742), .Z(n1744) );
  AND U2217 ( .A(n1745), .B(n1744), .Z(n1746) );
  AND U2218 ( .A(n1747), .B(n1746), .Z(n1766) );
  NANDN U2219 ( .A(y[384]), .B(x[384]), .Z(n2499) );
  NANDN U2220 ( .A(y[409]), .B(x[409]), .Z(n2521) );
  AND U2221 ( .A(n2499), .B(n2521), .Z(n1749) );
  NANDN U2222 ( .A(x[385]), .B(y[385]), .Z(n2500) );
  ANDN U2223 ( .B(x[382]), .A(y[382]), .Z(n2053) );
  ANDN U2224 ( .B(n2500), .A(n2053), .Z(n1748) );
  AND U2225 ( .A(n1749), .B(n1748), .Z(n1750) );
  ANDN U2226 ( .B(x[410]), .A(y[410]), .Z(n2520) );
  ANDN U2227 ( .B(n1750), .A(n2520), .Z(n1754) );
  NANDN U2228 ( .A(x[419]), .B(y[419]), .Z(n2043) );
  NANDN U2229 ( .A(y[398]), .B(x[398]), .Z(n1752) );
  NANDN U2230 ( .A(y[397]), .B(x[397]), .Z(n1751) );
  NAND U2231 ( .A(n1752), .B(n1751), .Z(n2511) );
  ANDN U2232 ( .B(n2043), .A(n2511), .Z(n1753) );
  AND U2233 ( .A(n1754), .B(n1753), .Z(n1755) );
  ANDN U2234 ( .B(x[463]), .A(y[463]), .Z(n2032) );
  ANDN U2235 ( .B(n1755), .A(n2032), .Z(n1759) );
  NANDN U2236 ( .A(x[418]), .B(y[418]), .Z(n2042) );
  NANDN U2237 ( .A(y[456]), .B(x[456]), .Z(n1757) );
  NANDN U2238 ( .A(y[455]), .B(x[455]), .Z(n1756) );
  NAND U2239 ( .A(n1757), .B(n1756), .Z(n2560) );
  ANDN U2240 ( .B(n2042), .A(n2560), .Z(n1758) );
  AND U2241 ( .A(n1759), .B(n1758), .Z(n1760) );
  NANDN U2242 ( .A(x[511]), .B(y[511]), .Z(n2609) );
  AND U2243 ( .A(n1760), .B(n2609), .Z(n1764) );
  NANDN U2244 ( .A(y[473]), .B(x[473]), .Z(n1762) );
  NANDN U2245 ( .A(y[474]), .B(x[474]), .Z(n1761) );
  AND U2246 ( .A(n1762), .B(n1761), .Z(n2577) );
  ANDN U2247 ( .B(x[464]), .A(y[464]), .Z(n2568) );
  ANDN U2248 ( .B(n2577), .A(n2568), .Z(n1763) );
  AND U2249 ( .A(n1764), .B(n1763), .Z(n1765) );
  AND U2250 ( .A(n1766), .B(n1765), .Z(n1784) );
  NANDN U2251 ( .A(y[178]), .B(x[178]), .Z(n1768) );
  NANDN U2252 ( .A(y[177]), .B(x[177]), .Z(n1767) );
  AND U2253 ( .A(n1768), .B(n1767), .Z(n2309) );
  NANDN U2254 ( .A(y[206]), .B(x[206]), .Z(n2334) );
  AND U2255 ( .A(n2309), .B(n2334), .Z(n1773) );
  NANDN U2256 ( .A(x[251]), .B(y[251]), .Z(n2372) );
  NANDN U2257 ( .A(y[253]), .B(x[253]), .Z(n2376) );
  AND U2258 ( .A(n2372), .B(n2376), .Z(n1770) );
  NANDN U2259 ( .A(x[249]), .B(y[249]), .Z(n2371) );
  ANDN U2260 ( .B(x[254]), .A(y[254]), .Z(n2379) );
  ANDN U2261 ( .B(n2371), .A(n2379), .Z(n1769) );
  AND U2262 ( .A(n1770), .B(n1769), .Z(n1771) );
  NANDN U2263 ( .A(x[195]), .B(y[195]), .Z(n2325) );
  AND U2264 ( .A(n1771), .B(n2325), .Z(n1772) );
  AND U2265 ( .A(n1773), .B(n1772), .Z(n1774) );
  NANDN U2266 ( .A(x[248]), .B(y[248]), .Z(n2370) );
  AND U2267 ( .A(n1774), .B(n2370), .Z(n1778) );
  NANDN U2268 ( .A(x[244]), .B(y[244]), .Z(n1776) );
  NANDN U2269 ( .A(x[245]), .B(y[245]), .Z(n1775) );
  AND U2270 ( .A(n1776), .B(n1775), .Z(n2368) );
  ANDN U2271 ( .B(x[205]), .A(y[205]), .Z(n2333) );
  ANDN U2272 ( .B(n2368), .A(n2333), .Z(n1777) );
  AND U2273 ( .A(n1778), .B(n1777), .Z(n1782) );
  NANDN U2274 ( .A(x[283]), .B(y[283]), .Z(n2408) );
  ANDN U2275 ( .B(x[256]), .A(y[256]), .Z(n2382) );
  ANDN U2276 ( .B(n2408), .A(n2382), .Z(n1780) );
  NANDN U2277 ( .A(y[257]), .B(x[257]), .Z(n2384) );
  ANDN U2278 ( .B(x[282]), .A(y[282]), .Z(n2084) );
  ANDN U2279 ( .B(n2384), .A(n2084), .Z(n1779) );
  AND U2280 ( .A(n1780), .B(n1779), .Z(n1781) );
  AND U2281 ( .A(n1782), .B(n1781), .Z(n1783) );
  AND U2282 ( .A(n1784), .B(n1783), .Z(n1832) );
  NANDN U2283 ( .A(y[458]), .B(x[458]), .Z(n1786) );
  NANDN U2284 ( .A(y[457]), .B(x[457]), .Z(n1785) );
  AND U2285 ( .A(n1786), .B(n1785), .Z(n2562) );
  NANDN U2286 ( .A(y[442]), .B(x[442]), .Z(n1788) );
  NANDN U2287 ( .A(y[441]), .B(x[441]), .Z(n1787) );
  NAND U2288 ( .A(n1788), .B(n1787), .Z(n2037) );
  ANDN U2289 ( .B(n2562), .A(n2037), .Z(n1794) );
  NANDN U2290 ( .A(x[447]), .B(y[447]), .Z(n1790) );
  NANDN U2291 ( .A(x[446]), .B(y[446]), .Z(n1789) );
  AND U2292 ( .A(n1790), .B(n1789), .Z(n2554) );
  NANDN U2293 ( .A(y[448]), .B(x[448]), .Z(n1792) );
  NANDN U2294 ( .A(y[447]), .B(x[447]), .Z(n1791) );
  NAND U2295 ( .A(n1792), .B(n1791), .Z(n2036) );
  ANDN U2296 ( .B(n2554), .A(n2036), .Z(n1793) );
  AND U2297 ( .A(n1794), .B(n1793), .Z(n1806) );
  NANDN U2298 ( .A(x[435]), .B(y[435]), .Z(n1796) );
  NANDN U2299 ( .A(x[434]), .B(y[434]), .Z(n1795) );
  AND U2300 ( .A(n1796), .B(n1795), .Z(n2543) );
  NANDN U2301 ( .A(y[438]), .B(x[438]), .Z(n1798) );
  NANDN U2302 ( .A(y[437]), .B(x[437]), .Z(n1797) );
  NAND U2303 ( .A(n1798), .B(n1797), .Z(n2545) );
  ANDN U2304 ( .B(n2543), .A(n2545), .Z(n1804) );
  NANDN U2305 ( .A(y[446]), .B(x[446]), .Z(n1800) );
  NANDN U2306 ( .A(y[445]), .B(x[445]), .Z(n1799) );
  AND U2307 ( .A(n1800), .B(n1799), .Z(n2553) );
  NANDN U2308 ( .A(y[436]), .B(x[436]), .Z(n1802) );
  NANDN U2309 ( .A(y[435]), .B(x[435]), .Z(n1801) );
  NAND U2310 ( .A(n1802), .B(n1801), .Z(n2039) );
  ANDN U2311 ( .B(n2553), .A(n2039), .Z(n1803) );
  AND U2312 ( .A(n1804), .B(n1803), .Z(n1805) );
  AND U2313 ( .A(n1806), .B(n1805), .Z(n1830) );
  NANDN U2314 ( .A(x[449]), .B(y[449]), .Z(n1808) );
  NANDN U2315 ( .A(x[448]), .B(y[448]), .Z(n1807) );
  AND U2316 ( .A(n1808), .B(n1807), .Z(n2555) );
  NANDN U2317 ( .A(y[460]), .B(x[460]), .Z(n1810) );
  NANDN U2318 ( .A(y[459]), .B(x[459]), .Z(n1809) );
  NAND U2319 ( .A(n1810), .B(n1809), .Z(n2033) );
  ANDN U2320 ( .B(n2555), .A(n2033), .Z(n1816) );
  NANDN U2321 ( .A(x[459]), .B(y[459]), .Z(n1812) );
  NANDN U2322 ( .A(x[458]), .B(y[458]), .Z(n1811) );
  AND U2323 ( .A(n1812), .B(n1811), .Z(n2564) );
  NANDN U2324 ( .A(y[450]), .B(x[450]), .Z(n1814) );
  NANDN U2325 ( .A(y[449]), .B(x[449]), .Z(n1813) );
  NAND U2326 ( .A(n1814), .B(n1813), .Z(n2556) );
  ANDN U2327 ( .B(n2564), .A(n2556), .Z(n1815) );
  AND U2328 ( .A(n1816), .B(n1815), .Z(n1828) );
  NANDN U2329 ( .A(x[427]), .B(y[427]), .Z(n1818) );
  NANDN U2330 ( .A(x[426]), .B(y[426]), .Z(n1817) );
  AND U2331 ( .A(n1818), .B(n1817), .Z(n2535) );
  NANDN U2332 ( .A(x[425]), .B(y[425]), .Z(n1820) );
  NANDN U2333 ( .A(x[424]), .B(y[424]), .Z(n1819) );
  AND U2334 ( .A(n1820), .B(n1819), .Z(n2533) );
  AND U2335 ( .A(n2535), .B(n2533), .Z(n1826) );
  NANDN U2336 ( .A(x[433]), .B(y[433]), .Z(n1822) );
  NANDN U2337 ( .A(x[432]), .B(y[432]), .Z(n1821) );
  AND U2338 ( .A(n1822), .B(n1821), .Z(n2541) );
  NANDN U2339 ( .A(y[426]), .B(x[426]), .Z(n1824) );
  NANDN U2340 ( .A(y[425]), .B(x[425]), .Z(n1823) );
  NAND U2341 ( .A(n1824), .B(n1823), .Z(n2534) );
  ANDN U2342 ( .B(n2541), .A(n2534), .Z(n1825) );
  AND U2343 ( .A(n1826), .B(n1825), .Z(n1827) );
  AND U2344 ( .A(n1828), .B(n1827), .Z(n1829) );
  AND U2345 ( .A(n1830), .B(n1829), .Z(n1831) );
  AND U2346 ( .A(n1832), .B(n1831), .Z(n1967) );
  NANDN U2347 ( .A(x[252]), .B(y[252]), .Z(n2374) );
  ANDN U2348 ( .B(x[251]), .A(y[251]), .Z(n2091) );
  ANDN U2349 ( .B(n2374), .A(n2091), .Z(n1833) );
  NANDN U2350 ( .A(x[250]), .B(y[250]), .Z(n2373) );
  AND U2351 ( .A(n1833), .B(n2373), .Z(n1836) );
  NANDN U2352 ( .A(x[258]), .B(y[258]), .Z(n2385) );
  ANDN U2353 ( .B(x[252]), .A(y[252]), .Z(n2375) );
  ANDN U2354 ( .B(n2385), .A(n2375), .Z(n1834) );
  NANDN U2355 ( .A(x[287]), .B(y[287]), .Z(n2082) );
  AND U2356 ( .A(n1834), .B(n2082), .Z(n1835) );
  AND U2357 ( .A(n1836), .B(n1835), .Z(n1838) );
  XNOR U2358 ( .A(x[255]), .B(y[255]), .Z(n1837) );
  AND U2359 ( .A(n1838), .B(n1837), .Z(n1839) );
  ANDN U2360 ( .B(x[0]), .A(y[0]), .Z(n2162) );
  ANDN U2361 ( .B(n1839), .A(n2162), .Z(n1843) );
  NANDN U2362 ( .A(x[3]), .B(y[3]), .Z(n2166) );
  NANDN U2363 ( .A(y[507]), .B(x[507]), .Z(n1841) );
  NANDN U2364 ( .A(y[508]), .B(x[508]), .Z(n1840) );
  NAND U2365 ( .A(n1841), .B(n1840), .Z(n2607) );
  ANDN U2366 ( .B(n2166), .A(n2607), .Z(n1842) );
  AND U2367 ( .A(n1843), .B(n1842), .Z(n1855) );
  NANDN U2368 ( .A(y[490]), .B(x[490]), .Z(n1845) );
  NANDN U2369 ( .A(y[489]), .B(x[489]), .Z(n1844) );
  AND U2370 ( .A(n1845), .B(n1844), .Z(n2592) );
  NANDN U2371 ( .A(y[486]), .B(x[486]), .Z(n1847) );
  NANDN U2372 ( .A(y[485]), .B(x[485]), .Z(n1846) );
  NAND U2373 ( .A(n1847), .B(n1846), .Z(n2027) );
  ANDN U2374 ( .B(n2592), .A(n2027), .Z(n1853) );
  NANDN U2375 ( .A(x[487]), .B(y[487]), .Z(n1849) );
  NANDN U2376 ( .A(x[486]), .B(y[486]), .Z(n1848) );
  AND U2377 ( .A(n1849), .B(n1848), .Z(n2588) );
  NANDN U2378 ( .A(y[492]), .B(x[492]), .Z(n1851) );
  NANDN U2379 ( .A(y[491]), .B(x[491]), .Z(n1850) );
  NAND U2380 ( .A(n1851), .B(n1850), .Z(n2026) );
  ANDN U2381 ( .B(n2588), .A(n2026), .Z(n1852) );
  AND U2382 ( .A(n1853), .B(n1852), .Z(n1854) );
  AND U2383 ( .A(n1855), .B(n1854), .Z(n1871) );
  NANDN U2384 ( .A(x[308]), .B(y[308]), .Z(n2074) );
  ANDN U2385 ( .B(x[264]), .A(y[264]), .Z(n2089) );
  ANDN U2386 ( .B(n2074), .A(n2089), .Z(n1857) );
  NANDN U2387 ( .A(y[292]), .B(x[292]), .Z(n2418) );
  ANDN U2388 ( .B(x[287]), .A(y[287]), .Z(n2412) );
  ANDN U2389 ( .B(n2418), .A(n2412), .Z(n1856) );
  AND U2390 ( .A(n1857), .B(n1856), .Z(n1869) );
  NANDN U2391 ( .A(x[479]), .B(y[479]), .Z(n1859) );
  NANDN U2392 ( .A(x[478]), .B(y[478]), .Z(n1858) );
  AND U2393 ( .A(n1859), .B(n1858), .Z(n2582) );
  NANDN U2394 ( .A(x[477]), .B(y[477]), .Z(n1861) );
  NANDN U2395 ( .A(x[476]), .B(y[476]), .Z(n1860) );
  AND U2396 ( .A(n1861), .B(n1860), .Z(n2580) );
  AND U2397 ( .A(n2582), .B(n2580), .Z(n1867) );
  NANDN U2398 ( .A(y[478]), .B(x[478]), .Z(n1863) );
  NANDN U2399 ( .A(y[477]), .B(x[477]), .Z(n1862) );
  AND U2400 ( .A(n1863), .B(n1862), .Z(n2581) );
  NANDN U2401 ( .A(y[480]), .B(x[480]), .Z(n1865) );
  NANDN U2402 ( .A(y[479]), .B(x[479]), .Z(n1864) );
  NAND U2403 ( .A(n1865), .B(n1864), .Z(n2029) );
  ANDN U2404 ( .B(n2581), .A(n2029), .Z(n1866) );
  AND U2405 ( .A(n1867), .B(n1866), .Z(n1868) );
  AND U2406 ( .A(n1869), .B(n1868), .Z(n1870) );
  AND U2407 ( .A(n1871), .B(n1870), .Z(n1883) );
  NANDN U2408 ( .A(y[476]), .B(x[476]), .Z(n1873) );
  NANDN U2409 ( .A(y[475]), .B(x[475]), .Z(n1872) );
  AND U2410 ( .A(n1873), .B(n1872), .Z(n2579) );
  NANDN U2411 ( .A(y[472]), .B(x[472]), .Z(n1875) );
  NANDN U2412 ( .A(y[471]), .B(x[471]), .Z(n1874) );
  NAND U2413 ( .A(n1875), .B(n1874), .Z(n2030) );
  ANDN U2414 ( .B(n2579), .A(n2030), .Z(n1881) );
  NANDN U2415 ( .A(x[469]), .B(y[469]), .Z(n1877) );
  NANDN U2416 ( .A(x[468]), .B(y[468]), .Z(n1876) );
  AND U2417 ( .A(n1877), .B(n1876), .Z(n2572) );
  NANDN U2418 ( .A(y[470]), .B(x[470]), .Z(n1879) );
  NANDN U2419 ( .A(y[469]), .B(x[469]), .Z(n1878) );
  NAND U2420 ( .A(n1879), .B(n1878), .Z(n2573) );
  ANDN U2421 ( .B(n2572), .A(n2573), .Z(n1880) );
  AND U2422 ( .A(n1881), .B(n1880), .Z(n1882) );
  AND U2423 ( .A(n1883), .B(n1882), .Z(n1917) );
  NANDN U2424 ( .A(x[503]), .B(y[503]), .Z(n1885) );
  NANDN U2425 ( .A(x[502]), .B(y[502]), .Z(n1884) );
  AND U2426 ( .A(n1885), .B(n1884), .Z(n2603) );
  NANDN U2427 ( .A(x[499]), .B(y[499]), .Z(n1887) );
  NANDN U2428 ( .A(x[498]), .B(y[498]), .Z(n1886) );
  AND U2429 ( .A(n1887), .B(n1886), .Z(n2598) );
  AND U2430 ( .A(n2603), .B(n2598), .Z(n1893) );
  NANDN U2431 ( .A(x[505]), .B(y[505]), .Z(n1889) );
  NANDN U2432 ( .A(x[504]), .B(y[504]), .Z(n1888) );
  AND U2433 ( .A(n1889), .B(n1888), .Z(n2604) );
  NANDN U2434 ( .A(y[502]), .B(x[502]), .Z(n1891) );
  NANDN U2435 ( .A(y[501]), .B(x[501]), .Z(n1890) );
  NAND U2436 ( .A(n1891), .B(n1890), .Z(n2023) );
  ANDN U2437 ( .B(n2604), .A(n2023), .Z(n1892) );
  AND U2438 ( .A(n1893), .B(n1892), .Z(n1896) );
  NANDN U2439 ( .A(x[491]), .B(y[491]), .Z(n1895) );
  NANDN U2440 ( .A(x[490]), .B(y[490]), .Z(n1894) );
  AND U2441 ( .A(n1895), .B(n1894), .Z(n2593) );
  AND U2442 ( .A(n1896), .B(n2593), .Z(n1903) );
  NANDN U2443 ( .A(x[295]), .B(y[295]), .Z(n2421) );
  ANDN U2444 ( .B(x[316]), .A(y[316]), .Z(n2438) );
  ANDN U2445 ( .B(n2421), .A(n2438), .Z(n1898) );
  NANDN U2446 ( .A(x[510]), .B(y[510]), .Z(n2610) );
  ANDN U2447 ( .B(x[511]), .A(y[511]), .Z(n2020) );
  ANDN U2448 ( .B(n2610), .A(n2020), .Z(n1897) );
  AND U2449 ( .A(n1898), .B(n1897), .Z(n1901) );
  NANDN U2450 ( .A(y[498]), .B(x[498]), .Z(n1900) );
  NANDN U2451 ( .A(y[497]), .B(x[497]), .Z(n1899) );
  NAND U2452 ( .A(n1900), .B(n1899), .Z(n2024) );
  ANDN U2453 ( .B(n1901), .A(n2024), .Z(n1902) );
  AND U2454 ( .A(n1903), .B(n1902), .Z(n1915) );
  NANDN U2455 ( .A(x[461]), .B(y[461]), .Z(n1905) );
  NANDN U2456 ( .A(x[460]), .B(y[460]), .Z(n1904) );
  AND U2457 ( .A(n1905), .B(n1904), .Z(n2565) );
  NANDN U2458 ( .A(y[468]), .B(x[468]), .Z(n1907) );
  NANDN U2459 ( .A(y[467]), .B(x[467]), .Z(n1906) );
  NAND U2460 ( .A(n1907), .B(n1906), .Z(n2031) );
  ANDN U2461 ( .B(n2565), .A(n2031), .Z(n1913) );
  NANDN U2462 ( .A(y[466]), .B(x[466]), .Z(n1909) );
  NANDN U2463 ( .A(y[465]), .B(x[465]), .Z(n1908) );
  AND U2464 ( .A(n1909), .B(n1908), .Z(n2570) );
  NANDN U2465 ( .A(y[462]), .B(x[462]), .Z(n1911) );
  NANDN U2466 ( .A(y[461]), .B(x[461]), .Z(n1910) );
  NAND U2467 ( .A(n1911), .B(n1910), .Z(n2566) );
  ANDN U2468 ( .B(n2570), .A(n2566), .Z(n1912) );
  AND U2469 ( .A(n1913), .B(n1912), .Z(n1914) );
  AND U2470 ( .A(n1915), .B(n1914), .Z(n1916) );
  AND U2471 ( .A(n1917), .B(n1916), .Z(n1965) );
  NANDN U2472 ( .A(x[415]), .B(y[415]), .Z(n1919) );
  NANDN U2473 ( .A(x[414]), .B(y[414]), .Z(n1918) );
  AND U2474 ( .A(n1919), .B(n1918), .Z(n2525) );
  NANDN U2475 ( .A(x[413]), .B(y[413]), .Z(n1921) );
  NANDN U2476 ( .A(x[412]), .B(y[412]), .Z(n1920) );
  AND U2477 ( .A(n1921), .B(n1920), .Z(n2524) );
  AND U2478 ( .A(n2525), .B(n2524), .Z(n1927) );
  NANDN U2479 ( .A(y[412]), .B(x[412]), .Z(n1923) );
  NANDN U2480 ( .A(y[411]), .B(x[411]), .Z(n1922) );
  AND U2481 ( .A(n1923), .B(n1922), .Z(n2523) );
  NANDN U2482 ( .A(y[406]), .B(x[406]), .Z(n1925) );
  NANDN U2483 ( .A(y[405]), .B(x[405]), .Z(n1924) );
  NAND U2484 ( .A(n1925), .B(n1924), .Z(n2047) );
  ANDN U2485 ( .B(n2523), .A(n2047), .Z(n1926) );
  AND U2486 ( .A(n1927), .B(n1926), .Z(n1939) );
  NANDN U2487 ( .A(x[405]), .B(y[405]), .Z(n1929) );
  NANDN U2488 ( .A(x[404]), .B(y[404]), .Z(n1928) );
  AND U2489 ( .A(n1929), .B(n1928), .Z(n2517) );
  NANDN U2490 ( .A(y[396]), .B(x[396]), .Z(n1931) );
  NANDN U2491 ( .A(y[395]), .B(x[395]), .Z(n1930) );
  NAND U2492 ( .A(n1931), .B(n1930), .Z(n2050) );
  ANDN U2493 ( .B(n2517), .A(n2050), .Z(n1937) );
  NANDN U2494 ( .A(y[404]), .B(x[404]), .Z(n1933) );
  NANDN U2495 ( .A(y[403]), .B(x[403]), .Z(n1932) );
  AND U2496 ( .A(n1933), .B(n1932), .Z(n2516) );
  NANDN U2497 ( .A(y[400]), .B(x[400]), .Z(n1935) );
  NANDN U2498 ( .A(y[399]), .B(x[399]), .Z(n1934) );
  NAND U2499 ( .A(n1935), .B(n1934), .Z(n2049) );
  ANDN U2500 ( .B(n2516), .A(n2049), .Z(n1936) );
  AND U2501 ( .A(n1937), .B(n1936), .Z(n1938) );
  AND U2502 ( .A(n1939), .B(n1938), .Z(n1963) );
  NANDN U2503 ( .A(y[422]), .B(x[422]), .Z(n1941) );
  NANDN U2504 ( .A(y[421]), .B(x[421]), .Z(n1940) );
  AND U2505 ( .A(n1941), .B(n1940), .Z(n2531) );
  NANDN U2506 ( .A(y[416]), .B(x[416]), .Z(n1943) );
  NANDN U2507 ( .A(y[415]), .B(x[415]), .Z(n1942) );
  NAND U2508 ( .A(n1943), .B(n1942), .Z(n2044) );
  ANDN U2509 ( .B(n2531), .A(n2044), .Z(n1949) );
  NANDN U2510 ( .A(x[421]), .B(y[421]), .Z(n1945) );
  NANDN U2511 ( .A(x[420]), .B(y[420]), .Z(n1944) );
  AND U2512 ( .A(n1945), .B(n1944), .Z(n2530) );
  NANDN U2513 ( .A(x[417]), .B(y[417]), .Z(n1947) );
  NANDN U2514 ( .A(x[416]), .B(y[416]), .Z(n1946) );
  AND U2515 ( .A(n1947), .B(n1946), .Z(n2527) );
  AND U2516 ( .A(n2530), .B(n2527), .Z(n1948) );
  AND U2517 ( .A(n1949), .B(n1948), .Z(n1961) );
  NANDN U2518 ( .A(x[403]), .B(y[403]), .Z(n1951) );
  NANDN U2519 ( .A(x[402]), .B(y[402]), .Z(n1950) );
  AND U2520 ( .A(n1951), .B(n1950), .Z(n2515) );
  NANDN U2521 ( .A(x[389]), .B(y[389]), .Z(n1953) );
  NANDN U2522 ( .A(x[388]), .B(y[388]), .Z(n1952) );
  AND U2523 ( .A(n1953), .B(n1952), .Z(n2505) );
  AND U2524 ( .A(n2515), .B(n2505), .Z(n1959) );
  NANDN U2525 ( .A(x[391]), .B(y[391]), .Z(n1955) );
  NANDN U2526 ( .A(x[390]), .B(y[390]), .Z(n1954) );
  AND U2527 ( .A(n1955), .B(n1954), .Z(n2506) );
  NANDN U2528 ( .A(y[392]), .B(x[392]), .Z(n1957) );
  NANDN U2529 ( .A(y[391]), .B(x[391]), .Z(n1956) );
  NAND U2530 ( .A(n1957), .B(n1956), .Z(n2507) );
  ANDN U2531 ( .B(n2506), .A(n2507), .Z(n1958) );
  AND U2532 ( .A(n1959), .B(n1958), .Z(n1960) );
  AND U2533 ( .A(n1961), .B(n1960), .Z(n1962) );
  AND U2534 ( .A(n1963), .B(n1962), .Z(n1964) );
  AND U2535 ( .A(n1965), .B(n1964), .Z(n1966) );
  AND U2536 ( .A(n1967), .B(n1966), .Z(n2015) );
  NANDN U2537 ( .A(y[337]), .B(x[337]), .Z(n1969) );
  NANDN U2538 ( .A(y[336]), .B(x[336]), .Z(n1968) );
  AND U2539 ( .A(n1969), .B(n1968), .Z(n2459) );
  NANDN U2540 ( .A(y[335]), .B(x[335]), .Z(n1971) );
  NANDN U2541 ( .A(y[334]), .B(x[334]), .Z(n1970) );
  NAND U2542 ( .A(n1971), .B(n1970), .Z(n2457) );
  ANDN U2543 ( .B(n2459), .A(n2457), .Z(n1977) );
  NANDN U2544 ( .A(x[342]), .B(y[342]), .Z(n1973) );
  NANDN U2545 ( .A(x[341]), .B(y[341]), .Z(n1972) );
  AND U2546 ( .A(n1973), .B(n1972), .Z(n2463) );
  NANDN U2547 ( .A(x[336]), .B(y[336]), .Z(n1975) );
  NANDN U2548 ( .A(x[335]), .B(y[335]), .Z(n1974) );
  AND U2549 ( .A(n1975), .B(n1974), .Z(n2458) );
  AND U2550 ( .A(n2463), .B(n2458), .Z(n1976) );
  AND U2551 ( .A(n1977), .B(n1976), .Z(n1989) );
  NANDN U2552 ( .A(x[332]), .B(y[332]), .Z(n1979) );
  NANDN U2553 ( .A(x[331]), .B(y[331]), .Z(n1978) );
  AND U2554 ( .A(n1979), .B(n1978), .Z(n2455) );
  NANDN U2555 ( .A(x[323]), .B(y[323]), .Z(n1981) );
  NANDN U2556 ( .A(x[322]), .B(y[322]), .Z(n1980) );
  AND U2557 ( .A(n1981), .B(n1980), .Z(n2446) );
  AND U2558 ( .A(n2455), .B(n2446), .Z(n1987) );
  NANDN U2559 ( .A(y[331]), .B(x[331]), .Z(n1983) );
  NANDN U2560 ( .A(y[330]), .B(x[330]), .Z(n1982) );
  AND U2561 ( .A(n1983), .B(n1982), .Z(n2453) );
  NANDN U2562 ( .A(y[326]), .B(x[326]), .Z(n1985) );
  NANDN U2563 ( .A(y[325]), .B(x[325]), .Z(n1984) );
  NAND U2564 ( .A(n1985), .B(n1984), .Z(n2070) );
  ANDN U2565 ( .B(n2453), .A(n2070), .Z(n1986) );
  AND U2566 ( .A(n1987), .B(n1986), .Z(n1988) );
  AND U2567 ( .A(n1989), .B(n1988), .Z(n2013) );
  NANDN U2568 ( .A(y[353]), .B(x[353]), .Z(n1991) );
  NANDN U2569 ( .A(y[352]), .B(x[352]), .Z(n1990) );
  AND U2570 ( .A(n1991), .B(n1990), .Z(n2471) );
  NANDN U2571 ( .A(y[341]), .B(x[341]), .Z(n1993) );
  NANDN U2572 ( .A(y[340]), .B(x[340]), .Z(n1992) );
  NAND U2573 ( .A(n1993), .B(n1992), .Z(n2462) );
  ANDN U2574 ( .B(n2471), .A(n2462), .Z(n1999) );
  NANDN U2575 ( .A(x[344]), .B(y[344]), .Z(n1995) );
  NANDN U2576 ( .A(x[343]), .B(y[343]), .Z(n1994) );
  AND U2577 ( .A(n1995), .B(n1994), .Z(n2464) );
  NANDN U2578 ( .A(y[343]), .B(x[343]), .Z(n1997) );
  NANDN U2579 ( .A(y[342]), .B(x[342]), .Z(n1996) );
  NAND U2580 ( .A(n1997), .B(n1996), .Z(n2066) );
  ANDN U2581 ( .B(n2464), .A(n2066), .Z(n1998) );
  AND U2582 ( .A(n1999), .B(n1998), .Z(n2011) );
  NANDN U2583 ( .A(x[321]), .B(y[321]), .Z(n2001) );
  NANDN U2584 ( .A(x[320]), .B(y[320]), .Z(n2000) );
  AND U2585 ( .A(n2001), .B(n2000), .Z(n2445) );
  NANDN U2586 ( .A(x[303]), .B(y[303]), .Z(n2003) );
  NANDN U2587 ( .A(x[302]), .B(y[302]), .Z(n2002) );
  AND U2588 ( .A(n2003), .B(n2002), .Z(n2426) );
  AND U2589 ( .A(n2445), .B(n2426), .Z(n2009) );
  NANDN U2590 ( .A(y[320]), .B(x[320]), .Z(n2005) );
  NANDN U2591 ( .A(y[319]), .B(x[319]), .Z(n2004) );
  AND U2592 ( .A(n2005), .B(n2004), .Z(n2444) );
  NANDN U2593 ( .A(y[322]), .B(x[322]), .Z(n2007) );
  NANDN U2594 ( .A(y[321]), .B(x[321]), .Z(n2006) );
  NAND U2595 ( .A(n2007), .B(n2006), .Z(n2071) );
  ANDN U2596 ( .B(n2444), .A(n2071), .Z(n2008) );
  AND U2597 ( .A(n2009), .B(n2008), .Z(n2010) );
  AND U2598 ( .A(n2011), .B(n2010), .Z(n2012) );
  AND U2599 ( .A(n2013), .B(n2012), .Z(n2014) );
  AND U2600 ( .A(n2015), .B(n2014), .Z(n2016) );
  AND U2601 ( .A(n2017), .B(n2016), .Z(n2018) );
  NAND U2602 ( .A(n2019), .B(n2018), .Z(n2611) );
  OR U2603 ( .A(n2611), .B(ebreg), .Z(n5) );
  IV U2604 ( .A(n2023), .Z(n2602) );
  IV U2605 ( .A(n2055), .Z(n2490) );
  IV U2606 ( .A(n2060), .Z(n2478) );
  IV U2607 ( .A(n2076), .Z(n2428) );
  IV U2608 ( .A(n2089), .Z(n2393) );
  IV U2609 ( .A(n2188), .Z(n2189) );
  IV U2610 ( .A(n2290), .Z(n2291) );
  IV U2611 ( .A(n2316), .Z(n2317) );
  IV U2612 ( .A(n2366), .Z(n2367) );
  IV U2613 ( .A(n2379), .Z(n2381) );
  ANDN U2614 ( .B(x[255]), .A(y[255]), .Z(n2380) );
  IV U2615 ( .A(n2549), .Z(n2550) );
  IV U2616 ( .A(n2589), .Z(n2590) );
endmodule

