
module sum_N1024_CC4 ( clk, rst, a, b, c );
  input [255:0] a;
  input [255:0] b;
  output [255:0] c;
  input clk, rst;
  wire   N514, N515, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801;
  wire   [1:0] carry_on;

  DFF \carry_on_reg[1]  ( .D(N515), .CLK(clk), .RST(rst), .Q(carry_on[1]) );
  DFF \carry_on_reg[0]  ( .D(N514), .CLK(clk), .RST(rst), .Q(carry_on[0]) );
  DFF \rc_reg[255]  ( .D(n1024), .CLK(clk), .RST(1'b0), .Q(c[255]) );
  DFF \rc_reg[254]  ( .D(n1023), .CLK(clk), .RST(1'b0), .Q(c[254]) );
  DFF \rc_reg[253]  ( .D(n1022), .CLK(clk), .RST(1'b0), .Q(c[253]) );
  DFF \rc_reg[252]  ( .D(n1021), .CLK(clk), .RST(1'b0), .Q(c[252]) );
  DFF \rc_reg[251]  ( .D(n1020), .CLK(clk), .RST(1'b0), .Q(c[251]) );
  DFF \rc_reg[250]  ( .D(n1019), .CLK(clk), .RST(1'b0), .Q(c[250]) );
  DFF \rc_reg[249]  ( .D(n1018), .CLK(clk), .RST(1'b0), .Q(c[249]) );
  DFF \rc_reg[248]  ( .D(n1017), .CLK(clk), .RST(1'b0), .Q(c[248]) );
  DFF \rc_reg[247]  ( .D(n1016), .CLK(clk), .RST(1'b0), .Q(c[247]) );
  DFF \rc_reg[246]  ( .D(n1015), .CLK(clk), .RST(1'b0), .Q(c[246]) );
  DFF \rc_reg[245]  ( .D(n1014), .CLK(clk), .RST(1'b0), .Q(c[245]) );
  DFF \rc_reg[244]  ( .D(n1013), .CLK(clk), .RST(1'b0), .Q(c[244]) );
  DFF \rc_reg[243]  ( .D(n1012), .CLK(clk), .RST(1'b0), .Q(c[243]) );
  DFF \rc_reg[242]  ( .D(n1011), .CLK(clk), .RST(1'b0), .Q(c[242]) );
  DFF \rc_reg[241]  ( .D(n1010), .CLK(clk), .RST(1'b0), .Q(c[241]) );
  DFF \rc_reg[240]  ( .D(n1009), .CLK(clk), .RST(1'b0), .Q(c[240]) );
  DFF \rc_reg[239]  ( .D(n1008), .CLK(clk), .RST(1'b0), .Q(c[239]) );
  DFF \rc_reg[238]  ( .D(n1007), .CLK(clk), .RST(1'b0), .Q(c[238]) );
  DFF \rc_reg[237]  ( .D(n1006), .CLK(clk), .RST(1'b0), .Q(c[237]) );
  DFF \rc_reg[236]  ( .D(n1005), .CLK(clk), .RST(1'b0), .Q(c[236]) );
  DFF \rc_reg[235]  ( .D(n1004), .CLK(clk), .RST(1'b0), .Q(c[235]) );
  DFF \rc_reg[234]  ( .D(n1003), .CLK(clk), .RST(1'b0), .Q(c[234]) );
  DFF \rc_reg[233]  ( .D(n1002), .CLK(clk), .RST(1'b0), .Q(c[233]) );
  DFF \rc_reg[232]  ( .D(n1001), .CLK(clk), .RST(1'b0), .Q(c[232]) );
  DFF \rc_reg[231]  ( .D(n1000), .CLK(clk), .RST(1'b0), .Q(c[231]) );
  DFF \rc_reg[230]  ( .D(n999), .CLK(clk), .RST(1'b0), .Q(c[230]) );
  DFF \rc_reg[229]  ( .D(n998), .CLK(clk), .RST(1'b0), .Q(c[229]) );
  DFF \rc_reg[228]  ( .D(n997), .CLK(clk), .RST(1'b0), .Q(c[228]) );
  DFF \rc_reg[227]  ( .D(n996), .CLK(clk), .RST(1'b0), .Q(c[227]) );
  DFF \rc_reg[226]  ( .D(n995), .CLK(clk), .RST(1'b0), .Q(c[226]) );
  DFF \rc_reg[225]  ( .D(n994), .CLK(clk), .RST(1'b0), .Q(c[225]) );
  DFF \rc_reg[224]  ( .D(n993), .CLK(clk), .RST(1'b0), .Q(c[224]) );
  DFF \rc_reg[223]  ( .D(n992), .CLK(clk), .RST(1'b0), .Q(c[223]) );
  DFF \rc_reg[222]  ( .D(n991), .CLK(clk), .RST(1'b0), .Q(c[222]) );
  DFF \rc_reg[221]  ( .D(n990), .CLK(clk), .RST(1'b0), .Q(c[221]) );
  DFF \rc_reg[220]  ( .D(n989), .CLK(clk), .RST(1'b0), .Q(c[220]) );
  DFF \rc_reg[219]  ( .D(n988), .CLK(clk), .RST(1'b0), .Q(c[219]) );
  DFF \rc_reg[218]  ( .D(n987), .CLK(clk), .RST(1'b0), .Q(c[218]) );
  DFF \rc_reg[217]  ( .D(n986), .CLK(clk), .RST(1'b0), .Q(c[217]) );
  DFF \rc_reg[216]  ( .D(n985), .CLK(clk), .RST(1'b0), .Q(c[216]) );
  DFF \rc_reg[215]  ( .D(n984), .CLK(clk), .RST(1'b0), .Q(c[215]) );
  DFF \rc_reg[214]  ( .D(n983), .CLK(clk), .RST(1'b0), .Q(c[214]) );
  DFF \rc_reg[213]  ( .D(n982), .CLK(clk), .RST(1'b0), .Q(c[213]) );
  DFF \rc_reg[212]  ( .D(n981), .CLK(clk), .RST(1'b0), .Q(c[212]) );
  DFF \rc_reg[211]  ( .D(n980), .CLK(clk), .RST(1'b0), .Q(c[211]) );
  DFF \rc_reg[210]  ( .D(n979), .CLK(clk), .RST(1'b0), .Q(c[210]) );
  DFF \rc_reg[209]  ( .D(n978), .CLK(clk), .RST(1'b0), .Q(c[209]) );
  DFF \rc_reg[208]  ( .D(n977), .CLK(clk), .RST(1'b0), .Q(c[208]) );
  DFF \rc_reg[207]  ( .D(n976), .CLK(clk), .RST(1'b0), .Q(c[207]) );
  DFF \rc_reg[206]  ( .D(n975), .CLK(clk), .RST(1'b0), .Q(c[206]) );
  DFF \rc_reg[205]  ( .D(n974), .CLK(clk), .RST(1'b0), .Q(c[205]) );
  DFF \rc_reg[204]  ( .D(n973), .CLK(clk), .RST(1'b0), .Q(c[204]) );
  DFF \rc_reg[203]  ( .D(n972), .CLK(clk), .RST(1'b0), .Q(c[203]) );
  DFF \rc_reg[202]  ( .D(n971), .CLK(clk), .RST(1'b0), .Q(c[202]) );
  DFF \rc_reg[201]  ( .D(n970), .CLK(clk), .RST(1'b0), .Q(c[201]) );
  DFF \rc_reg[200]  ( .D(n969), .CLK(clk), .RST(1'b0), .Q(c[200]) );
  DFF \rc_reg[199]  ( .D(n968), .CLK(clk), .RST(1'b0), .Q(c[199]) );
  DFF \rc_reg[198]  ( .D(n967), .CLK(clk), .RST(1'b0), .Q(c[198]) );
  DFF \rc_reg[197]  ( .D(n966), .CLK(clk), .RST(1'b0), .Q(c[197]) );
  DFF \rc_reg[196]  ( .D(n965), .CLK(clk), .RST(1'b0), .Q(c[196]) );
  DFF \rc_reg[195]  ( .D(n964), .CLK(clk), .RST(1'b0), .Q(c[195]) );
  DFF \rc_reg[194]  ( .D(n963), .CLK(clk), .RST(1'b0), .Q(c[194]) );
  DFF \rc_reg[193]  ( .D(n962), .CLK(clk), .RST(1'b0), .Q(c[193]) );
  DFF \rc_reg[192]  ( .D(n961), .CLK(clk), .RST(1'b0), .Q(c[192]) );
  DFF \rc_reg[191]  ( .D(n960), .CLK(clk), .RST(1'b0), .Q(c[191]) );
  DFF \rc_reg[190]  ( .D(n959), .CLK(clk), .RST(1'b0), .Q(c[190]) );
  DFF \rc_reg[189]  ( .D(n958), .CLK(clk), .RST(1'b0), .Q(c[189]) );
  DFF \rc_reg[188]  ( .D(n957), .CLK(clk), .RST(1'b0), .Q(c[188]) );
  DFF \rc_reg[187]  ( .D(n956), .CLK(clk), .RST(1'b0), .Q(c[187]) );
  DFF \rc_reg[186]  ( .D(n955), .CLK(clk), .RST(1'b0), .Q(c[186]) );
  DFF \rc_reg[185]  ( .D(n954), .CLK(clk), .RST(1'b0), .Q(c[185]) );
  DFF \rc_reg[184]  ( .D(n953), .CLK(clk), .RST(1'b0), .Q(c[184]) );
  DFF \rc_reg[183]  ( .D(n952), .CLK(clk), .RST(1'b0), .Q(c[183]) );
  DFF \rc_reg[182]  ( .D(n951), .CLK(clk), .RST(1'b0), .Q(c[182]) );
  DFF \rc_reg[181]  ( .D(n950), .CLK(clk), .RST(1'b0), .Q(c[181]) );
  DFF \rc_reg[180]  ( .D(n949), .CLK(clk), .RST(1'b0), .Q(c[180]) );
  DFF \rc_reg[179]  ( .D(n948), .CLK(clk), .RST(1'b0), .Q(c[179]) );
  DFF \rc_reg[178]  ( .D(n947), .CLK(clk), .RST(1'b0), .Q(c[178]) );
  DFF \rc_reg[177]  ( .D(n946), .CLK(clk), .RST(1'b0), .Q(c[177]) );
  DFF \rc_reg[176]  ( .D(n945), .CLK(clk), .RST(1'b0), .Q(c[176]) );
  DFF \rc_reg[175]  ( .D(n944), .CLK(clk), .RST(1'b0), .Q(c[175]) );
  DFF \rc_reg[174]  ( .D(n943), .CLK(clk), .RST(1'b0), .Q(c[174]) );
  DFF \rc_reg[173]  ( .D(n942), .CLK(clk), .RST(1'b0), .Q(c[173]) );
  DFF \rc_reg[172]  ( .D(n941), .CLK(clk), .RST(1'b0), .Q(c[172]) );
  DFF \rc_reg[171]  ( .D(n940), .CLK(clk), .RST(1'b0), .Q(c[171]) );
  DFF \rc_reg[170]  ( .D(n939), .CLK(clk), .RST(1'b0), .Q(c[170]) );
  DFF \rc_reg[169]  ( .D(n938), .CLK(clk), .RST(1'b0), .Q(c[169]) );
  DFF \rc_reg[168]  ( .D(n937), .CLK(clk), .RST(1'b0), .Q(c[168]) );
  DFF \rc_reg[167]  ( .D(n936), .CLK(clk), .RST(1'b0), .Q(c[167]) );
  DFF \rc_reg[166]  ( .D(n935), .CLK(clk), .RST(1'b0), .Q(c[166]) );
  DFF \rc_reg[165]  ( .D(n934), .CLK(clk), .RST(1'b0), .Q(c[165]) );
  DFF \rc_reg[164]  ( .D(n933), .CLK(clk), .RST(1'b0), .Q(c[164]) );
  DFF \rc_reg[163]  ( .D(n932), .CLK(clk), .RST(1'b0), .Q(c[163]) );
  DFF \rc_reg[162]  ( .D(n931), .CLK(clk), .RST(1'b0), .Q(c[162]) );
  DFF \rc_reg[161]  ( .D(n930), .CLK(clk), .RST(1'b0), .Q(c[161]) );
  DFF \rc_reg[160]  ( .D(n929), .CLK(clk), .RST(1'b0), .Q(c[160]) );
  DFF \rc_reg[159]  ( .D(n928), .CLK(clk), .RST(1'b0), .Q(c[159]) );
  DFF \rc_reg[158]  ( .D(n927), .CLK(clk), .RST(1'b0), .Q(c[158]) );
  DFF \rc_reg[157]  ( .D(n926), .CLK(clk), .RST(1'b0), .Q(c[157]) );
  DFF \rc_reg[156]  ( .D(n925), .CLK(clk), .RST(1'b0), .Q(c[156]) );
  DFF \rc_reg[155]  ( .D(n924), .CLK(clk), .RST(1'b0), .Q(c[155]) );
  DFF \rc_reg[154]  ( .D(n923), .CLK(clk), .RST(1'b0), .Q(c[154]) );
  DFF \rc_reg[153]  ( .D(n922), .CLK(clk), .RST(1'b0), .Q(c[153]) );
  DFF \rc_reg[152]  ( .D(n921), .CLK(clk), .RST(1'b0), .Q(c[152]) );
  DFF \rc_reg[151]  ( .D(n920), .CLK(clk), .RST(1'b0), .Q(c[151]) );
  DFF \rc_reg[150]  ( .D(n919), .CLK(clk), .RST(1'b0), .Q(c[150]) );
  DFF \rc_reg[149]  ( .D(n918), .CLK(clk), .RST(1'b0), .Q(c[149]) );
  DFF \rc_reg[148]  ( .D(n917), .CLK(clk), .RST(1'b0), .Q(c[148]) );
  DFF \rc_reg[147]  ( .D(n916), .CLK(clk), .RST(1'b0), .Q(c[147]) );
  DFF \rc_reg[146]  ( .D(n915), .CLK(clk), .RST(1'b0), .Q(c[146]) );
  DFF \rc_reg[145]  ( .D(n914), .CLK(clk), .RST(1'b0), .Q(c[145]) );
  DFF \rc_reg[144]  ( .D(n913), .CLK(clk), .RST(1'b0), .Q(c[144]) );
  DFF \rc_reg[143]  ( .D(n912), .CLK(clk), .RST(1'b0), .Q(c[143]) );
  DFF \rc_reg[142]  ( .D(n911), .CLK(clk), .RST(1'b0), .Q(c[142]) );
  DFF \rc_reg[141]  ( .D(n910), .CLK(clk), .RST(1'b0), .Q(c[141]) );
  DFF \rc_reg[140]  ( .D(n909), .CLK(clk), .RST(1'b0), .Q(c[140]) );
  DFF \rc_reg[139]  ( .D(n908), .CLK(clk), .RST(1'b0), .Q(c[139]) );
  DFF \rc_reg[138]  ( .D(n907), .CLK(clk), .RST(1'b0), .Q(c[138]) );
  DFF \rc_reg[137]  ( .D(n906), .CLK(clk), .RST(1'b0), .Q(c[137]) );
  DFF \rc_reg[136]  ( .D(n905), .CLK(clk), .RST(1'b0), .Q(c[136]) );
  DFF \rc_reg[135]  ( .D(n904), .CLK(clk), .RST(1'b0), .Q(c[135]) );
  DFF \rc_reg[134]  ( .D(n903), .CLK(clk), .RST(1'b0), .Q(c[134]) );
  DFF \rc_reg[133]  ( .D(n902), .CLK(clk), .RST(1'b0), .Q(c[133]) );
  DFF \rc_reg[132]  ( .D(n901), .CLK(clk), .RST(1'b0), .Q(c[132]) );
  DFF \rc_reg[131]  ( .D(n900), .CLK(clk), .RST(1'b0), .Q(c[131]) );
  DFF \rc_reg[130]  ( .D(n899), .CLK(clk), .RST(1'b0), .Q(c[130]) );
  DFF \rc_reg[129]  ( .D(n898), .CLK(clk), .RST(1'b0), .Q(c[129]) );
  DFF \rc_reg[128]  ( .D(n897), .CLK(clk), .RST(1'b0), .Q(c[128]) );
  DFF \rc_reg[127]  ( .D(n896), .CLK(clk), .RST(1'b0), .Q(c[127]) );
  DFF \rc_reg[126]  ( .D(n895), .CLK(clk), .RST(1'b0), .Q(c[126]) );
  DFF \rc_reg[125]  ( .D(n894), .CLK(clk), .RST(1'b0), .Q(c[125]) );
  DFF \rc_reg[124]  ( .D(n893), .CLK(clk), .RST(1'b0), .Q(c[124]) );
  DFF \rc_reg[123]  ( .D(n892), .CLK(clk), .RST(1'b0), .Q(c[123]) );
  DFF \rc_reg[122]  ( .D(n891), .CLK(clk), .RST(1'b0), .Q(c[122]) );
  DFF \rc_reg[121]  ( .D(n890), .CLK(clk), .RST(1'b0), .Q(c[121]) );
  DFF \rc_reg[120]  ( .D(n889), .CLK(clk), .RST(1'b0), .Q(c[120]) );
  DFF \rc_reg[119]  ( .D(n888), .CLK(clk), .RST(1'b0), .Q(c[119]) );
  DFF \rc_reg[118]  ( .D(n887), .CLK(clk), .RST(1'b0), .Q(c[118]) );
  DFF \rc_reg[117]  ( .D(n886), .CLK(clk), .RST(1'b0), .Q(c[117]) );
  DFF \rc_reg[116]  ( .D(n885), .CLK(clk), .RST(1'b0), .Q(c[116]) );
  DFF \rc_reg[115]  ( .D(n884), .CLK(clk), .RST(1'b0), .Q(c[115]) );
  DFF \rc_reg[114]  ( .D(n883), .CLK(clk), .RST(1'b0), .Q(c[114]) );
  DFF \rc_reg[113]  ( .D(n882), .CLK(clk), .RST(1'b0), .Q(c[113]) );
  DFF \rc_reg[112]  ( .D(n881), .CLK(clk), .RST(1'b0), .Q(c[112]) );
  DFF \rc_reg[111]  ( .D(n880), .CLK(clk), .RST(1'b0), .Q(c[111]) );
  DFF \rc_reg[110]  ( .D(n879), .CLK(clk), .RST(1'b0), .Q(c[110]) );
  DFF \rc_reg[109]  ( .D(n878), .CLK(clk), .RST(1'b0), .Q(c[109]) );
  DFF \rc_reg[108]  ( .D(n877), .CLK(clk), .RST(1'b0), .Q(c[108]) );
  DFF \rc_reg[107]  ( .D(n876), .CLK(clk), .RST(1'b0), .Q(c[107]) );
  DFF \rc_reg[106]  ( .D(n875), .CLK(clk), .RST(1'b0), .Q(c[106]) );
  DFF \rc_reg[105]  ( .D(n874), .CLK(clk), .RST(1'b0), .Q(c[105]) );
  DFF \rc_reg[104]  ( .D(n873), .CLK(clk), .RST(1'b0), .Q(c[104]) );
  DFF \rc_reg[103]  ( .D(n872), .CLK(clk), .RST(1'b0), .Q(c[103]) );
  DFF \rc_reg[102]  ( .D(n871), .CLK(clk), .RST(1'b0), .Q(c[102]) );
  DFF \rc_reg[101]  ( .D(n870), .CLK(clk), .RST(1'b0), .Q(c[101]) );
  DFF \rc_reg[100]  ( .D(n869), .CLK(clk), .RST(1'b0), .Q(c[100]) );
  DFF \rc_reg[99]  ( .D(n868), .CLK(clk), .RST(1'b0), .Q(c[99]) );
  DFF \rc_reg[98]  ( .D(n867), .CLK(clk), .RST(1'b0), .Q(c[98]) );
  DFF \rc_reg[97]  ( .D(n866), .CLK(clk), .RST(1'b0), .Q(c[97]) );
  DFF \rc_reg[96]  ( .D(n865), .CLK(clk), .RST(1'b0), .Q(c[96]) );
  DFF \rc_reg[95]  ( .D(n864), .CLK(clk), .RST(1'b0), .Q(c[95]) );
  DFF \rc_reg[94]  ( .D(n863), .CLK(clk), .RST(1'b0), .Q(c[94]) );
  DFF \rc_reg[93]  ( .D(n862), .CLK(clk), .RST(1'b0), .Q(c[93]) );
  DFF \rc_reg[92]  ( .D(n861), .CLK(clk), .RST(1'b0), .Q(c[92]) );
  DFF \rc_reg[91]  ( .D(n860), .CLK(clk), .RST(1'b0), .Q(c[91]) );
  DFF \rc_reg[90]  ( .D(n859), .CLK(clk), .RST(1'b0), .Q(c[90]) );
  DFF \rc_reg[89]  ( .D(n858), .CLK(clk), .RST(1'b0), .Q(c[89]) );
  DFF \rc_reg[88]  ( .D(n857), .CLK(clk), .RST(1'b0), .Q(c[88]) );
  DFF \rc_reg[87]  ( .D(n856), .CLK(clk), .RST(1'b0), .Q(c[87]) );
  DFF \rc_reg[86]  ( .D(n855), .CLK(clk), .RST(1'b0), .Q(c[86]) );
  DFF \rc_reg[85]  ( .D(n854), .CLK(clk), .RST(1'b0), .Q(c[85]) );
  DFF \rc_reg[84]  ( .D(n853), .CLK(clk), .RST(1'b0), .Q(c[84]) );
  DFF \rc_reg[83]  ( .D(n852), .CLK(clk), .RST(1'b0), .Q(c[83]) );
  DFF \rc_reg[82]  ( .D(n851), .CLK(clk), .RST(1'b0), .Q(c[82]) );
  DFF \rc_reg[81]  ( .D(n850), .CLK(clk), .RST(1'b0), .Q(c[81]) );
  DFF \rc_reg[80]  ( .D(n849), .CLK(clk), .RST(1'b0), .Q(c[80]) );
  DFF \rc_reg[79]  ( .D(n848), .CLK(clk), .RST(1'b0), .Q(c[79]) );
  DFF \rc_reg[78]  ( .D(n847), .CLK(clk), .RST(1'b0), .Q(c[78]) );
  DFF \rc_reg[77]  ( .D(n846), .CLK(clk), .RST(1'b0), .Q(c[77]) );
  DFF \rc_reg[76]  ( .D(n845), .CLK(clk), .RST(1'b0), .Q(c[76]) );
  DFF \rc_reg[75]  ( .D(n844), .CLK(clk), .RST(1'b0), .Q(c[75]) );
  DFF \rc_reg[74]  ( .D(n843), .CLK(clk), .RST(1'b0), .Q(c[74]) );
  DFF \rc_reg[73]  ( .D(n842), .CLK(clk), .RST(1'b0), .Q(c[73]) );
  DFF \rc_reg[72]  ( .D(n841), .CLK(clk), .RST(1'b0), .Q(c[72]) );
  DFF \rc_reg[71]  ( .D(n840), .CLK(clk), .RST(1'b0), .Q(c[71]) );
  DFF \rc_reg[70]  ( .D(n839), .CLK(clk), .RST(1'b0), .Q(c[70]) );
  DFF \rc_reg[69]  ( .D(n838), .CLK(clk), .RST(1'b0), .Q(c[69]) );
  DFF \rc_reg[68]  ( .D(n837), .CLK(clk), .RST(1'b0), .Q(c[68]) );
  DFF \rc_reg[67]  ( .D(n836), .CLK(clk), .RST(1'b0), .Q(c[67]) );
  DFF \rc_reg[66]  ( .D(n835), .CLK(clk), .RST(1'b0), .Q(c[66]) );
  DFF \rc_reg[65]  ( .D(n834), .CLK(clk), .RST(1'b0), .Q(c[65]) );
  DFF \rc_reg[64]  ( .D(n833), .CLK(clk), .RST(1'b0), .Q(c[64]) );
  DFF \rc_reg[63]  ( .D(n832), .CLK(clk), .RST(1'b0), .Q(c[63]) );
  DFF \rc_reg[62]  ( .D(n831), .CLK(clk), .RST(1'b0), .Q(c[62]) );
  DFF \rc_reg[61]  ( .D(n830), .CLK(clk), .RST(1'b0), .Q(c[61]) );
  DFF \rc_reg[60]  ( .D(n829), .CLK(clk), .RST(1'b0), .Q(c[60]) );
  DFF \rc_reg[59]  ( .D(n828), .CLK(clk), .RST(1'b0), .Q(c[59]) );
  DFF \rc_reg[58]  ( .D(n827), .CLK(clk), .RST(1'b0), .Q(c[58]) );
  DFF \rc_reg[57]  ( .D(n826), .CLK(clk), .RST(1'b0), .Q(c[57]) );
  DFF \rc_reg[56]  ( .D(n825), .CLK(clk), .RST(1'b0), .Q(c[56]) );
  DFF \rc_reg[55]  ( .D(n824), .CLK(clk), .RST(1'b0), .Q(c[55]) );
  DFF \rc_reg[54]  ( .D(n823), .CLK(clk), .RST(1'b0), .Q(c[54]) );
  DFF \rc_reg[53]  ( .D(n822), .CLK(clk), .RST(1'b0), .Q(c[53]) );
  DFF \rc_reg[52]  ( .D(n821), .CLK(clk), .RST(1'b0), .Q(c[52]) );
  DFF \rc_reg[51]  ( .D(n820), .CLK(clk), .RST(1'b0), .Q(c[51]) );
  DFF \rc_reg[50]  ( .D(n819), .CLK(clk), .RST(1'b0), .Q(c[50]) );
  DFF \rc_reg[49]  ( .D(n818), .CLK(clk), .RST(1'b0), .Q(c[49]) );
  DFF \rc_reg[48]  ( .D(n817), .CLK(clk), .RST(1'b0), .Q(c[48]) );
  DFF \rc_reg[47]  ( .D(n816), .CLK(clk), .RST(1'b0), .Q(c[47]) );
  DFF \rc_reg[46]  ( .D(n815), .CLK(clk), .RST(1'b0), .Q(c[46]) );
  DFF \rc_reg[45]  ( .D(n814), .CLK(clk), .RST(1'b0), .Q(c[45]) );
  DFF \rc_reg[44]  ( .D(n813), .CLK(clk), .RST(1'b0), .Q(c[44]) );
  DFF \rc_reg[43]  ( .D(n812), .CLK(clk), .RST(1'b0), .Q(c[43]) );
  DFF \rc_reg[42]  ( .D(n811), .CLK(clk), .RST(1'b0), .Q(c[42]) );
  DFF \rc_reg[41]  ( .D(n810), .CLK(clk), .RST(1'b0), .Q(c[41]) );
  DFF \rc_reg[40]  ( .D(n809), .CLK(clk), .RST(1'b0), .Q(c[40]) );
  DFF \rc_reg[39]  ( .D(n808), .CLK(clk), .RST(1'b0), .Q(c[39]) );
  DFF \rc_reg[38]  ( .D(n807), .CLK(clk), .RST(1'b0), .Q(c[38]) );
  DFF \rc_reg[37]  ( .D(n806), .CLK(clk), .RST(1'b0), .Q(c[37]) );
  DFF \rc_reg[36]  ( .D(n805), .CLK(clk), .RST(1'b0), .Q(c[36]) );
  DFF \rc_reg[35]  ( .D(n804), .CLK(clk), .RST(1'b0), .Q(c[35]) );
  DFF \rc_reg[34]  ( .D(n803), .CLK(clk), .RST(1'b0), .Q(c[34]) );
  DFF \rc_reg[33]  ( .D(n802), .CLK(clk), .RST(1'b0), .Q(c[33]) );
  DFF \rc_reg[32]  ( .D(n801), .CLK(clk), .RST(1'b0), .Q(c[32]) );
  DFF \rc_reg[31]  ( .D(n800), .CLK(clk), .RST(1'b0), .Q(c[31]) );
  DFF \rc_reg[30]  ( .D(n799), .CLK(clk), .RST(1'b0), .Q(c[30]) );
  DFF \rc_reg[29]  ( .D(n798), .CLK(clk), .RST(1'b0), .Q(c[29]) );
  DFF \rc_reg[28]  ( .D(n797), .CLK(clk), .RST(1'b0), .Q(c[28]) );
  DFF \rc_reg[27]  ( .D(n796), .CLK(clk), .RST(1'b0), .Q(c[27]) );
  DFF \rc_reg[26]  ( .D(n795), .CLK(clk), .RST(1'b0), .Q(c[26]) );
  DFF \rc_reg[25]  ( .D(n794), .CLK(clk), .RST(1'b0), .Q(c[25]) );
  DFF \rc_reg[24]  ( .D(n793), .CLK(clk), .RST(1'b0), .Q(c[24]) );
  DFF \rc_reg[23]  ( .D(n792), .CLK(clk), .RST(1'b0), .Q(c[23]) );
  DFF \rc_reg[22]  ( .D(n791), .CLK(clk), .RST(1'b0), .Q(c[22]) );
  DFF \rc_reg[21]  ( .D(n790), .CLK(clk), .RST(1'b0), .Q(c[21]) );
  DFF \rc_reg[20]  ( .D(n789), .CLK(clk), .RST(1'b0), .Q(c[20]) );
  DFF \rc_reg[19]  ( .D(n788), .CLK(clk), .RST(1'b0), .Q(c[19]) );
  DFF \rc_reg[18]  ( .D(n787), .CLK(clk), .RST(1'b0), .Q(c[18]) );
  DFF \rc_reg[17]  ( .D(n786), .CLK(clk), .RST(1'b0), .Q(c[17]) );
  DFF \rc_reg[16]  ( .D(n785), .CLK(clk), .RST(1'b0), .Q(c[16]) );
  DFF \rc_reg[15]  ( .D(n784), .CLK(clk), .RST(1'b0), .Q(c[15]) );
  DFF \rc_reg[14]  ( .D(n783), .CLK(clk), .RST(1'b0), .Q(c[14]) );
  DFF \rc_reg[13]  ( .D(n782), .CLK(clk), .RST(1'b0), .Q(c[13]) );
  DFF \rc_reg[12]  ( .D(n781), .CLK(clk), .RST(1'b0), .Q(c[12]) );
  DFF \rc_reg[11]  ( .D(n780), .CLK(clk), .RST(1'b0), .Q(c[11]) );
  DFF \rc_reg[10]  ( .D(n779), .CLK(clk), .RST(1'b0), .Q(c[10]) );
  DFF \rc_reg[9]  ( .D(n778), .CLK(clk), .RST(1'b0), .Q(c[9]) );
  DFF \rc_reg[8]  ( .D(n777), .CLK(clk), .RST(1'b0), .Q(c[8]) );
  DFF \rc_reg[7]  ( .D(n776), .CLK(clk), .RST(1'b0), .Q(c[7]) );
  DFF \rc_reg[6]  ( .D(n775), .CLK(clk), .RST(1'b0), .Q(c[6]) );
  DFF \rc_reg[5]  ( .D(n774), .CLK(clk), .RST(1'b0), .Q(c[5]) );
  DFF \rc_reg[4]  ( .D(n773), .CLK(clk), .RST(1'b0), .Q(c[4]) );
  DFF \rc_reg[3]  ( .D(n772), .CLK(clk), .RST(1'b0), .Q(c[3]) );
  DFF \rc_reg[2]  ( .D(n771), .CLK(clk), .RST(1'b0), .Q(c[2]) );
  DFF \rc_reg[1]  ( .D(n770), .CLK(clk), .RST(1'b0), .Q(c[1]) );
  DFF \rc_reg[0]  ( .D(n769), .CLK(clk), .RST(1'b0), .Q(c[0]) );
  NANDN U1027 ( .A(n1994), .B(n1995), .Z(n1025) );
  NANDN U1028 ( .A(n3343), .B(n3342), .Z(n1026) );
  AND U1029 ( .A(n1025), .B(n1026), .Z(n1027) );
  NAND U1030 ( .A(n3348), .B(n3347), .Z(n1028) );
  NANDN U1031 ( .A(n1027), .B(n1996), .Z(n1029) );
  AND U1032 ( .A(n1028), .B(n1029), .Z(n1997) );
  XOR U1033 ( .A(n1089), .B(n1088), .Z(n2572) );
  XOR U1034 ( .A(n1113), .B(n1112), .Z(n2592) );
  XOR U1035 ( .A(n1137), .B(n1136), .Z(n2612) );
  XOR U1036 ( .A(n1177), .B(n1176), .Z(n2647) );
  XOR U1037 ( .A(n1217), .B(n1216), .Z(n2682) );
  XOR U1038 ( .A(n1241), .B(n1240), .Z(n2702) );
  XOR U1039 ( .A(n1265), .B(n1264), .Z(n2722) );
  XOR U1040 ( .A(n1289), .B(n1288), .Z(n2742) );
  XOR U1041 ( .A(n1313), .B(n1312), .Z(n2762) );
  XOR U1042 ( .A(n1337), .B(n1336), .Z(n2782) );
  XOR U1043 ( .A(n1361), .B(n1360), .Z(n2802) );
  XOR U1044 ( .A(n1385), .B(n1384), .Z(n2822) );
  XOR U1045 ( .A(n1409), .B(n1408), .Z(n2842) );
  XOR U1046 ( .A(n1433), .B(n1432), .Z(n2862) );
  XOR U1047 ( .A(n1457), .B(n1456), .Z(n2882) );
  XOR U1048 ( .A(n1481), .B(n1480), .Z(n2902) );
  XOR U1049 ( .A(n1505), .B(n1504), .Z(n2922) );
  XOR U1050 ( .A(n1601), .B(n1600), .Z(n3007) );
  XOR U1051 ( .A(n1625), .B(n1624), .Z(n3027) );
  XOR U1052 ( .A(n1649), .B(n1648), .Z(n3047) );
  XOR U1053 ( .A(n1673), .B(n1672), .Z(n3067) );
  XOR U1054 ( .A(n1697), .B(n1696), .Z(n3087) );
  XOR U1055 ( .A(n1721), .B(n1720), .Z(n3107) );
  XOR U1056 ( .A(n1745), .B(n1744), .Z(n3127) );
  XOR U1057 ( .A(n1785), .B(n1784), .Z(n3162) );
  XOR U1058 ( .A(n1809), .B(n1808), .Z(n3182) );
  XOR U1059 ( .A(n1833), .B(n1832), .Z(n3202) );
  XOR U1060 ( .A(n1857), .B(n1856), .Z(n3222) );
  XOR U1061 ( .A(n1881), .B(n1880), .Z(n3242) );
  XOR U1062 ( .A(n1905), .B(n1904), .Z(n3262) );
  XOR U1063 ( .A(n1973), .B(n1972), .Z(n3322) );
  XOR U1064 ( .A(n2016), .B(n2015), .Z(n3367) );
  XOR U1065 ( .A(n2040), .B(n2039), .Z(n3387) );
  XOR U1066 ( .A(n2064), .B(n2063), .Z(n3407) );
  XOR U1067 ( .A(n2088), .B(n2087), .Z(n3427) );
  OR U1068 ( .A(n2117), .B(n2118), .Z(n1030) );
  ANDN U1069 ( .B(n1030), .A(n2120), .Z(n3458) );
  XOR U1070 ( .A(n2155), .B(n2154), .Z(n3487) );
  XOR U1071 ( .A(n2179), .B(n2178), .Z(n3507) );
  XOR U1072 ( .A(n2231), .B(n2230), .Z(n3552) );
  XOR U1073 ( .A(n2255), .B(n2254), .Z(n3572) );
  XOR U1074 ( .A(n2279), .B(n2278), .Z(n3592) );
  XOR U1075 ( .A(n2319), .B(n2318), .Z(n3627) );
  XOR U1076 ( .A(n2343), .B(n2342), .Z(n3647) );
  XOR U1077 ( .A(n2367), .B(n2366), .Z(n3667) );
  XOR U1078 ( .A(n2391), .B(n2390), .Z(n3687) );
  XOR U1079 ( .A(n2431), .B(n2430), .Z(n3722) );
  XOR U1080 ( .A(n2455), .B(n2454), .Z(n3742) );
  XOR U1081 ( .A(n2479), .B(n2478), .Z(n3762) );
  XOR U1082 ( .A(n2503), .B(n2502), .Z(n3782) );
  NAND U1083 ( .A(n3353), .B(n3352), .Z(n1031) );
  NAND U1084 ( .A(n1999), .B(n1998), .Z(n1032) );
  NAND U1085 ( .A(n1031), .B(n1032), .Z(n1033) );
  ANDN U1086 ( .B(n1033), .A(n2001), .Z(n2003) );
  XOR U1087 ( .A(n1059), .B(n1060), .Z(n2548) );
  XOR U1088 ( .A(n1077), .B(n1076), .Z(n2562) );
  XOR U1089 ( .A(n1101), .B(n1100), .Z(n2582) );
  XOR U1090 ( .A(n1125), .B(n1124), .Z(n2602) );
  XOR U1091 ( .A(n1149), .B(n1148), .Z(n2622) );
  XOR U1092 ( .A(n1189), .B(n1188), .Z(n2657) );
  XOR U1093 ( .A(n1229), .B(n1228), .Z(n2692) );
  XOR U1094 ( .A(n1253), .B(n1252), .Z(n2712) );
  XOR U1095 ( .A(n1277), .B(n1276), .Z(n2732) );
  XOR U1096 ( .A(n1301), .B(n1300), .Z(n2752) );
  XOR U1097 ( .A(n1325), .B(n1324), .Z(n2772) );
  XOR U1098 ( .A(n1349), .B(n1348), .Z(n2792) );
  XOR U1099 ( .A(n1373), .B(n1372), .Z(n2812) );
  XOR U1100 ( .A(n1397), .B(n1396), .Z(n2832) );
  XOR U1101 ( .A(n1421), .B(n1420), .Z(n2852) );
  XOR U1102 ( .A(n1445), .B(n1444), .Z(n2872) );
  XOR U1103 ( .A(n1469), .B(n1468), .Z(n2892) );
  XOR U1104 ( .A(n1493), .B(n1492), .Z(n2912) );
  XOR U1105 ( .A(n1517), .B(n1516), .Z(n2932) );
  XOR U1106 ( .A(n1545), .B(n1544), .Z(n2957) );
  XOR U1107 ( .A(n1573), .B(n1572), .Z(n2982) );
  XOR U1108 ( .A(n1613), .B(n1612), .Z(n3017) );
  XOR U1109 ( .A(n1637), .B(n1636), .Z(n3037) );
  XOR U1110 ( .A(n1661), .B(n1660), .Z(n3057) );
  XOR U1111 ( .A(n1685), .B(n1684), .Z(n3077) );
  XOR U1112 ( .A(n1709), .B(n1708), .Z(n3097) );
  XOR U1113 ( .A(n1733), .B(n1732), .Z(n3117) );
  XOR U1114 ( .A(n1757), .B(n1756), .Z(n3137) );
  XOR U1115 ( .A(n1797), .B(n1796), .Z(n3172) );
  XOR U1116 ( .A(n1821), .B(n1820), .Z(n3192) );
  XOR U1117 ( .A(n1845), .B(n1844), .Z(n3212) );
  XOR U1118 ( .A(n1869), .B(n1868), .Z(n3232) );
  XOR U1119 ( .A(n1893), .B(n1892), .Z(n3252) );
  XOR U1120 ( .A(n1917), .B(n1916), .Z(n3272) );
  XOR U1121 ( .A(n1945), .B(n1944), .Z(n3297) );
  XOR U1122 ( .A(n1985), .B(n1984), .Z(n3332) );
  XOR U1123 ( .A(n2028), .B(n2027), .Z(n3377) );
  XOR U1124 ( .A(n2052), .B(n2051), .Z(n3397) );
  XOR U1125 ( .A(n2076), .B(n2075), .Z(n3417) );
  XOR U1126 ( .A(n2100), .B(n2099), .Z(n3437) );
  XOR U1127 ( .A(n2127), .B(n2126), .Z(n3462) );
  XOR U1128 ( .A(n2167), .B(n2166), .Z(n3497) );
  XOR U1129 ( .A(n2191), .B(n2190), .Z(n3517) );
  XOR U1130 ( .A(n2219), .B(n2218), .Z(n3542) );
  XOR U1131 ( .A(n2243), .B(n2242), .Z(n3562) );
  XOR U1132 ( .A(n2267), .B(n2266), .Z(n3582) );
  XOR U1133 ( .A(n2291), .B(n2290), .Z(n3602) );
  XOR U1134 ( .A(n2331), .B(n2330), .Z(n3637) );
  XOR U1135 ( .A(n2355), .B(n2354), .Z(n3657) );
  XOR U1136 ( .A(n2379), .B(n2378), .Z(n3677) );
  XOR U1137 ( .A(n2403), .B(n2402), .Z(n3697) );
  XOR U1138 ( .A(n2443), .B(n2442), .Z(n3732) );
  XOR U1139 ( .A(n2467), .B(n2466), .Z(n3752) );
  XOR U1140 ( .A(n2491), .B(n2490), .Z(n3772) );
  XOR U1141 ( .A(n2513), .B(n2514), .Z(n3792) );
  AND U1142 ( .A(a[255]), .B(b[255]), .Z(n2522) );
  NAND U1143 ( .A(a[254]), .B(b[254]), .Z(n2518) );
  NAND U1144 ( .A(a[253]), .B(b[253]), .Z(n2513) );
  NAND U1145 ( .A(a[186]), .B(b[186]), .Z(n2117) );
  NAND U1146 ( .A(a[167]), .B(b[167]), .Z(n2005) );
  NAND U1147 ( .A(a[165]), .B(b[165]), .Z(n1998) );
  NAND U1148 ( .A(a[164]), .B(b[164]), .Z(n1996) );
  AND U1149 ( .A(a[163]), .B(b[163]), .Z(n1994) );
  NAND U1150 ( .A(a[153]), .B(b[153]), .Z(n1934) );
  NAND U1151 ( .A(a[126]), .B(b[126]), .Z(n1774) );
  NAND U1152 ( .A(a[85]), .B(b[85]), .Z(n1534) );
  NAND U1153 ( .A(a[23]), .B(b[23]), .Z(n1166) );
  AND U1154 ( .A(a[4]), .B(b[4]), .Z(n1059) );
  AND U1155 ( .A(a[3]), .B(b[3]), .Z(n1052) );
  AND U1156 ( .A(a[2]), .B(b[2]), .Z(n1048) );
  XNOR U1157 ( .A(a[1]), .B(b[1]), .Z(n1036) );
  XNOR U1158 ( .A(carry_on[1]), .B(n1036), .Z(n2528) );
  NAND U1159 ( .A(a[0]), .B(b[0]), .Z(n1035) );
  XOR U1160 ( .A(a[0]), .B(b[0]), .Z(n2523) );
  NAND U1161 ( .A(n2523), .B(carry_on[0]), .Z(n1034) );
  NAND U1162 ( .A(n1035), .B(n1034), .Z(n2527) );
  NAND U1163 ( .A(n2528), .B(n2527), .Z(n1038) );
  ANDN U1164 ( .B(carry_on[1]), .A(n1036), .Z(n1039) );
  ANDN U1165 ( .B(n1038), .A(n1039), .Z(n1037) );
  NAND U1166 ( .A(a[1]), .B(b[1]), .Z(n1040) );
  NAND U1167 ( .A(n1037), .B(n1040), .Z(n1044) );
  XNOR U1168 ( .A(n1040), .B(n1038), .Z(n1042) );
  NAND U1169 ( .A(n1040), .B(n1039), .Z(n1041) );
  NAND U1170 ( .A(n1042), .B(n1041), .Z(n2533) );
  XNOR U1171 ( .A(a[2]), .B(b[2]), .Z(n2532) );
  NAND U1172 ( .A(n2533), .B(n2532), .Z(n1043) );
  NAND U1173 ( .A(n1044), .B(n1043), .Z(n1049) );
  ANDN U1174 ( .B(n1048), .A(n1049), .Z(n1045) );
  XNOR U1175 ( .A(n1052), .B(n1045), .Z(n1047) );
  XNOR U1176 ( .A(n1048), .B(n1049), .Z(n2537) );
  XOR U1177 ( .A(a[3]), .B(b[3]), .Z(n2538) );
  NAND U1178 ( .A(n2537), .B(n2538), .Z(n1046) );
  NAND U1179 ( .A(n1047), .B(n1046), .Z(n2543) );
  XNOR U1180 ( .A(a[4]), .B(b[4]), .Z(n2542) );
  NAND U1181 ( .A(n2543), .B(n2542), .Z(n1055) );
  ANDN U1182 ( .B(n1049), .A(n1048), .Z(n1051) );
  ANDN U1183 ( .B(n2537), .A(n2538), .Z(n1050) );
  OR U1184 ( .A(n1051), .B(n1050), .Z(n1053) );
  ANDN U1185 ( .B(n1053), .A(n1052), .Z(n1054) );
  ANDN U1186 ( .B(n1055), .A(n1054), .Z(n1060) );
  NOR U1187 ( .A(n1059), .B(n1060), .Z(n1057) );
  XNOR U1188 ( .A(a[5]), .B(b[5]), .Z(n2547) );
  NAND U1189 ( .A(n2548), .B(n2547), .Z(n1056) );
  NANDN U1190 ( .A(n1057), .B(n1056), .Z(n1058) );
  AND U1191 ( .A(a[5]), .B(b[5]), .Z(n1062) );
  ANDN U1192 ( .B(n1058), .A(n1062), .Z(n1064) );
  AND U1193 ( .A(n1060), .B(n1059), .Z(n1061) );
  NAND U1194 ( .A(n1062), .B(n1061), .Z(n1067) );
  ANDN U1195 ( .B(n1067), .A(n1064), .Z(n2553) );
  XNOR U1196 ( .A(a[6]), .B(b[6]), .Z(n2552) );
  AND U1197 ( .A(n2553), .B(n2552), .Z(n1063) );
  OR U1198 ( .A(n1064), .B(n1063), .Z(n1065) );
  NAND U1199 ( .A(a[6]), .B(b[6]), .Z(n1066) );
  AND U1200 ( .A(n1065), .B(n1066), .Z(n1070) );
  OR U1201 ( .A(n1067), .B(n1066), .Z(n1068) );
  ANDN U1202 ( .B(n1068), .A(n1070), .Z(n2558) );
  XNOR U1203 ( .A(a[7]), .B(b[7]), .Z(n2557) );
  NAND U1204 ( .A(n2558), .B(n2557), .Z(n1069) );
  NANDN U1205 ( .A(n1070), .B(n1069), .Z(n1076) );
  NAND U1206 ( .A(a[7]), .B(b[7]), .Z(n1077) );
  AND U1207 ( .A(n1076), .B(n1077), .Z(n1072) );
  XOR U1208 ( .A(a[8]), .B(b[8]), .Z(n2563) );
  ANDN U1209 ( .B(n2562), .A(n2563), .Z(n1071) );
  OR U1210 ( .A(n1072), .B(n1071), .Z(n1073) );
  AND U1211 ( .A(a[8]), .B(b[8]), .Z(n1075) );
  ANDN U1212 ( .B(n1073), .A(n1075), .Z(n1082) );
  NOR U1213 ( .A(n1077), .B(n1076), .Z(n1074) );
  XNOR U1214 ( .A(n1075), .B(n1074), .Z(n1080) );
  XOR U1215 ( .A(n1077), .B(n1076), .Z(n1078) );
  NAND U1216 ( .A(n1078), .B(n2563), .Z(n1079) );
  NAND U1217 ( .A(n1080), .B(n1079), .Z(n2568) );
  XNOR U1218 ( .A(a[9]), .B(b[9]), .Z(n2567) );
  NAND U1219 ( .A(n2568), .B(n2567), .Z(n1081) );
  NANDN U1220 ( .A(n1082), .B(n1081), .Z(n1088) );
  NAND U1221 ( .A(a[9]), .B(b[9]), .Z(n1089) );
  AND U1222 ( .A(n1088), .B(n1089), .Z(n1084) );
  XOR U1223 ( .A(a[10]), .B(b[10]), .Z(n2573) );
  ANDN U1224 ( .B(n2572), .A(n2573), .Z(n1083) );
  OR U1225 ( .A(n1084), .B(n1083), .Z(n1085) );
  AND U1226 ( .A(a[10]), .B(b[10]), .Z(n1087) );
  ANDN U1227 ( .B(n1085), .A(n1087), .Z(n1094) );
  NOR U1228 ( .A(n1089), .B(n1088), .Z(n1086) );
  XNOR U1229 ( .A(n1087), .B(n1086), .Z(n1092) );
  XOR U1230 ( .A(n1089), .B(n1088), .Z(n1090) );
  NAND U1231 ( .A(n1090), .B(n2573), .Z(n1091) );
  NAND U1232 ( .A(n1092), .B(n1091), .Z(n2578) );
  XNOR U1233 ( .A(a[11]), .B(b[11]), .Z(n2577) );
  NAND U1234 ( .A(n2578), .B(n2577), .Z(n1093) );
  NANDN U1235 ( .A(n1094), .B(n1093), .Z(n1100) );
  NAND U1236 ( .A(a[11]), .B(b[11]), .Z(n1101) );
  AND U1237 ( .A(n1100), .B(n1101), .Z(n1096) );
  XOR U1238 ( .A(a[12]), .B(b[12]), .Z(n2583) );
  ANDN U1239 ( .B(n2582), .A(n2583), .Z(n1095) );
  OR U1240 ( .A(n1096), .B(n1095), .Z(n1097) );
  AND U1241 ( .A(a[12]), .B(b[12]), .Z(n1099) );
  ANDN U1242 ( .B(n1097), .A(n1099), .Z(n1106) );
  NOR U1243 ( .A(n1101), .B(n1100), .Z(n1098) );
  XNOR U1244 ( .A(n1099), .B(n1098), .Z(n1104) );
  XOR U1245 ( .A(n1101), .B(n1100), .Z(n1102) );
  NAND U1246 ( .A(n1102), .B(n2583), .Z(n1103) );
  NAND U1247 ( .A(n1104), .B(n1103), .Z(n2588) );
  XNOR U1248 ( .A(a[13]), .B(b[13]), .Z(n2587) );
  NAND U1249 ( .A(n2588), .B(n2587), .Z(n1105) );
  NANDN U1250 ( .A(n1106), .B(n1105), .Z(n1112) );
  NAND U1251 ( .A(a[13]), .B(b[13]), .Z(n1113) );
  AND U1252 ( .A(n1112), .B(n1113), .Z(n1108) );
  XOR U1253 ( .A(a[14]), .B(b[14]), .Z(n2593) );
  ANDN U1254 ( .B(n2592), .A(n2593), .Z(n1107) );
  OR U1255 ( .A(n1108), .B(n1107), .Z(n1109) );
  AND U1256 ( .A(a[14]), .B(b[14]), .Z(n1111) );
  ANDN U1257 ( .B(n1109), .A(n1111), .Z(n1118) );
  NOR U1258 ( .A(n1113), .B(n1112), .Z(n1110) );
  XNOR U1259 ( .A(n1111), .B(n1110), .Z(n1116) );
  XOR U1260 ( .A(n1113), .B(n1112), .Z(n1114) );
  NAND U1261 ( .A(n1114), .B(n2593), .Z(n1115) );
  NAND U1262 ( .A(n1116), .B(n1115), .Z(n2598) );
  XNOR U1263 ( .A(a[15]), .B(b[15]), .Z(n2597) );
  NAND U1264 ( .A(n2598), .B(n2597), .Z(n1117) );
  NANDN U1265 ( .A(n1118), .B(n1117), .Z(n1124) );
  NAND U1266 ( .A(a[15]), .B(b[15]), .Z(n1125) );
  AND U1267 ( .A(n1124), .B(n1125), .Z(n1120) );
  XOR U1268 ( .A(a[16]), .B(b[16]), .Z(n2603) );
  ANDN U1269 ( .B(n2602), .A(n2603), .Z(n1119) );
  OR U1270 ( .A(n1120), .B(n1119), .Z(n1121) );
  AND U1271 ( .A(a[16]), .B(b[16]), .Z(n1123) );
  ANDN U1272 ( .B(n1121), .A(n1123), .Z(n1130) );
  NOR U1273 ( .A(n1125), .B(n1124), .Z(n1122) );
  XNOR U1274 ( .A(n1123), .B(n1122), .Z(n1128) );
  XOR U1275 ( .A(n1125), .B(n1124), .Z(n1126) );
  NAND U1276 ( .A(n1126), .B(n2603), .Z(n1127) );
  NAND U1277 ( .A(n1128), .B(n1127), .Z(n2608) );
  XNOR U1278 ( .A(a[17]), .B(b[17]), .Z(n2607) );
  NAND U1279 ( .A(n2608), .B(n2607), .Z(n1129) );
  NANDN U1280 ( .A(n1130), .B(n1129), .Z(n1136) );
  NAND U1281 ( .A(a[17]), .B(b[17]), .Z(n1137) );
  AND U1282 ( .A(n1136), .B(n1137), .Z(n1132) );
  XOR U1283 ( .A(a[18]), .B(b[18]), .Z(n2613) );
  ANDN U1284 ( .B(n2612), .A(n2613), .Z(n1131) );
  OR U1285 ( .A(n1132), .B(n1131), .Z(n1133) );
  AND U1286 ( .A(a[18]), .B(b[18]), .Z(n1135) );
  ANDN U1287 ( .B(n1133), .A(n1135), .Z(n1142) );
  NOR U1288 ( .A(n1137), .B(n1136), .Z(n1134) );
  XNOR U1289 ( .A(n1135), .B(n1134), .Z(n1140) );
  XOR U1290 ( .A(n1137), .B(n1136), .Z(n1138) );
  NAND U1291 ( .A(n1138), .B(n2613), .Z(n1139) );
  NAND U1292 ( .A(n1140), .B(n1139), .Z(n2618) );
  XNOR U1293 ( .A(a[19]), .B(b[19]), .Z(n2617) );
  NAND U1294 ( .A(n2618), .B(n2617), .Z(n1141) );
  NANDN U1295 ( .A(n1142), .B(n1141), .Z(n1148) );
  NAND U1296 ( .A(a[19]), .B(b[19]), .Z(n1149) );
  AND U1297 ( .A(n1148), .B(n1149), .Z(n1144) );
  XOR U1298 ( .A(a[20]), .B(b[20]), .Z(n2623) );
  ANDN U1299 ( .B(n2622), .A(n2623), .Z(n1143) );
  OR U1300 ( .A(n1144), .B(n1143), .Z(n1145) );
  AND U1301 ( .A(a[20]), .B(b[20]), .Z(n1147) );
  ANDN U1302 ( .B(n1145), .A(n1147), .Z(n1154) );
  NOR U1303 ( .A(n1149), .B(n1148), .Z(n1146) );
  XNOR U1304 ( .A(n1147), .B(n1146), .Z(n1152) );
  XOR U1305 ( .A(n1149), .B(n1148), .Z(n1150) );
  NAND U1306 ( .A(n1150), .B(n2623), .Z(n1151) );
  NAND U1307 ( .A(n1152), .B(n1151), .Z(n2628) );
  XNOR U1308 ( .A(a[21]), .B(b[21]), .Z(n2627) );
  NAND U1309 ( .A(n2628), .B(n2627), .Z(n1153) );
  NANDN U1310 ( .A(n1154), .B(n1153), .Z(n1155) );
  IV U1311 ( .A(n1155), .Z(n1159) );
  AND U1312 ( .A(a[21]), .B(b[21]), .Z(n1160) );
  NOR U1313 ( .A(n1159), .B(n1160), .Z(n1157) );
  XNOR U1314 ( .A(n1160), .B(n1155), .Z(n2633) );
  XNOR U1315 ( .A(a[22]), .B(b[22]), .Z(n2632) );
  AND U1316 ( .A(n2633), .B(n2632), .Z(n1156) );
  OR U1317 ( .A(n1157), .B(n1156), .Z(n1158) );
  AND U1318 ( .A(a[22]), .B(b[22]), .Z(n1162) );
  ANDN U1319 ( .B(n1158), .A(n1162), .Z(n1164) );
  AND U1320 ( .A(n1160), .B(n1159), .Z(n1161) );
  NAND U1321 ( .A(n1162), .B(n1161), .Z(n1167) );
  ANDN U1322 ( .B(n1167), .A(n1164), .Z(n2638) );
  XNOR U1323 ( .A(a[23]), .B(b[23]), .Z(n2637) );
  AND U1324 ( .A(n2638), .B(n2637), .Z(n1163) );
  OR U1325 ( .A(n1164), .B(n1163), .Z(n1165) );
  AND U1326 ( .A(n1166), .B(n1165), .Z(n1170) );
  OR U1327 ( .A(n1167), .B(n1166), .Z(n1168) );
  ANDN U1328 ( .B(n1168), .A(n1170), .Z(n2643) );
  XNOR U1329 ( .A(a[24]), .B(b[24]), .Z(n2642) );
  NAND U1330 ( .A(n2643), .B(n2642), .Z(n1169) );
  NANDN U1331 ( .A(n1170), .B(n1169), .Z(n1176) );
  NAND U1332 ( .A(a[24]), .B(b[24]), .Z(n1177) );
  AND U1333 ( .A(n1176), .B(n1177), .Z(n1172) );
  XOR U1334 ( .A(a[25]), .B(b[25]), .Z(n2648) );
  ANDN U1335 ( .B(n2647), .A(n2648), .Z(n1171) );
  OR U1336 ( .A(n1172), .B(n1171), .Z(n1173) );
  AND U1337 ( .A(a[25]), .B(b[25]), .Z(n1175) );
  ANDN U1338 ( .B(n1173), .A(n1175), .Z(n1182) );
  NOR U1339 ( .A(n1177), .B(n1176), .Z(n1174) );
  XNOR U1340 ( .A(n1175), .B(n1174), .Z(n1180) );
  XOR U1341 ( .A(n1177), .B(n1176), .Z(n1178) );
  NAND U1342 ( .A(n1178), .B(n2648), .Z(n1179) );
  NAND U1343 ( .A(n1180), .B(n1179), .Z(n2653) );
  XNOR U1344 ( .A(a[26]), .B(b[26]), .Z(n2652) );
  NAND U1345 ( .A(n2653), .B(n2652), .Z(n1181) );
  NANDN U1346 ( .A(n1182), .B(n1181), .Z(n1188) );
  NAND U1347 ( .A(a[26]), .B(b[26]), .Z(n1189) );
  AND U1348 ( .A(n1188), .B(n1189), .Z(n1184) );
  XOR U1349 ( .A(a[27]), .B(b[27]), .Z(n2658) );
  ANDN U1350 ( .B(n2657), .A(n2658), .Z(n1183) );
  OR U1351 ( .A(n1184), .B(n1183), .Z(n1185) );
  AND U1352 ( .A(a[27]), .B(b[27]), .Z(n1187) );
  ANDN U1353 ( .B(n1185), .A(n1187), .Z(n1194) );
  NOR U1354 ( .A(n1189), .B(n1188), .Z(n1186) );
  XNOR U1355 ( .A(n1187), .B(n1186), .Z(n1192) );
  XOR U1356 ( .A(n1189), .B(n1188), .Z(n1190) );
  NAND U1357 ( .A(n1190), .B(n2658), .Z(n1191) );
  NAND U1358 ( .A(n1192), .B(n1191), .Z(n2663) );
  XNOR U1359 ( .A(a[28]), .B(b[28]), .Z(n2662) );
  NAND U1360 ( .A(n2663), .B(n2662), .Z(n1193) );
  NANDN U1361 ( .A(n1194), .B(n1193), .Z(n1195) );
  IV U1362 ( .A(n1195), .Z(n1199) );
  AND U1363 ( .A(a[28]), .B(b[28]), .Z(n1200) );
  NOR U1364 ( .A(n1199), .B(n1200), .Z(n1197) );
  XNOR U1365 ( .A(n1200), .B(n1195), .Z(n2668) );
  XNOR U1366 ( .A(a[29]), .B(b[29]), .Z(n2667) );
  AND U1367 ( .A(n2668), .B(n2667), .Z(n1196) );
  OR U1368 ( .A(n1197), .B(n1196), .Z(n1198) );
  AND U1369 ( .A(a[29]), .B(b[29]), .Z(n1202) );
  ANDN U1370 ( .B(n1198), .A(n1202), .Z(n1204) );
  AND U1371 ( .A(n1200), .B(n1199), .Z(n1201) );
  NAND U1372 ( .A(n1202), .B(n1201), .Z(n1207) );
  ANDN U1373 ( .B(n1207), .A(n1204), .Z(n2673) );
  XNOR U1374 ( .A(a[30]), .B(b[30]), .Z(n2672) );
  AND U1375 ( .A(n2673), .B(n2672), .Z(n1203) );
  OR U1376 ( .A(n1204), .B(n1203), .Z(n1205) );
  AND U1377 ( .A(a[30]), .B(b[30]), .Z(n1206) );
  ANDN U1378 ( .B(n1205), .A(n1206), .Z(n1210) );
  NANDN U1379 ( .A(n1207), .B(n1206), .Z(n1208) );
  ANDN U1380 ( .B(n1208), .A(n1210), .Z(n2678) );
  XNOR U1381 ( .A(a[31]), .B(b[31]), .Z(n2677) );
  NAND U1382 ( .A(n2678), .B(n2677), .Z(n1209) );
  NANDN U1383 ( .A(n1210), .B(n1209), .Z(n1216) );
  NAND U1384 ( .A(a[31]), .B(b[31]), .Z(n1217) );
  AND U1385 ( .A(n1216), .B(n1217), .Z(n1212) );
  XOR U1386 ( .A(a[32]), .B(b[32]), .Z(n2683) );
  ANDN U1387 ( .B(n2682), .A(n2683), .Z(n1211) );
  OR U1388 ( .A(n1212), .B(n1211), .Z(n1213) );
  AND U1389 ( .A(a[32]), .B(b[32]), .Z(n1215) );
  ANDN U1390 ( .B(n1213), .A(n1215), .Z(n1222) );
  NOR U1391 ( .A(n1217), .B(n1216), .Z(n1214) );
  XNOR U1392 ( .A(n1215), .B(n1214), .Z(n1220) );
  XOR U1393 ( .A(n1217), .B(n1216), .Z(n1218) );
  NAND U1394 ( .A(n1218), .B(n2683), .Z(n1219) );
  NAND U1395 ( .A(n1220), .B(n1219), .Z(n2688) );
  XNOR U1396 ( .A(a[33]), .B(b[33]), .Z(n2687) );
  NAND U1397 ( .A(n2688), .B(n2687), .Z(n1221) );
  NANDN U1398 ( .A(n1222), .B(n1221), .Z(n1228) );
  NAND U1399 ( .A(a[33]), .B(b[33]), .Z(n1229) );
  AND U1400 ( .A(n1228), .B(n1229), .Z(n1224) );
  XOR U1401 ( .A(a[34]), .B(b[34]), .Z(n2693) );
  ANDN U1402 ( .B(n2692), .A(n2693), .Z(n1223) );
  OR U1403 ( .A(n1224), .B(n1223), .Z(n1225) );
  AND U1404 ( .A(a[34]), .B(b[34]), .Z(n1227) );
  ANDN U1405 ( .B(n1225), .A(n1227), .Z(n1234) );
  NOR U1406 ( .A(n1229), .B(n1228), .Z(n1226) );
  XNOR U1407 ( .A(n1227), .B(n1226), .Z(n1232) );
  XOR U1408 ( .A(n1229), .B(n1228), .Z(n1230) );
  NAND U1409 ( .A(n1230), .B(n2693), .Z(n1231) );
  NAND U1410 ( .A(n1232), .B(n1231), .Z(n2698) );
  XNOR U1411 ( .A(a[35]), .B(b[35]), .Z(n2697) );
  NAND U1412 ( .A(n2698), .B(n2697), .Z(n1233) );
  NANDN U1413 ( .A(n1234), .B(n1233), .Z(n1240) );
  NAND U1414 ( .A(a[35]), .B(b[35]), .Z(n1241) );
  AND U1415 ( .A(n1240), .B(n1241), .Z(n1236) );
  XOR U1416 ( .A(a[36]), .B(b[36]), .Z(n2703) );
  ANDN U1417 ( .B(n2702), .A(n2703), .Z(n1235) );
  OR U1418 ( .A(n1236), .B(n1235), .Z(n1237) );
  AND U1419 ( .A(a[36]), .B(b[36]), .Z(n1239) );
  ANDN U1420 ( .B(n1237), .A(n1239), .Z(n1246) );
  NOR U1421 ( .A(n1241), .B(n1240), .Z(n1238) );
  XNOR U1422 ( .A(n1239), .B(n1238), .Z(n1244) );
  XOR U1423 ( .A(n1241), .B(n1240), .Z(n1242) );
  NAND U1424 ( .A(n1242), .B(n2703), .Z(n1243) );
  NAND U1425 ( .A(n1244), .B(n1243), .Z(n2708) );
  XNOR U1426 ( .A(a[37]), .B(b[37]), .Z(n2707) );
  NAND U1427 ( .A(n2708), .B(n2707), .Z(n1245) );
  NANDN U1428 ( .A(n1246), .B(n1245), .Z(n1252) );
  NAND U1429 ( .A(a[37]), .B(b[37]), .Z(n1253) );
  AND U1430 ( .A(n1252), .B(n1253), .Z(n1248) );
  XOR U1431 ( .A(a[38]), .B(b[38]), .Z(n2713) );
  ANDN U1432 ( .B(n2712), .A(n2713), .Z(n1247) );
  OR U1433 ( .A(n1248), .B(n1247), .Z(n1249) );
  AND U1434 ( .A(a[38]), .B(b[38]), .Z(n1251) );
  ANDN U1435 ( .B(n1249), .A(n1251), .Z(n1258) );
  NOR U1436 ( .A(n1253), .B(n1252), .Z(n1250) );
  XNOR U1437 ( .A(n1251), .B(n1250), .Z(n1256) );
  XOR U1438 ( .A(n1253), .B(n1252), .Z(n1254) );
  NAND U1439 ( .A(n1254), .B(n2713), .Z(n1255) );
  NAND U1440 ( .A(n1256), .B(n1255), .Z(n2718) );
  XNOR U1441 ( .A(a[39]), .B(b[39]), .Z(n2717) );
  NAND U1442 ( .A(n2718), .B(n2717), .Z(n1257) );
  NANDN U1443 ( .A(n1258), .B(n1257), .Z(n1264) );
  NAND U1444 ( .A(a[39]), .B(b[39]), .Z(n1265) );
  AND U1445 ( .A(n1264), .B(n1265), .Z(n1260) );
  XOR U1446 ( .A(a[40]), .B(b[40]), .Z(n2723) );
  ANDN U1447 ( .B(n2722), .A(n2723), .Z(n1259) );
  OR U1448 ( .A(n1260), .B(n1259), .Z(n1261) );
  AND U1449 ( .A(a[40]), .B(b[40]), .Z(n1263) );
  ANDN U1450 ( .B(n1261), .A(n1263), .Z(n1270) );
  NOR U1451 ( .A(n1265), .B(n1264), .Z(n1262) );
  XNOR U1452 ( .A(n1263), .B(n1262), .Z(n1268) );
  XOR U1453 ( .A(n1265), .B(n1264), .Z(n1266) );
  NAND U1454 ( .A(n1266), .B(n2723), .Z(n1267) );
  NAND U1455 ( .A(n1268), .B(n1267), .Z(n2728) );
  XNOR U1456 ( .A(a[41]), .B(b[41]), .Z(n2727) );
  NAND U1457 ( .A(n2728), .B(n2727), .Z(n1269) );
  NANDN U1458 ( .A(n1270), .B(n1269), .Z(n1276) );
  NAND U1459 ( .A(a[41]), .B(b[41]), .Z(n1277) );
  AND U1460 ( .A(n1276), .B(n1277), .Z(n1272) );
  XOR U1461 ( .A(a[42]), .B(b[42]), .Z(n2733) );
  ANDN U1462 ( .B(n2732), .A(n2733), .Z(n1271) );
  OR U1463 ( .A(n1272), .B(n1271), .Z(n1273) );
  AND U1464 ( .A(a[42]), .B(b[42]), .Z(n1275) );
  ANDN U1465 ( .B(n1273), .A(n1275), .Z(n1282) );
  NOR U1466 ( .A(n1277), .B(n1276), .Z(n1274) );
  XNOR U1467 ( .A(n1275), .B(n1274), .Z(n1280) );
  XOR U1468 ( .A(n1277), .B(n1276), .Z(n1278) );
  NAND U1469 ( .A(n1278), .B(n2733), .Z(n1279) );
  NAND U1470 ( .A(n1280), .B(n1279), .Z(n2738) );
  XNOR U1471 ( .A(a[43]), .B(b[43]), .Z(n2737) );
  NAND U1472 ( .A(n2738), .B(n2737), .Z(n1281) );
  NANDN U1473 ( .A(n1282), .B(n1281), .Z(n1288) );
  NAND U1474 ( .A(a[43]), .B(b[43]), .Z(n1289) );
  AND U1475 ( .A(n1288), .B(n1289), .Z(n1284) );
  XOR U1476 ( .A(a[44]), .B(b[44]), .Z(n2743) );
  ANDN U1477 ( .B(n2742), .A(n2743), .Z(n1283) );
  OR U1478 ( .A(n1284), .B(n1283), .Z(n1285) );
  AND U1479 ( .A(a[44]), .B(b[44]), .Z(n1287) );
  ANDN U1480 ( .B(n1285), .A(n1287), .Z(n1294) );
  NOR U1481 ( .A(n1289), .B(n1288), .Z(n1286) );
  XNOR U1482 ( .A(n1287), .B(n1286), .Z(n1292) );
  XOR U1483 ( .A(n1289), .B(n1288), .Z(n1290) );
  NAND U1484 ( .A(n1290), .B(n2743), .Z(n1291) );
  NAND U1485 ( .A(n1292), .B(n1291), .Z(n2748) );
  XNOR U1486 ( .A(a[45]), .B(b[45]), .Z(n2747) );
  NAND U1487 ( .A(n2748), .B(n2747), .Z(n1293) );
  NANDN U1488 ( .A(n1294), .B(n1293), .Z(n1300) );
  NAND U1489 ( .A(a[45]), .B(b[45]), .Z(n1301) );
  AND U1490 ( .A(n1300), .B(n1301), .Z(n1296) );
  XOR U1491 ( .A(a[46]), .B(b[46]), .Z(n2753) );
  ANDN U1492 ( .B(n2752), .A(n2753), .Z(n1295) );
  OR U1493 ( .A(n1296), .B(n1295), .Z(n1297) );
  AND U1494 ( .A(a[46]), .B(b[46]), .Z(n1299) );
  ANDN U1495 ( .B(n1297), .A(n1299), .Z(n1306) );
  NOR U1496 ( .A(n1301), .B(n1300), .Z(n1298) );
  XNOR U1497 ( .A(n1299), .B(n1298), .Z(n1304) );
  XOR U1498 ( .A(n1301), .B(n1300), .Z(n1302) );
  NAND U1499 ( .A(n1302), .B(n2753), .Z(n1303) );
  NAND U1500 ( .A(n1304), .B(n1303), .Z(n2758) );
  XNOR U1501 ( .A(a[47]), .B(b[47]), .Z(n2757) );
  NAND U1502 ( .A(n2758), .B(n2757), .Z(n1305) );
  NANDN U1503 ( .A(n1306), .B(n1305), .Z(n1312) );
  NAND U1504 ( .A(a[47]), .B(b[47]), .Z(n1313) );
  AND U1505 ( .A(n1312), .B(n1313), .Z(n1308) );
  XOR U1506 ( .A(a[48]), .B(b[48]), .Z(n2763) );
  ANDN U1507 ( .B(n2762), .A(n2763), .Z(n1307) );
  OR U1508 ( .A(n1308), .B(n1307), .Z(n1309) );
  AND U1509 ( .A(a[48]), .B(b[48]), .Z(n1311) );
  ANDN U1510 ( .B(n1309), .A(n1311), .Z(n1318) );
  NOR U1511 ( .A(n1313), .B(n1312), .Z(n1310) );
  XNOR U1512 ( .A(n1311), .B(n1310), .Z(n1316) );
  XOR U1513 ( .A(n1313), .B(n1312), .Z(n1314) );
  NAND U1514 ( .A(n1314), .B(n2763), .Z(n1315) );
  NAND U1515 ( .A(n1316), .B(n1315), .Z(n2768) );
  XNOR U1516 ( .A(a[49]), .B(b[49]), .Z(n2767) );
  NAND U1517 ( .A(n2768), .B(n2767), .Z(n1317) );
  NANDN U1518 ( .A(n1318), .B(n1317), .Z(n1324) );
  NAND U1519 ( .A(a[49]), .B(b[49]), .Z(n1325) );
  AND U1520 ( .A(n1324), .B(n1325), .Z(n1320) );
  XOR U1521 ( .A(a[50]), .B(b[50]), .Z(n2773) );
  ANDN U1522 ( .B(n2772), .A(n2773), .Z(n1319) );
  OR U1523 ( .A(n1320), .B(n1319), .Z(n1321) );
  AND U1524 ( .A(a[50]), .B(b[50]), .Z(n1323) );
  ANDN U1525 ( .B(n1321), .A(n1323), .Z(n1330) );
  NOR U1526 ( .A(n1325), .B(n1324), .Z(n1322) );
  XNOR U1527 ( .A(n1323), .B(n1322), .Z(n1328) );
  XOR U1528 ( .A(n1325), .B(n1324), .Z(n1326) );
  NAND U1529 ( .A(n1326), .B(n2773), .Z(n1327) );
  NAND U1530 ( .A(n1328), .B(n1327), .Z(n2778) );
  XNOR U1531 ( .A(a[51]), .B(b[51]), .Z(n2777) );
  NAND U1532 ( .A(n2778), .B(n2777), .Z(n1329) );
  NANDN U1533 ( .A(n1330), .B(n1329), .Z(n1336) );
  NAND U1534 ( .A(a[51]), .B(b[51]), .Z(n1337) );
  AND U1535 ( .A(n1336), .B(n1337), .Z(n1332) );
  XOR U1536 ( .A(a[52]), .B(b[52]), .Z(n2783) );
  ANDN U1537 ( .B(n2782), .A(n2783), .Z(n1331) );
  OR U1538 ( .A(n1332), .B(n1331), .Z(n1333) );
  AND U1539 ( .A(a[52]), .B(b[52]), .Z(n1335) );
  ANDN U1540 ( .B(n1333), .A(n1335), .Z(n1342) );
  NOR U1541 ( .A(n1337), .B(n1336), .Z(n1334) );
  XNOR U1542 ( .A(n1335), .B(n1334), .Z(n1340) );
  XOR U1543 ( .A(n1337), .B(n1336), .Z(n1338) );
  NAND U1544 ( .A(n1338), .B(n2783), .Z(n1339) );
  NAND U1545 ( .A(n1340), .B(n1339), .Z(n2788) );
  XNOR U1546 ( .A(a[53]), .B(b[53]), .Z(n2787) );
  NAND U1547 ( .A(n2788), .B(n2787), .Z(n1341) );
  NANDN U1548 ( .A(n1342), .B(n1341), .Z(n1348) );
  NAND U1549 ( .A(a[53]), .B(b[53]), .Z(n1349) );
  AND U1550 ( .A(n1348), .B(n1349), .Z(n1344) );
  XOR U1551 ( .A(a[54]), .B(b[54]), .Z(n2793) );
  ANDN U1552 ( .B(n2792), .A(n2793), .Z(n1343) );
  OR U1553 ( .A(n1344), .B(n1343), .Z(n1345) );
  AND U1554 ( .A(a[54]), .B(b[54]), .Z(n1347) );
  ANDN U1555 ( .B(n1345), .A(n1347), .Z(n1354) );
  NOR U1556 ( .A(n1349), .B(n1348), .Z(n1346) );
  XNOR U1557 ( .A(n1347), .B(n1346), .Z(n1352) );
  XOR U1558 ( .A(n1349), .B(n1348), .Z(n1350) );
  NAND U1559 ( .A(n1350), .B(n2793), .Z(n1351) );
  NAND U1560 ( .A(n1352), .B(n1351), .Z(n2798) );
  XNOR U1561 ( .A(a[55]), .B(b[55]), .Z(n2797) );
  NAND U1562 ( .A(n2798), .B(n2797), .Z(n1353) );
  NANDN U1563 ( .A(n1354), .B(n1353), .Z(n1360) );
  NAND U1564 ( .A(a[55]), .B(b[55]), .Z(n1361) );
  AND U1565 ( .A(n1360), .B(n1361), .Z(n1356) );
  XOR U1566 ( .A(a[56]), .B(b[56]), .Z(n2803) );
  ANDN U1567 ( .B(n2802), .A(n2803), .Z(n1355) );
  OR U1568 ( .A(n1356), .B(n1355), .Z(n1357) );
  AND U1569 ( .A(a[56]), .B(b[56]), .Z(n1359) );
  ANDN U1570 ( .B(n1357), .A(n1359), .Z(n1366) );
  NOR U1571 ( .A(n1361), .B(n1360), .Z(n1358) );
  XNOR U1572 ( .A(n1359), .B(n1358), .Z(n1364) );
  XOR U1573 ( .A(n1361), .B(n1360), .Z(n1362) );
  NAND U1574 ( .A(n1362), .B(n2803), .Z(n1363) );
  NAND U1575 ( .A(n1364), .B(n1363), .Z(n2808) );
  XNOR U1576 ( .A(a[57]), .B(b[57]), .Z(n2807) );
  NAND U1577 ( .A(n2808), .B(n2807), .Z(n1365) );
  NANDN U1578 ( .A(n1366), .B(n1365), .Z(n1372) );
  NAND U1579 ( .A(a[57]), .B(b[57]), .Z(n1373) );
  AND U1580 ( .A(n1372), .B(n1373), .Z(n1368) );
  XOR U1581 ( .A(a[58]), .B(b[58]), .Z(n2813) );
  ANDN U1582 ( .B(n2812), .A(n2813), .Z(n1367) );
  OR U1583 ( .A(n1368), .B(n1367), .Z(n1369) );
  AND U1584 ( .A(a[58]), .B(b[58]), .Z(n1371) );
  ANDN U1585 ( .B(n1369), .A(n1371), .Z(n1378) );
  NOR U1586 ( .A(n1373), .B(n1372), .Z(n1370) );
  XNOR U1587 ( .A(n1371), .B(n1370), .Z(n1376) );
  XOR U1588 ( .A(n1373), .B(n1372), .Z(n1374) );
  NAND U1589 ( .A(n1374), .B(n2813), .Z(n1375) );
  NAND U1590 ( .A(n1376), .B(n1375), .Z(n2818) );
  XNOR U1591 ( .A(a[59]), .B(b[59]), .Z(n2817) );
  NAND U1592 ( .A(n2818), .B(n2817), .Z(n1377) );
  NANDN U1593 ( .A(n1378), .B(n1377), .Z(n1384) );
  NAND U1594 ( .A(a[59]), .B(b[59]), .Z(n1385) );
  AND U1595 ( .A(n1384), .B(n1385), .Z(n1380) );
  XOR U1596 ( .A(a[60]), .B(b[60]), .Z(n2823) );
  ANDN U1597 ( .B(n2822), .A(n2823), .Z(n1379) );
  OR U1598 ( .A(n1380), .B(n1379), .Z(n1381) );
  AND U1599 ( .A(a[60]), .B(b[60]), .Z(n1383) );
  ANDN U1600 ( .B(n1381), .A(n1383), .Z(n1390) );
  NOR U1601 ( .A(n1385), .B(n1384), .Z(n1382) );
  XNOR U1602 ( .A(n1383), .B(n1382), .Z(n1388) );
  XOR U1603 ( .A(n1385), .B(n1384), .Z(n1386) );
  NAND U1604 ( .A(n1386), .B(n2823), .Z(n1387) );
  NAND U1605 ( .A(n1388), .B(n1387), .Z(n2828) );
  XNOR U1606 ( .A(a[61]), .B(b[61]), .Z(n2827) );
  NAND U1607 ( .A(n2828), .B(n2827), .Z(n1389) );
  NANDN U1608 ( .A(n1390), .B(n1389), .Z(n1396) );
  NAND U1609 ( .A(a[61]), .B(b[61]), .Z(n1397) );
  AND U1610 ( .A(n1396), .B(n1397), .Z(n1392) );
  XOR U1611 ( .A(a[62]), .B(b[62]), .Z(n2833) );
  ANDN U1612 ( .B(n2832), .A(n2833), .Z(n1391) );
  OR U1613 ( .A(n1392), .B(n1391), .Z(n1393) );
  AND U1614 ( .A(a[62]), .B(b[62]), .Z(n1395) );
  ANDN U1615 ( .B(n1393), .A(n1395), .Z(n1402) );
  NOR U1616 ( .A(n1397), .B(n1396), .Z(n1394) );
  XNOR U1617 ( .A(n1395), .B(n1394), .Z(n1400) );
  XOR U1618 ( .A(n1397), .B(n1396), .Z(n1398) );
  NAND U1619 ( .A(n1398), .B(n2833), .Z(n1399) );
  NAND U1620 ( .A(n1400), .B(n1399), .Z(n2838) );
  XNOR U1621 ( .A(a[63]), .B(b[63]), .Z(n2837) );
  NAND U1622 ( .A(n2838), .B(n2837), .Z(n1401) );
  NANDN U1623 ( .A(n1402), .B(n1401), .Z(n1408) );
  NAND U1624 ( .A(a[63]), .B(b[63]), .Z(n1409) );
  AND U1625 ( .A(n1408), .B(n1409), .Z(n1404) );
  XOR U1626 ( .A(a[64]), .B(b[64]), .Z(n2843) );
  ANDN U1627 ( .B(n2842), .A(n2843), .Z(n1403) );
  OR U1628 ( .A(n1404), .B(n1403), .Z(n1405) );
  AND U1629 ( .A(a[64]), .B(b[64]), .Z(n1407) );
  ANDN U1630 ( .B(n1405), .A(n1407), .Z(n1414) );
  NOR U1631 ( .A(n1409), .B(n1408), .Z(n1406) );
  XNOR U1632 ( .A(n1407), .B(n1406), .Z(n1412) );
  XOR U1633 ( .A(n1409), .B(n1408), .Z(n1410) );
  NAND U1634 ( .A(n1410), .B(n2843), .Z(n1411) );
  NAND U1635 ( .A(n1412), .B(n1411), .Z(n2848) );
  XNOR U1636 ( .A(a[65]), .B(b[65]), .Z(n2847) );
  NAND U1637 ( .A(n2848), .B(n2847), .Z(n1413) );
  NANDN U1638 ( .A(n1414), .B(n1413), .Z(n1420) );
  NAND U1639 ( .A(a[65]), .B(b[65]), .Z(n1421) );
  AND U1640 ( .A(n1420), .B(n1421), .Z(n1416) );
  XOR U1641 ( .A(a[66]), .B(b[66]), .Z(n2853) );
  ANDN U1642 ( .B(n2852), .A(n2853), .Z(n1415) );
  OR U1643 ( .A(n1416), .B(n1415), .Z(n1417) );
  AND U1644 ( .A(a[66]), .B(b[66]), .Z(n1419) );
  ANDN U1645 ( .B(n1417), .A(n1419), .Z(n1426) );
  NOR U1646 ( .A(n1421), .B(n1420), .Z(n1418) );
  XNOR U1647 ( .A(n1419), .B(n1418), .Z(n1424) );
  XOR U1648 ( .A(n1421), .B(n1420), .Z(n1422) );
  NAND U1649 ( .A(n1422), .B(n2853), .Z(n1423) );
  NAND U1650 ( .A(n1424), .B(n1423), .Z(n2858) );
  XNOR U1651 ( .A(a[67]), .B(b[67]), .Z(n2857) );
  NAND U1652 ( .A(n2858), .B(n2857), .Z(n1425) );
  NANDN U1653 ( .A(n1426), .B(n1425), .Z(n1432) );
  NAND U1654 ( .A(a[67]), .B(b[67]), .Z(n1433) );
  AND U1655 ( .A(n1432), .B(n1433), .Z(n1428) );
  XOR U1656 ( .A(a[68]), .B(b[68]), .Z(n2863) );
  ANDN U1657 ( .B(n2862), .A(n2863), .Z(n1427) );
  OR U1658 ( .A(n1428), .B(n1427), .Z(n1429) );
  AND U1659 ( .A(a[68]), .B(b[68]), .Z(n1431) );
  ANDN U1660 ( .B(n1429), .A(n1431), .Z(n1438) );
  NOR U1661 ( .A(n1433), .B(n1432), .Z(n1430) );
  XNOR U1662 ( .A(n1431), .B(n1430), .Z(n1436) );
  XOR U1663 ( .A(n1433), .B(n1432), .Z(n1434) );
  NAND U1664 ( .A(n1434), .B(n2863), .Z(n1435) );
  NAND U1665 ( .A(n1436), .B(n1435), .Z(n2868) );
  XNOR U1666 ( .A(a[69]), .B(b[69]), .Z(n2867) );
  NAND U1667 ( .A(n2868), .B(n2867), .Z(n1437) );
  NANDN U1668 ( .A(n1438), .B(n1437), .Z(n1444) );
  NAND U1669 ( .A(a[69]), .B(b[69]), .Z(n1445) );
  AND U1670 ( .A(n1444), .B(n1445), .Z(n1440) );
  XOR U1671 ( .A(a[70]), .B(b[70]), .Z(n2873) );
  ANDN U1672 ( .B(n2872), .A(n2873), .Z(n1439) );
  OR U1673 ( .A(n1440), .B(n1439), .Z(n1441) );
  AND U1674 ( .A(a[70]), .B(b[70]), .Z(n1443) );
  ANDN U1675 ( .B(n1441), .A(n1443), .Z(n1450) );
  NOR U1676 ( .A(n1445), .B(n1444), .Z(n1442) );
  XNOR U1677 ( .A(n1443), .B(n1442), .Z(n1448) );
  XOR U1678 ( .A(n1445), .B(n1444), .Z(n1446) );
  NAND U1679 ( .A(n1446), .B(n2873), .Z(n1447) );
  NAND U1680 ( .A(n1448), .B(n1447), .Z(n2878) );
  XNOR U1681 ( .A(a[71]), .B(b[71]), .Z(n2877) );
  NAND U1682 ( .A(n2878), .B(n2877), .Z(n1449) );
  NANDN U1683 ( .A(n1450), .B(n1449), .Z(n1456) );
  NAND U1684 ( .A(a[71]), .B(b[71]), .Z(n1457) );
  AND U1685 ( .A(n1456), .B(n1457), .Z(n1452) );
  XOR U1686 ( .A(a[72]), .B(b[72]), .Z(n2883) );
  ANDN U1687 ( .B(n2882), .A(n2883), .Z(n1451) );
  OR U1688 ( .A(n1452), .B(n1451), .Z(n1453) );
  AND U1689 ( .A(a[72]), .B(b[72]), .Z(n1455) );
  ANDN U1690 ( .B(n1453), .A(n1455), .Z(n1462) );
  NOR U1691 ( .A(n1457), .B(n1456), .Z(n1454) );
  XNOR U1692 ( .A(n1455), .B(n1454), .Z(n1460) );
  XOR U1693 ( .A(n1457), .B(n1456), .Z(n1458) );
  NAND U1694 ( .A(n1458), .B(n2883), .Z(n1459) );
  NAND U1695 ( .A(n1460), .B(n1459), .Z(n2888) );
  XNOR U1696 ( .A(a[73]), .B(b[73]), .Z(n2887) );
  NAND U1697 ( .A(n2888), .B(n2887), .Z(n1461) );
  NANDN U1698 ( .A(n1462), .B(n1461), .Z(n1468) );
  NAND U1699 ( .A(a[73]), .B(b[73]), .Z(n1469) );
  AND U1700 ( .A(n1468), .B(n1469), .Z(n1464) );
  XOR U1701 ( .A(a[74]), .B(b[74]), .Z(n2893) );
  ANDN U1702 ( .B(n2892), .A(n2893), .Z(n1463) );
  OR U1703 ( .A(n1464), .B(n1463), .Z(n1465) );
  AND U1704 ( .A(a[74]), .B(b[74]), .Z(n1467) );
  ANDN U1705 ( .B(n1465), .A(n1467), .Z(n1474) );
  NOR U1706 ( .A(n1469), .B(n1468), .Z(n1466) );
  XNOR U1707 ( .A(n1467), .B(n1466), .Z(n1472) );
  XOR U1708 ( .A(n1469), .B(n1468), .Z(n1470) );
  NAND U1709 ( .A(n1470), .B(n2893), .Z(n1471) );
  NAND U1710 ( .A(n1472), .B(n1471), .Z(n2898) );
  XNOR U1711 ( .A(a[75]), .B(b[75]), .Z(n2897) );
  NAND U1712 ( .A(n2898), .B(n2897), .Z(n1473) );
  NANDN U1713 ( .A(n1474), .B(n1473), .Z(n1480) );
  NAND U1714 ( .A(a[75]), .B(b[75]), .Z(n1481) );
  AND U1715 ( .A(n1480), .B(n1481), .Z(n1476) );
  XOR U1716 ( .A(a[76]), .B(b[76]), .Z(n2903) );
  ANDN U1717 ( .B(n2902), .A(n2903), .Z(n1475) );
  OR U1718 ( .A(n1476), .B(n1475), .Z(n1477) );
  AND U1719 ( .A(a[76]), .B(b[76]), .Z(n1479) );
  ANDN U1720 ( .B(n1477), .A(n1479), .Z(n1486) );
  NOR U1721 ( .A(n1481), .B(n1480), .Z(n1478) );
  XNOR U1722 ( .A(n1479), .B(n1478), .Z(n1484) );
  XOR U1723 ( .A(n1481), .B(n1480), .Z(n1482) );
  NAND U1724 ( .A(n1482), .B(n2903), .Z(n1483) );
  NAND U1725 ( .A(n1484), .B(n1483), .Z(n2908) );
  XNOR U1726 ( .A(a[77]), .B(b[77]), .Z(n2907) );
  NAND U1727 ( .A(n2908), .B(n2907), .Z(n1485) );
  NANDN U1728 ( .A(n1486), .B(n1485), .Z(n1492) );
  NAND U1729 ( .A(a[77]), .B(b[77]), .Z(n1493) );
  AND U1730 ( .A(n1492), .B(n1493), .Z(n1488) );
  XOR U1731 ( .A(a[78]), .B(b[78]), .Z(n2913) );
  ANDN U1732 ( .B(n2912), .A(n2913), .Z(n1487) );
  OR U1733 ( .A(n1488), .B(n1487), .Z(n1489) );
  AND U1734 ( .A(a[78]), .B(b[78]), .Z(n1491) );
  ANDN U1735 ( .B(n1489), .A(n1491), .Z(n1498) );
  NOR U1736 ( .A(n1493), .B(n1492), .Z(n1490) );
  XNOR U1737 ( .A(n1491), .B(n1490), .Z(n1496) );
  XOR U1738 ( .A(n1493), .B(n1492), .Z(n1494) );
  NAND U1739 ( .A(n1494), .B(n2913), .Z(n1495) );
  NAND U1740 ( .A(n1496), .B(n1495), .Z(n2918) );
  XNOR U1741 ( .A(a[79]), .B(b[79]), .Z(n2917) );
  NAND U1742 ( .A(n2918), .B(n2917), .Z(n1497) );
  NANDN U1743 ( .A(n1498), .B(n1497), .Z(n1504) );
  NAND U1744 ( .A(a[79]), .B(b[79]), .Z(n1505) );
  AND U1745 ( .A(n1504), .B(n1505), .Z(n1500) );
  XOR U1746 ( .A(a[80]), .B(b[80]), .Z(n2923) );
  ANDN U1747 ( .B(n2922), .A(n2923), .Z(n1499) );
  OR U1748 ( .A(n1500), .B(n1499), .Z(n1501) );
  AND U1749 ( .A(a[80]), .B(b[80]), .Z(n1503) );
  ANDN U1750 ( .B(n1501), .A(n1503), .Z(n1510) );
  NOR U1751 ( .A(n1505), .B(n1504), .Z(n1502) );
  XNOR U1752 ( .A(n1503), .B(n1502), .Z(n1508) );
  XOR U1753 ( .A(n1505), .B(n1504), .Z(n1506) );
  NAND U1754 ( .A(n1506), .B(n2923), .Z(n1507) );
  NAND U1755 ( .A(n1508), .B(n1507), .Z(n2928) );
  XNOR U1756 ( .A(a[81]), .B(b[81]), .Z(n2927) );
  NAND U1757 ( .A(n2928), .B(n2927), .Z(n1509) );
  NANDN U1758 ( .A(n1510), .B(n1509), .Z(n1516) );
  NAND U1759 ( .A(a[81]), .B(b[81]), .Z(n1517) );
  AND U1760 ( .A(n1516), .B(n1517), .Z(n1512) );
  XOR U1761 ( .A(a[82]), .B(b[82]), .Z(n2933) );
  ANDN U1762 ( .B(n2932), .A(n2933), .Z(n1511) );
  OR U1763 ( .A(n1512), .B(n1511), .Z(n1513) );
  AND U1764 ( .A(a[82]), .B(b[82]), .Z(n1515) );
  ANDN U1765 ( .B(n1513), .A(n1515), .Z(n1522) );
  NOR U1766 ( .A(n1517), .B(n1516), .Z(n1514) );
  XNOR U1767 ( .A(n1515), .B(n1514), .Z(n1520) );
  XOR U1768 ( .A(n1517), .B(n1516), .Z(n1518) );
  NAND U1769 ( .A(n1518), .B(n2933), .Z(n1519) );
  NAND U1770 ( .A(n1520), .B(n1519), .Z(n2938) );
  XNOR U1771 ( .A(a[83]), .B(b[83]), .Z(n2937) );
  NAND U1772 ( .A(n2938), .B(n2937), .Z(n1521) );
  NANDN U1773 ( .A(n1522), .B(n1521), .Z(n1523) );
  IV U1774 ( .A(n1523), .Z(n1527) );
  AND U1775 ( .A(a[83]), .B(b[83]), .Z(n1528) );
  NOR U1776 ( .A(n1527), .B(n1528), .Z(n1525) );
  XNOR U1777 ( .A(n1528), .B(n1523), .Z(n2943) );
  XNOR U1778 ( .A(a[84]), .B(b[84]), .Z(n2942) );
  AND U1779 ( .A(n2943), .B(n2942), .Z(n1524) );
  OR U1780 ( .A(n1525), .B(n1524), .Z(n1526) );
  AND U1781 ( .A(a[84]), .B(b[84]), .Z(n1530) );
  ANDN U1782 ( .B(n1526), .A(n1530), .Z(n1532) );
  AND U1783 ( .A(n1528), .B(n1527), .Z(n1529) );
  NAND U1784 ( .A(n1530), .B(n1529), .Z(n1535) );
  ANDN U1785 ( .B(n1535), .A(n1532), .Z(n2948) );
  XNOR U1786 ( .A(a[85]), .B(b[85]), .Z(n2947) );
  AND U1787 ( .A(n2948), .B(n2947), .Z(n1531) );
  OR U1788 ( .A(n1532), .B(n1531), .Z(n1533) );
  AND U1789 ( .A(n1534), .B(n1533), .Z(n1538) );
  OR U1790 ( .A(n1535), .B(n1534), .Z(n1536) );
  ANDN U1791 ( .B(n1536), .A(n1538), .Z(n2953) );
  XNOR U1792 ( .A(a[86]), .B(b[86]), .Z(n2952) );
  NAND U1793 ( .A(n2953), .B(n2952), .Z(n1537) );
  NANDN U1794 ( .A(n1538), .B(n1537), .Z(n1544) );
  NAND U1795 ( .A(a[86]), .B(b[86]), .Z(n1545) );
  AND U1796 ( .A(n1544), .B(n1545), .Z(n1540) );
  XOR U1797 ( .A(a[87]), .B(b[87]), .Z(n2958) );
  ANDN U1798 ( .B(n2957), .A(n2958), .Z(n1539) );
  OR U1799 ( .A(n1540), .B(n1539), .Z(n1541) );
  AND U1800 ( .A(a[87]), .B(b[87]), .Z(n1543) );
  ANDN U1801 ( .B(n1541), .A(n1543), .Z(n1550) );
  NOR U1802 ( .A(n1545), .B(n1544), .Z(n1542) );
  XNOR U1803 ( .A(n1543), .B(n1542), .Z(n1548) );
  XOR U1804 ( .A(n1545), .B(n1544), .Z(n1546) );
  NAND U1805 ( .A(n1546), .B(n2958), .Z(n1547) );
  NAND U1806 ( .A(n1548), .B(n1547), .Z(n2963) );
  XNOR U1807 ( .A(a[88]), .B(b[88]), .Z(n2962) );
  NAND U1808 ( .A(n2963), .B(n2962), .Z(n1549) );
  NANDN U1809 ( .A(n1550), .B(n1549), .Z(n1551) );
  IV U1810 ( .A(n1551), .Z(n1555) );
  AND U1811 ( .A(a[88]), .B(b[88]), .Z(n1556) );
  NOR U1812 ( .A(n1555), .B(n1556), .Z(n1553) );
  XNOR U1813 ( .A(n1556), .B(n1551), .Z(n2968) );
  XNOR U1814 ( .A(a[89]), .B(b[89]), .Z(n2967) );
  AND U1815 ( .A(n2968), .B(n2967), .Z(n1552) );
  OR U1816 ( .A(n1553), .B(n1552), .Z(n1554) );
  AND U1817 ( .A(a[89]), .B(b[89]), .Z(n1558) );
  ANDN U1818 ( .B(n1554), .A(n1558), .Z(n1560) );
  AND U1819 ( .A(n1556), .B(n1555), .Z(n1557) );
  NAND U1820 ( .A(n1558), .B(n1557), .Z(n1563) );
  ANDN U1821 ( .B(n1563), .A(n1560), .Z(n2973) );
  XNOR U1822 ( .A(a[90]), .B(b[90]), .Z(n2972) );
  AND U1823 ( .A(n2973), .B(n2972), .Z(n1559) );
  OR U1824 ( .A(n1560), .B(n1559), .Z(n1561) );
  AND U1825 ( .A(a[90]), .B(b[90]), .Z(n1562) );
  ANDN U1826 ( .B(n1561), .A(n1562), .Z(n1566) );
  NANDN U1827 ( .A(n1563), .B(n1562), .Z(n1564) );
  ANDN U1828 ( .B(n1564), .A(n1566), .Z(n2978) );
  XNOR U1829 ( .A(a[91]), .B(b[91]), .Z(n2977) );
  NAND U1830 ( .A(n2978), .B(n2977), .Z(n1565) );
  NANDN U1831 ( .A(n1566), .B(n1565), .Z(n1572) );
  NAND U1832 ( .A(a[91]), .B(b[91]), .Z(n1573) );
  AND U1833 ( .A(n1572), .B(n1573), .Z(n1568) );
  XOR U1834 ( .A(a[92]), .B(b[92]), .Z(n2983) );
  ANDN U1835 ( .B(n2982), .A(n2983), .Z(n1567) );
  OR U1836 ( .A(n1568), .B(n1567), .Z(n1569) );
  AND U1837 ( .A(a[92]), .B(b[92]), .Z(n1571) );
  ANDN U1838 ( .B(n1569), .A(n1571), .Z(n1578) );
  NOR U1839 ( .A(n1573), .B(n1572), .Z(n1570) );
  XNOR U1840 ( .A(n1571), .B(n1570), .Z(n1576) );
  XOR U1841 ( .A(n1573), .B(n1572), .Z(n1574) );
  NAND U1842 ( .A(n1574), .B(n2983), .Z(n1575) );
  NAND U1843 ( .A(n1576), .B(n1575), .Z(n2988) );
  XNOR U1844 ( .A(a[93]), .B(b[93]), .Z(n2987) );
  NAND U1845 ( .A(n2988), .B(n2987), .Z(n1577) );
  NANDN U1846 ( .A(n1578), .B(n1577), .Z(n1579) );
  IV U1847 ( .A(n1579), .Z(n1583) );
  AND U1848 ( .A(a[93]), .B(b[93]), .Z(n1584) );
  NOR U1849 ( .A(n1583), .B(n1584), .Z(n1581) );
  XNOR U1850 ( .A(n1584), .B(n1579), .Z(n2993) );
  XNOR U1851 ( .A(a[94]), .B(b[94]), .Z(n2992) );
  AND U1852 ( .A(n2993), .B(n2992), .Z(n1580) );
  OR U1853 ( .A(n1581), .B(n1580), .Z(n1582) );
  AND U1854 ( .A(a[94]), .B(b[94]), .Z(n1586) );
  ANDN U1855 ( .B(n1582), .A(n1586), .Z(n1588) );
  AND U1856 ( .A(n1584), .B(n1583), .Z(n1585) );
  NAND U1857 ( .A(n1586), .B(n1585), .Z(n1591) );
  ANDN U1858 ( .B(n1591), .A(n1588), .Z(n2998) );
  XNOR U1859 ( .A(a[95]), .B(b[95]), .Z(n2997) );
  AND U1860 ( .A(n2998), .B(n2997), .Z(n1587) );
  OR U1861 ( .A(n1588), .B(n1587), .Z(n1589) );
  AND U1862 ( .A(a[95]), .B(b[95]), .Z(n1590) );
  ANDN U1863 ( .B(n1589), .A(n1590), .Z(n1594) );
  NANDN U1864 ( .A(n1591), .B(n1590), .Z(n1592) );
  ANDN U1865 ( .B(n1592), .A(n1594), .Z(n3003) );
  XNOR U1866 ( .A(a[96]), .B(b[96]), .Z(n3002) );
  NAND U1867 ( .A(n3003), .B(n3002), .Z(n1593) );
  NANDN U1868 ( .A(n1594), .B(n1593), .Z(n1600) );
  NAND U1869 ( .A(a[96]), .B(b[96]), .Z(n1601) );
  AND U1870 ( .A(n1600), .B(n1601), .Z(n1596) );
  XOR U1871 ( .A(a[97]), .B(b[97]), .Z(n3008) );
  ANDN U1872 ( .B(n3007), .A(n3008), .Z(n1595) );
  OR U1873 ( .A(n1596), .B(n1595), .Z(n1597) );
  AND U1874 ( .A(a[97]), .B(b[97]), .Z(n1599) );
  ANDN U1875 ( .B(n1597), .A(n1599), .Z(n1606) );
  NOR U1876 ( .A(n1601), .B(n1600), .Z(n1598) );
  XNOR U1877 ( .A(n1599), .B(n1598), .Z(n1604) );
  XOR U1878 ( .A(n1601), .B(n1600), .Z(n1602) );
  NAND U1879 ( .A(n1602), .B(n3008), .Z(n1603) );
  NAND U1880 ( .A(n1604), .B(n1603), .Z(n3013) );
  XNOR U1881 ( .A(a[98]), .B(b[98]), .Z(n3012) );
  NAND U1882 ( .A(n3013), .B(n3012), .Z(n1605) );
  NANDN U1883 ( .A(n1606), .B(n1605), .Z(n1612) );
  NAND U1884 ( .A(a[98]), .B(b[98]), .Z(n1613) );
  AND U1885 ( .A(n1612), .B(n1613), .Z(n1608) );
  XOR U1886 ( .A(a[99]), .B(b[99]), .Z(n3018) );
  ANDN U1887 ( .B(n3017), .A(n3018), .Z(n1607) );
  OR U1888 ( .A(n1608), .B(n1607), .Z(n1609) );
  AND U1889 ( .A(a[99]), .B(b[99]), .Z(n1611) );
  ANDN U1890 ( .B(n1609), .A(n1611), .Z(n1618) );
  NOR U1891 ( .A(n1613), .B(n1612), .Z(n1610) );
  XNOR U1892 ( .A(n1611), .B(n1610), .Z(n1616) );
  XOR U1893 ( .A(n1613), .B(n1612), .Z(n1614) );
  NAND U1894 ( .A(n1614), .B(n3018), .Z(n1615) );
  NAND U1895 ( .A(n1616), .B(n1615), .Z(n3023) );
  XNOR U1896 ( .A(a[100]), .B(b[100]), .Z(n3022) );
  NAND U1897 ( .A(n3023), .B(n3022), .Z(n1617) );
  NANDN U1898 ( .A(n1618), .B(n1617), .Z(n1624) );
  NAND U1899 ( .A(a[100]), .B(b[100]), .Z(n1625) );
  AND U1900 ( .A(n1624), .B(n1625), .Z(n1620) );
  XOR U1901 ( .A(a[101]), .B(b[101]), .Z(n3028) );
  ANDN U1902 ( .B(n3027), .A(n3028), .Z(n1619) );
  OR U1903 ( .A(n1620), .B(n1619), .Z(n1621) );
  AND U1904 ( .A(a[101]), .B(b[101]), .Z(n1623) );
  ANDN U1905 ( .B(n1621), .A(n1623), .Z(n1630) );
  NOR U1906 ( .A(n1625), .B(n1624), .Z(n1622) );
  XNOR U1907 ( .A(n1623), .B(n1622), .Z(n1628) );
  XOR U1908 ( .A(n1625), .B(n1624), .Z(n1626) );
  NAND U1909 ( .A(n1626), .B(n3028), .Z(n1627) );
  NAND U1910 ( .A(n1628), .B(n1627), .Z(n3033) );
  XNOR U1911 ( .A(a[102]), .B(b[102]), .Z(n3032) );
  NAND U1912 ( .A(n3033), .B(n3032), .Z(n1629) );
  NANDN U1913 ( .A(n1630), .B(n1629), .Z(n1636) );
  NAND U1914 ( .A(a[102]), .B(b[102]), .Z(n1637) );
  AND U1915 ( .A(n1636), .B(n1637), .Z(n1632) );
  XOR U1916 ( .A(a[103]), .B(b[103]), .Z(n3038) );
  ANDN U1917 ( .B(n3037), .A(n3038), .Z(n1631) );
  OR U1918 ( .A(n1632), .B(n1631), .Z(n1633) );
  AND U1919 ( .A(a[103]), .B(b[103]), .Z(n1635) );
  ANDN U1920 ( .B(n1633), .A(n1635), .Z(n1642) );
  NOR U1921 ( .A(n1637), .B(n1636), .Z(n1634) );
  XNOR U1922 ( .A(n1635), .B(n1634), .Z(n1640) );
  XOR U1923 ( .A(n1637), .B(n1636), .Z(n1638) );
  NAND U1924 ( .A(n1638), .B(n3038), .Z(n1639) );
  NAND U1925 ( .A(n1640), .B(n1639), .Z(n3043) );
  XNOR U1926 ( .A(a[104]), .B(b[104]), .Z(n3042) );
  NAND U1927 ( .A(n3043), .B(n3042), .Z(n1641) );
  NANDN U1928 ( .A(n1642), .B(n1641), .Z(n1648) );
  NAND U1929 ( .A(a[104]), .B(b[104]), .Z(n1649) );
  AND U1930 ( .A(n1648), .B(n1649), .Z(n1644) );
  XOR U1931 ( .A(a[105]), .B(b[105]), .Z(n3048) );
  ANDN U1932 ( .B(n3047), .A(n3048), .Z(n1643) );
  OR U1933 ( .A(n1644), .B(n1643), .Z(n1645) );
  AND U1934 ( .A(a[105]), .B(b[105]), .Z(n1647) );
  ANDN U1935 ( .B(n1645), .A(n1647), .Z(n1654) );
  NOR U1936 ( .A(n1649), .B(n1648), .Z(n1646) );
  XNOR U1937 ( .A(n1647), .B(n1646), .Z(n1652) );
  XOR U1938 ( .A(n1649), .B(n1648), .Z(n1650) );
  NAND U1939 ( .A(n1650), .B(n3048), .Z(n1651) );
  NAND U1940 ( .A(n1652), .B(n1651), .Z(n3053) );
  XNOR U1941 ( .A(a[106]), .B(b[106]), .Z(n3052) );
  NAND U1942 ( .A(n3053), .B(n3052), .Z(n1653) );
  NANDN U1943 ( .A(n1654), .B(n1653), .Z(n1660) );
  NAND U1944 ( .A(a[106]), .B(b[106]), .Z(n1661) );
  AND U1945 ( .A(n1660), .B(n1661), .Z(n1656) );
  XOR U1946 ( .A(a[107]), .B(b[107]), .Z(n3058) );
  ANDN U1947 ( .B(n3057), .A(n3058), .Z(n1655) );
  OR U1948 ( .A(n1656), .B(n1655), .Z(n1657) );
  AND U1949 ( .A(a[107]), .B(b[107]), .Z(n1659) );
  ANDN U1950 ( .B(n1657), .A(n1659), .Z(n1666) );
  NOR U1951 ( .A(n1661), .B(n1660), .Z(n1658) );
  XNOR U1952 ( .A(n1659), .B(n1658), .Z(n1664) );
  XOR U1953 ( .A(n1661), .B(n1660), .Z(n1662) );
  NAND U1954 ( .A(n1662), .B(n3058), .Z(n1663) );
  NAND U1955 ( .A(n1664), .B(n1663), .Z(n3063) );
  XNOR U1956 ( .A(a[108]), .B(b[108]), .Z(n3062) );
  NAND U1957 ( .A(n3063), .B(n3062), .Z(n1665) );
  NANDN U1958 ( .A(n1666), .B(n1665), .Z(n1672) );
  NAND U1959 ( .A(a[108]), .B(b[108]), .Z(n1673) );
  AND U1960 ( .A(n1672), .B(n1673), .Z(n1668) );
  XOR U1961 ( .A(a[109]), .B(b[109]), .Z(n3068) );
  ANDN U1962 ( .B(n3067), .A(n3068), .Z(n1667) );
  OR U1963 ( .A(n1668), .B(n1667), .Z(n1669) );
  AND U1964 ( .A(a[109]), .B(b[109]), .Z(n1671) );
  ANDN U1965 ( .B(n1669), .A(n1671), .Z(n1678) );
  NOR U1966 ( .A(n1673), .B(n1672), .Z(n1670) );
  XNOR U1967 ( .A(n1671), .B(n1670), .Z(n1676) );
  XOR U1968 ( .A(n1673), .B(n1672), .Z(n1674) );
  NAND U1969 ( .A(n1674), .B(n3068), .Z(n1675) );
  NAND U1970 ( .A(n1676), .B(n1675), .Z(n3073) );
  XNOR U1971 ( .A(a[110]), .B(b[110]), .Z(n3072) );
  NAND U1972 ( .A(n3073), .B(n3072), .Z(n1677) );
  NANDN U1973 ( .A(n1678), .B(n1677), .Z(n1684) );
  NAND U1974 ( .A(a[110]), .B(b[110]), .Z(n1685) );
  AND U1975 ( .A(n1684), .B(n1685), .Z(n1680) );
  XOR U1976 ( .A(a[111]), .B(b[111]), .Z(n3078) );
  ANDN U1977 ( .B(n3077), .A(n3078), .Z(n1679) );
  OR U1978 ( .A(n1680), .B(n1679), .Z(n1681) );
  AND U1979 ( .A(a[111]), .B(b[111]), .Z(n1683) );
  ANDN U1980 ( .B(n1681), .A(n1683), .Z(n1690) );
  NOR U1981 ( .A(n1685), .B(n1684), .Z(n1682) );
  XNOR U1982 ( .A(n1683), .B(n1682), .Z(n1688) );
  XOR U1983 ( .A(n1685), .B(n1684), .Z(n1686) );
  NAND U1984 ( .A(n1686), .B(n3078), .Z(n1687) );
  NAND U1985 ( .A(n1688), .B(n1687), .Z(n3083) );
  XNOR U1986 ( .A(a[112]), .B(b[112]), .Z(n3082) );
  NAND U1987 ( .A(n3083), .B(n3082), .Z(n1689) );
  NANDN U1988 ( .A(n1690), .B(n1689), .Z(n1696) );
  NAND U1989 ( .A(a[112]), .B(b[112]), .Z(n1697) );
  AND U1990 ( .A(n1696), .B(n1697), .Z(n1692) );
  XOR U1991 ( .A(a[113]), .B(b[113]), .Z(n3088) );
  ANDN U1992 ( .B(n3087), .A(n3088), .Z(n1691) );
  OR U1993 ( .A(n1692), .B(n1691), .Z(n1693) );
  AND U1994 ( .A(a[113]), .B(b[113]), .Z(n1695) );
  ANDN U1995 ( .B(n1693), .A(n1695), .Z(n1702) );
  NOR U1996 ( .A(n1697), .B(n1696), .Z(n1694) );
  XNOR U1997 ( .A(n1695), .B(n1694), .Z(n1700) );
  XOR U1998 ( .A(n1697), .B(n1696), .Z(n1698) );
  NAND U1999 ( .A(n1698), .B(n3088), .Z(n1699) );
  NAND U2000 ( .A(n1700), .B(n1699), .Z(n3093) );
  XNOR U2001 ( .A(a[114]), .B(b[114]), .Z(n3092) );
  NAND U2002 ( .A(n3093), .B(n3092), .Z(n1701) );
  NANDN U2003 ( .A(n1702), .B(n1701), .Z(n1708) );
  NAND U2004 ( .A(a[114]), .B(b[114]), .Z(n1709) );
  AND U2005 ( .A(n1708), .B(n1709), .Z(n1704) );
  XOR U2006 ( .A(a[115]), .B(b[115]), .Z(n3098) );
  ANDN U2007 ( .B(n3097), .A(n3098), .Z(n1703) );
  OR U2008 ( .A(n1704), .B(n1703), .Z(n1705) );
  AND U2009 ( .A(a[115]), .B(b[115]), .Z(n1707) );
  ANDN U2010 ( .B(n1705), .A(n1707), .Z(n1714) );
  NOR U2011 ( .A(n1709), .B(n1708), .Z(n1706) );
  XNOR U2012 ( .A(n1707), .B(n1706), .Z(n1712) );
  XOR U2013 ( .A(n1709), .B(n1708), .Z(n1710) );
  NAND U2014 ( .A(n1710), .B(n3098), .Z(n1711) );
  NAND U2015 ( .A(n1712), .B(n1711), .Z(n3103) );
  XNOR U2016 ( .A(a[116]), .B(b[116]), .Z(n3102) );
  NAND U2017 ( .A(n3103), .B(n3102), .Z(n1713) );
  NANDN U2018 ( .A(n1714), .B(n1713), .Z(n1720) );
  NAND U2019 ( .A(a[116]), .B(b[116]), .Z(n1721) );
  AND U2020 ( .A(n1720), .B(n1721), .Z(n1716) );
  XOR U2021 ( .A(a[117]), .B(b[117]), .Z(n3108) );
  ANDN U2022 ( .B(n3107), .A(n3108), .Z(n1715) );
  OR U2023 ( .A(n1716), .B(n1715), .Z(n1717) );
  AND U2024 ( .A(a[117]), .B(b[117]), .Z(n1719) );
  ANDN U2025 ( .B(n1717), .A(n1719), .Z(n1726) );
  NOR U2026 ( .A(n1721), .B(n1720), .Z(n1718) );
  XNOR U2027 ( .A(n1719), .B(n1718), .Z(n1724) );
  XOR U2028 ( .A(n1721), .B(n1720), .Z(n1722) );
  NAND U2029 ( .A(n1722), .B(n3108), .Z(n1723) );
  NAND U2030 ( .A(n1724), .B(n1723), .Z(n3113) );
  XNOR U2031 ( .A(a[118]), .B(b[118]), .Z(n3112) );
  NAND U2032 ( .A(n3113), .B(n3112), .Z(n1725) );
  NANDN U2033 ( .A(n1726), .B(n1725), .Z(n1732) );
  NAND U2034 ( .A(a[118]), .B(b[118]), .Z(n1733) );
  AND U2035 ( .A(n1732), .B(n1733), .Z(n1728) );
  XOR U2036 ( .A(a[119]), .B(b[119]), .Z(n3118) );
  ANDN U2037 ( .B(n3117), .A(n3118), .Z(n1727) );
  OR U2038 ( .A(n1728), .B(n1727), .Z(n1729) );
  AND U2039 ( .A(a[119]), .B(b[119]), .Z(n1731) );
  ANDN U2040 ( .B(n1729), .A(n1731), .Z(n1738) );
  NOR U2041 ( .A(n1733), .B(n1732), .Z(n1730) );
  XNOR U2042 ( .A(n1731), .B(n1730), .Z(n1736) );
  XOR U2043 ( .A(n1733), .B(n1732), .Z(n1734) );
  NAND U2044 ( .A(n1734), .B(n3118), .Z(n1735) );
  NAND U2045 ( .A(n1736), .B(n1735), .Z(n3123) );
  XNOR U2046 ( .A(a[120]), .B(b[120]), .Z(n3122) );
  NAND U2047 ( .A(n3123), .B(n3122), .Z(n1737) );
  NANDN U2048 ( .A(n1738), .B(n1737), .Z(n1744) );
  NAND U2049 ( .A(a[120]), .B(b[120]), .Z(n1745) );
  AND U2050 ( .A(n1744), .B(n1745), .Z(n1740) );
  XOR U2051 ( .A(a[121]), .B(b[121]), .Z(n3128) );
  ANDN U2052 ( .B(n3127), .A(n3128), .Z(n1739) );
  OR U2053 ( .A(n1740), .B(n1739), .Z(n1741) );
  AND U2054 ( .A(a[121]), .B(b[121]), .Z(n1743) );
  ANDN U2055 ( .B(n1741), .A(n1743), .Z(n1750) );
  NOR U2056 ( .A(n1745), .B(n1744), .Z(n1742) );
  XNOR U2057 ( .A(n1743), .B(n1742), .Z(n1748) );
  XOR U2058 ( .A(n1745), .B(n1744), .Z(n1746) );
  NAND U2059 ( .A(n1746), .B(n3128), .Z(n1747) );
  NAND U2060 ( .A(n1748), .B(n1747), .Z(n3133) );
  XNOR U2061 ( .A(a[122]), .B(b[122]), .Z(n3132) );
  NAND U2062 ( .A(n3133), .B(n3132), .Z(n1749) );
  NANDN U2063 ( .A(n1750), .B(n1749), .Z(n1756) );
  NAND U2064 ( .A(a[122]), .B(b[122]), .Z(n1757) );
  AND U2065 ( .A(n1756), .B(n1757), .Z(n1752) );
  XOR U2066 ( .A(a[123]), .B(b[123]), .Z(n3138) );
  ANDN U2067 ( .B(n3137), .A(n3138), .Z(n1751) );
  OR U2068 ( .A(n1752), .B(n1751), .Z(n1753) );
  AND U2069 ( .A(a[123]), .B(b[123]), .Z(n1755) );
  ANDN U2070 ( .B(n1753), .A(n1755), .Z(n1762) );
  NOR U2071 ( .A(n1757), .B(n1756), .Z(n1754) );
  XNOR U2072 ( .A(n1755), .B(n1754), .Z(n1760) );
  XOR U2073 ( .A(n1757), .B(n1756), .Z(n1758) );
  NAND U2074 ( .A(n1758), .B(n3138), .Z(n1759) );
  NAND U2075 ( .A(n1760), .B(n1759), .Z(n3143) );
  XNOR U2076 ( .A(a[124]), .B(b[124]), .Z(n3142) );
  NAND U2077 ( .A(n3143), .B(n3142), .Z(n1761) );
  NANDN U2078 ( .A(n1762), .B(n1761), .Z(n1763) );
  IV U2079 ( .A(n1763), .Z(n1767) );
  AND U2080 ( .A(a[124]), .B(b[124]), .Z(n1768) );
  NOR U2081 ( .A(n1767), .B(n1768), .Z(n1765) );
  XNOR U2082 ( .A(n1768), .B(n1763), .Z(n3148) );
  XNOR U2083 ( .A(a[125]), .B(b[125]), .Z(n3147) );
  AND U2084 ( .A(n3148), .B(n3147), .Z(n1764) );
  OR U2085 ( .A(n1765), .B(n1764), .Z(n1766) );
  AND U2086 ( .A(a[125]), .B(b[125]), .Z(n1770) );
  ANDN U2087 ( .B(n1766), .A(n1770), .Z(n1772) );
  AND U2088 ( .A(n1768), .B(n1767), .Z(n1769) );
  NAND U2089 ( .A(n1770), .B(n1769), .Z(n1775) );
  ANDN U2090 ( .B(n1775), .A(n1772), .Z(n3153) );
  XNOR U2091 ( .A(a[126]), .B(b[126]), .Z(n3152) );
  AND U2092 ( .A(n3153), .B(n3152), .Z(n1771) );
  OR U2093 ( .A(n1772), .B(n1771), .Z(n1773) );
  AND U2094 ( .A(n1774), .B(n1773), .Z(n1778) );
  OR U2095 ( .A(n1775), .B(n1774), .Z(n1776) );
  ANDN U2096 ( .B(n1776), .A(n1778), .Z(n3158) );
  XNOR U2097 ( .A(a[127]), .B(b[127]), .Z(n3157) );
  NAND U2098 ( .A(n3158), .B(n3157), .Z(n1777) );
  NANDN U2099 ( .A(n1778), .B(n1777), .Z(n1784) );
  NAND U2100 ( .A(a[127]), .B(b[127]), .Z(n1785) );
  AND U2101 ( .A(n1784), .B(n1785), .Z(n1780) );
  XOR U2102 ( .A(a[128]), .B(b[128]), .Z(n3163) );
  ANDN U2103 ( .B(n3162), .A(n3163), .Z(n1779) );
  OR U2104 ( .A(n1780), .B(n1779), .Z(n1781) );
  AND U2105 ( .A(a[128]), .B(b[128]), .Z(n1783) );
  ANDN U2106 ( .B(n1781), .A(n1783), .Z(n1790) );
  NOR U2107 ( .A(n1785), .B(n1784), .Z(n1782) );
  XNOR U2108 ( .A(n1783), .B(n1782), .Z(n1788) );
  XOR U2109 ( .A(n1785), .B(n1784), .Z(n1786) );
  NAND U2110 ( .A(n1786), .B(n3163), .Z(n1787) );
  NAND U2111 ( .A(n1788), .B(n1787), .Z(n3168) );
  XNOR U2112 ( .A(a[129]), .B(b[129]), .Z(n3167) );
  NAND U2113 ( .A(n3168), .B(n3167), .Z(n1789) );
  NANDN U2114 ( .A(n1790), .B(n1789), .Z(n1796) );
  NAND U2115 ( .A(a[129]), .B(b[129]), .Z(n1797) );
  AND U2116 ( .A(n1796), .B(n1797), .Z(n1792) );
  XOR U2117 ( .A(a[130]), .B(b[130]), .Z(n3173) );
  ANDN U2118 ( .B(n3172), .A(n3173), .Z(n1791) );
  OR U2119 ( .A(n1792), .B(n1791), .Z(n1793) );
  AND U2120 ( .A(a[130]), .B(b[130]), .Z(n1795) );
  ANDN U2121 ( .B(n1793), .A(n1795), .Z(n1802) );
  NOR U2122 ( .A(n1797), .B(n1796), .Z(n1794) );
  XNOR U2123 ( .A(n1795), .B(n1794), .Z(n1800) );
  XOR U2124 ( .A(n1797), .B(n1796), .Z(n1798) );
  NAND U2125 ( .A(n1798), .B(n3173), .Z(n1799) );
  NAND U2126 ( .A(n1800), .B(n1799), .Z(n3178) );
  XNOR U2127 ( .A(a[131]), .B(b[131]), .Z(n3177) );
  NAND U2128 ( .A(n3178), .B(n3177), .Z(n1801) );
  NANDN U2129 ( .A(n1802), .B(n1801), .Z(n1808) );
  NAND U2130 ( .A(a[131]), .B(b[131]), .Z(n1809) );
  AND U2131 ( .A(n1808), .B(n1809), .Z(n1804) );
  XOR U2132 ( .A(a[132]), .B(b[132]), .Z(n3183) );
  ANDN U2133 ( .B(n3182), .A(n3183), .Z(n1803) );
  OR U2134 ( .A(n1804), .B(n1803), .Z(n1805) );
  AND U2135 ( .A(a[132]), .B(b[132]), .Z(n1807) );
  ANDN U2136 ( .B(n1805), .A(n1807), .Z(n1814) );
  NOR U2137 ( .A(n1809), .B(n1808), .Z(n1806) );
  XNOR U2138 ( .A(n1807), .B(n1806), .Z(n1812) );
  XOR U2139 ( .A(n1809), .B(n1808), .Z(n1810) );
  NAND U2140 ( .A(n1810), .B(n3183), .Z(n1811) );
  NAND U2141 ( .A(n1812), .B(n1811), .Z(n3188) );
  XNOR U2142 ( .A(a[133]), .B(b[133]), .Z(n3187) );
  NAND U2143 ( .A(n3188), .B(n3187), .Z(n1813) );
  NANDN U2144 ( .A(n1814), .B(n1813), .Z(n1820) );
  NAND U2145 ( .A(a[133]), .B(b[133]), .Z(n1821) );
  AND U2146 ( .A(n1820), .B(n1821), .Z(n1816) );
  XOR U2147 ( .A(a[134]), .B(b[134]), .Z(n3193) );
  ANDN U2148 ( .B(n3192), .A(n3193), .Z(n1815) );
  OR U2149 ( .A(n1816), .B(n1815), .Z(n1817) );
  AND U2150 ( .A(a[134]), .B(b[134]), .Z(n1819) );
  ANDN U2151 ( .B(n1817), .A(n1819), .Z(n1826) );
  NOR U2152 ( .A(n1821), .B(n1820), .Z(n1818) );
  XNOR U2153 ( .A(n1819), .B(n1818), .Z(n1824) );
  XOR U2154 ( .A(n1821), .B(n1820), .Z(n1822) );
  NAND U2155 ( .A(n1822), .B(n3193), .Z(n1823) );
  NAND U2156 ( .A(n1824), .B(n1823), .Z(n3198) );
  XNOR U2157 ( .A(a[135]), .B(b[135]), .Z(n3197) );
  NAND U2158 ( .A(n3198), .B(n3197), .Z(n1825) );
  NANDN U2159 ( .A(n1826), .B(n1825), .Z(n1832) );
  NAND U2160 ( .A(a[135]), .B(b[135]), .Z(n1833) );
  AND U2161 ( .A(n1832), .B(n1833), .Z(n1828) );
  XOR U2162 ( .A(a[136]), .B(b[136]), .Z(n3203) );
  ANDN U2163 ( .B(n3202), .A(n3203), .Z(n1827) );
  OR U2164 ( .A(n1828), .B(n1827), .Z(n1829) );
  AND U2165 ( .A(a[136]), .B(b[136]), .Z(n1831) );
  ANDN U2166 ( .B(n1829), .A(n1831), .Z(n1838) );
  NOR U2167 ( .A(n1833), .B(n1832), .Z(n1830) );
  XNOR U2168 ( .A(n1831), .B(n1830), .Z(n1836) );
  XOR U2169 ( .A(n1833), .B(n1832), .Z(n1834) );
  NAND U2170 ( .A(n1834), .B(n3203), .Z(n1835) );
  NAND U2171 ( .A(n1836), .B(n1835), .Z(n3208) );
  XNOR U2172 ( .A(a[137]), .B(b[137]), .Z(n3207) );
  NAND U2173 ( .A(n3208), .B(n3207), .Z(n1837) );
  NANDN U2174 ( .A(n1838), .B(n1837), .Z(n1844) );
  NAND U2175 ( .A(a[137]), .B(b[137]), .Z(n1845) );
  AND U2176 ( .A(n1844), .B(n1845), .Z(n1840) );
  XOR U2177 ( .A(a[138]), .B(b[138]), .Z(n3213) );
  ANDN U2178 ( .B(n3212), .A(n3213), .Z(n1839) );
  OR U2179 ( .A(n1840), .B(n1839), .Z(n1841) );
  AND U2180 ( .A(a[138]), .B(b[138]), .Z(n1843) );
  ANDN U2181 ( .B(n1841), .A(n1843), .Z(n1850) );
  NOR U2182 ( .A(n1845), .B(n1844), .Z(n1842) );
  XNOR U2183 ( .A(n1843), .B(n1842), .Z(n1848) );
  XOR U2184 ( .A(n1845), .B(n1844), .Z(n1846) );
  NAND U2185 ( .A(n1846), .B(n3213), .Z(n1847) );
  NAND U2186 ( .A(n1848), .B(n1847), .Z(n3218) );
  XNOR U2187 ( .A(a[139]), .B(b[139]), .Z(n3217) );
  NAND U2188 ( .A(n3218), .B(n3217), .Z(n1849) );
  NANDN U2189 ( .A(n1850), .B(n1849), .Z(n1856) );
  NAND U2190 ( .A(a[139]), .B(b[139]), .Z(n1857) );
  AND U2191 ( .A(n1856), .B(n1857), .Z(n1852) );
  XOR U2192 ( .A(a[140]), .B(b[140]), .Z(n3223) );
  ANDN U2193 ( .B(n3222), .A(n3223), .Z(n1851) );
  OR U2194 ( .A(n1852), .B(n1851), .Z(n1853) );
  AND U2195 ( .A(a[140]), .B(b[140]), .Z(n1855) );
  ANDN U2196 ( .B(n1853), .A(n1855), .Z(n1862) );
  NOR U2197 ( .A(n1857), .B(n1856), .Z(n1854) );
  XNOR U2198 ( .A(n1855), .B(n1854), .Z(n1860) );
  XOR U2199 ( .A(n1857), .B(n1856), .Z(n1858) );
  NAND U2200 ( .A(n1858), .B(n3223), .Z(n1859) );
  NAND U2201 ( .A(n1860), .B(n1859), .Z(n3228) );
  XNOR U2202 ( .A(a[141]), .B(b[141]), .Z(n3227) );
  NAND U2203 ( .A(n3228), .B(n3227), .Z(n1861) );
  NANDN U2204 ( .A(n1862), .B(n1861), .Z(n1868) );
  NAND U2205 ( .A(a[141]), .B(b[141]), .Z(n1869) );
  AND U2206 ( .A(n1868), .B(n1869), .Z(n1864) );
  XOR U2207 ( .A(a[142]), .B(b[142]), .Z(n3233) );
  ANDN U2208 ( .B(n3232), .A(n3233), .Z(n1863) );
  OR U2209 ( .A(n1864), .B(n1863), .Z(n1865) );
  AND U2210 ( .A(a[142]), .B(b[142]), .Z(n1867) );
  ANDN U2211 ( .B(n1865), .A(n1867), .Z(n1874) );
  NOR U2212 ( .A(n1869), .B(n1868), .Z(n1866) );
  XNOR U2213 ( .A(n1867), .B(n1866), .Z(n1872) );
  XOR U2214 ( .A(n1869), .B(n1868), .Z(n1870) );
  NAND U2215 ( .A(n1870), .B(n3233), .Z(n1871) );
  NAND U2216 ( .A(n1872), .B(n1871), .Z(n3238) );
  XNOR U2217 ( .A(a[143]), .B(b[143]), .Z(n3237) );
  NAND U2218 ( .A(n3238), .B(n3237), .Z(n1873) );
  NANDN U2219 ( .A(n1874), .B(n1873), .Z(n1880) );
  NAND U2220 ( .A(a[143]), .B(b[143]), .Z(n1881) );
  AND U2221 ( .A(n1880), .B(n1881), .Z(n1876) );
  XOR U2222 ( .A(a[144]), .B(b[144]), .Z(n3243) );
  ANDN U2223 ( .B(n3242), .A(n3243), .Z(n1875) );
  OR U2224 ( .A(n1876), .B(n1875), .Z(n1877) );
  AND U2225 ( .A(a[144]), .B(b[144]), .Z(n1879) );
  ANDN U2226 ( .B(n1877), .A(n1879), .Z(n1886) );
  NOR U2227 ( .A(n1881), .B(n1880), .Z(n1878) );
  XNOR U2228 ( .A(n1879), .B(n1878), .Z(n1884) );
  XOR U2229 ( .A(n1881), .B(n1880), .Z(n1882) );
  NAND U2230 ( .A(n1882), .B(n3243), .Z(n1883) );
  NAND U2231 ( .A(n1884), .B(n1883), .Z(n3248) );
  XNOR U2232 ( .A(a[145]), .B(b[145]), .Z(n3247) );
  NAND U2233 ( .A(n3248), .B(n3247), .Z(n1885) );
  NANDN U2234 ( .A(n1886), .B(n1885), .Z(n1892) );
  NAND U2235 ( .A(a[145]), .B(b[145]), .Z(n1893) );
  AND U2236 ( .A(n1892), .B(n1893), .Z(n1888) );
  XOR U2237 ( .A(a[146]), .B(b[146]), .Z(n3253) );
  ANDN U2238 ( .B(n3252), .A(n3253), .Z(n1887) );
  OR U2239 ( .A(n1888), .B(n1887), .Z(n1889) );
  AND U2240 ( .A(a[146]), .B(b[146]), .Z(n1891) );
  ANDN U2241 ( .B(n1889), .A(n1891), .Z(n1898) );
  NOR U2242 ( .A(n1893), .B(n1892), .Z(n1890) );
  XNOR U2243 ( .A(n1891), .B(n1890), .Z(n1896) );
  XOR U2244 ( .A(n1893), .B(n1892), .Z(n1894) );
  NAND U2245 ( .A(n1894), .B(n3253), .Z(n1895) );
  NAND U2246 ( .A(n1896), .B(n1895), .Z(n3258) );
  XNOR U2247 ( .A(a[147]), .B(b[147]), .Z(n3257) );
  NAND U2248 ( .A(n3258), .B(n3257), .Z(n1897) );
  NANDN U2249 ( .A(n1898), .B(n1897), .Z(n1904) );
  NAND U2250 ( .A(a[147]), .B(b[147]), .Z(n1905) );
  AND U2251 ( .A(n1904), .B(n1905), .Z(n1900) );
  XOR U2252 ( .A(a[148]), .B(b[148]), .Z(n3263) );
  ANDN U2253 ( .B(n3262), .A(n3263), .Z(n1899) );
  OR U2254 ( .A(n1900), .B(n1899), .Z(n1901) );
  AND U2255 ( .A(a[148]), .B(b[148]), .Z(n1903) );
  ANDN U2256 ( .B(n1901), .A(n1903), .Z(n1910) );
  NOR U2257 ( .A(n1905), .B(n1904), .Z(n1902) );
  XNOR U2258 ( .A(n1903), .B(n1902), .Z(n1908) );
  XOR U2259 ( .A(n1905), .B(n1904), .Z(n1906) );
  NAND U2260 ( .A(n1906), .B(n3263), .Z(n1907) );
  NAND U2261 ( .A(n1908), .B(n1907), .Z(n3268) );
  XNOR U2262 ( .A(a[149]), .B(b[149]), .Z(n3267) );
  NAND U2263 ( .A(n3268), .B(n3267), .Z(n1909) );
  NANDN U2264 ( .A(n1910), .B(n1909), .Z(n1916) );
  NAND U2265 ( .A(a[149]), .B(b[149]), .Z(n1917) );
  AND U2266 ( .A(n1916), .B(n1917), .Z(n1912) );
  XOR U2267 ( .A(a[150]), .B(b[150]), .Z(n3273) );
  ANDN U2268 ( .B(n3272), .A(n3273), .Z(n1911) );
  OR U2269 ( .A(n1912), .B(n1911), .Z(n1913) );
  AND U2270 ( .A(a[150]), .B(b[150]), .Z(n1915) );
  ANDN U2271 ( .B(n1913), .A(n1915), .Z(n1922) );
  NOR U2272 ( .A(n1917), .B(n1916), .Z(n1914) );
  XNOR U2273 ( .A(n1915), .B(n1914), .Z(n1920) );
  XOR U2274 ( .A(n1917), .B(n1916), .Z(n1918) );
  NAND U2275 ( .A(n1918), .B(n3273), .Z(n1919) );
  NAND U2276 ( .A(n1920), .B(n1919), .Z(n3278) );
  XNOR U2277 ( .A(a[151]), .B(b[151]), .Z(n3277) );
  NAND U2278 ( .A(n3278), .B(n3277), .Z(n1921) );
  NANDN U2279 ( .A(n1922), .B(n1921), .Z(n1923) );
  IV U2280 ( .A(n1923), .Z(n1927) );
  AND U2281 ( .A(a[151]), .B(b[151]), .Z(n1928) );
  NOR U2282 ( .A(n1927), .B(n1928), .Z(n1925) );
  XNOR U2283 ( .A(n1928), .B(n1923), .Z(n3283) );
  XNOR U2284 ( .A(a[152]), .B(b[152]), .Z(n3282) );
  AND U2285 ( .A(n3283), .B(n3282), .Z(n1924) );
  OR U2286 ( .A(n1925), .B(n1924), .Z(n1926) );
  AND U2287 ( .A(a[152]), .B(b[152]), .Z(n1930) );
  ANDN U2288 ( .B(n1926), .A(n1930), .Z(n1932) );
  AND U2289 ( .A(n1928), .B(n1927), .Z(n1929) );
  NAND U2290 ( .A(n1930), .B(n1929), .Z(n1935) );
  ANDN U2291 ( .B(n1935), .A(n1932), .Z(n3288) );
  XNOR U2292 ( .A(a[153]), .B(b[153]), .Z(n3287) );
  AND U2293 ( .A(n3288), .B(n3287), .Z(n1931) );
  OR U2294 ( .A(n1932), .B(n1931), .Z(n1933) );
  AND U2295 ( .A(n1934), .B(n1933), .Z(n1938) );
  OR U2296 ( .A(n1935), .B(n1934), .Z(n1936) );
  ANDN U2297 ( .B(n1936), .A(n1938), .Z(n3293) );
  XNOR U2298 ( .A(a[154]), .B(b[154]), .Z(n3292) );
  NAND U2299 ( .A(n3293), .B(n3292), .Z(n1937) );
  NANDN U2300 ( .A(n1938), .B(n1937), .Z(n1944) );
  NAND U2301 ( .A(a[154]), .B(b[154]), .Z(n1945) );
  AND U2302 ( .A(n1944), .B(n1945), .Z(n1940) );
  XOR U2303 ( .A(a[155]), .B(b[155]), .Z(n3298) );
  ANDN U2304 ( .B(n3297), .A(n3298), .Z(n1939) );
  OR U2305 ( .A(n1940), .B(n1939), .Z(n1941) );
  AND U2306 ( .A(a[155]), .B(b[155]), .Z(n1943) );
  ANDN U2307 ( .B(n1941), .A(n1943), .Z(n1950) );
  NOR U2308 ( .A(n1945), .B(n1944), .Z(n1942) );
  XNOR U2309 ( .A(n1943), .B(n1942), .Z(n1948) );
  XOR U2310 ( .A(n1945), .B(n1944), .Z(n1946) );
  NAND U2311 ( .A(n1946), .B(n3298), .Z(n1947) );
  NAND U2312 ( .A(n1948), .B(n1947), .Z(n3303) );
  XNOR U2313 ( .A(a[156]), .B(b[156]), .Z(n3302) );
  NAND U2314 ( .A(n3303), .B(n3302), .Z(n1949) );
  NANDN U2315 ( .A(n1950), .B(n1949), .Z(n1951) );
  IV U2316 ( .A(n1951), .Z(n1955) );
  AND U2317 ( .A(a[156]), .B(b[156]), .Z(n1956) );
  NOR U2318 ( .A(n1955), .B(n1956), .Z(n1953) );
  XNOR U2319 ( .A(n1956), .B(n1951), .Z(n3308) );
  XNOR U2320 ( .A(a[157]), .B(b[157]), .Z(n3307) );
  AND U2321 ( .A(n3308), .B(n3307), .Z(n1952) );
  OR U2322 ( .A(n1953), .B(n1952), .Z(n1954) );
  AND U2323 ( .A(a[157]), .B(b[157]), .Z(n1958) );
  ANDN U2324 ( .B(n1954), .A(n1958), .Z(n1960) );
  AND U2325 ( .A(n1956), .B(n1955), .Z(n1957) );
  NAND U2326 ( .A(n1958), .B(n1957), .Z(n1963) );
  ANDN U2327 ( .B(n1963), .A(n1960), .Z(n3313) );
  XNOR U2328 ( .A(a[158]), .B(b[158]), .Z(n3312) );
  AND U2329 ( .A(n3313), .B(n3312), .Z(n1959) );
  OR U2330 ( .A(n1960), .B(n1959), .Z(n1961) );
  AND U2331 ( .A(a[158]), .B(b[158]), .Z(n1962) );
  ANDN U2332 ( .B(n1961), .A(n1962), .Z(n1966) );
  NANDN U2333 ( .A(n1963), .B(n1962), .Z(n1964) );
  ANDN U2334 ( .B(n1964), .A(n1966), .Z(n3318) );
  XNOR U2335 ( .A(a[159]), .B(b[159]), .Z(n3317) );
  NAND U2336 ( .A(n3318), .B(n3317), .Z(n1965) );
  NANDN U2337 ( .A(n1966), .B(n1965), .Z(n1972) );
  NAND U2338 ( .A(a[159]), .B(b[159]), .Z(n1973) );
  AND U2339 ( .A(n1972), .B(n1973), .Z(n1968) );
  XOR U2340 ( .A(a[160]), .B(b[160]), .Z(n3323) );
  ANDN U2341 ( .B(n3322), .A(n3323), .Z(n1967) );
  OR U2342 ( .A(n1968), .B(n1967), .Z(n1969) );
  AND U2343 ( .A(a[160]), .B(b[160]), .Z(n1971) );
  ANDN U2344 ( .B(n1969), .A(n1971), .Z(n1978) );
  NOR U2345 ( .A(n1973), .B(n1972), .Z(n1970) );
  XNOR U2346 ( .A(n1971), .B(n1970), .Z(n1976) );
  XOR U2347 ( .A(n1973), .B(n1972), .Z(n1974) );
  NAND U2348 ( .A(n1974), .B(n3323), .Z(n1975) );
  NAND U2349 ( .A(n1976), .B(n1975), .Z(n3328) );
  XNOR U2350 ( .A(a[161]), .B(b[161]), .Z(n3327) );
  NAND U2351 ( .A(n3328), .B(n3327), .Z(n1977) );
  NANDN U2352 ( .A(n1978), .B(n1977), .Z(n1984) );
  NAND U2353 ( .A(a[161]), .B(b[161]), .Z(n1985) );
  AND U2354 ( .A(n1984), .B(n1985), .Z(n1980) );
  XOR U2355 ( .A(a[162]), .B(b[162]), .Z(n3333) );
  ANDN U2356 ( .B(n3332), .A(n3333), .Z(n1979) );
  OR U2357 ( .A(n1980), .B(n1979), .Z(n1981) );
  AND U2358 ( .A(a[162]), .B(b[162]), .Z(n1983) );
  ANDN U2359 ( .B(n1981), .A(n1983), .Z(n1990) );
  NOR U2360 ( .A(n1985), .B(n1984), .Z(n1982) );
  XNOR U2361 ( .A(n1983), .B(n1982), .Z(n1988) );
  XOR U2362 ( .A(n1985), .B(n1984), .Z(n1986) );
  NAND U2363 ( .A(n1986), .B(n3333), .Z(n1987) );
  NAND U2364 ( .A(n1988), .B(n1987), .Z(n3338) );
  XNOR U2365 ( .A(a[163]), .B(b[163]), .Z(n3337) );
  NAND U2366 ( .A(n3338), .B(n3337), .Z(n1989) );
  NANDN U2367 ( .A(n1990), .B(n1989), .Z(n1995) );
  ANDN U2368 ( .B(n1994), .A(n1995), .Z(n1991) );
  XOR U2369 ( .A(n1996), .B(n1991), .Z(n1993) );
  XOR U2370 ( .A(a[164]), .B(b[164]), .Z(n3343) );
  XNOR U2371 ( .A(n1994), .B(n1995), .Z(n3342) );
  NAND U2372 ( .A(n3343), .B(n3342), .Z(n1992) );
  NAND U2373 ( .A(n1993), .B(n1992), .Z(n3348) );
  XNOR U2374 ( .A(a[165]), .B(b[165]), .Z(n3347) );
  IV U2375 ( .A(n1997), .Z(n1999) );
  XNOR U2376 ( .A(n1998), .B(n1997), .Z(n3353) );
  XNOR U2377 ( .A(a[166]), .B(b[166]), .Z(n3352) );
  AND U2378 ( .A(a[166]), .B(b[166]), .Z(n2001) );
  NOR U2379 ( .A(n1999), .B(n1998), .Z(n2000) );
  NAND U2380 ( .A(n2001), .B(n2000), .Z(n2006) );
  ANDN U2381 ( .B(n2006), .A(n2003), .Z(n3358) );
  XNOR U2382 ( .A(a[167]), .B(b[167]), .Z(n3357) );
  NAND U2383 ( .A(n3358), .B(n3357), .Z(n2002) );
  NANDN U2384 ( .A(n2003), .B(n2002), .Z(n2004) );
  AND U2385 ( .A(n2005), .B(n2004), .Z(n2009) );
  OR U2386 ( .A(n2006), .B(n2005), .Z(n2007) );
  ANDN U2387 ( .B(n2007), .A(n2009), .Z(n3363) );
  XNOR U2388 ( .A(a[168]), .B(b[168]), .Z(n3362) );
  NAND U2389 ( .A(n3363), .B(n3362), .Z(n2008) );
  NANDN U2390 ( .A(n2009), .B(n2008), .Z(n2015) );
  NAND U2391 ( .A(a[168]), .B(b[168]), .Z(n2016) );
  AND U2392 ( .A(n2015), .B(n2016), .Z(n2011) );
  XOR U2393 ( .A(a[169]), .B(b[169]), .Z(n3368) );
  ANDN U2394 ( .B(n3367), .A(n3368), .Z(n2010) );
  OR U2395 ( .A(n2011), .B(n2010), .Z(n2012) );
  AND U2396 ( .A(a[169]), .B(b[169]), .Z(n2014) );
  ANDN U2397 ( .B(n2012), .A(n2014), .Z(n2021) );
  NOR U2398 ( .A(n2016), .B(n2015), .Z(n2013) );
  XNOR U2399 ( .A(n2014), .B(n2013), .Z(n2019) );
  XOR U2400 ( .A(n2016), .B(n2015), .Z(n2017) );
  NAND U2401 ( .A(n2017), .B(n3368), .Z(n2018) );
  NAND U2402 ( .A(n2019), .B(n2018), .Z(n3373) );
  XNOR U2403 ( .A(a[170]), .B(b[170]), .Z(n3372) );
  NAND U2404 ( .A(n3373), .B(n3372), .Z(n2020) );
  NANDN U2405 ( .A(n2021), .B(n2020), .Z(n2027) );
  NAND U2406 ( .A(a[170]), .B(b[170]), .Z(n2028) );
  AND U2407 ( .A(n2027), .B(n2028), .Z(n2023) );
  XOR U2408 ( .A(a[171]), .B(b[171]), .Z(n3378) );
  ANDN U2409 ( .B(n3377), .A(n3378), .Z(n2022) );
  OR U2410 ( .A(n2023), .B(n2022), .Z(n2024) );
  AND U2411 ( .A(a[171]), .B(b[171]), .Z(n2026) );
  ANDN U2412 ( .B(n2024), .A(n2026), .Z(n2033) );
  NOR U2413 ( .A(n2028), .B(n2027), .Z(n2025) );
  XNOR U2414 ( .A(n2026), .B(n2025), .Z(n2031) );
  XOR U2415 ( .A(n2028), .B(n2027), .Z(n2029) );
  NAND U2416 ( .A(n2029), .B(n3378), .Z(n2030) );
  NAND U2417 ( .A(n2031), .B(n2030), .Z(n3383) );
  XNOR U2418 ( .A(a[172]), .B(b[172]), .Z(n3382) );
  NAND U2419 ( .A(n3383), .B(n3382), .Z(n2032) );
  NANDN U2420 ( .A(n2033), .B(n2032), .Z(n2039) );
  NAND U2421 ( .A(a[172]), .B(b[172]), .Z(n2040) );
  AND U2422 ( .A(n2039), .B(n2040), .Z(n2035) );
  XOR U2423 ( .A(a[173]), .B(b[173]), .Z(n3388) );
  ANDN U2424 ( .B(n3387), .A(n3388), .Z(n2034) );
  OR U2425 ( .A(n2035), .B(n2034), .Z(n2036) );
  AND U2426 ( .A(a[173]), .B(b[173]), .Z(n2038) );
  ANDN U2427 ( .B(n2036), .A(n2038), .Z(n2045) );
  NOR U2428 ( .A(n2040), .B(n2039), .Z(n2037) );
  XNOR U2429 ( .A(n2038), .B(n2037), .Z(n2043) );
  XOR U2430 ( .A(n2040), .B(n2039), .Z(n2041) );
  NAND U2431 ( .A(n2041), .B(n3388), .Z(n2042) );
  NAND U2432 ( .A(n2043), .B(n2042), .Z(n3393) );
  XNOR U2433 ( .A(a[174]), .B(b[174]), .Z(n3392) );
  NAND U2434 ( .A(n3393), .B(n3392), .Z(n2044) );
  NANDN U2435 ( .A(n2045), .B(n2044), .Z(n2051) );
  NAND U2436 ( .A(a[174]), .B(b[174]), .Z(n2052) );
  AND U2437 ( .A(n2051), .B(n2052), .Z(n2047) );
  XOR U2438 ( .A(a[175]), .B(b[175]), .Z(n3398) );
  ANDN U2439 ( .B(n3397), .A(n3398), .Z(n2046) );
  OR U2440 ( .A(n2047), .B(n2046), .Z(n2048) );
  AND U2441 ( .A(a[175]), .B(b[175]), .Z(n2050) );
  ANDN U2442 ( .B(n2048), .A(n2050), .Z(n2057) );
  NOR U2443 ( .A(n2052), .B(n2051), .Z(n2049) );
  XNOR U2444 ( .A(n2050), .B(n2049), .Z(n2055) );
  XOR U2445 ( .A(n2052), .B(n2051), .Z(n2053) );
  NAND U2446 ( .A(n2053), .B(n3398), .Z(n2054) );
  NAND U2447 ( .A(n2055), .B(n2054), .Z(n3403) );
  XNOR U2448 ( .A(a[176]), .B(b[176]), .Z(n3402) );
  NAND U2449 ( .A(n3403), .B(n3402), .Z(n2056) );
  NANDN U2450 ( .A(n2057), .B(n2056), .Z(n2063) );
  NAND U2451 ( .A(a[176]), .B(b[176]), .Z(n2064) );
  AND U2452 ( .A(n2063), .B(n2064), .Z(n2059) );
  XOR U2453 ( .A(a[177]), .B(b[177]), .Z(n3408) );
  ANDN U2454 ( .B(n3407), .A(n3408), .Z(n2058) );
  OR U2455 ( .A(n2059), .B(n2058), .Z(n2060) );
  AND U2456 ( .A(a[177]), .B(b[177]), .Z(n2062) );
  ANDN U2457 ( .B(n2060), .A(n2062), .Z(n2069) );
  NOR U2458 ( .A(n2064), .B(n2063), .Z(n2061) );
  XNOR U2459 ( .A(n2062), .B(n2061), .Z(n2067) );
  XOR U2460 ( .A(n2064), .B(n2063), .Z(n2065) );
  NAND U2461 ( .A(n2065), .B(n3408), .Z(n2066) );
  NAND U2462 ( .A(n2067), .B(n2066), .Z(n3413) );
  XNOR U2463 ( .A(a[178]), .B(b[178]), .Z(n3412) );
  NAND U2464 ( .A(n3413), .B(n3412), .Z(n2068) );
  NANDN U2465 ( .A(n2069), .B(n2068), .Z(n2075) );
  NAND U2466 ( .A(a[178]), .B(b[178]), .Z(n2076) );
  AND U2467 ( .A(n2075), .B(n2076), .Z(n2071) );
  XOR U2468 ( .A(a[179]), .B(b[179]), .Z(n3418) );
  ANDN U2469 ( .B(n3417), .A(n3418), .Z(n2070) );
  OR U2470 ( .A(n2071), .B(n2070), .Z(n2072) );
  AND U2471 ( .A(a[179]), .B(b[179]), .Z(n2074) );
  ANDN U2472 ( .B(n2072), .A(n2074), .Z(n2081) );
  NOR U2473 ( .A(n2076), .B(n2075), .Z(n2073) );
  XNOR U2474 ( .A(n2074), .B(n2073), .Z(n2079) );
  XOR U2475 ( .A(n2076), .B(n2075), .Z(n2077) );
  NAND U2476 ( .A(n2077), .B(n3418), .Z(n2078) );
  NAND U2477 ( .A(n2079), .B(n2078), .Z(n3423) );
  XNOR U2478 ( .A(a[180]), .B(b[180]), .Z(n3422) );
  NAND U2479 ( .A(n3423), .B(n3422), .Z(n2080) );
  NANDN U2480 ( .A(n2081), .B(n2080), .Z(n2087) );
  NAND U2481 ( .A(a[180]), .B(b[180]), .Z(n2088) );
  AND U2482 ( .A(n2087), .B(n2088), .Z(n2083) );
  XOR U2483 ( .A(a[181]), .B(b[181]), .Z(n3428) );
  ANDN U2484 ( .B(n3427), .A(n3428), .Z(n2082) );
  OR U2485 ( .A(n2083), .B(n2082), .Z(n2084) );
  AND U2486 ( .A(a[181]), .B(b[181]), .Z(n2086) );
  ANDN U2487 ( .B(n2084), .A(n2086), .Z(n2093) );
  NOR U2488 ( .A(n2088), .B(n2087), .Z(n2085) );
  XNOR U2489 ( .A(n2086), .B(n2085), .Z(n2091) );
  XOR U2490 ( .A(n2088), .B(n2087), .Z(n2089) );
  NAND U2491 ( .A(n2089), .B(n3428), .Z(n2090) );
  NAND U2492 ( .A(n2091), .B(n2090), .Z(n3433) );
  XNOR U2493 ( .A(a[182]), .B(b[182]), .Z(n3432) );
  NAND U2494 ( .A(n3433), .B(n3432), .Z(n2092) );
  NANDN U2495 ( .A(n2093), .B(n2092), .Z(n2099) );
  NAND U2496 ( .A(a[182]), .B(b[182]), .Z(n2100) );
  AND U2497 ( .A(n2099), .B(n2100), .Z(n2095) );
  XOR U2498 ( .A(a[183]), .B(b[183]), .Z(n3438) );
  ANDN U2499 ( .B(n3437), .A(n3438), .Z(n2094) );
  OR U2500 ( .A(n2095), .B(n2094), .Z(n2096) );
  AND U2501 ( .A(a[183]), .B(b[183]), .Z(n2098) );
  ANDN U2502 ( .B(n2096), .A(n2098), .Z(n2105) );
  NOR U2503 ( .A(n2100), .B(n2099), .Z(n2097) );
  XNOR U2504 ( .A(n2098), .B(n2097), .Z(n2103) );
  XOR U2505 ( .A(n2100), .B(n2099), .Z(n2101) );
  NAND U2506 ( .A(n2101), .B(n3438), .Z(n2102) );
  NAND U2507 ( .A(n2103), .B(n2102), .Z(n3443) );
  XNOR U2508 ( .A(a[184]), .B(b[184]), .Z(n3442) );
  NAND U2509 ( .A(n3443), .B(n3442), .Z(n2104) );
  NANDN U2510 ( .A(n2105), .B(n2104), .Z(n2106) );
  IV U2511 ( .A(n2106), .Z(n2110) );
  AND U2512 ( .A(a[184]), .B(b[184]), .Z(n2111) );
  NOR U2513 ( .A(n2110), .B(n2111), .Z(n2108) );
  XNOR U2514 ( .A(n2111), .B(n2106), .Z(n3448) );
  XNOR U2515 ( .A(a[185]), .B(b[185]), .Z(n3447) );
  AND U2516 ( .A(n3448), .B(n3447), .Z(n2107) );
  OR U2517 ( .A(n2108), .B(n2107), .Z(n2109) );
  AND U2518 ( .A(a[185]), .B(b[185]), .Z(n2113) );
  ANDN U2519 ( .B(n2109), .A(n2113), .Z(n2115) );
  AND U2520 ( .A(n2111), .B(n2110), .Z(n2112) );
  NAND U2521 ( .A(n2113), .B(n2112), .Z(n2118) );
  ANDN U2522 ( .B(n2118), .A(n2115), .Z(n3453) );
  XNOR U2523 ( .A(a[186]), .B(b[186]), .Z(n3452) );
  AND U2524 ( .A(n3453), .B(n3452), .Z(n2114) );
  OR U2525 ( .A(n2115), .B(n2114), .Z(n2116) );
  AND U2526 ( .A(n2117), .B(n2116), .Z(n2120) );
  XNOR U2527 ( .A(a[187]), .B(b[187]), .Z(n3457) );
  NAND U2528 ( .A(n3458), .B(n3457), .Z(n2119) );
  NANDN U2529 ( .A(n2120), .B(n2119), .Z(n2126) );
  NAND U2530 ( .A(a[187]), .B(b[187]), .Z(n2127) );
  AND U2531 ( .A(n2126), .B(n2127), .Z(n2122) );
  XOR U2532 ( .A(a[188]), .B(b[188]), .Z(n3463) );
  ANDN U2533 ( .B(n3462), .A(n3463), .Z(n2121) );
  OR U2534 ( .A(n2122), .B(n2121), .Z(n2123) );
  AND U2535 ( .A(a[188]), .B(b[188]), .Z(n2125) );
  ANDN U2536 ( .B(n2123), .A(n2125), .Z(n2132) );
  NOR U2537 ( .A(n2127), .B(n2126), .Z(n2124) );
  XNOR U2538 ( .A(n2125), .B(n2124), .Z(n2130) );
  XOR U2539 ( .A(n2127), .B(n2126), .Z(n2128) );
  NAND U2540 ( .A(n2128), .B(n3463), .Z(n2129) );
  NAND U2541 ( .A(n2130), .B(n2129), .Z(n3468) );
  XNOR U2542 ( .A(a[189]), .B(b[189]), .Z(n3467) );
  NAND U2543 ( .A(n3468), .B(n3467), .Z(n2131) );
  NANDN U2544 ( .A(n2132), .B(n2131), .Z(n2133) );
  IV U2545 ( .A(n2133), .Z(n2137) );
  AND U2546 ( .A(a[189]), .B(b[189]), .Z(n2138) );
  NOR U2547 ( .A(n2137), .B(n2138), .Z(n2135) );
  XNOR U2548 ( .A(n2138), .B(n2133), .Z(n3473) );
  XNOR U2549 ( .A(a[190]), .B(b[190]), .Z(n3472) );
  AND U2550 ( .A(n3473), .B(n3472), .Z(n2134) );
  OR U2551 ( .A(n2135), .B(n2134), .Z(n2136) );
  AND U2552 ( .A(a[190]), .B(b[190]), .Z(n2140) );
  ANDN U2553 ( .B(n2136), .A(n2140), .Z(n2142) );
  AND U2554 ( .A(n2138), .B(n2137), .Z(n2139) );
  NAND U2555 ( .A(n2140), .B(n2139), .Z(n2145) );
  ANDN U2556 ( .B(n2145), .A(n2142), .Z(n3478) );
  XNOR U2557 ( .A(a[191]), .B(b[191]), .Z(n3477) );
  AND U2558 ( .A(n3478), .B(n3477), .Z(n2141) );
  OR U2559 ( .A(n2142), .B(n2141), .Z(n2143) );
  AND U2560 ( .A(a[191]), .B(b[191]), .Z(n2144) );
  ANDN U2561 ( .B(n2143), .A(n2144), .Z(n2148) );
  NANDN U2562 ( .A(n2145), .B(n2144), .Z(n2146) );
  ANDN U2563 ( .B(n2146), .A(n2148), .Z(n3483) );
  XNOR U2564 ( .A(a[192]), .B(b[192]), .Z(n3482) );
  NAND U2565 ( .A(n3483), .B(n3482), .Z(n2147) );
  NANDN U2566 ( .A(n2148), .B(n2147), .Z(n2154) );
  NAND U2567 ( .A(a[192]), .B(b[192]), .Z(n2155) );
  AND U2568 ( .A(n2154), .B(n2155), .Z(n2150) );
  XOR U2569 ( .A(a[193]), .B(b[193]), .Z(n3488) );
  ANDN U2570 ( .B(n3487), .A(n3488), .Z(n2149) );
  OR U2571 ( .A(n2150), .B(n2149), .Z(n2151) );
  AND U2572 ( .A(a[193]), .B(b[193]), .Z(n2153) );
  ANDN U2573 ( .B(n2151), .A(n2153), .Z(n2160) );
  NOR U2574 ( .A(n2155), .B(n2154), .Z(n2152) );
  XNOR U2575 ( .A(n2153), .B(n2152), .Z(n2158) );
  XOR U2576 ( .A(n2155), .B(n2154), .Z(n2156) );
  NAND U2577 ( .A(n2156), .B(n3488), .Z(n2157) );
  NAND U2578 ( .A(n2158), .B(n2157), .Z(n3493) );
  XNOR U2579 ( .A(a[194]), .B(b[194]), .Z(n3492) );
  NAND U2580 ( .A(n3493), .B(n3492), .Z(n2159) );
  NANDN U2581 ( .A(n2160), .B(n2159), .Z(n2166) );
  NAND U2582 ( .A(a[194]), .B(b[194]), .Z(n2167) );
  AND U2583 ( .A(n2166), .B(n2167), .Z(n2162) );
  XOR U2584 ( .A(a[195]), .B(b[195]), .Z(n3498) );
  ANDN U2585 ( .B(n3497), .A(n3498), .Z(n2161) );
  OR U2586 ( .A(n2162), .B(n2161), .Z(n2163) );
  AND U2587 ( .A(a[195]), .B(b[195]), .Z(n2165) );
  ANDN U2588 ( .B(n2163), .A(n2165), .Z(n2172) );
  NOR U2589 ( .A(n2167), .B(n2166), .Z(n2164) );
  XNOR U2590 ( .A(n2165), .B(n2164), .Z(n2170) );
  XOR U2591 ( .A(n2167), .B(n2166), .Z(n2168) );
  NAND U2592 ( .A(n2168), .B(n3498), .Z(n2169) );
  NAND U2593 ( .A(n2170), .B(n2169), .Z(n3503) );
  XNOR U2594 ( .A(a[196]), .B(b[196]), .Z(n3502) );
  NAND U2595 ( .A(n3503), .B(n3502), .Z(n2171) );
  NANDN U2596 ( .A(n2172), .B(n2171), .Z(n2178) );
  NAND U2597 ( .A(a[196]), .B(b[196]), .Z(n2179) );
  AND U2598 ( .A(n2178), .B(n2179), .Z(n2174) );
  XOR U2599 ( .A(a[197]), .B(b[197]), .Z(n3508) );
  ANDN U2600 ( .B(n3507), .A(n3508), .Z(n2173) );
  OR U2601 ( .A(n2174), .B(n2173), .Z(n2175) );
  AND U2602 ( .A(a[197]), .B(b[197]), .Z(n2177) );
  ANDN U2603 ( .B(n2175), .A(n2177), .Z(n2184) );
  NOR U2604 ( .A(n2179), .B(n2178), .Z(n2176) );
  XNOR U2605 ( .A(n2177), .B(n2176), .Z(n2182) );
  XOR U2606 ( .A(n2179), .B(n2178), .Z(n2180) );
  NAND U2607 ( .A(n2180), .B(n3508), .Z(n2181) );
  NAND U2608 ( .A(n2182), .B(n2181), .Z(n3513) );
  XNOR U2609 ( .A(a[198]), .B(b[198]), .Z(n3512) );
  NAND U2610 ( .A(n3513), .B(n3512), .Z(n2183) );
  NANDN U2611 ( .A(n2184), .B(n2183), .Z(n2190) );
  NAND U2612 ( .A(a[198]), .B(b[198]), .Z(n2191) );
  AND U2613 ( .A(n2190), .B(n2191), .Z(n2186) );
  XOR U2614 ( .A(a[199]), .B(b[199]), .Z(n3518) );
  ANDN U2615 ( .B(n3517), .A(n3518), .Z(n2185) );
  OR U2616 ( .A(n2186), .B(n2185), .Z(n2187) );
  AND U2617 ( .A(a[199]), .B(b[199]), .Z(n2189) );
  ANDN U2618 ( .B(n2187), .A(n2189), .Z(n2196) );
  NOR U2619 ( .A(n2191), .B(n2190), .Z(n2188) );
  XNOR U2620 ( .A(n2189), .B(n2188), .Z(n2194) );
  XOR U2621 ( .A(n2191), .B(n2190), .Z(n2192) );
  NAND U2622 ( .A(n2192), .B(n3518), .Z(n2193) );
  NAND U2623 ( .A(n2194), .B(n2193), .Z(n3523) );
  XNOR U2624 ( .A(a[200]), .B(b[200]), .Z(n3522) );
  NAND U2625 ( .A(n3523), .B(n3522), .Z(n2195) );
  NANDN U2626 ( .A(n2196), .B(n2195), .Z(n2197) );
  IV U2627 ( .A(n2197), .Z(n2201) );
  AND U2628 ( .A(a[200]), .B(b[200]), .Z(n2202) );
  NOR U2629 ( .A(n2201), .B(n2202), .Z(n2199) );
  XNOR U2630 ( .A(n2202), .B(n2197), .Z(n3528) );
  XNOR U2631 ( .A(a[201]), .B(b[201]), .Z(n3527) );
  AND U2632 ( .A(n3528), .B(n3527), .Z(n2198) );
  OR U2633 ( .A(n2199), .B(n2198), .Z(n2200) );
  AND U2634 ( .A(a[201]), .B(b[201]), .Z(n2204) );
  ANDN U2635 ( .B(n2200), .A(n2204), .Z(n2206) );
  AND U2636 ( .A(n2202), .B(n2201), .Z(n2203) );
  NAND U2637 ( .A(n2204), .B(n2203), .Z(n2209) );
  ANDN U2638 ( .B(n2209), .A(n2206), .Z(n3533) );
  XNOR U2639 ( .A(a[202]), .B(b[202]), .Z(n3532) );
  AND U2640 ( .A(n3533), .B(n3532), .Z(n2205) );
  OR U2641 ( .A(n2206), .B(n2205), .Z(n2207) );
  AND U2642 ( .A(a[202]), .B(b[202]), .Z(n2208) );
  ANDN U2643 ( .B(n2207), .A(n2208), .Z(n2212) );
  NANDN U2644 ( .A(n2209), .B(n2208), .Z(n2210) );
  ANDN U2645 ( .B(n2210), .A(n2212), .Z(n3538) );
  XNOR U2646 ( .A(a[203]), .B(b[203]), .Z(n3537) );
  NAND U2647 ( .A(n3538), .B(n3537), .Z(n2211) );
  NANDN U2648 ( .A(n2212), .B(n2211), .Z(n2218) );
  NAND U2649 ( .A(a[203]), .B(b[203]), .Z(n2219) );
  AND U2650 ( .A(n2218), .B(n2219), .Z(n2214) );
  XOR U2651 ( .A(a[204]), .B(b[204]), .Z(n3543) );
  ANDN U2652 ( .B(n3542), .A(n3543), .Z(n2213) );
  OR U2653 ( .A(n2214), .B(n2213), .Z(n2215) );
  AND U2654 ( .A(a[204]), .B(b[204]), .Z(n2217) );
  ANDN U2655 ( .B(n2215), .A(n2217), .Z(n2224) );
  NOR U2656 ( .A(n2219), .B(n2218), .Z(n2216) );
  XNOR U2657 ( .A(n2217), .B(n2216), .Z(n2222) );
  XOR U2658 ( .A(n2219), .B(n2218), .Z(n2220) );
  NAND U2659 ( .A(n2220), .B(n3543), .Z(n2221) );
  NAND U2660 ( .A(n2222), .B(n2221), .Z(n3548) );
  XNOR U2661 ( .A(a[205]), .B(b[205]), .Z(n3547) );
  NAND U2662 ( .A(n3548), .B(n3547), .Z(n2223) );
  NANDN U2663 ( .A(n2224), .B(n2223), .Z(n2230) );
  NAND U2664 ( .A(a[205]), .B(b[205]), .Z(n2231) );
  AND U2665 ( .A(n2230), .B(n2231), .Z(n2226) );
  XOR U2666 ( .A(a[206]), .B(b[206]), .Z(n3553) );
  ANDN U2667 ( .B(n3552), .A(n3553), .Z(n2225) );
  OR U2668 ( .A(n2226), .B(n2225), .Z(n2227) );
  AND U2669 ( .A(a[206]), .B(b[206]), .Z(n2229) );
  ANDN U2670 ( .B(n2227), .A(n2229), .Z(n2236) );
  NOR U2671 ( .A(n2231), .B(n2230), .Z(n2228) );
  XNOR U2672 ( .A(n2229), .B(n2228), .Z(n2234) );
  XOR U2673 ( .A(n2231), .B(n2230), .Z(n2232) );
  NAND U2674 ( .A(n2232), .B(n3553), .Z(n2233) );
  NAND U2675 ( .A(n2234), .B(n2233), .Z(n3558) );
  XNOR U2676 ( .A(a[207]), .B(b[207]), .Z(n3557) );
  NAND U2677 ( .A(n3558), .B(n3557), .Z(n2235) );
  NANDN U2678 ( .A(n2236), .B(n2235), .Z(n2242) );
  NAND U2679 ( .A(a[207]), .B(b[207]), .Z(n2243) );
  AND U2680 ( .A(n2242), .B(n2243), .Z(n2238) );
  XOR U2681 ( .A(a[208]), .B(b[208]), .Z(n3563) );
  ANDN U2682 ( .B(n3562), .A(n3563), .Z(n2237) );
  OR U2683 ( .A(n2238), .B(n2237), .Z(n2239) );
  AND U2684 ( .A(a[208]), .B(b[208]), .Z(n2241) );
  ANDN U2685 ( .B(n2239), .A(n2241), .Z(n2248) );
  NOR U2686 ( .A(n2243), .B(n2242), .Z(n2240) );
  XNOR U2687 ( .A(n2241), .B(n2240), .Z(n2246) );
  XOR U2688 ( .A(n2243), .B(n2242), .Z(n2244) );
  NAND U2689 ( .A(n2244), .B(n3563), .Z(n2245) );
  NAND U2690 ( .A(n2246), .B(n2245), .Z(n3568) );
  XNOR U2691 ( .A(a[209]), .B(b[209]), .Z(n3567) );
  NAND U2692 ( .A(n3568), .B(n3567), .Z(n2247) );
  NANDN U2693 ( .A(n2248), .B(n2247), .Z(n2254) );
  NAND U2694 ( .A(a[209]), .B(b[209]), .Z(n2255) );
  AND U2695 ( .A(n2254), .B(n2255), .Z(n2250) );
  XOR U2696 ( .A(a[210]), .B(b[210]), .Z(n3573) );
  ANDN U2697 ( .B(n3572), .A(n3573), .Z(n2249) );
  OR U2698 ( .A(n2250), .B(n2249), .Z(n2251) );
  AND U2699 ( .A(a[210]), .B(b[210]), .Z(n2253) );
  ANDN U2700 ( .B(n2251), .A(n2253), .Z(n2260) );
  NOR U2701 ( .A(n2255), .B(n2254), .Z(n2252) );
  XNOR U2702 ( .A(n2253), .B(n2252), .Z(n2258) );
  XOR U2703 ( .A(n2255), .B(n2254), .Z(n2256) );
  NAND U2704 ( .A(n2256), .B(n3573), .Z(n2257) );
  NAND U2705 ( .A(n2258), .B(n2257), .Z(n3578) );
  XNOR U2706 ( .A(a[211]), .B(b[211]), .Z(n3577) );
  NAND U2707 ( .A(n3578), .B(n3577), .Z(n2259) );
  NANDN U2708 ( .A(n2260), .B(n2259), .Z(n2266) );
  NAND U2709 ( .A(a[211]), .B(b[211]), .Z(n2267) );
  AND U2710 ( .A(n2266), .B(n2267), .Z(n2262) );
  XOR U2711 ( .A(a[212]), .B(b[212]), .Z(n3583) );
  ANDN U2712 ( .B(n3582), .A(n3583), .Z(n2261) );
  OR U2713 ( .A(n2262), .B(n2261), .Z(n2263) );
  AND U2714 ( .A(a[212]), .B(b[212]), .Z(n2265) );
  ANDN U2715 ( .B(n2263), .A(n2265), .Z(n2272) );
  NOR U2716 ( .A(n2267), .B(n2266), .Z(n2264) );
  XNOR U2717 ( .A(n2265), .B(n2264), .Z(n2270) );
  XOR U2718 ( .A(n2267), .B(n2266), .Z(n2268) );
  NAND U2719 ( .A(n2268), .B(n3583), .Z(n2269) );
  NAND U2720 ( .A(n2270), .B(n2269), .Z(n3588) );
  XNOR U2721 ( .A(a[213]), .B(b[213]), .Z(n3587) );
  NAND U2722 ( .A(n3588), .B(n3587), .Z(n2271) );
  NANDN U2723 ( .A(n2272), .B(n2271), .Z(n2278) );
  NAND U2724 ( .A(a[213]), .B(b[213]), .Z(n2279) );
  AND U2725 ( .A(n2278), .B(n2279), .Z(n2274) );
  XOR U2726 ( .A(a[214]), .B(b[214]), .Z(n3593) );
  ANDN U2727 ( .B(n3592), .A(n3593), .Z(n2273) );
  OR U2728 ( .A(n2274), .B(n2273), .Z(n2275) );
  AND U2729 ( .A(a[214]), .B(b[214]), .Z(n2277) );
  ANDN U2730 ( .B(n2275), .A(n2277), .Z(n2284) );
  NOR U2731 ( .A(n2279), .B(n2278), .Z(n2276) );
  XNOR U2732 ( .A(n2277), .B(n2276), .Z(n2282) );
  XOR U2733 ( .A(n2279), .B(n2278), .Z(n2280) );
  NAND U2734 ( .A(n2280), .B(n3593), .Z(n2281) );
  NAND U2735 ( .A(n2282), .B(n2281), .Z(n3598) );
  XNOR U2736 ( .A(a[215]), .B(b[215]), .Z(n3597) );
  NAND U2737 ( .A(n3598), .B(n3597), .Z(n2283) );
  NANDN U2738 ( .A(n2284), .B(n2283), .Z(n2290) );
  NAND U2739 ( .A(a[215]), .B(b[215]), .Z(n2291) );
  AND U2740 ( .A(n2290), .B(n2291), .Z(n2286) );
  XOR U2741 ( .A(a[216]), .B(b[216]), .Z(n3603) );
  ANDN U2742 ( .B(n3602), .A(n3603), .Z(n2285) );
  OR U2743 ( .A(n2286), .B(n2285), .Z(n2287) );
  AND U2744 ( .A(a[216]), .B(b[216]), .Z(n2289) );
  ANDN U2745 ( .B(n2287), .A(n2289), .Z(n2296) );
  NOR U2746 ( .A(n2291), .B(n2290), .Z(n2288) );
  XNOR U2747 ( .A(n2289), .B(n2288), .Z(n2294) );
  XOR U2748 ( .A(n2291), .B(n2290), .Z(n2292) );
  NAND U2749 ( .A(n2292), .B(n3603), .Z(n2293) );
  NAND U2750 ( .A(n2294), .B(n2293), .Z(n3608) );
  XNOR U2751 ( .A(a[217]), .B(b[217]), .Z(n3607) );
  NAND U2752 ( .A(n3608), .B(n3607), .Z(n2295) );
  NANDN U2753 ( .A(n2296), .B(n2295), .Z(n2297) );
  IV U2754 ( .A(n2297), .Z(n2301) );
  AND U2755 ( .A(a[217]), .B(b[217]), .Z(n2302) );
  NOR U2756 ( .A(n2301), .B(n2302), .Z(n2299) );
  XNOR U2757 ( .A(n2302), .B(n2297), .Z(n3613) );
  XNOR U2758 ( .A(a[218]), .B(b[218]), .Z(n3612) );
  AND U2759 ( .A(n3613), .B(n3612), .Z(n2298) );
  OR U2760 ( .A(n2299), .B(n2298), .Z(n2300) );
  AND U2761 ( .A(a[218]), .B(b[218]), .Z(n2304) );
  ANDN U2762 ( .B(n2300), .A(n2304), .Z(n2306) );
  AND U2763 ( .A(n2302), .B(n2301), .Z(n2303) );
  NAND U2764 ( .A(n2304), .B(n2303), .Z(n2309) );
  ANDN U2765 ( .B(n2309), .A(n2306), .Z(n3618) );
  XNOR U2766 ( .A(a[219]), .B(b[219]), .Z(n3617) );
  AND U2767 ( .A(n3618), .B(n3617), .Z(n2305) );
  OR U2768 ( .A(n2306), .B(n2305), .Z(n2307) );
  AND U2769 ( .A(a[219]), .B(b[219]), .Z(n2308) );
  ANDN U2770 ( .B(n2307), .A(n2308), .Z(n2312) );
  NANDN U2771 ( .A(n2309), .B(n2308), .Z(n2310) );
  ANDN U2772 ( .B(n2310), .A(n2312), .Z(n3623) );
  XNOR U2773 ( .A(a[220]), .B(b[220]), .Z(n3622) );
  NAND U2774 ( .A(n3623), .B(n3622), .Z(n2311) );
  NANDN U2775 ( .A(n2312), .B(n2311), .Z(n2318) );
  NAND U2776 ( .A(a[220]), .B(b[220]), .Z(n2319) );
  AND U2777 ( .A(n2318), .B(n2319), .Z(n2314) );
  XOR U2778 ( .A(a[221]), .B(b[221]), .Z(n3628) );
  ANDN U2779 ( .B(n3627), .A(n3628), .Z(n2313) );
  OR U2780 ( .A(n2314), .B(n2313), .Z(n2315) );
  AND U2781 ( .A(a[221]), .B(b[221]), .Z(n2317) );
  ANDN U2782 ( .B(n2315), .A(n2317), .Z(n2324) );
  NOR U2783 ( .A(n2319), .B(n2318), .Z(n2316) );
  XNOR U2784 ( .A(n2317), .B(n2316), .Z(n2322) );
  XOR U2785 ( .A(n2319), .B(n2318), .Z(n2320) );
  NAND U2786 ( .A(n2320), .B(n3628), .Z(n2321) );
  NAND U2787 ( .A(n2322), .B(n2321), .Z(n3633) );
  XNOR U2788 ( .A(a[222]), .B(b[222]), .Z(n3632) );
  NAND U2789 ( .A(n3633), .B(n3632), .Z(n2323) );
  NANDN U2790 ( .A(n2324), .B(n2323), .Z(n2330) );
  NAND U2791 ( .A(a[222]), .B(b[222]), .Z(n2331) );
  AND U2792 ( .A(n2330), .B(n2331), .Z(n2326) );
  XOR U2793 ( .A(a[223]), .B(b[223]), .Z(n3638) );
  ANDN U2794 ( .B(n3637), .A(n3638), .Z(n2325) );
  OR U2795 ( .A(n2326), .B(n2325), .Z(n2327) );
  AND U2796 ( .A(a[223]), .B(b[223]), .Z(n2329) );
  ANDN U2797 ( .B(n2327), .A(n2329), .Z(n2336) );
  NOR U2798 ( .A(n2331), .B(n2330), .Z(n2328) );
  XNOR U2799 ( .A(n2329), .B(n2328), .Z(n2334) );
  XOR U2800 ( .A(n2331), .B(n2330), .Z(n2332) );
  NAND U2801 ( .A(n2332), .B(n3638), .Z(n2333) );
  NAND U2802 ( .A(n2334), .B(n2333), .Z(n3643) );
  XNOR U2803 ( .A(a[224]), .B(b[224]), .Z(n3642) );
  NAND U2804 ( .A(n3643), .B(n3642), .Z(n2335) );
  NANDN U2805 ( .A(n2336), .B(n2335), .Z(n2342) );
  NAND U2806 ( .A(a[224]), .B(b[224]), .Z(n2343) );
  AND U2807 ( .A(n2342), .B(n2343), .Z(n2338) );
  XOR U2808 ( .A(a[225]), .B(b[225]), .Z(n3648) );
  ANDN U2809 ( .B(n3647), .A(n3648), .Z(n2337) );
  OR U2810 ( .A(n2338), .B(n2337), .Z(n2339) );
  AND U2811 ( .A(a[225]), .B(b[225]), .Z(n2341) );
  ANDN U2812 ( .B(n2339), .A(n2341), .Z(n2348) );
  NOR U2813 ( .A(n2343), .B(n2342), .Z(n2340) );
  XNOR U2814 ( .A(n2341), .B(n2340), .Z(n2346) );
  XOR U2815 ( .A(n2343), .B(n2342), .Z(n2344) );
  NAND U2816 ( .A(n2344), .B(n3648), .Z(n2345) );
  NAND U2817 ( .A(n2346), .B(n2345), .Z(n3653) );
  XNOR U2818 ( .A(a[226]), .B(b[226]), .Z(n3652) );
  NAND U2819 ( .A(n3653), .B(n3652), .Z(n2347) );
  NANDN U2820 ( .A(n2348), .B(n2347), .Z(n2354) );
  NAND U2821 ( .A(a[226]), .B(b[226]), .Z(n2355) );
  AND U2822 ( .A(n2354), .B(n2355), .Z(n2350) );
  XOR U2823 ( .A(a[227]), .B(b[227]), .Z(n3658) );
  ANDN U2824 ( .B(n3657), .A(n3658), .Z(n2349) );
  OR U2825 ( .A(n2350), .B(n2349), .Z(n2351) );
  AND U2826 ( .A(a[227]), .B(b[227]), .Z(n2353) );
  ANDN U2827 ( .B(n2351), .A(n2353), .Z(n2360) );
  NOR U2828 ( .A(n2355), .B(n2354), .Z(n2352) );
  XNOR U2829 ( .A(n2353), .B(n2352), .Z(n2358) );
  XOR U2830 ( .A(n2355), .B(n2354), .Z(n2356) );
  NAND U2831 ( .A(n2356), .B(n3658), .Z(n2357) );
  NAND U2832 ( .A(n2358), .B(n2357), .Z(n3663) );
  XNOR U2833 ( .A(a[228]), .B(b[228]), .Z(n3662) );
  NAND U2834 ( .A(n3663), .B(n3662), .Z(n2359) );
  NANDN U2835 ( .A(n2360), .B(n2359), .Z(n2366) );
  NAND U2836 ( .A(a[228]), .B(b[228]), .Z(n2367) );
  AND U2837 ( .A(n2366), .B(n2367), .Z(n2362) );
  XOR U2838 ( .A(a[229]), .B(b[229]), .Z(n3668) );
  ANDN U2839 ( .B(n3667), .A(n3668), .Z(n2361) );
  OR U2840 ( .A(n2362), .B(n2361), .Z(n2363) );
  AND U2841 ( .A(a[229]), .B(b[229]), .Z(n2365) );
  ANDN U2842 ( .B(n2363), .A(n2365), .Z(n2372) );
  NOR U2843 ( .A(n2367), .B(n2366), .Z(n2364) );
  XNOR U2844 ( .A(n2365), .B(n2364), .Z(n2370) );
  XOR U2845 ( .A(n2367), .B(n2366), .Z(n2368) );
  NAND U2846 ( .A(n2368), .B(n3668), .Z(n2369) );
  NAND U2847 ( .A(n2370), .B(n2369), .Z(n3673) );
  XNOR U2848 ( .A(a[230]), .B(b[230]), .Z(n3672) );
  NAND U2849 ( .A(n3673), .B(n3672), .Z(n2371) );
  NANDN U2850 ( .A(n2372), .B(n2371), .Z(n2378) );
  NAND U2851 ( .A(a[230]), .B(b[230]), .Z(n2379) );
  AND U2852 ( .A(n2378), .B(n2379), .Z(n2374) );
  XOR U2853 ( .A(a[231]), .B(b[231]), .Z(n3678) );
  ANDN U2854 ( .B(n3677), .A(n3678), .Z(n2373) );
  OR U2855 ( .A(n2374), .B(n2373), .Z(n2375) );
  AND U2856 ( .A(a[231]), .B(b[231]), .Z(n2377) );
  ANDN U2857 ( .B(n2375), .A(n2377), .Z(n2384) );
  NOR U2858 ( .A(n2379), .B(n2378), .Z(n2376) );
  XNOR U2859 ( .A(n2377), .B(n2376), .Z(n2382) );
  XOR U2860 ( .A(n2379), .B(n2378), .Z(n2380) );
  NAND U2861 ( .A(n2380), .B(n3678), .Z(n2381) );
  NAND U2862 ( .A(n2382), .B(n2381), .Z(n3683) );
  XNOR U2863 ( .A(a[232]), .B(b[232]), .Z(n3682) );
  NAND U2864 ( .A(n3683), .B(n3682), .Z(n2383) );
  NANDN U2865 ( .A(n2384), .B(n2383), .Z(n2390) );
  NAND U2866 ( .A(a[232]), .B(b[232]), .Z(n2391) );
  AND U2867 ( .A(n2390), .B(n2391), .Z(n2386) );
  XOR U2868 ( .A(a[233]), .B(b[233]), .Z(n3688) );
  ANDN U2869 ( .B(n3687), .A(n3688), .Z(n2385) );
  OR U2870 ( .A(n2386), .B(n2385), .Z(n2387) );
  AND U2871 ( .A(a[233]), .B(b[233]), .Z(n2389) );
  ANDN U2872 ( .B(n2387), .A(n2389), .Z(n2396) );
  NOR U2873 ( .A(n2391), .B(n2390), .Z(n2388) );
  XNOR U2874 ( .A(n2389), .B(n2388), .Z(n2394) );
  XOR U2875 ( .A(n2391), .B(n2390), .Z(n2392) );
  NAND U2876 ( .A(n2392), .B(n3688), .Z(n2393) );
  NAND U2877 ( .A(n2394), .B(n2393), .Z(n3693) );
  XNOR U2878 ( .A(a[234]), .B(b[234]), .Z(n3692) );
  NAND U2879 ( .A(n3693), .B(n3692), .Z(n2395) );
  NANDN U2880 ( .A(n2396), .B(n2395), .Z(n2402) );
  NAND U2881 ( .A(a[234]), .B(b[234]), .Z(n2403) );
  AND U2882 ( .A(n2402), .B(n2403), .Z(n2398) );
  XOR U2883 ( .A(a[235]), .B(b[235]), .Z(n3698) );
  ANDN U2884 ( .B(n3697), .A(n3698), .Z(n2397) );
  OR U2885 ( .A(n2398), .B(n2397), .Z(n2399) );
  AND U2886 ( .A(a[235]), .B(b[235]), .Z(n2401) );
  ANDN U2887 ( .B(n2399), .A(n2401), .Z(n2408) );
  NOR U2888 ( .A(n2403), .B(n2402), .Z(n2400) );
  XNOR U2889 ( .A(n2401), .B(n2400), .Z(n2406) );
  XOR U2890 ( .A(n2403), .B(n2402), .Z(n2404) );
  NAND U2891 ( .A(n2404), .B(n3698), .Z(n2405) );
  NAND U2892 ( .A(n2406), .B(n2405), .Z(n3703) );
  XNOR U2893 ( .A(a[236]), .B(b[236]), .Z(n3702) );
  NAND U2894 ( .A(n3703), .B(n3702), .Z(n2407) );
  NANDN U2895 ( .A(n2408), .B(n2407), .Z(n2409) );
  IV U2896 ( .A(n2409), .Z(n2413) );
  AND U2897 ( .A(a[236]), .B(b[236]), .Z(n2414) );
  NOR U2898 ( .A(n2413), .B(n2414), .Z(n2411) );
  XNOR U2899 ( .A(n2414), .B(n2409), .Z(n3708) );
  XNOR U2900 ( .A(a[237]), .B(b[237]), .Z(n3707) );
  AND U2901 ( .A(n3708), .B(n3707), .Z(n2410) );
  OR U2902 ( .A(n2411), .B(n2410), .Z(n2412) );
  AND U2903 ( .A(a[237]), .B(b[237]), .Z(n2416) );
  ANDN U2904 ( .B(n2412), .A(n2416), .Z(n2418) );
  AND U2905 ( .A(n2414), .B(n2413), .Z(n2415) );
  NAND U2906 ( .A(n2416), .B(n2415), .Z(n2421) );
  ANDN U2907 ( .B(n2421), .A(n2418), .Z(n3713) );
  XNOR U2908 ( .A(a[238]), .B(b[238]), .Z(n3712) );
  AND U2909 ( .A(n3713), .B(n3712), .Z(n2417) );
  OR U2910 ( .A(n2418), .B(n2417), .Z(n2419) );
  AND U2911 ( .A(a[238]), .B(b[238]), .Z(n2420) );
  ANDN U2912 ( .B(n2419), .A(n2420), .Z(n2424) );
  NANDN U2913 ( .A(n2421), .B(n2420), .Z(n2422) );
  ANDN U2914 ( .B(n2422), .A(n2424), .Z(n3718) );
  XNOR U2915 ( .A(a[239]), .B(b[239]), .Z(n3717) );
  NAND U2916 ( .A(n3718), .B(n3717), .Z(n2423) );
  NANDN U2917 ( .A(n2424), .B(n2423), .Z(n2430) );
  NAND U2918 ( .A(a[239]), .B(b[239]), .Z(n2431) );
  AND U2919 ( .A(n2430), .B(n2431), .Z(n2426) );
  XOR U2920 ( .A(a[240]), .B(b[240]), .Z(n3723) );
  ANDN U2921 ( .B(n3722), .A(n3723), .Z(n2425) );
  OR U2922 ( .A(n2426), .B(n2425), .Z(n2427) );
  AND U2923 ( .A(a[240]), .B(b[240]), .Z(n2429) );
  ANDN U2924 ( .B(n2427), .A(n2429), .Z(n2436) );
  NOR U2925 ( .A(n2431), .B(n2430), .Z(n2428) );
  XNOR U2926 ( .A(n2429), .B(n2428), .Z(n2434) );
  XOR U2927 ( .A(n2431), .B(n2430), .Z(n2432) );
  NAND U2928 ( .A(n2432), .B(n3723), .Z(n2433) );
  NAND U2929 ( .A(n2434), .B(n2433), .Z(n3728) );
  XNOR U2930 ( .A(a[241]), .B(b[241]), .Z(n3727) );
  NAND U2931 ( .A(n3728), .B(n3727), .Z(n2435) );
  NANDN U2932 ( .A(n2436), .B(n2435), .Z(n2442) );
  NAND U2933 ( .A(a[241]), .B(b[241]), .Z(n2443) );
  AND U2934 ( .A(n2442), .B(n2443), .Z(n2438) );
  XOR U2935 ( .A(a[242]), .B(b[242]), .Z(n3733) );
  ANDN U2936 ( .B(n3732), .A(n3733), .Z(n2437) );
  OR U2937 ( .A(n2438), .B(n2437), .Z(n2439) );
  AND U2938 ( .A(a[242]), .B(b[242]), .Z(n2441) );
  ANDN U2939 ( .B(n2439), .A(n2441), .Z(n2448) );
  NOR U2940 ( .A(n2443), .B(n2442), .Z(n2440) );
  XNOR U2941 ( .A(n2441), .B(n2440), .Z(n2446) );
  XOR U2942 ( .A(n2443), .B(n2442), .Z(n2444) );
  NAND U2943 ( .A(n2444), .B(n3733), .Z(n2445) );
  NAND U2944 ( .A(n2446), .B(n2445), .Z(n3738) );
  XNOR U2945 ( .A(a[243]), .B(b[243]), .Z(n3737) );
  NAND U2946 ( .A(n3738), .B(n3737), .Z(n2447) );
  NANDN U2947 ( .A(n2448), .B(n2447), .Z(n2454) );
  NAND U2948 ( .A(a[243]), .B(b[243]), .Z(n2455) );
  AND U2949 ( .A(n2454), .B(n2455), .Z(n2450) );
  XOR U2950 ( .A(a[244]), .B(b[244]), .Z(n3743) );
  ANDN U2951 ( .B(n3742), .A(n3743), .Z(n2449) );
  OR U2952 ( .A(n2450), .B(n2449), .Z(n2451) );
  AND U2953 ( .A(a[244]), .B(b[244]), .Z(n2453) );
  ANDN U2954 ( .B(n2451), .A(n2453), .Z(n2460) );
  NOR U2955 ( .A(n2455), .B(n2454), .Z(n2452) );
  XNOR U2956 ( .A(n2453), .B(n2452), .Z(n2458) );
  XOR U2957 ( .A(n2455), .B(n2454), .Z(n2456) );
  NAND U2958 ( .A(n2456), .B(n3743), .Z(n2457) );
  NAND U2959 ( .A(n2458), .B(n2457), .Z(n3748) );
  XNOR U2960 ( .A(a[245]), .B(b[245]), .Z(n3747) );
  NAND U2961 ( .A(n3748), .B(n3747), .Z(n2459) );
  NANDN U2962 ( .A(n2460), .B(n2459), .Z(n2466) );
  NAND U2963 ( .A(a[245]), .B(b[245]), .Z(n2467) );
  AND U2964 ( .A(n2466), .B(n2467), .Z(n2462) );
  XOR U2965 ( .A(a[246]), .B(b[246]), .Z(n3753) );
  ANDN U2966 ( .B(n3752), .A(n3753), .Z(n2461) );
  OR U2967 ( .A(n2462), .B(n2461), .Z(n2463) );
  AND U2968 ( .A(a[246]), .B(b[246]), .Z(n2465) );
  ANDN U2969 ( .B(n2463), .A(n2465), .Z(n2472) );
  NOR U2970 ( .A(n2467), .B(n2466), .Z(n2464) );
  XNOR U2971 ( .A(n2465), .B(n2464), .Z(n2470) );
  XOR U2972 ( .A(n2467), .B(n2466), .Z(n2468) );
  NAND U2973 ( .A(n2468), .B(n3753), .Z(n2469) );
  NAND U2974 ( .A(n2470), .B(n2469), .Z(n3758) );
  XNOR U2975 ( .A(a[247]), .B(b[247]), .Z(n3757) );
  NAND U2976 ( .A(n3758), .B(n3757), .Z(n2471) );
  NANDN U2977 ( .A(n2472), .B(n2471), .Z(n2478) );
  NAND U2978 ( .A(a[247]), .B(b[247]), .Z(n2479) );
  AND U2979 ( .A(n2478), .B(n2479), .Z(n2474) );
  XOR U2980 ( .A(a[248]), .B(b[248]), .Z(n3763) );
  ANDN U2981 ( .B(n3762), .A(n3763), .Z(n2473) );
  OR U2982 ( .A(n2474), .B(n2473), .Z(n2475) );
  AND U2983 ( .A(a[248]), .B(b[248]), .Z(n2477) );
  ANDN U2984 ( .B(n2475), .A(n2477), .Z(n2484) );
  NOR U2985 ( .A(n2479), .B(n2478), .Z(n2476) );
  XNOR U2986 ( .A(n2477), .B(n2476), .Z(n2482) );
  XOR U2987 ( .A(n2479), .B(n2478), .Z(n2480) );
  NAND U2988 ( .A(n2480), .B(n3763), .Z(n2481) );
  NAND U2989 ( .A(n2482), .B(n2481), .Z(n3768) );
  XNOR U2990 ( .A(a[249]), .B(b[249]), .Z(n3767) );
  NAND U2991 ( .A(n3768), .B(n3767), .Z(n2483) );
  NANDN U2992 ( .A(n2484), .B(n2483), .Z(n2490) );
  NAND U2993 ( .A(a[249]), .B(b[249]), .Z(n2491) );
  AND U2994 ( .A(n2490), .B(n2491), .Z(n2486) );
  XOR U2995 ( .A(a[250]), .B(b[250]), .Z(n3773) );
  ANDN U2996 ( .B(n3772), .A(n3773), .Z(n2485) );
  OR U2997 ( .A(n2486), .B(n2485), .Z(n2487) );
  AND U2998 ( .A(a[250]), .B(b[250]), .Z(n2489) );
  ANDN U2999 ( .B(n2487), .A(n2489), .Z(n2496) );
  NOR U3000 ( .A(n2491), .B(n2490), .Z(n2488) );
  XNOR U3001 ( .A(n2489), .B(n2488), .Z(n2494) );
  XOR U3002 ( .A(n2491), .B(n2490), .Z(n2492) );
  NAND U3003 ( .A(n2492), .B(n3773), .Z(n2493) );
  NAND U3004 ( .A(n2494), .B(n2493), .Z(n3778) );
  XNOR U3005 ( .A(a[251]), .B(b[251]), .Z(n3777) );
  NAND U3006 ( .A(n3778), .B(n3777), .Z(n2495) );
  NANDN U3007 ( .A(n2496), .B(n2495), .Z(n2502) );
  NAND U3008 ( .A(a[251]), .B(b[251]), .Z(n2503) );
  AND U3009 ( .A(n2502), .B(n2503), .Z(n2498) );
  XOR U3010 ( .A(a[252]), .B(b[252]), .Z(n3783) );
  ANDN U3011 ( .B(n3782), .A(n3783), .Z(n2497) );
  OR U3012 ( .A(n2498), .B(n2497), .Z(n2499) );
  AND U3013 ( .A(a[252]), .B(b[252]), .Z(n2501) );
  ANDN U3014 ( .B(n2499), .A(n2501), .Z(n2508) );
  NOR U3015 ( .A(n2503), .B(n2502), .Z(n2500) );
  XNOR U3016 ( .A(n2501), .B(n2500), .Z(n2506) );
  XOR U3017 ( .A(n2503), .B(n2502), .Z(n2504) );
  NAND U3018 ( .A(n2504), .B(n3783), .Z(n2505) );
  NAND U3019 ( .A(n2506), .B(n2505), .Z(n3788) );
  XNOR U3020 ( .A(a[253]), .B(b[253]), .Z(n3787) );
  NAND U3021 ( .A(n3788), .B(n3787), .Z(n2507) );
  NANDN U3022 ( .A(n2508), .B(n2507), .Z(n2514) );
  NOR U3023 ( .A(n2513), .B(n2514), .Z(n2509) );
  XOR U3024 ( .A(n2518), .B(n2509), .Z(n2512) );
  XNOR U3025 ( .A(a[254]), .B(b[254]), .Z(n3793) );
  XOR U3026 ( .A(n2513), .B(n2514), .Z(n2510) );
  NANDN U3027 ( .A(n3793), .B(n2510), .Z(n2511) );
  NAND U3028 ( .A(n2512), .B(n2511), .Z(n3798) );
  XNOR U3029 ( .A(a[255]), .B(b[255]), .Z(n3797) );
  NAND U3030 ( .A(n3798), .B(n3797), .Z(n2520) );
  AND U3031 ( .A(n2514), .B(n2513), .Z(n2516) );
  AND U3032 ( .A(n3792), .B(n3793), .Z(n2515) );
  OR U3033 ( .A(n2516), .B(n2515), .Z(n2517) );
  AND U3034 ( .A(n2518), .B(n2517), .Z(n2519) );
  ANDN U3035 ( .B(n2520), .A(n2519), .Z(n2521) );
  XOR U3036 ( .A(n2522), .B(n2521), .Z(N514) );
  AND U3037 ( .A(n2522), .B(n2521), .Z(N515) );
  NAND U3039 ( .A(c[0]), .B(rst), .Z(n2526) );
  XOR U3040 ( .A(n2523), .B(carry_on[0]), .Z(n2524) );
  NANDN U3041 ( .A(rst), .B(n2524), .Z(n2525) );
  NAND U3042 ( .A(n2526), .B(n2525), .Z(n769) );
  NAND U3043 ( .A(c[1]), .B(rst), .Z(n2531) );
  XOR U3044 ( .A(n2528), .B(n2527), .Z(n2529) );
  NANDN U3045 ( .A(rst), .B(n2529), .Z(n2530) );
  NAND U3046 ( .A(n2531), .B(n2530), .Z(n770) );
  NAND U3047 ( .A(c[2]), .B(rst), .Z(n2536) );
  XNOR U3048 ( .A(n2533), .B(n2532), .Z(n2534) );
  NANDN U3049 ( .A(rst), .B(n2534), .Z(n2535) );
  NAND U3050 ( .A(n2536), .B(n2535), .Z(n771) );
  NAND U3051 ( .A(c[3]), .B(rst), .Z(n2541) );
  XOR U3052 ( .A(n2538), .B(n2537), .Z(n2539) );
  NANDN U3053 ( .A(rst), .B(n2539), .Z(n2540) );
  NAND U3054 ( .A(n2541), .B(n2540), .Z(n772) );
  NAND U3055 ( .A(c[4]), .B(rst), .Z(n2546) );
  XNOR U3056 ( .A(n2543), .B(n2542), .Z(n2544) );
  NANDN U3057 ( .A(rst), .B(n2544), .Z(n2545) );
  NAND U3058 ( .A(n2546), .B(n2545), .Z(n773) );
  NAND U3059 ( .A(c[5]), .B(rst), .Z(n2551) );
  XNOR U3060 ( .A(n2548), .B(n2547), .Z(n2549) );
  NANDN U3061 ( .A(rst), .B(n2549), .Z(n2550) );
  NAND U3062 ( .A(n2551), .B(n2550), .Z(n774) );
  NAND U3063 ( .A(c[6]), .B(rst), .Z(n2556) );
  XNOR U3064 ( .A(n2553), .B(n2552), .Z(n2554) );
  NANDN U3065 ( .A(rst), .B(n2554), .Z(n2555) );
  NAND U3066 ( .A(n2556), .B(n2555), .Z(n775) );
  NAND U3067 ( .A(c[7]), .B(rst), .Z(n2561) );
  XNOR U3068 ( .A(n2558), .B(n2557), .Z(n2559) );
  NANDN U3069 ( .A(rst), .B(n2559), .Z(n2560) );
  NAND U3070 ( .A(n2561), .B(n2560), .Z(n776) );
  NAND U3071 ( .A(c[8]), .B(rst), .Z(n2566) );
  XOR U3072 ( .A(n2563), .B(n2562), .Z(n2564) );
  NANDN U3073 ( .A(rst), .B(n2564), .Z(n2565) );
  NAND U3074 ( .A(n2566), .B(n2565), .Z(n777) );
  NAND U3075 ( .A(c[9]), .B(rst), .Z(n2571) );
  XNOR U3076 ( .A(n2568), .B(n2567), .Z(n2569) );
  NANDN U3077 ( .A(rst), .B(n2569), .Z(n2570) );
  NAND U3078 ( .A(n2571), .B(n2570), .Z(n778) );
  NAND U3079 ( .A(c[10]), .B(rst), .Z(n2576) );
  XOR U3080 ( .A(n2573), .B(n2572), .Z(n2574) );
  NANDN U3081 ( .A(rst), .B(n2574), .Z(n2575) );
  NAND U3082 ( .A(n2576), .B(n2575), .Z(n779) );
  NAND U3083 ( .A(c[11]), .B(rst), .Z(n2581) );
  XNOR U3084 ( .A(n2578), .B(n2577), .Z(n2579) );
  NANDN U3085 ( .A(rst), .B(n2579), .Z(n2580) );
  NAND U3086 ( .A(n2581), .B(n2580), .Z(n780) );
  NAND U3087 ( .A(c[12]), .B(rst), .Z(n2586) );
  XOR U3088 ( .A(n2583), .B(n2582), .Z(n2584) );
  NANDN U3089 ( .A(rst), .B(n2584), .Z(n2585) );
  NAND U3090 ( .A(n2586), .B(n2585), .Z(n781) );
  NAND U3091 ( .A(c[13]), .B(rst), .Z(n2591) );
  XNOR U3092 ( .A(n2588), .B(n2587), .Z(n2589) );
  NANDN U3093 ( .A(rst), .B(n2589), .Z(n2590) );
  NAND U3094 ( .A(n2591), .B(n2590), .Z(n782) );
  NAND U3095 ( .A(c[14]), .B(rst), .Z(n2596) );
  XOR U3096 ( .A(n2593), .B(n2592), .Z(n2594) );
  NANDN U3097 ( .A(rst), .B(n2594), .Z(n2595) );
  NAND U3098 ( .A(n2596), .B(n2595), .Z(n783) );
  NAND U3099 ( .A(c[15]), .B(rst), .Z(n2601) );
  XNOR U3100 ( .A(n2598), .B(n2597), .Z(n2599) );
  NANDN U3101 ( .A(rst), .B(n2599), .Z(n2600) );
  NAND U3102 ( .A(n2601), .B(n2600), .Z(n784) );
  NAND U3103 ( .A(c[16]), .B(rst), .Z(n2606) );
  XOR U3104 ( .A(n2603), .B(n2602), .Z(n2604) );
  NANDN U3105 ( .A(rst), .B(n2604), .Z(n2605) );
  NAND U3106 ( .A(n2606), .B(n2605), .Z(n785) );
  NAND U3107 ( .A(c[17]), .B(rst), .Z(n2611) );
  XNOR U3108 ( .A(n2608), .B(n2607), .Z(n2609) );
  NANDN U3109 ( .A(rst), .B(n2609), .Z(n2610) );
  NAND U3110 ( .A(n2611), .B(n2610), .Z(n786) );
  NAND U3111 ( .A(c[18]), .B(rst), .Z(n2616) );
  XOR U3112 ( .A(n2613), .B(n2612), .Z(n2614) );
  NANDN U3113 ( .A(rst), .B(n2614), .Z(n2615) );
  NAND U3114 ( .A(n2616), .B(n2615), .Z(n787) );
  NAND U3115 ( .A(c[19]), .B(rst), .Z(n2621) );
  XNOR U3116 ( .A(n2618), .B(n2617), .Z(n2619) );
  NANDN U3117 ( .A(rst), .B(n2619), .Z(n2620) );
  NAND U3118 ( .A(n2621), .B(n2620), .Z(n788) );
  NAND U3119 ( .A(c[20]), .B(rst), .Z(n2626) );
  XOR U3120 ( .A(n2623), .B(n2622), .Z(n2624) );
  NANDN U3121 ( .A(rst), .B(n2624), .Z(n2625) );
  NAND U3122 ( .A(n2626), .B(n2625), .Z(n789) );
  NAND U3123 ( .A(c[21]), .B(rst), .Z(n2631) );
  XNOR U3124 ( .A(n2628), .B(n2627), .Z(n2629) );
  NANDN U3125 ( .A(rst), .B(n2629), .Z(n2630) );
  NAND U3126 ( .A(n2631), .B(n2630), .Z(n790) );
  NAND U3127 ( .A(c[22]), .B(rst), .Z(n2636) );
  XNOR U3128 ( .A(n2633), .B(n2632), .Z(n2634) );
  NANDN U3129 ( .A(rst), .B(n2634), .Z(n2635) );
  NAND U3130 ( .A(n2636), .B(n2635), .Z(n791) );
  NAND U3131 ( .A(c[23]), .B(rst), .Z(n2641) );
  XNOR U3132 ( .A(n2638), .B(n2637), .Z(n2639) );
  NANDN U3133 ( .A(rst), .B(n2639), .Z(n2640) );
  NAND U3134 ( .A(n2641), .B(n2640), .Z(n792) );
  NAND U3135 ( .A(c[24]), .B(rst), .Z(n2646) );
  XNOR U3136 ( .A(n2643), .B(n2642), .Z(n2644) );
  NANDN U3137 ( .A(rst), .B(n2644), .Z(n2645) );
  NAND U3138 ( .A(n2646), .B(n2645), .Z(n793) );
  NAND U3139 ( .A(c[25]), .B(rst), .Z(n2651) );
  XOR U3140 ( .A(n2648), .B(n2647), .Z(n2649) );
  NANDN U3141 ( .A(rst), .B(n2649), .Z(n2650) );
  NAND U3142 ( .A(n2651), .B(n2650), .Z(n794) );
  NAND U3143 ( .A(c[26]), .B(rst), .Z(n2656) );
  XNOR U3144 ( .A(n2653), .B(n2652), .Z(n2654) );
  NANDN U3145 ( .A(rst), .B(n2654), .Z(n2655) );
  NAND U3146 ( .A(n2656), .B(n2655), .Z(n795) );
  NAND U3147 ( .A(c[27]), .B(rst), .Z(n2661) );
  XOR U3148 ( .A(n2658), .B(n2657), .Z(n2659) );
  NANDN U3149 ( .A(rst), .B(n2659), .Z(n2660) );
  NAND U3150 ( .A(n2661), .B(n2660), .Z(n796) );
  NAND U3151 ( .A(c[28]), .B(rst), .Z(n2666) );
  XNOR U3152 ( .A(n2663), .B(n2662), .Z(n2664) );
  NANDN U3153 ( .A(rst), .B(n2664), .Z(n2665) );
  NAND U3154 ( .A(n2666), .B(n2665), .Z(n797) );
  NAND U3155 ( .A(c[29]), .B(rst), .Z(n2671) );
  XNOR U3156 ( .A(n2668), .B(n2667), .Z(n2669) );
  NANDN U3157 ( .A(rst), .B(n2669), .Z(n2670) );
  NAND U3158 ( .A(n2671), .B(n2670), .Z(n798) );
  NAND U3159 ( .A(c[30]), .B(rst), .Z(n2676) );
  XNOR U3160 ( .A(n2673), .B(n2672), .Z(n2674) );
  NANDN U3161 ( .A(rst), .B(n2674), .Z(n2675) );
  NAND U3162 ( .A(n2676), .B(n2675), .Z(n799) );
  NAND U3163 ( .A(c[31]), .B(rst), .Z(n2681) );
  XNOR U3164 ( .A(n2678), .B(n2677), .Z(n2679) );
  NANDN U3165 ( .A(rst), .B(n2679), .Z(n2680) );
  NAND U3166 ( .A(n2681), .B(n2680), .Z(n800) );
  NAND U3167 ( .A(c[32]), .B(rst), .Z(n2686) );
  XOR U3168 ( .A(n2683), .B(n2682), .Z(n2684) );
  NANDN U3169 ( .A(rst), .B(n2684), .Z(n2685) );
  NAND U3170 ( .A(n2686), .B(n2685), .Z(n801) );
  NAND U3171 ( .A(c[33]), .B(rst), .Z(n2691) );
  XNOR U3172 ( .A(n2688), .B(n2687), .Z(n2689) );
  NANDN U3173 ( .A(rst), .B(n2689), .Z(n2690) );
  NAND U3174 ( .A(n2691), .B(n2690), .Z(n802) );
  NAND U3175 ( .A(c[34]), .B(rst), .Z(n2696) );
  XOR U3176 ( .A(n2693), .B(n2692), .Z(n2694) );
  NANDN U3177 ( .A(rst), .B(n2694), .Z(n2695) );
  NAND U3178 ( .A(n2696), .B(n2695), .Z(n803) );
  NAND U3179 ( .A(c[35]), .B(rst), .Z(n2701) );
  XNOR U3180 ( .A(n2698), .B(n2697), .Z(n2699) );
  NANDN U3181 ( .A(rst), .B(n2699), .Z(n2700) );
  NAND U3182 ( .A(n2701), .B(n2700), .Z(n804) );
  NAND U3183 ( .A(c[36]), .B(rst), .Z(n2706) );
  XOR U3184 ( .A(n2703), .B(n2702), .Z(n2704) );
  NANDN U3185 ( .A(rst), .B(n2704), .Z(n2705) );
  NAND U3186 ( .A(n2706), .B(n2705), .Z(n805) );
  NAND U3187 ( .A(c[37]), .B(rst), .Z(n2711) );
  XNOR U3188 ( .A(n2708), .B(n2707), .Z(n2709) );
  NANDN U3189 ( .A(rst), .B(n2709), .Z(n2710) );
  NAND U3190 ( .A(n2711), .B(n2710), .Z(n806) );
  NAND U3191 ( .A(c[38]), .B(rst), .Z(n2716) );
  XOR U3192 ( .A(n2713), .B(n2712), .Z(n2714) );
  NANDN U3193 ( .A(rst), .B(n2714), .Z(n2715) );
  NAND U3194 ( .A(n2716), .B(n2715), .Z(n807) );
  NAND U3195 ( .A(c[39]), .B(rst), .Z(n2721) );
  XNOR U3196 ( .A(n2718), .B(n2717), .Z(n2719) );
  NANDN U3197 ( .A(rst), .B(n2719), .Z(n2720) );
  NAND U3198 ( .A(n2721), .B(n2720), .Z(n808) );
  NAND U3199 ( .A(c[40]), .B(rst), .Z(n2726) );
  XOR U3200 ( .A(n2723), .B(n2722), .Z(n2724) );
  NANDN U3201 ( .A(rst), .B(n2724), .Z(n2725) );
  NAND U3202 ( .A(n2726), .B(n2725), .Z(n809) );
  NAND U3203 ( .A(c[41]), .B(rst), .Z(n2731) );
  XNOR U3204 ( .A(n2728), .B(n2727), .Z(n2729) );
  NANDN U3205 ( .A(rst), .B(n2729), .Z(n2730) );
  NAND U3206 ( .A(n2731), .B(n2730), .Z(n810) );
  NAND U3207 ( .A(c[42]), .B(rst), .Z(n2736) );
  XOR U3208 ( .A(n2733), .B(n2732), .Z(n2734) );
  NANDN U3209 ( .A(rst), .B(n2734), .Z(n2735) );
  NAND U3210 ( .A(n2736), .B(n2735), .Z(n811) );
  NAND U3211 ( .A(c[43]), .B(rst), .Z(n2741) );
  XNOR U3212 ( .A(n2738), .B(n2737), .Z(n2739) );
  NANDN U3213 ( .A(rst), .B(n2739), .Z(n2740) );
  NAND U3214 ( .A(n2741), .B(n2740), .Z(n812) );
  NAND U3215 ( .A(c[44]), .B(rst), .Z(n2746) );
  XOR U3216 ( .A(n2743), .B(n2742), .Z(n2744) );
  NANDN U3217 ( .A(rst), .B(n2744), .Z(n2745) );
  NAND U3218 ( .A(n2746), .B(n2745), .Z(n813) );
  NAND U3219 ( .A(c[45]), .B(rst), .Z(n2751) );
  XNOR U3220 ( .A(n2748), .B(n2747), .Z(n2749) );
  NANDN U3221 ( .A(rst), .B(n2749), .Z(n2750) );
  NAND U3222 ( .A(n2751), .B(n2750), .Z(n814) );
  NAND U3223 ( .A(c[46]), .B(rst), .Z(n2756) );
  XOR U3224 ( .A(n2753), .B(n2752), .Z(n2754) );
  NANDN U3225 ( .A(rst), .B(n2754), .Z(n2755) );
  NAND U3226 ( .A(n2756), .B(n2755), .Z(n815) );
  NAND U3227 ( .A(c[47]), .B(rst), .Z(n2761) );
  XNOR U3228 ( .A(n2758), .B(n2757), .Z(n2759) );
  NANDN U3229 ( .A(rst), .B(n2759), .Z(n2760) );
  NAND U3230 ( .A(n2761), .B(n2760), .Z(n816) );
  NAND U3231 ( .A(c[48]), .B(rst), .Z(n2766) );
  XOR U3232 ( .A(n2763), .B(n2762), .Z(n2764) );
  NANDN U3233 ( .A(rst), .B(n2764), .Z(n2765) );
  NAND U3234 ( .A(n2766), .B(n2765), .Z(n817) );
  NAND U3235 ( .A(c[49]), .B(rst), .Z(n2771) );
  XNOR U3236 ( .A(n2768), .B(n2767), .Z(n2769) );
  NANDN U3237 ( .A(rst), .B(n2769), .Z(n2770) );
  NAND U3238 ( .A(n2771), .B(n2770), .Z(n818) );
  NAND U3239 ( .A(c[50]), .B(rst), .Z(n2776) );
  XOR U3240 ( .A(n2773), .B(n2772), .Z(n2774) );
  NANDN U3241 ( .A(rst), .B(n2774), .Z(n2775) );
  NAND U3242 ( .A(n2776), .B(n2775), .Z(n819) );
  NAND U3243 ( .A(c[51]), .B(rst), .Z(n2781) );
  XNOR U3244 ( .A(n2778), .B(n2777), .Z(n2779) );
  NANDN U3245 ( .A(rst), .B(n2779), .Z(n2780) );
  NAND U3246 ( .A(n2781), .B(n2780), .Z(n820) );
  NAND U3247 ( .A(c[52]), .B(rst), .Z(n2786) );
  XOR U3248 ( .A(n2783), .B(n2782), .Z(n2784) );
  NANDN U3249 ( .A(rst), .B(n2784), .Z(n2785) );
  NAND U3250 ( .A(n2786), .B(n2785), .Z(n821) );
  NAND U3251 ( .A(c[53]), .B(rst), .Z(n2791) );
  XNOR U3252 ( .A(n2788), .B(n2787), .Z(n2789) );
  NANDN U3253 ( .A(rst), .B(n2789), .Z(n2790) );
  NAND U3254 ( .A(n2791), .B(n2790), .Z(n822) );
  NAND U3255 ( .A(c[54]), .B(rst), .Z(n2796) );
  XOR U3256 ( .A(n2793), .B(n2792), .Z(n2794) );
  NANDN U3257 ( .A(rst), .B(n2794), .Z(n2795) );
  NAND U3258 ( .A(n2796), .B(n2795), .Z(n823) );
  NAND U3259 ( .A(c[55]), .B(rst), .Z(n2801) );
  XNOR U3260 ( .A(n2798), .B(n2797), .Z(n2799) );
  NANDN U3261 ( .A(rst), .B(n2799), .Z(n2800) );
  NAND U3262 ( .A(n2801), .B(n2800), .Z(n824) );
  NAND U3263 ( .A(c[56]), .B(rst), .Z(n2806) );
  XOR U3264 ( .A(n2803), .B(n2802), .Z(n2804) );
  NANDN U3265 ( .A(rst), .B(n2804), .Z(n2805) );
  NAND U3266 ( .A(n2806), .B(n2805), .Z(n825) );
  NAND U3267 ( .A(c[57]), .B(rst), .Z(n2811) );
  XNOR U3268 ( .A(n2808), .B(n2807), .Z(n2809) );
  NANDN U3269 ( .A(rst), .B(n2809), .Z(n2810) );
  NAND U3270 ( .A(n2811), .B(n2810), .Z(n826) );
  NAND U3271 ( .A(c[58]), .B(rst), .Z(n2816) );
  XOR U3272 ( .A(n2813), .B(n2812), .Z(n2814) );
  NANDN U3273 ( .A(rst), .B(n2814), .Z(n2815) );
  NAND U3274 ( .A(n2816), .B(n2815), .Z(n827) );
  NAND U3275 ( .A(c[59]), .B(rst), .Z(n2821) );
  XNOR U3276 ( .A(n2818), .B(n2817), .Z(n2819) );
  NANDN U3277 ( .A(rst), .B(n2819), .Z(n2820) );
  NAND U3278 ( .A(n2821), .B(n2820), .Z(n828) );
  NAND U3279 ( .A(c[60]), .B(rst), .Z(n2826) );
  XOR U3280 ( .A(n2823), .B(n2822), .Z(n2824) );
  NANDN U3281 ( .A(rst), .B(n2824), .Z(n2825) );
  NAND U3282 ( .A(n2826), .B(n2825), .Z(n829) );
  NAND U3283 ( .A(c[61]), .B(rst), .Z(n2831) );
  XNOR U3284 ( .A(n2828), .B(n2827), .Z(n2829) );
  NANDN U3285 ( .A(rst), .B(n2829), .Z(n2830) );
  NAND U3286 ( .A(n2831), .B(n2830), .Z(n830) );
  NAND U3287 ( .A(c[62]), .B(rst), .Z(n2836) );
  XOR U3288 ( .A(n2833), .B(n2832), .Z(n2834) );
  NANDN U3289 ( .A(rst), .B(n2834), .Z(n2835) );
  NAND U3290 ( .A(n2836), .B(n2835), .Z(n831) );
  NAND U3291 ( .A(c[63]), .B(rst), .Z(n2841) );
  XNOR U3292 ( .A(n2838), .B(n2837), .Z(n2839) );
  NANDN U3293 ( .A(rst), .B(n2839), .Z(n2840) );
  NAND U3294 ( .A(n2841), .B(n2840), .Z(n832) );
  NAND U3295 ( .A(c[64]), .B(rst), .Z(n2846) );
  XOR U3296 ( .A(n2843), .B(n2842), .Z(n2844) );
  NANDN U3297 ( .A(rst), .B(n2844), .Z(n2845) );
  NAND U3298 ( .A(n2846), .B(n2845), .Z(n833) );
  NAND U3299 ( .A(c[65]), .B(rst), .Z(n2851) );
  XNOR U3300 ( .A(n2848), .B(n2847), .Z(n2849) );
  NANDN U3301 ( .A(rst), .B(n2849), .Z(n2850) );
  NAND U3302 ( .A(n2851), .B(n2850), .Z(n834) );
  NAND U3303 ( .A(c[66]), .B(rst), .Z(n2856) );
  XOR U3304 ( .A(n2853), .B(n2852), .Z(n2854) );
  NANDN U3305 ( .A(rst), .B(n2854), .Z(n2855) );
  NAND U3306 ( .A(n2856), .B(n2855), .Z(n835) );
  NAND U3307 ( .A(c[67]), .B(rst), .Z(n2861) );
  XNOR U3308 ( .A(n2858), .B(n2857), .Z(n2859) );
  NANDN U3309 ( .A(rst), .B(n2859), .Z(n2860) );
  NAND U3310 ( .A(n2861), .B(n2860), .Z(n836) );
  NAND U3311 ( .A(c[68]), .B(rst), .Z(n2866) );
  XOR U3312 ( .A(n2863), .B(n2862), .Z(n2864) );
  NANDN U3313 ( .A(rst), .B(n2864), .Z(n2865) );
  NAND U3314 ( .A(n2866), .B(n2865), .Z(n837) );
  NAND U3315 ( .A(c[69]), .B(rst), .Z(n2871) );
  XNOR U3316 ( .A(n2868), .B(n2867), .Z(n2869) );
  NANDN U3317 ( .A(rst), .B(n2869), .Z(n2870) );
  NAND U3318 ( .A(n2871), .B(n2870), .Z(n838) );
  NAND U3319 ( .A(c[70]), .B(rst), .Z(n2876) );
  XOR U3320 ( .A(n2873), .B(n2872), .Z(n2874) );
  NANDN U3321 ( .A(rst), .B(n2874), .Z(n2875) );
  NAND U3322 ( .A(n2876), .B(n2875), .Z(n839) );
  NAND U3323 ( .A(c[71]), .B(rst), .Z(n2881) );
  XNOR U3324 ( .A(n2878), .B(n2877), .Z(n2879) );
  NANDN U3325 ( .A(rst), .B(n2879), .Z(n2880) );
  NAND U3326 ( .A(n2881), .B(n2880), .Z(n840) );
  NAND U3327 ( .A(c[72]), .B(rst), .Z(n2886) );
  XOR U3328 ( .A(n2883), .B(n2882), .Z(n2884) );
  NANDN U3329 ( .A(rst), .B(n2884), .Z(n2885) );
  NAND U3330 ( .A(n2886), .B(n2885), .Z(n841) );
  NAND U3331 ( .A(c[73]), .B(rst), .Z(n2891) );
  XNOR U3332 ( .A(n2888), .B(n2887), .Z(n2889) );
  NANDN U3333 ( .A(rst), .B(n2889), .Z(n2890) );
  NAND U3334 ( .A(n2891), .B(n2890), .Z(n842) );
  NAND U3335 ( .A(c[74]), .B(rst), .Z(n2896) );
  XOR U3336 ( .A(n2893), .B(n2892), .Z(n2894) );
  NANDN U3337 ( .A(rst), .B(n2894), .Z(n2895) );
  NAND U3338 ( .A(n2896), .B(n2895), .Z(n843) );
  NAND U3339 ( .A(c[75]), .B(rst), .Z(n2901) );
  XNOR U3340 ( .A(n2898), .B(n2897), .Z(n2899) );
  NANDN U3341 ( .A(rst), .B(n2899), .Z(n2900) );
  NAND U3342 ( .A(n2901), .B(n2900), .Z(n844) );
  NAND U3343 ( .A(c[76]), .B(rst), .Z(n2906) );
  XOR U3344 ( .A(n2903), .B(n2902), .Z(n2904) );
  NANDN U3345 ( .A(rst), .B(n2904), .Z(n2905) );
  NAND U3346 ( .A(n2906), .B(n2905), .Z(n845) );
  NAND U3347 ( .A(c[77]), .B(rst), .Z(n2911) );
  XNOR U3348 ( .A(n2908), .B(n2907), .Z(n2909) );
  NANDN U3349 ( .A(rst), .B(n2909), .Z(n2910) );
  NAND U3350 ( .A(n2911), .B(n2910), .Z(n846) );
  NAND U3351 ( .A(c[78]), .B(rst), .Z(n2916) );
  XOR U3352 ( .A(n2913), .B(n2912), .Z(n2914) );
  NANDN U3353 ( .A(rst), .B(n2914), .Z(n2915) );
  NAND U3354 ( .A(n2916), .B(n2915), .Z(n847) );
  NAND U3355 ( .A(c[79]), .B(rst), .Z(n2921) );
  XNOR U3356 ( .A(n2918), .B(n2917), .Z(n2919) );
  NANDN U3357 ( .A(rst), .B(n2919), .Z(n2920) );
  NAND U3358 ( .A(n2921), .B(n2920), .Z(n848) );
  NAND U3359 ( .A(c[80]), .B(rst), .Z(n2926) );
  XOR U3360 ( .A(n2923), .B(n2922), .Z(n2924) );
  NANDN U3361 ( .A(rst), .B(n2924), .Z(n2925) );
  NAND U3362 ( .A(n2926), .B(n2925), .Z(n849) );
  NAND U3363 ( .A(c[81]), .B(rst), .Z(n2931) );
  XNOR U3364 ( .A(n2928), .B(n2927), .Z(n2929) );
  NANDN U3365 ( .A(rst), .B(n2929), .Z(n2930) );
  NAND U3366 ( .A(n2931), .B(n2930), .Z(n850) );
  NAND U3367 ( .A(c[82]), .B(rst), .Z(n2936) );
  XOR U3368 ( .A(n2933), .B(n2932), .Z(n2934) );
  NANDN U3369 ( .A(rst), .B(n2934), .Z(n2935) );
  NAND U3370 ( .A(n2936), .B(n2935), .Z(n851) );
  NAND U3371 ( .A(c[83]), .B(rst), .Z(n2941) );
  XNOR U3372 ( .A(n2938), .B(n2937), .Z(n2939) );
  NANDN U3373 ( .A(rst), .B(n2939), .Z(n2940) );
  NAND U3374 ( .A(n2941), .B(n2940), .Z(n852) );
  NAND U3375 ( .A(c[84]), .B(rst), .Z(n2946) );
  XNOR U3376 ( .A(n2943), .B(n2942), .Z(n2944) );
  NANDN U3377 ( .A(rst), .B(n2944), .Z(n2945) );
  NAND U3378 ( .A(n2946), .B(n2945), .Z(n853) );
  NAND U3379 ( .A(c[85]), .B(rst), .Z(n2951) );
  XNOR U3380 ( .A(n2948), .B(n2947), .Z(n2949) );
  NANDN U3381 ( .A(rst), .B(n2949), .Z(n2950) );
  NAND U3382 ( .A(n2951), .B(n2950), .Z(n854) );
  NAND U3383 ( .A(c[86]), .B(rst), .Z(n2956) );
  XNOR U3384 ( .A(n2953), .B(n2952), .Z(n2954) );
  NANDN U3385 ( .A(rst), .B(n2954), .Z(n2955) );
  NAND U3386 ( .A(n2956), .B(n2955), .Z(n855) );
  NAND U3387 ( .A(c[87]), .B(rst), .Z(n2961) );
  XOR U3388 ( .A(n2958), .B(n2957), .Z(n2959) );
  NANDN U3389 ( .A(rst), .B(n2959), .Z(n2960) );
  NAND U3390 ( .A(n2961), .B(n2960), .Z(n856) );
  NAND U3391 ( .A(c[88]), .B(rst), .Z(n2966) );
  XNOR U3392 ( .A(n2963), .B(n2962), .Z(n2964) );
  NANDN U3393 ( .A(rst), .B(n2964), .Z(n2965) );
  NAND U3394 ( .A(n2966), .B(n2965), .Z(n857) );
  NAND U3395 ( .A(c[89]), .B(rst), .Z(n2971) );
  XNOR U3396 ( .A(n2968), .B(n2967), .Z(n2969) );
  NANDN U3397 ( .A(rst), .B(n2969), .Z(n2970) );
  NAND U3398 ( .A(n2971), .B(n2970), .Z(n858) );
  NAND U3399 ( .A(c[90]), .B(rst), .Z(n2976) );
  XNOR U3400 ( .A(n2973), .B(n2972), .Z(n2974) );
  NANDN U3401 ( .A(rst), .B(n2974), .Z(n2975) );
  NAND U3402 ( .A(n2976), .B(n2975), .Z(n859) );
  NAND U3403 ( .A(c[91]), .B(rst), .Z(n2981) );
  XNOR U3404 ( .A(n2978), .B(n2977), .Z(n2979) );
  NANDN U3405 ( .A(rst), .B(n2979), .Z(n2980) );
  NAND U3406 ( .A(n2981), .B(n2980), .Z(n860) );
  NAND U3407 ( .A(c[92]), .B(rst), .Z(n2986) );
  XOR U3408 ( .A(n2983), .B(n2982), .Z(n2984) );
  NANDN U3409 ( .A(rst), .B(n2984), .Z(n2985) );
  NAND U3410 ( .A(n2986), .B(n2985), .Z(n861) );
  NAND U3411 ( .A(c[93]), .B(rst), .Z(n2991) );
  XNOR U3412 ( .A(n2988), .B(n2987), .Z(n2989) );
  NANDN U3413 ( .A(rst), .B(n2989), .Z(n2990) );
  NAND U3414 ( .A(n2991), .B(n2990), .Z(n862) );
  NAND U3415 ( .A(c[94]), .B(rst), .Z(n2996) );
  XNOR U3416 ( .A(n2993), .B(n2992), .Z(n2994) );
  NANDN U3417 ( .A(rst), .B(n2994), .Z(n2995) );
  NAND U3418 ( .A(n2996), .B(n2995), .Z(n863) );
  NAND U3419 ( .A(c[95]), .B(rst), .Z(n3001) );
  XNOR U3420 ( .A(n2998), .B(n2997), .Z(n2999) );
  NANDN U3421 ( .A(rst), .B(n2999), .Z(n3000) );
  NAND U3422 ( .A(n3001), .B(n3000), .Z(n864) );
  NAND U3423 ( .A(c[96]), .B(rst), .Z(n3006) );
  XNOR U3424 ( .A(n3003), .B(n3002), .Z(n3004) );
  NANDN U3425 ( .A(rst), .B(n3004), .Z(n3005) );
  NAND U3426 ( .A(n3006), .B(n3005), .Z(n865) );
  NAND U3427 ( .A(c[97]), .B(rst), .Z(n3011) );
  XOR U3428 ( .A(n3008), .B(n3007), .Z(n3009) );
  NANDN U3429 ( .A(rst), .B(n3009), .Z(n3010) );
  NAND U3430 ( .A(n3011), .B(n3010), .Z(n866) );
  NAND U3431 ( .A(c[98]), .B(rst), .Z(n3016) );
  XNOR U3432 ( .A(n3013), .B(n3012), .Z(n3014) );
  NANDN U3433 ( .A(rst), .B(n3014), .Z(n3015) );
  NAND U3434 ( .A(n3016), .B(n3015), .Z(n867) );
  NAND U3435 ( .A(c[99]), .B(rst), .Z(n3021) );
  XOR U3436 ( .A(n3018), .B(n3017), .Z(n3019) );
  NANDN U3437 ( .A(rst), .B(n3019), .Z(n3020) );
  NAND U3438 ( .A(n3021), .B(n3020), .Z(n868) );
  NAND U3439 ( .A(c[100]), .B(rst), .Z(n3026) );
  XNOR U3440 ( .A(n3023), .B(n3022), .Z(n3024) );
  NANDN U3441 ( .A(rst), .B(n3024), .Z(n3025) );
  NAND U3442 ( .A(n3026), .B(n3025), .Z(n869) );
  NAND U3443 ( .A(c[101]), .B(rst), .Z(n3031) );
  XOR U3444 ( .A(n3028), .B(n3027), .Z(n3029) );
  NANDN U3445 ( .A(rst), .B(n3029), .Z(n3030) );
  NAND U3446 ( .A(n3031), .B(n3030), .Z(n870) );
  NAND U3447 ( .A(c[102]), .B(rst), .Z(n3036) );
  XNOR U3448 ( .A(n3033), .B(n3032), .Z(n3034) );
  NANDN U3449 ( .A(rst), .B(n3034), .Z(n3035) );
  NAND U3450 ( .A(n3036), .B(n3035), .Z(n871) );
  NAND U3451 ( .A(c[103]), .B(rst), .Z(n3041) );
  XOR U3452 ( .A(n3038), .B(n3037), .Z(n3039) );
  NANDN U3453 ( .A(rst), .B(n3039), .Z(n3040) );
  NAND U3454 ( .A(n3041), .B(n3040), .Z(n872) );
  NAND U3455 ( .A(c[104]), .B(rst), .Z(n3046) );
  XNOR U3456 ( .A(n3043), .B(n3042), .Z(n3044) );
  NANDN U3457 ( .A(rst), .B(n3044), .Z(n3045) );
  NAND U3458 ( .A(n3046), .B(n3045), .Z(n873) );
  NAND U3459 ( .A(c[105]), .B(rst), .Z(n3051) );
  XOR U3460 ( .A(n3048), .B(n3047), .Z(n3049) );
  NANDN U3461 ( .A(rst), .B(n3049), .Z(n3050) );
  NAND U3462 ( .A(n3051), .B(n3050), .Z(n874) );
  NAND U3463 ( .A(c[106]), .B(rst), .Z(n3056) );
  XNOR U3464 ( .A(n3053), .B(n3052), .Z(n3054) );
  NANDN U3465 ( .A(rst), .B(n3054), .Z(n3055) );
  NAND U3466 ( .A(n3056), .B(n3055), .Z(n875) );
  NAND U3467 ( .A(c[107]), .B(rst), .Z(n3061) );
  XOR U3468 ( .A(n3058), .B(n3057), .Z(n3059) );
  NANDN U3469 ( .A(rst), .B(n3059), .Z(n3060) );
  NAND U3470 ( .A(n3061), .B(n3060), .Z(n876) );
  NAND U3471 ( .A(c[108]), .B(rst), .Z(n3066) );
  XNOR U3472 ( .A(n3063), .B(n3062), .Z(n3064) );
  NANDN U3473 ( .A(rst), .B(n3064), .Z(n3065) );
  NAND U3474 ( .A(n3066), .B(n3065), .Z(n877) );
  NAND U3475 ( .A(c[109]), .B(rst), .Z(n3071) );
  XOR U3476 ( .A(n3068), .B(n3067), .Z(n3069) );
  NANDN U3477 ( .A(rst), .B(n3069), .Z(n3070) );
  NAND U3478 ( .A(n3071), .B(n3070), .Z(n878) );
  NAND U3479 ( .A(c[110]), .B(rst), .Z(n3076) );
  XNOR U3480 ( .A(n3073), .B(n3072), .Z(n3074) );
  NANDN U3481 ( .A(rst), .B(n3074), .Z(n3075) );
  NAND U3482 ( .A(n3076), .B(n3075), .Z(n879) );
  NAND U3483 ( .A(c[111]), .B(rst), .Z(n3081) );
  XOR U3484 ( .A(n3078), .B(n3077), .Z(n3079) );
  NANDN U3485 ( .A(rst), .B(n3079), .Z(n3080) );
  NAND U3486 ( .A(n3081), .B(n3080), .Z(n880) );
  NAND U3487 ( .A(c[112]), .B(rst), .Z(n3086) );
  XNOR U3488 ( .A(n3083), .B(n3082), .Z(n3084) );
  NANDN U3489 ( .A(rst), .B(n3084), .Z(n3085) );
  NAND U3490 ( .A(n3086), .B(n3085), .Z(n881) );
  NAND U3491 ( .A(c[113]), .B(rst), .Z(n3091) );
  XOR U3492 ( .A(n3088), .B(n3087), .Z(n3089) );
  NANDN U3493 ( .A(rst), .B(n3089), .Z(n3090) );
  NAND U3494 ( .A(n3091), .B(n3090), .Z(n882) );
  NAND U3495 ( .A(c[114]), .B(rst), .Z(n3096) );
  XNOR U3496 ( .A(n3093), .B(n3092), .Z(n3094) );
  NANDN U3497 ( .A(rst), .B(n3094), .Z(n3095) );
  NAND U3498 ( .A(n3096), .B(n3095), .Z(n883) );
  NAND U3499 ( .A(c[115]), .B(rst), .Z(n3101) );
  XOR U3500 ( .A(n3098), .B(n3097), .Z(n3099) );
  NANDN U3501 ( .A(rst), .B(n3099), .Z(n3100) );
  NAND U3502 ( .A(n3101), .B(n3100), .Z(n884) );
  NAND U3503 ( .A(c[116]), .B(rst), .Z(n3106) );
  XNOR U3504 ( .A(n3103), .B(n3102), .Z(n3104) );
  NANDN U3505 ( .A(rst), .B(n3104), .Z(n3105) );
  NAND U3506 ( .A(n3106), .B(n3105), .Z(n885) );
  NAND U3507 ( .A(c[117]), .B(rst), .Z(n3111) );
  XOR U3508 ( .A(n3108), .B(n3107), .Z(n3109) );
  NANDN U3509 ( .A(rst), .B(n3109), .Z(n3110) );
  NAND U3510 ( .A(n3111), .B(n3110), .Z(n886) );
  NAND U3511 ( .A(c[118]), .B(rst), .Z(n3116) );
  XNOR U3512 ( .A(n3113), .B(n3112), .Z(n3114) );
  NANDN U3513 ( .A(rst), .B(n3114), .Z(n3115) );
  NAND U3514 ( .A(n3116), .B(n3115), .Z(n887) );
  NAND U3515 ( .A(c[119]), .B(rst), .Z(n3121) );
  XOR U3516 ( .A(n3118), .B(n3117), .Z(n3119) );
  NANDN U3517 ( .A(rst), .B(n3119), .Z(n3120) );
  NAND U3518 ( .A(n3121), .B(n3120), .Z(n888) );
  NAND U3519 ( .A(c[120]), .B(rst), .Z(n3126) );
  XNOR U3520 ( .A(n3123), .B(n3122), .Z(n3124) );
  NANDN U3521 ( .A(rst), .B(n3124), .Z(n3125) );
  NAND U3522 ( .A(n3126), .B(n3125), .Z(n889) );
  NAND U3523 ( .A(c[121]), .B(rst), .Z(n3131) );
  XOR U3524 ( .A(n3128), .B(n3127), .Z(n3129) );
  NANDN U3525 ( .A(rst), .B(n3129), .Z(n3130) );
  NAND U3526 ( .A(n3131), .B(n3130), .Z(n890) );
  NAND U3527 ( .A(c[122]), .B(rst), .Z(n3136) );
  XNOR U3528 ( .A(n3133), .B(n3132), .Z(n3134) );
  NANDN U3529 ( .A(rst), .B(n3134), .Z(n3135) );
  NAND U3530 ( .A(n3136), .B(n3135), .Z(n891) );
  NAND U3531 ( .A(c[123]), .B(rst), .Z(n3141) );
  XOR U3532 ( .A(n3138), .B(n3137), .Z(n3139) );
  NANDN U3533 ( .A(rst), .B(n3139), .Z(n3140) );
  NAND U3534 ( .A(n3141), .B(n3140), .Z(n892) );
  NAND U3535 ( .A(c[124]), .B(rst), .Z(n3146) );
  XNOR U3536 ( .A(n3143), .B(n3142), .Z(n3144) );
  NANDN U3537 ( .A(rst), .B(n3144), .Z(n3145) );
  NAND U3538 ( .A(n3146), .B(n3145), .Z(n893) );
  NAND U3539 ( .A(c[125]), .B(rst), .Z(n3151) );
  XNOR U3540 ( .A(n3148), .B(n3147), .Z(n3149) );
  NANDN U3541 ( .A(rst), .B(n3149), .Z(n3150) );
  NAND U3542 ( .A(n3151), .B(n3150), .Z(n894) );
  NAND U3543 ( .A(c[126]), .B(rst), .Z(n3156) );
  XNOR U3544 ( .A(n3153), .B(n3152), .Z(n3154) );
  NANDN U3545 ( .A(rst), .B(n3154), .Z(n3155) );
  NAND U3546 ( .A(n3156), .B(n3155), .Z(n895) );
  NAND U3547 ( .A(c[127]), .B(rst), .Z(n3161) );
  XNOR U3548 ( .A(n3158), .B(n3157), .Z(n3159) );
  NANDN U3549 ( .A(rst), .B(n3159), .Z(n3160) );
  NAND U3550 ( .A(n3161), .B(n3160), .Z(n896) );
  NAND U3551 ( .A(c[128]), .B(rst), .Z(n3166) );
  XOR U3552 ( .A(n3163), .B(n3162), .Z(n3164) );
  NANDN U3553 ( .A(rst), .B(n3164), .Z(n3165) );
  NAND U3554 ( .A(n3166), .B(n3165), .Z(n897) );
  NAND U3555 ( .A(c[129]), .B(rst), .Z(n3171) );
  XNOR U3556 ( .A(n3168), .B(n3167), .Z(n3169) );
  NANDN U3557 ( .A(rst), .B(n3169), .Z(n3170) );
  NAND U3558 ( .A(n3171), .B(n3170), .Z(n898) );
  NAND U3559 ( .A(c[130]), .B(rst), .Z(n3176) );
  XOR U3560 ( .A(n3173), .B(n3172), .Z(n3174) );
  NANDN U3561 ( .A(rst), .B(n3174), .Z(n3175) );
  NAND U3562 ( .A(n3176), .B(n3175), .Z(n899) );
  NAND U3563 ( .A(c[131]), .B(rst), .Z(n3181) );
  XNOR U3564 ( .A(n3178), .B(n3177), .Z(n3179) );
  NANDN U3565 ( .A(rst), .B(n3179), .Z(n3180) );
  NAND U3566 ( .A(n3181), .B(n3180), .Z(n900) );
  NAND U3567 ( .A(c[132]), .B(rst), .Z(n3186) );
  XOR U3568 ( .A(n3183), .B(n3182), .Z(n3184) );
  NANDN U3569 ( .A(rst), .B(n3184), .Z(n3185) );
  NAND U3570 ( .A(n3186), .B(n3185), .Z(n901) );
  NAND U3571 ( .A(c[133]), .B(rst), .Z(n3191) );
  XNOR U3572 ( .A(n3188), .B(n3187), .Z(n3189) );
  NANDN U3573 ( .A(rst), .B(n3189), .Z(n3190) );
  NAND U3574 ( .A(n3191), .B(n3190), .Z(n902) );
  NAND U3575 ( .A(c[134]), .B(rst), .Z(n3196) );
  XOR U3576 ( .A(n3193), .B(n3192), .Z(n3194) );
  NANDN U3577 ( .A(rst), .B(n3194), .Z(n3195) );
  NAND U3578 ( .A(n3196), .B(n3195), .Z(n903) );
  NAND U3579 ( .A(c[135]), .B(rst), .Z(n3201) );
  XNOR U3580 ( .A(n3198), .B(n3197), .Z(n3199) );
  NANDN U3581 ( .A(rst), .B(n3199), .Z(n3200) );
  NAND U3582 ( .A(n3201), .B(n3200), .Z(n904) );
  NAND U3583 ( .A(c[136]), .B(rst), .Z(n3206) );
  XOR U3584 ( .A(n3203), .B(n3202), .Z(n3204) );
  NANDN U3585 ( .A(rst), .B(n3204), .Z(n3205) );
  NAND U3586 ( .A(n3206), .B(n3205), .Z(n905) );
  NAND U3587 ( .A(c[137]), .B(rst), .Z(n3211) );
  XNOR U3588 ( .A(n3208), .B(n3207), .Z(n3209) );
  NANDN U3589 ( .A(rst), .B(n3209), .Z(n3210) );
  NAND U3590 ( .A(n3211), .B(n3210), .Z(n906) );
  NAND U3591 ( .A(c[138]), .B(rst), .Z(n3216) );
  XOR U3592 ( .A(n3213), .B(n3212), .Z(n3214) );
  NANDN U3593 ( .A(rst), .B(n3214), .Z(n3215) );
  NAND U3594 ( .A(n3216), .B(n3215), .Z(n907) );
  NAND U3595 ( .A(c[139]), .B(rst), .Z(n3221) );
  XNOR U3596 ( .A(n3218), .B(n3217), .Z(n3219) );
  NANDN U3597 ( .A(rst), .B(n3219), .Z(n3220) );
  NAND U3598 ( .A(n3221), .B(n3220), .Z(n908) );
  NAND U3599 ( .A(c[140]), .B(rst), .Z(n3226) );
  XOR U3600 ( .A(n3223), .B(n3222), .Z(n3224) );
  NANDN U3601 ( .A(rst), .B(n3224), .Z(n3225) );
  NAND U3602 ( .A(n3226), .B(n3225), .Z(n909) );
  NAND U3603 ( .A(c[141]), .B(rst), .Z(n3231) );
  XNOR U3604 ( .A(n3228), .B(n3227), .Z(n3229) );
  NANDN U3605 ( .A(rst), .B(n3229), .Z(n3230) );
  NAND U3606 ( .A(n3231), .B(n3230), .Z(n910) );
  NAND U3607 ( .A(c[142]), .B(rst), .Z(n3236) );
  XOR U3608 ( .A(n3233), .B(n3232), .Z(n3234) );
  NANDN U3609 ( .A(rst), .B(n3234), .Z(n3235) );
  NAND U3610 ( .A(n3236), .B(n3235), .Z(n911) );
  NAND U3611 ( .A(c[143]), .B(rst), .Z(n3241) );
  XNOR U3612 ( .A(n3238), .B(n3237), .Z(n3239) );
  NANDN U3613 ( .A(rst), .B(n3239), .Z(n3240) );
  NAND U3614 ( .A(n3241), .B(n3240), .Z(n912) );
  NAND U3615 ( .A(c[144]), .B(rst), .Z(n3246) );
  XOR U3616 ( .A(n3243), .B(n3242), .Z(n3244) );
  NANDN U3617 ( .A(rst), .B(n3244), .Z(n3245) );
  NAND U3618 ( .A(n3246), .B(n3245), .Z(n913) );
  NAND U3619 ( .A(c[145]), .B(rst), .Z(n3251) );
  XNOR U3620 ( .A(n3248), .B(n3247), .Z(n3249) );
  NANDN U3621 ( .A(rst), .B(n3249), .Z(n3250) );
  NAND U3622 ( .A(n3251), .B(n3250), .Z(n914) );
  NAND U3623 ( .A(c[146]), .B(rst), .Z(n3256) );
  XOR U3624 ( .A(n3253), .B(n3252), .Z(n3254) );
  NANDN U3625 ( .A(rst), .B(n3254), .Z(n3255) );
  NAND U3626 ( .A(n3256), .B(n3255), .Z(n915) );
  NAND U3627 ( .A(c[147]), .B(rst), .Z(n3261) );
  XNOR U3628 ( .A(n3258), .B(n3257), .Z(n3259) );
  NANDN U3629 ( .A(rst), .B(n3259), .Z(n3260) );
  NAND U3630 ( .A(n3261), .B(n3260), .Z(n916) );
  NAND U3631 ( .A(c[148]), .B(rst), .Z(n3266) );
  XOR U3632 ( .A(n3263), .B(n3262), .Z(n3264) );
  NANDN U3633 ( .A(rst), .B(n3264), .Z(n3265) );
  NAND U3634 ( .A(n3266), .B(n3265), .Z(n917) );
  NAND U3635 ( .A(c[149]), .B(rst), .Z(n3271) );
  XNOR U3636 ( .A(n3268), .B(n3267), .Z(n3269) );
  NANDN U3637 ( .A(rst), .B(n3269), .Z(n3270) );
  NAND U3638 ( .A(n3271), .B(n3270), .Z(n918) );
  NAND U3639 ( .A(c[150]), .B(rst), .Z(n3276) );
  XOR U3640 ( .A(n3273), .B(n3272), .Z(n3274) );
  NANDN U3641 ( .A(rst), .B(n3274), .Z(n3275) );
  NAND U3642 ( .A(n3276), .B(n3275), .Z(n919) );
  NAND U3643 ( .A(c[151]), .B(rst), .Z(n3281) );
  XNOR U3644 ( .A(n3278), .B(n3277), .Z(n3279) );
  NANDN U3645 ( .A(rst), .B(n3279), .Z(n3280) );
  NAND U3646 ( .A(n3281), .B(n3280), .Z(n920) );
  NAND U3647 ( .A(c[152]), .B(rst), .Z(n3286) );
  XNOR U3648 ( .A(n3283), .B(n3282), .Z(n3284) );
  NANDN U3649 ( .A(rst), .B(n3284), .Z(n3285) );
  NAND U3650 ( .A(n3286), .B(n3285), .Z(n921) );
  NAND U3651 ( .A(c[153]), .B(rst), .Z(n3291) );
  XNOR U3652 ( .A(n3288), .B(n3287), .Z(n3289) );
  NANDN U3653 ( .A(rst), .B(n3289), .Z(n3290) );
  NAND U3654 ( .A(n3291), .B(n3290), .Z(n922) );
  NAND U3655 ( .A(c[154]), .B(rst), .Z(n3296) );
  XNOR U3656 ( .A(n3293), .B(n3292), .Z(n3294) );
  NANDN U3657 ( .A(rst), .B(n3294), .Z(n3295) );
  NAND U3658 ( .A(n3296), .B(n3295), .Z(n923) );
  NAND U3659 ( .A(c[155]), .B(rst), .Z(n3301) );
  XOR U3660 ( .A(n3298), .B(n3297), .Z(n3299) );
  NANDN U3661 ( .A(rst), .B(n3299), .Z(n3300) );
  NAND U3662 ( .A(n3301), .B(n3300), .Z(n924) );
  NAND U3663 ( .A(c[156]), .B(rst), .Z(n3306) );
  XNOR U3664 ( .A(n3303), .B(n3302), .Z(n3304) );
  NANDN U3665 ( .A(rst), .B(n3304), .Z(n3305) );
  NAND U3666 ( .A(n3306), .B(n3305), .Z(n925) );
  NAND U3667 ( .A(c[157]), .B(rst), .Z(n3311) );
  XNOR U3668 ( .A(n3308), .B(n3307), .Z(n3309) );
  NANDN U3669 ( .A(rst), .B(n3309), .Z(n3310) );
  NAND U3670 ( .A(n3311), .B(n3310), .Z(n926) );
  NAND U3671 ( .A(c[158]), .B(rst), .Z(n3316) );
  XNOR U3672 ( .A(n3313), .B(n3312), .Z(n3314) );
  NANDN U3673 ( .A(rst), .B(n3314), .Z(n3315) );
  NAND U3674 ( .A(n3316), .B(n3315), .Z(n927) );
  NAND U3675 ( .A(c[159]), .B(rst), .Z(n3321) );
  XNOR U3676 ( .A(n3318), .B(n3317), .Z(n3319) );
  NANDN U3677 ( .A(rst), .B(n3319), .Z(n3320) );
  NAND U3678 ( .A(n3321), .B(n3320), .Z(n928) );
  NAND U3679 ( .A(c[160]), .B(rst), .Z(n3326) );
  XOR U3680 ( .A(n3323), .B(n3322), .Z(n3324) );
  NANDN U3681 ( .A(rst), .B(n3324), .Z(n3325) );
  NAND U3682 ( .A(n3326), .B(n3325), .Z(n929) );
  NAND U3683 ( .A(c[161]), .B(rst), .Z(n3331) );
  XNOR U3684 ( .A(n3328), .B(n3327), .Z(n3329) );
  NANDN U3685 ( .A(rst), .B(n3329), .Z(n3330) );
  NAND U3686 ( .A(n3331), .B(n3330), .Z(n930) );
  NAND U3687 ( .A(c[162]), .B(rst), .Z(n3336) );
  XOR U3688 ( .A(n3333), .B(n3332), .Z(n3334) );
  NANDN U3689 ( .A(rst), .B(n3334), .Z(n3335) );
  NAND U3690 ( .A(n3336), .B(n3335), .Z(n931) );
  NAND U3691 ( .A(c[163]), .B(rst), .Z(n3341) );
  XNOR U3692 ( .A(n3338), .B(n3337), .Z(n3339) );
  NANDN U3693 ( .A(rst), .B(n3339), .Z(n3340) );
  NAND U3694 ( .A(n3341), .B(n3340), .Z(n932) );
  NAND U3695 ( .A(c[164]), .B(rst), .Z(n3346) );
  XOR U3696 ( .A(n3343), .B(n3342), .Z(n3344) );
  NANDN U3697 ( .A(rst), .B(n3344), .Z(n3345) );
  NAND U3698 ( .A(n3346), .B(n3345), .Z(n933) );
  NAND U3699 ( .A(c[165]), .B(rst), .Z(n3351) );
  XNOR U3700 ( .A(n3348), .B(n3347), .Z(n3349) );
  NANDN U3701 ( .A(rst), .B(n3349), .Z(n3350) );
  NAND U3702 ( .A(n3351), .B(n3350), .Z(n934) );
  NAND U3703 ( .A(c[166]), .B(rst), .Z(n3356) );
  XNOR U3704 ( .A(n3353), .B(n3352), .Z(n3354) );
  NANDN U3705 ( .A(rst), .B(n3354), .Z(n3355) );
  NAND U3706 ( .A(n3356), .B(n3355), .Z(n935) );
  NAND U3707 ( .A(c[167]), .B(rst), .Z(n3361) );
  XNOR U3708 ( .A(n3358), .B(n3357), .Z(n3359) );
  NANDN U3709 ( .A(rst), .B(n3359), .Z(n3360) );
  NAND U3710 ( .A(n3361), .B(n3360), .Z(n936) );
  NAND U3711 ( .A(c[168]), .B(rst), .Z(n3366) );
  XNOR U3712 ( .A(n3363), .B(n3362), .Z(n3364) );
  NANDN U3713 ( .A(rst), .B(n3364), .Z(n3365) );
  NAND U3714 ( .A(n3366), .B(n3365), .Z(n937) );
  NAND U3715 ( .A(c[169]), .B(rst), .Z(n3371) );
  XOR U3716 ( .A(n3368), .B(n3367), .Z(n3369) );
  NANDN U3717 ( .A(rst), .B(n3369), .Z(n3370) );
  NAND U3718 ( .A(n3371), .B(n3370), .Z(n938) );
  NAND U3719 ( .A(c[170]), .B(rst), .Z(n3376) );
  XNOR U3720 ( .A(n3373), .B(n3372), .Z(n3374) );
  NANDN U3721 ( .A(rst), .B(n3374), .Z(n3375) );
  NAND U3722 ( .A(n3376), .B(n3375), .Z(n939) );
  NAND U3723 ( .A(c[171]), .B(rst), .Z(n3381) );
  XOR U3724 ( .A(n3378), .B(n3377), .Z(n3379) );
  NANDN U3725 ( .A(rst), .B(n3379), .Z(n3380) );
  NAND U3726 ( .A(n3381), .B(n3380), .Z(n940) );
  NAND U3727 ( .A(c[172]), .B(rst), .Z(n3386) );
  XNOR U3728 ( .A(n3383), .B(n3382), .Z(n3384) );
  NANDN U3729 ( .A(rst), .B(n3384), .Z(n3385) );
  NAND U3730 ( .A(n3386), .B(n3385), .Z(n941) );
  NAND U3731 ( .A(c[173]), .B(rst), .Z(n3391) );
  XOR U3732 ( .A(n3388), .B(n3387), .Z(n3389) );
  NANDN U3733 ( .A(rst), .B(n3389), .Z(n3390) );
  NAND U3734 ( .A(n3391), .B(n3390), .Z(n942) );
  NAND U3735 ( .A(c[174]), .B(rst), .Z(n3396) );
  XNOR U3736 ( .A(n3393), .B(n3392), .Z(n3394) );
  NANDN U3737 ( .A(rst), .B(n3394), .Z(n3395) );
  NAND U3738 ( .A(n3396), .B(n3395), .Z(n943) );
  NAND U3739 ( .A(c[175]), .B(rst), .Z(n3401) );
  XOR U3740 ( .A(n3398), .B(n3397), .Z(n3399) );
  NANDN U3741 ( .A(rst), .B(n3399), .Z(n3400) );
  NAND U3742 ( .A(n3401), .B(n3400), .Z(n944) );
  NAND U3743 ( .A(c[176]), .B(rst), .Z(n3406) );
  XNOR U3744 ( .A(n3403), .B(n3402), .Z(n3404) );
  NANDN U3745 ( .A(rst), .B(n3404), .Z(n3405) );
  NAND U3746 ( .A(n3406), .B(n3405), .Z(n945) );
  NAND U3747 ( .A(c[177]), .B(rst), .Z(n3411) );
  XOR U3748 ( .A(n3408), .B(n3407), .Z(n3409) );
  NANDN U3749 ( .A(rst), .B(n3409), .Z(n3410) );
  NAND U3750 ( .A(n3411), .B(n3410), .Z(n946) );
  NAND U3751 ( .A(c[178]), .B(rst), .Z(n3416) );
  XNOR U3752 ( .A(n3413), .B(n3412), .Z(n3414) );
  NANDN U3753 ( .A(rst), .B(n3414), .Z(n3415) );
  NAND U3754 ( .A(n3416), .B(n3415), .Z(n947) );
  NAND U3755 ( .A(c[179]), .B(rst), .Z(n3421) );
  XOR U3756 ( .A(n3418), .B(n3417), .Z(n3419) );
  NANDN U3757 ( .A(rst), .B(n3419), .Z(n3420) );
  NAND U3758 ( .A(n3421), .B(n3420), .Z(n948) );
  NAND U3759 ( .A(c[180]), .B(rst), .Z(n3426) );
  XNOR U3760 ( .A(n3423), .B(n3422), .Z(n3424) );
  NANDN U3761 ( .A(rst), .B(n3424), .Z(n3425) );
  NAND U3762 ( .A(n3426), .B(n3425), .Z(n949) );
  NAND U3763 ( .A(c[181]), .B(rst), .Z(n3431) );
  XOR U3764 ( .A(n3428), .B(n3427), .Z(n3429) );
  NANDN U3765 ( .A(rst), .B(n3429), .Z(n3430) );
  NAND U3766 ( .A(n3431), .B(n3430), .Z(n950) );
  NAND U3767 ( .A(c[182]), .B(rst), .Z(n3436) );
  XNOR U3768 ( .A(n3433), .B(n3432), .Z(n3434) );
  NANDN U3769 ( .A(rst), .B(n3434), .Z(n3435) );
  NAND U3770 ( .A(n3436), .B(n3435), .Z(n951) );
  NAND U3771 ( .A(c[183]), .B(rst), .Z(n3441) );
  XOR U3772 ( .A(n3438), .B(n3437), .Z(n3439) );
  NANDN U3773 ( .A(rst), .B(n3439), .Z(n3440) );
  NAND U3774 ( .A(n3441), .B(n3440), .Z(n952) );
  NAND U3775 ( .A(c[184]), .B(rst), .Z(n3446) );
  XNOR U3776 ( .A(n3443), .B(n3442), .Z(n3444) );
  NANDN U3777 ( .A(rst), .B(n3444), .Z(n3445) );
  NAND U3778 ( .A(n3446), .B(n3445), .Z(n953) );
  NAND U3779 ( .A(c[185]), .B(rst), .Z(n3451) );
  XNOR U3780 ( .A(n3448), .B(n3447), .Z(n3449) );
  NANDN U3781 ( .A(rst), .B(n3449), .Z(n3450) );
  NAND U3782 ( .A(n3451), .B(n3450), .Z(n954) );
  NAND U3783 ( .A(c[186]), .B(rst), .Z(n3456) );
  XNOR U3784 ( .A(n3453), .B(n3452), .Z(n3454) );
  NANDN U3785 ( .A(rst), .B(n3454), .Z(n3455) );
  NAND U3786 ( .A(n3456), .B(n3455), .Z(n955) );
  NAND U3787 ( .A(c[187]), .B(rst), .Z(n3461) );
  XNOR U3788 ( .A(n3458), .B(n3457), .Z(n3459) );
  NANDN U3789 ( .A(rst), .B(n3459), .Z(n3460) );
  NAND U3790 ( .A(n3461), .B(n3460), .Z(n956) );
  NAND U3791 ( .A(c[188]), .B(rst), .Z(n3466) );
  XOR U3792 ( .A(n3463), .B(n3462), .Z(n3464) );
  NANDN U3793 ( .A(rst), .B(n3464), .Z(n3465) );
  NAND U3794 ( .A(n3466), .B(n3465), .Z(n957) );
  NAND U3795 ( .A(c[189]), .B(rst), .Z(n3471) );
  XNOR U3796 ( .A(n3468), .B(n3467), .Z(n3469) );
  NANDN U3797 ( .A(rst), .B(n3469), .Z(n3470) );
  NAND U3798 ( .A(n3471), .B(n3470), .Z(n958) );
  NAND U3799 ( .A(c[190]), .B(rst), .Z(n3476) );
  XNOR U3800 ( .A(n3473), .B(n3472), .Z(n3474) );
  NANDN U3801 ( .A(rst), .B(n3474), .Z(n3475) );
  NAND U3802 ( .A(n3476), .B(n3475), .Z(n959) );
  NAND U3803 ( .A(c[191]), .B(rst), .Z(n3481) );
  XNOR U3804 ( .A(n3478), .B(n3477), .Z(n3479) );
  NANDN U3805 ( .A(rst), .B(n3479), .Z(n3480) );
  NAND U3806 ( .A(n3481), .B(n3480), .Z(n960) );
  NAND U3807 ( .A(c[192]), .B(rst), .Z(n3486) );
  XNOR U3808 ( .A(n3483), .B(n3482), .Z(n3484) );
  NANDN U3809 ( .A(rst), .B(n3484), .Z(n3485) );
  NAND U3810 ( .A(n3486), .B(n3485), .Z(n961) );
  NAND U3811 ( .A(c[193]), .B(rst), .Z(n3491) );
  XOR U3812 ( .A(n3488), .B(n3487), .Z(n3489) );
  NANDN U3813 ( .A(rst), .B(n3489), .Z(n3490) );
  NAND U3814 ( .A(n3491), .B(n3490), .Z(n962) );
  NAND U3815 ( .A(c[194]), .B(rst), .Z(n3496) );
  XNOR U3816 ( .A(n3493), .B(n3492), .Z(n3494) );
  NANDN U3817 ( .A(rst), .B(n3494), .Z(n3495) );
  NAND U3818 ( .A(n3496), .B(n3495), .Z(n963) );
  NAND U3819 ( .A(c[195]), .B(rst), .Z(n3501) );
  XOR U3820 ( .A(n3498), .B(n3497), .Z(n3499) );
  NANDN U3821 ( .A(rst), .B(n3499), .Z(n3500) );
  NAND U3822 ( .A(n3501), .B(n3500), .Z(n964) );
  NAND U3823 ( .A(c[196]), .B(rst), .Z(n3506) );
  XNOR U3824 ( .A(n3503), .B(n3502), .Z(n3504) );
  NANDN U3825 ( .A(rst), .B(n3504), .Z(n3505) );
  NAND U3826 ( .A(n3506), .B(n3505), .Z(n965) );
  NAND U3827 ( .A(c[197]), .B(rst), .Z(n3511) );
  XOR U3828 ( .A(n3508), .B(n3507), .Z(n3509) );
  NANDN U3829 ( .A(rst), .B(n3509), .Z(n3510) );
  NAND U3830 ( .A(n3511), .B(n3510), .Z(n966) );
  NAND U3831 ( .A(c[198]), .B(rst), .Z(n3516) );
  XNOR U3832 ( .A(n3513), .B(n3512), .Z(n3514) );
  NANDN U3833 ( .A(rst), .B(n3514), .Z(n3515) );
  NAND U3834 ( .A(n3516), .B(n3515), .Z(n967) );
  NAND U3835 ( .A(c[199]), .B(rst), .Z(n3521) );
  XOR U3836 ( .A(n3518), .B(n3517), .Z(n3519) );
  NANDN U3837 ( .A(rst), .B(n3519), .Z(n3520) );
  NAND U3838 ( .A(n3521), .B(n3520), .Z(n968) );
  NAND U3839 ( .A(c[200]), .B(rst), .Z(n3526) );
  XNOR U3840 ( .A(n3523), .B(n3522), .Z(n3524) );
  NANDN U3841 ( .A(rst), .B(n3524), .Z(n3525) );
  NAND U3842 ( .A(n3526), .B(n3525), .Z(n969) );
  NAND U3843 ( .A(c[201]), .B(rst), .Z(n3531) );
  XNOR U3844 ( .A(n3528), .B(n3527), .Z(n3529) );
  NANDN U3845 ( .A(rst), .B(n3529), .Z(n3530) );
  NAND U3846 ( .A(n3531), .B(n3530), .Z(n970) );
  NAND U3847 ( .A(c[202]), .B(rst), .Z(n3536) );
  XNOR U3848 ( .A(n3533), .B(n3532), .Z(n3534) );
  NANDN U3849 ( .A(rst), .B(n3534), .Z(n3535) );
  NAND U3850 ( .A(n3536), .B(n3535), .Z(n971) );
  NAND U3851 ( .A(c[203]), .B(rst), .Z(n3541) );
  XNOR U3852 ( .A(n3538), .B(n3537), .Z(n3539) );
  NANDN U3853 ( .A(rst), .B(n3539), .Z(n3540) );
  NAND U3854 ( .A(n3541), .B(n3540), .Z(n972) );
  NAND U3855 ( .A(c[204]), .B(rst), .Z(n3546) );
  XOR U3856 ( .A(n3543), .B(n3542), .Z(n3544) );
  NANDN U3857 ( .A(rst), .B(n3544), .Z(n3545) );
  NAND U3858 ( .A(n3546), .B(n3545), .Z(n973) );
  NAND U3859 ( .A(c[205]), .B(rst), .Z(n3551) );
  XNOR U3860 ( .A(n3548), .B(n3547), .Z(n3549) );
  NANDN U3861 ( .A(rst), .B(n3549), .Z(n3550) );
  NAND U3862 ( .A(n3551), .B(n3550), .Z(n974) );
  NAND U3863 ( .A(c[206]), .B(rst), .Z(n3556) );
  XOR U3864 ( .A(n3553), .B(n3552), .Z(n3554) );
  NANDN U3865 ( .A(rst), .B(n3554), .Z(n3555) );
  NAND U3866 ( .A(n3556), .B(n3555), .Z(n975) );
  NAND U3867 ( .A(c[207]), .B(rst), .Z(n3561) );
  XNOR U3868 ( .A(n3558), .B(n3557), .Z(n3559) );
  NANDN U3869 ( .A(rst), .B(n3559), .Z(n3560) );
  NAND U3870 ( .A(n3561), .B(n3560), .Z(n976) );
  NAND U3871 ( .A(c[208]), .B(rst), .Z(n3566) );
  XOR U3872 ( .A(n3563), .B(n3562), .Z(n3564) );
  NANDN U3873 ( .A(rst), .B(n3564), .Z(n3565) );
  NAND U3874 ( .A(n3566), .B(n3565), .Z(n977) );
  NAND U3875 ( .A(c[209]), .B(rst), .Z(n3571) );
  XNOR U3876 ( .A(n3568), .B(n3567), .Z(n3569) );
  NANDN U3877 ( .A(rst), .B(n3569), .Z(n3570) );
  NAND U3878 ( .A(n3571), .B(n3570), .Z(n978) );
  NAND U3879 ( .A(c[210]), .B(rst), .Z(n3576) );
  XOR U3880 ( .A(n3573), .B(n3572), .Z(n3574) );
  NANDN U3881 ( .A(rst), .B(n3574), .Z(n3575) );
  NAND U3882 ( .A(n3576), .B(n3575), .Z(n979) );
  NAND U3883 ( .A(c[211]), .B(rst), .Z(n3581) );
  XNOR U3884 ( .A(n3578), .B(n3577), .Z(n3579) );
  NANDN U3885 ( .A(rst), .B(n3579), .Z(n3580) );
  NAND U3886 ( .A(n3581), .B(n3580), .Z(n980) );
  NAND U3887 ( .A(c[212]), .B(rst), .Z(n3586) );
  XOR U3888 ( .A(n3583), .B(n3582), .Z(n3584) );
  NANDN U3889 ( .A(rst), .B(n3584), .Z(n3585) );
  NAND U3890 ( .A(n3586), .B(n3585), .Z(n981) );
  NAND U3891 ( .A(c[213]), .B(rst), .Z(n3591) );
  XNOR U3892 ( .A(n3588), .B(n3587), .Z(n3589) );
  NANDN U3893 ( .A(rst), .B(n3589), .Z(n3590) );
  NAND U3894 ( .A(n3591), .B(n3590), .Z(n982) );
  NAND U3895 ( .A(c[214]), .B(rst), .Z(n3596) );
  XOR U3896 ( .A(n3593), .B(n3592), .Z(n3594) );
  NANDN U3897 ( .A(rst), .B(n3594), .Z(n3595) );
  NAND U3898 ( .A(n3596), .B(n3595), .Z(n983) );
  NAND U3899 ( .A(c[215]), .B(rst), .Z(n3601) );
  XNOR U3900 ( .A(n3598), .B(n3597), .Z(n3599) );
  NANDN U3901 ( .A(rst), .B(n3599), .Z(n3600) );
  NAND U3902 ( .A(n3601), .B(n3600), .Z(n984) );
  NAND U3903 ( .A(c[216]), .B(rst), .Z(n3606) );
  XOR U3904 ( .A(n3603), .B(n3602), .Z(n3604) );
  NANDN U3905 ( .A(rst), .B(n3604), .Z(n3605) );
  NAND U3906 ( .A(n3606), .B(n3605), .Z(n985) );
  NAND U3907 ( .A(c[217]), .B(rst), .Z(n3611) );
  XNOR U3908 ( .A(n3608), .B(n3607), .Z(n3609) );
  NANDN U3909 ( .A(rst), .B(n3609), .Z(n3610) );
  NAND U3910 ( .A(n3611), .B(n3610), .Z(n986) );
  NAND U3911 ( .A(c[218]), .B(rst), .Z(n3616) );
  XNOR U3912 ( .A(n3613), .B(n3612), .Z(n3614) );
  NANDN U3913 ( .A(rst), .B(n3614), .Z(n3615) );
  NAND U3914 ( .A(n3616), .B(n3615), .Z(n987) );
  NAND U3915 ( .A(c[219]), .B(rst), .Z(n3621) );
  XNOR U3916 ( .A(n3618), .B(n3617), .Z(n3619) );
  NANDN U3917 ( .A(rst), .B(n3619), .Z(n3620) );
  NAND U3918 ( .A(n3621), .B(n3620), .Z(n988) );
  NAND U3919 ( .A(c[220]), .B(rst), .Z(n3626) );
  XNOR U3920 ( .A(n3623), .B(n3622), .Z(n3624) );
  NANDN U3921 ( .A(rst), .B(n3624), .Z(n3625) );
  NAND U3922 ( .A(n3626), .B(n3625), .Z(n989) );
  NAND U3923 ( .A(c[221]), .B(rst), .Z(n3631) );
  XOR U3924 ( .A(n3628), .B(n3627), .Z(n3629) );
  NANDN U3925 ( .A(rst), .B(n3629), .Z(n3630) );
  NAND U3926 ( .A(n3631), .B(n3630), .Z(n990) );
  NAND U3927 ( .A(c[222]), .B(rst), .Z(n3636) );
  XNOR U3928 ( .A(n3633), .B(n3632), .Z(n3634) );
  NANDN U3929 ( .A(rst), .B(n3634), .Z(n3635) );
  NAND U3930 ( .A(n3636), .B(n3635), .Z(n991) );
  NAND U3931 ( .A(c[223]), .B(rst), .Z(n3641) );
  XOR U3932 ( .A(n3638), .B(n3637), .Z(n3639) );
  NANDN U3933 ( .A(rst), .B(n3639), .Z(n3640) );
  NAND U3934 ( .A(n3641), .B(n3640), .Z(n992) );
  NAND U3935 ( .A(c[224]), .B(rst), .Z(n3646) );
  XNOR U3936 ( .A(n3643), .B(n3642), .Z(n3644) );
  NANDN U3937 ( .A(rst), .B(n3644), .Z(n3645) );
  NAND U3938 ( .A(n3646), .B(n3645), .Z(n993) );
  NAND U3939 ( .A(c[225]), .B(rst), .Z(n3651) );
  XOR U3940 ( .A(n3648), .B(n3647), .Z(n3649) );
  NANDN U3941 ( .A(rst), .B(n3649), .Z(n3650) );
  NAND U3942 ( .A(n3651), .B(n3650), .Z(n994) );
  NAND U3943 ( .A(c[226]), .B(rst), .Z(n3656) );
  XNOR U3944 ( .A(n3653), .B(n3652), .Z(n3654) );
  NANDN U3945 ( .A(rst), .B(n3654), .Z(n3655) );
  NAND U3946 ( .A(n3656), .B(n3655), .Z(n995) );
  NAND U3947 ( .A(c[227]), .B(rst), .Z(n3661) );
  XOR U3948 ( .A(n3658), .B(n3657), .Z(n3659) );
  NANDN U3949 ( .A(rst), .B(n3659), .Z(n3660) );
  NAND U3950 ( .A(n3661), .B(n3660), .Z(n996) );
  NAND U3951 ( .A(c[228]), .B(rst), .Z(n3666) );
  XNOR U3952 ( .A(n3663), .B(n3662), .Z(n3664) );
  NANDN U3953 ( .A(rst), .B(n3664), .Z(n3665) );
  NAND U3954 ( .A(n3666), .B(n3665), .Z(n997) );
  NAND U3955 ( .A(c[229]), .B(rst), .Z(n3671) );
  XOR U3956 ( .A(n3668), .B(n3667), .Z(n3669) );
  NANDN U3957 ( .A(rst), .B(n3669), .Z(n3670) );
  NAND U3958 ( .A(n3671), .B(n3670), .Z(n998) );
  NAND U3959 ( .A(c[230]), .B(rst), .Z(n3676) );
  XNOR U3960 ( .A(n3673), .B(n3672), .Z(n3674) );
  NANDN U3961 ( .A(rst), .B(n3674), .Z(n3675) );
  NAND U3962 ( .A(n3676), .B(n3675), .Z(n999) );
  NAND U3963 ( .A(c[231]), .B(rst), .Z(n3681) );
  XOR U3964 ( .A(n3678), .B(n3677), .Z(n3679) );
  NANDN U3965 ( .A(rst), .B(n3679), .Z(n3680) );
  NAND U3966 ( .A(n3681), .B(n3680), .Z(n1000) );
  NAND U3967 ( .A(c[232]), .B(rst), .Z(n3686) );
  XNOR U3968 ( .A(n3683), .B(n3682), .Z(n3684) );
  NANDN U3969 ( .A(rst), .B(n3684), .Z(n3685) );
  NAND U3970 ( .A(n3686), .B(n3685), .Z(n1001) );
  NAND U3971 ( .A(c[233]), .B(rst), .Z(n3691) );
  XOR U3972 ( .A(n3688), .B(n3687), .Z(n3689) );
  NANDN U3973 ( .A(rst), .B(n3689), .Z(n3690) );
  NAND U3974 ( .A(n3691), .B(n3690), .Z(n1002) );
  NAND U3975 ( .A(c[234]), .B(rst), .Z(n3696) );
  XNOR U3976 ( .A(n3693), .B(n3692), .Z(n3694) );
  NANDN U3977 ( .A(rst), .B(n3694), .Z(n3695) );
  NAND U3978 ( .A(n3696), .B(n3695), .Z(n1003) );
  NAND U3979 ( .A(c[235]), .B(rst), .Z(n3701) );
  XOR U3980 ( .A(n3698), .B(n3697), .Z(n3699) );
  NANDN U3981 ( .A(rst), .B(n3699), .Z(n3700) );
  NAND U3982 ( .A(n3701), .B(n3700), .Z(n1004) );
  NAND U3983 ( .A(c[236]), .B(rst), .Z(n3706) );
  XNOR U3984 ( .A(n3703), .B(n3702), .Z(n3704) );
  NANDN U3985 ( .A(rst), .B(n3704), .Z(n3705) );
  NAND U3986 ( .A(n3706), .B(n3705), .Z(n1005) );
  NAND U3987 ( .A(c[237]), .B(rst), .Z(n3711) );
  XNOR U3988 ( .A(n3708), .B(n3707), .Z(n3709) );
  NANDN U3989 ( .A(rst), .B(n3709), .Z(n3710) );
  NAND U3990 ( .A(n3711), .B(n3710), .Z(n1006) );
  NAND U3991 ( .A(c[238]), .B(rst), .Z(n3716) );
  XNOR U3992 ( .A(n3713), .B(n3712), .Z(n3714) );
  NANDN U3993 ( .A(rst), .B(n3714), .Z(n3715) );
  NAND U3994 ( .A(n3716), .B(n3715), .Z(n1007) );
  NAND U3995 ( .A(c[239]), .B(rst), .Z(n3721) );
  XNOR U3996 ( .A(n3718), .B(n3717), .Z(n3719) );
  NANDN U3997 ( .A(rst), .B(n3719), .Z(n3720) );
  NAND U3998 ( .A(n3721), .B(n3720), .Z(n1008) );
  NAND U3999 ( .A(c[240]), .B(rst), .Z(n3726) );
  XOR U4000 ( .A(n3723), .B(n3722), .Z(n3724) );
  NANDN U4001 ( .A(rst), .B(n3724), .Z(n3725) );
  NAND U4002 ( .A(n3726), .B(n3725), .Z(n1009) );
  NAND U4003 ( .A(c[241]), .B(rst), .Z(n3731) );
  XNOR U4004 ( .A(n3728), .B(n3727), .Z(n3729) );
  NANDN U4005 ( .A(rst), .B(n3729), .Z(n3730) );
  NAND U4006 ( .A(n3731), .B(n3730), .Z(n1010) );
  NAND U4007 ( .A(c[242]), .B(rst), .Z(n3736) );
  XOR U4008 ( .A(n3733), .B(n3732), .Z(n3734) );
  NANDN U4009 ( .A(rst), .B(n3734), .Z(n3735) );
  NAND U4010 ( .A(n3736), .B(n3735), .Z(n1011) );
  NAND U4011 ( .A(c[243]), .B(rst), .Z(n3741) );
  XNOR U4012 ( .A(n3738), .B(n3737), .Z(n3739) );
  NANDN U4013 ( .A(rst), .B(n3739), .Z(n3740) );
  NAND U4014 ( .A(n3741), .B(n3740), .Z(n1012) );
  NAND U4015 ( .A(c[244]), .B(rst), .Z(n3746) );
  XOR U4016 ( .A(n3743), .B(n3742), .Z(n3744) );
  NANDN U4017 ( .A(rst), .B(n3744), .Z(n3745) );
  NAND U4018 ( .A(n3746), .B(n3745), .Z(n1013) );
  NAND U4019 ( .A(c[245]), .B(rst), .Z(n3751) );
  XNOR U4020 ( .A(n3748), .B(n3747), .Z(n3749) );
  NANDN U4021 ( .A(rst), .B(n3749), .Z(n3750) );
  NAND U4022 ( .A(n3751), .B(n3750), .Z(n1014) );
  NAND U4023 ( .A(c[246]), .B(rst), .Z(n3756) );
  XOR U4024 ( .A(n3753), .B(n3752), .Z(n3754) );
  NANDN U4025 ( .A(rst), .B(n3754), .Z(n3755) );
  NAND U4026 ( .A(n3756), .B(n3755), .Z(n1015) );
  NAND U4027 ( .A(c[247]), .B(rst), .Z(n3761) );
  XNOR U4028 ( .A(n3758), .B(n3757), .Z(n3759) );
  NANDN U4029 ( .A(rst), .B(n3759), .Z(n3760) );
  NAND U4030 ( .A(n3761), .B(n3760), .Z(n1016) );
  NAND U4031 ( .A(c[248]), .B(rst), .Z(n3766) );
  XOR U4032 ( .A(n3763), .B(n3762), .Z(n3764) );
  NANDN U4033 ( .A(rst), .B(n3764), .Z(n3765) );
  NAND U4034 ( .A(n3766), .B(n3765), .Z(n1017) );
  NAND U4035 ( .A(c[249]), .B(rst), .Z(n3771) );
  XNOR U4036 ( .A(n3768), .B(n3767), .Z(n3769) );
  NANDN U4037 ( .A(rst), .B(n3769), .Z(n3770) );
  NAND U4038 ( .A(n3771), .B(n3770), .Z(n1018) );
  NAND U4039 ( .A(c[250]), .B(rst), .Z(n3776) );
  XOR U4040 ( .A(n3773), .B(n3772), .Z(n3774) );
  NANDN U4041 ( .A(rst), .B(n3774), .Z(n3775) );
  NAND U4042 ( .A(n3776), .B(n3775), .Z(n1019) );
  NAND U4043 ( .A(c[251]), .B(rst), .Z(n3781) );
  XNOR U4044 ( .A(n3778), .B(n3777), .Z(n3779) );
  NANDN U4045 ( .A(rst), .B(n3779), .Z(n3780) );
  NAND U4046 ( .A(n3781), .B(n3780), .Z(n1020) );
  NAND U4047 ( .A(c[252]), .B(rst), .Z(n3786) );
  XOR U4048 ( .A(n3783), .B(n3782), .Z(n3784) );
  NANDN U4049 ( .A(rst), .B(n3784), .Z(n3785) );
  NAND U4050 ( .A(n3786), .B(n3785), .Z(n1021) );
  NAND U4051 ( .A(c[253]), .B(rst), .Z(n3791) );
  XNOR U4052 ( .A(n3788), .B(n3787), .Z(n3789) );
  NANDN U4053 ( .A(rst), .B(n3789), .Z(n3790) );
  NAND U4054 ( .A(n3791), .B(n3790), .Z(n1022) );
  NAND U4055 ( .A(c[254]), .B(rst), .Z(n3796) );
  XNOR U4056 ( .A(n3793), .B(n3792), .Z(n3794) );
  NANDN U4057 ( .A(rst), .B(n3794), .Z(n3795) );
  NAND U4058 ( .A(n3796), .B(n3795), .Z(n1023) );
  NAND U4059 ( .A(c[255]), .B(rst), .Z(n3801) );
  XNOR U4060 ( .A(n3798), .B(n3797), .Z(n3799) );
  NANDN U4061 ( .A(rst), .B(n3799), .Z(n3800) );
  NAND U4062 ( .A(n3801), .B(n3800), .Z(n1024) );
endmodule

