
module FA_6945 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_6946 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6947 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6948 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6949 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6950 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6951 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6952 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6953 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6954 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6955 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6956 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6957 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6958 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6959 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6960 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6961 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6962 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6963 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6964 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6965 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6966 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6967 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6968 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6969 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6970 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6971 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6972 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6973 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6974 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6975 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_221 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;


  FA_6975 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_6974 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_6973 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_6972 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_6971 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_6970 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_6969 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_6968 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_6967 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_6966 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_6965 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_6964 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_6963 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_6962 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_6961 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_6960 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_6959 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_6958 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_6957 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_6956 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_6955 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_6954 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_6953 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_6952 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_6951 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_6950 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_6949 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_6948 \FAINST[28].FA_  ( .A(1'b0), .B(B[28]), .CI(1'b0), .S(S[28]) );
  FA_6947 \FAINST[29].FA_  ( .A(1'b0), .B(B[29]), .CI(1'b0), .S(S[29]) );
  FA_6946 \FAINST[30].FA_  ( .A(1'b0), .B(B[30]), .CI(1'b0), .S(S[30]) );
  FA_6945 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(1'b0), .S(S[31]) );
endmodule


module FA_6977 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_6978 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_6979 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6980 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6981 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6982 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6983 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6984 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6985 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6986 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6987 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6988 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6989 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6990 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6991 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6992 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6993 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6994 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6995 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6996 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6997 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6998 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6999 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7000 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7001 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7002 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7003 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7004 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7005 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7006 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7007 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_222 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;
  wire   \C[31] ;

  FA_7007 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_7006 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_7005 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_7004 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_7003 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_7002 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_7001 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_7000 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_6999 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_6998 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_6997 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_6996 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_6995 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_6994 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_6993 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_6992 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_6991 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_6990 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_6989 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_6988 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_6987 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_6986 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_6985 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_6984 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_6983 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_6982 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_6981 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_6980 \FAINST[28].FA_  ( .A(1'b0), .B(B[28]), .CI(1'b0), .S(S[28]) );
  FA_6979 \FAINST[29].FA_  ( .A(1'b0), .B(B[29]), .CI(1'b0), .S(S[29]) );
  FA_6978 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(1'b0), .S(S[30]), .CO(
        \C[31] ) );
  FA_6977 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(\C[31] ), .S(S[31]) );
endmodule


module FA_7009 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_7010 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7011 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_7012 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7013 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7014 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7015 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7016 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7017 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7018 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7019 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7020 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7021 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7022 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7023 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7024 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7025 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7026 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7027 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7028 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7029 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7030 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7031 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7032 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7033 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7034 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7035 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7036 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7037 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7038 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7039 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_223 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_7039 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_7038 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_7037 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_7036 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_7035 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_7034 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_7033 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_7032 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_7031 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_7030 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_7029 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_7028 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_7027 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_7026 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_7025 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_7024 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_7023 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_7022 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_7021 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_7020 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_7019 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_7018 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_7017 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_7016 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_7015 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_7014 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_7013 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_7012 \FAINST[28].FA_  ( .A(1'b0), .B(B[28]), .CI(1'b0), .S(S[28]) );
  FA_7011 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(1'b0), .S(S[29]), .CO(
        C[30]) );
  FA_7010 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_7009 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_7041 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_7042 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7043 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7044 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_7045 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7046 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7047 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7048 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7049 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7050 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7051 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7052 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7053 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7054 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7055 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7056 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7057 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7058 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7059 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7060 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7061 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7062 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7063 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7064 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7065 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7066 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7067 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7068 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7069 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7070 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7071 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_224 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_7071 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_7070 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_7069 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_7068 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_7067 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_7066 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_7065 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_7064 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_7063 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_7062 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_7061 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_7060 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_7059 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_7058 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_7057 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_7056 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_7055 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_7054 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_7053 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_7052 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_7051 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_7050 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_7049 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_7048 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_7047 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_7046 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_7045 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_7044 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(1'b0), .S(S[28]), .CO(
        C[29]) );
  FA_7043 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_7042 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_7041 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_7073 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_7074 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7075 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7076 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7077 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_7078 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7079 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7080 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7081 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7082 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7083 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7084 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7085 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7086 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7087 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7088 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7089 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7090 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7091 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7092 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7093 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7094 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7095 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7096 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7097 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7098 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7099 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_225 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_7103 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_7102 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_7101 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_7100 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_7099 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_7098 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_7097 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_7096 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_7095 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_7094 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_7093 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_7092 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_7091 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_7090 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_7089 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_7088 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_7087 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_7086 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_7085 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_7084 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_7083 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_7082 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_7081 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_7080 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_7079 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_7078 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_7077 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(1'b0), .S(S[27]), .CO(
        C[28]) );
  FA_7076 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_7075 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_7074 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_7073 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_7105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_7106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_7111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7120 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_226 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_7135 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_7134 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_7133 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_7132 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_7131 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_7130 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_7129 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_7128 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_7127 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_7126 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_7125 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_7124 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_7123 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_7122 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_7121 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_7120 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_7119 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_7118 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_7117 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_7116 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_7115 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_7114 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_7113 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_7112 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_7111 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_7110 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(1'b0), .S(S[26]), .CO(
        C[27]) );
  FA_7109 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_7108 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_7107 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_7106 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_7105 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_7137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_7138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_7144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7152 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_227 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_7167 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_7166 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_7165 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_7164 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_7163 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_7162 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_7161 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_7160 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_7159 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_7158 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_7157 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_7156 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_7155 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_7154 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_7153 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_7152 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_7151 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_7150 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_7149 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_7148 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_7147 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_7146 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_7145 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_7144 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_7143 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(1'b0), .S(S[25]), .CO(
        C[26]) );
  FA_7142 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_7141 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_7140 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_7139 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_7138 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_7137 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_7169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_7170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_7177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7184 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_228 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_7199 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_7198 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_7197 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_7196 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_7195 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_7194 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_7193 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_7192 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_7191 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_7190 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_7189 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_7188 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_7187 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_7186 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_7185 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_7184 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_7183 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_7182 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_7181 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_7180 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_7179 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_7178 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_7177 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_7176 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(1'b0), .S(S[24]), .CO(
        C[25]) );
  FA_7175 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_7174 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_7173 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_7172 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_7171 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_7170 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_7169 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_7201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_7202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_7210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7216 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_229 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_7231 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_7230 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_7229 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_7228 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_7227 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_7226 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_7225 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_7224 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_7223 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_7222 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_7221 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_7220 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_7219 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_7218 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_7217 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_7216 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_7215 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_7214 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_7213 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_7212 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_7211 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_7210 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_7209 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(1'b0), .S(S[23]), .CO(
        C[24]) );
  FA_7208 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_7207 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_7206 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_7205 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_7204 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_7203 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_7202 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_7201 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_7233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_7234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_7243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7248 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_230 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_7263 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_7262 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_7261 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_7260 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_7259 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_7258 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_7257 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_7256 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_7255 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_7254 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_7253 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_7252 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_7251 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_7250 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_7249 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_7248 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_7247 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_7246 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_7245 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_7244 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_7243 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_7242 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(1'b0), .S(S[22]), .CO(
        C[23]) );
  FA_7241 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_7240 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_7239 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_7238 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_7237 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_7236 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_7235 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_7234 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_7233 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_7265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_7266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_7276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7280 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_231 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_7295 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_7294 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_7293 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_7292 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_7291 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_7290 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_7289 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_7288 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_7287 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_7286 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_7285 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_7284 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_7283 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_7282 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_7281 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_7280 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_7279 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_7278 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_7277 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_7276 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_7275 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(1'b0), .S(S[21]), .CO(
        C[22]) );
  FA_7274 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_7273 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_7272 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_7271 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_7270 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_7269 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_7268 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_7267 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_7266 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_7265 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_7297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_7298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_7309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7312 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_232 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_7327 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_7326 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_7325 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_7324 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_7323 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_7322 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_7321 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_7320 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_7319 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_7318 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_7317 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_7316 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_7315 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_7314 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_7313 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_7312 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_7311 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_7310 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_7309 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_7308 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(1'b0), .S(S[20]), .CO(
        C[21]) );
  FA_7307 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_7306 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_7305 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_7304 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_7303 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_7302 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_7301 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_7300 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_7299 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_7298 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_7297 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_7329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_7330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_7342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7344 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_233 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_7359 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_7358 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_7357 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_7356 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_7355 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_7354 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_7353 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_7352 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_7351 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_7350 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_7349 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_7348 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_7347 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_7346 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_7345 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_7344 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_7343 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_7342 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_7341 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(1'b0), .S(S[19]), .CO(
        C[20]) );
  FA_7340 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_7339 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_7338 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_7337 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_7336 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_7335 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_7334 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_7333 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_7332 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_7331 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_7330 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_7329 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_7361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_7362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_7375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7376 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_234 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_7391 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_7390 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_7389 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_7388 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_7387 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_7386 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_7385 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_7384 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_7383 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_7382 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_7381 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_7380 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_7379 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_7378 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_7377 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_7376 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_7375 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_7374 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(1'b0), .S(S[18]), .CO(
        C[19]) );
  FA_7373 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_7372 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_7371 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_7370 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_7369 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_7368 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_7367 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_7366 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_7365 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_7364 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_7363 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_7362 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_7361 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_7393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_7394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_7408 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_235 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_7423 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_7422 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_7421 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_7420 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_7419 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_7418 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_7417 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_7416 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_7415 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_7414 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_7413 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_7412 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_7411 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_7410 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_7409 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_7408 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_7407 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(1'b0), .S(S[17]), .CO(
        C[18]) );
  FA_7406 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_7405 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_7404 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_7403 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_7402 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_7401 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_7400 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_7399 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_7398 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_7397 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_7396 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_7395 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_7394 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_7393 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_7425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_7426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7440 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_7441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_236 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_7455 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_7454 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_7453 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_7452 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_7451 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_7450 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_7449 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_7448 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_7447 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_7446 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_7445 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_7444 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_7443 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_7442 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_7441 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_7440 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(1'b0), .S(S[16]), .CO(
        C[17]) );
  FA_7439 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_7438 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_7437 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_7436 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_7435 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_7434 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_7433 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_7432 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_7431 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_7430 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_7429 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_7428 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_7427 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_7426 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_7425 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_7457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_7458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7472 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_7474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_237 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_7487 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_7486 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_7485 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_7484 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_7483 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_7482 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_7481 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_7480 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_7479 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_7478 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_7477 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_7476 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_7475 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_7474 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_7473 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(1'b0), .S(S[15]), .CO(
        C[16]) );
  FA_7472 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_7471 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_7470 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_7469 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_7468 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_7467 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_7466 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_7465 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_7464 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_7463 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_7462 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_7461 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_7460 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_7459 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_7458 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_7457 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_7489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_7490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7504 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_7507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7512 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7513 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7514 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7515 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7516 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7517 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7518 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7519 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_238 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_7519 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_7518 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_7517 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_7516 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_7515 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_7514 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_7513 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_7512 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_7511 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_7510 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_7509 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_7508 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_7507 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_7506 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(1'b0), .S(S[14]), .CO(
        C[15]) );
  FA_7505 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_7504 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_7503 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_7502 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_7501 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_7500 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_7499 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_7498 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_7497 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_7496 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_7495 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_7494 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_7493 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_7492 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_7491 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_7490 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_7489 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_7521 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_7522 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7523 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7524 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7525 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7526 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7527 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7528 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7529 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7530 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7531 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7532 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7533 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7534 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7535 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7536 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7537 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7538 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7539 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_7540 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7541 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7542 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7543 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7544 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7545 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7546 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7547 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7548 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7549 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7550 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7551 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_239 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_7551 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_7550 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_7549 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_7548 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_7547 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_7546 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_7545 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_7544 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_7543 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_7542 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_7541 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_7540 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_7539 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(1'b0), .S(S[13]), .CO(
        C[14]) );
  FA_7538 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_7537 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_7536 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_7535 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_7534 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_7533 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_7532 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_7531 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_7530 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_7529 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_7528 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_7527 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_7526 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_7525 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_7524 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_7523 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_7522 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_7521 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_7553 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_7554 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7555 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7556 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7557 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7558 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7559 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7560 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7561 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7562 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7563 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7564 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7565 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7566 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7567 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7568 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7569 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7570 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7571 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7572 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_7573 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7574 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7575 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7576 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7577 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7578 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7579 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7580 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7581 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7582 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7583 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_240 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_7583 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_7582 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_7581 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_7580 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_7579 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_7578 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_7577 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_7576 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_7575 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_7574 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_7573 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_7572 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(1'b0), .S(S[12]), .CO(
        C[13]) );
  FA_7571 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_7570 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_7569 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_7568 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_7567 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_7566 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_7565 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_7564 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_7563 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_7562 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_7561 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_7560 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_7559 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_7558 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_7557 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_7556 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_7555 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_7554 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_7553 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_7585 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_7586 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7587 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7588 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7589 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7590 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7591 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7592 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7593 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7594 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7595 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7596 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7597 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7598 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7599 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7600 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7601 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7602 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7603 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7604 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7605 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_7606 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7607 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7608 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7609 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7610 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7611 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7612 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7613 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7614 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7615 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_241 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_7615 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_7614 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_7613 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_7612 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_7611 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_7610 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_7609 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_7608 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_7607 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_7606 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_7605 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(1'b0), .S(S[11]), .CO(
        C[12]) );
  FA_7604 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_7603 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_7602 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_7601 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_7600 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_7599 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_7598 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_7597 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_7596 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_7595 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_7594 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_7593 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_7592 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_7591 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_7590 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_7589 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_7588 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_7587 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_7586 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_7585 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_7617 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_7618 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7619 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7620 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7621 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7622 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7623 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7624 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7625 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7626 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7627 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7628 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7629 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7630 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7631 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7632 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7633 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7634 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7635 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7636 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7637 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7638 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_7639 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7640 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7641 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7642 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7643 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7644 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7645 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7646 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7647 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_242 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_7647 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_7646 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_7645 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_7644 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_7643 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_7642 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_7641 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_7640 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_7639 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_7638 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(1'b0), .S(S[10]), .CO(
        C[11]) );
  FA_7637 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_7636 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_7635 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_7634 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_7633 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_7632 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_7631 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_7630 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_7629 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_7628 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_7627 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_7626 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_7625 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_7624 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_7623 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_7622 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_7621 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_7620 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_7619 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_7618 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_7617 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_7649 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_7650 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7651 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7652 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7653 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7654 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7655 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7656 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7657 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7658 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7659 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7660 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7661 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7662 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7663 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7664 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7665 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7666 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7667 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7668 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7669 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7670 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7671 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_7672 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7673 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7674 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7675 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7676 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7677 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7678 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7679 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_243 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_7679 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_7678 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_7677 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_7676 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_7675 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_7674 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_7673 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_7672 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_7671 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(1'b0), .S(S[9]), .CO(C[10]) );
  FA_7670 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_7669 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_7668 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_7667 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_7666 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_7665 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_7664 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_7663 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_7662 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_7661 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_7660 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_7659 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_7658 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_7657 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_7656 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_7655 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_7654 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_7653 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_7652 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_7651 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_7650 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_7649 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_7681 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_7682 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7683 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7684 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7685 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7686 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7687 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7688 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7689 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7690 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7691 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7692 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7693 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7694 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7695 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7696 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7697 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7698 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7699 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7700 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7701 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7702 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7703 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7704 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_7705 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7706 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7707 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7708 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7709 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7710 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7711 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_244 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_7711 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_7710 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_7709 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_7708 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_7707 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_7706 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_7705 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_7704 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(1'b0), .S(S[8]), .CO(C[9])
         );
  FA_7703 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_7702 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_7701 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_7700 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_7699 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_7698 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_7697 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_7696 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_7695 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_7694 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_7693 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_7692 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_7691 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_7690 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_7689 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_7688 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_7687 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_7686 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_7685 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_7684 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_7683 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_7682 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_7681 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_7713 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_7714 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7715 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7716 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7717 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7718 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7719 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7720 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7721 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7722 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7723 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7724 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7725 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7726 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7727 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7728 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7729 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7730 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7731 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7732 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7733 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7734 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7735 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7736 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7737 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_7738 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7739 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7740 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7741 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7742 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7743 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_245 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_7743 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_7742 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_7741 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_7740 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_7739 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_7738 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_7737 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(1'b0), .S(S[7]), .CO(C[8])
         );
  FA_7736 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_7735 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_7734 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_7733 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_7732 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_7731 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_7730 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_7729 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_7728 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_7727 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_7726 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_7725 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_7724 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_7723 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_7722 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_7721 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_7720 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_7719 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_7718 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_7717 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_7716 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_7715 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_7714 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_7713 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_7745 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_7746 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7747 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7748 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7749 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7750 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7751 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7752 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7753 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7754 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7755 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7756 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7757 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7758 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7759 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7760 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7761 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7762 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7763 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7764 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7765 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7766 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7767 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7768 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7769 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7770 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_7771 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7772 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7773 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7774 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7775 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_246 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_7775 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_7774 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_7773 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_7772 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_7771 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_7770 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(1'b0), .S(S[6]), .CO(C[7])
         );
  FA_7769 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_7768 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_7767 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_7766 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_7765 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_7764 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_7763 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_7762 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_7761 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_7760 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_7759 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_7758 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_7757 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_7756 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_7755 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_7754 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_7753 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_7752 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_7751 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_7750 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_7749 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_7748 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_7747 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_7746 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_7745 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_7777 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_7778 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7779 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7780 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7781 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7782 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7783 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7784 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7785 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7786 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7787 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7788 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7789 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7790 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7791 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7792 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7793 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7794 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7795 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7796 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7797 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7798 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7799 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7800 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7801 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7802 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7803 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_7804 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7805 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7806 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7807 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_247 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_7807 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_7806 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_7805 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_7804 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_7803 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(1'b0), .S(S[5]), .CO(C[6])
         );
  FA_7802 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_7801 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_7800 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_7799 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_7798 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_7797 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_7796 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_7795 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_7794 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_7793 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_7792 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_7791 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_7790 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_7789 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_7788 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_7787 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_7786 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_7785 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_7784 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_7783 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_7782 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_7781 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_7780 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_7779 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_7778 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_7777 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_7809 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_7810 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7811 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7812 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7813 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7814 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7815 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7816 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7817 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7818 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7819 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7820 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7821 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7822 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7823 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7824 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7825 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7826 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7827 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7828 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7829 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7830 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7831 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7832 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7833 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7834 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7835 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7836 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_7837 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7838 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7839 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_248 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_7839 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_7838 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_7837 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_7836 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(1'b0), .S(S[4]), .CO(C[5])
         );
  FA_7835 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_7834 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_7833 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_7832 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_7831 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_7830 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_7829 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_7828 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_7827 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_7826 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_7825 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_7824 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_7823 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_7822 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_7821 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_7820 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_7819 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_7818 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_7817 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_7816 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_7815 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_7814 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_7813 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_7812 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_7811 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_7810 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_7809 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_7841 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_7842 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7843 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7844 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7845 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7846 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7847 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7848 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7849 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7850 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7851 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7852 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7853 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7854 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7855 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7856 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7857 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7858 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7859 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7860 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7861 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7862 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7863 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7864 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7865 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7866 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7867 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7868 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7869 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_7870 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7871 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_249 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_7871 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_7870 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_7869 \FAINST[3].FA_  ( .A(A[3]), .B(B[3]), .CI(1'b0), .S(S[3]), .CO(C[4])
         );
  FA_7868 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_7867 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_7866 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_7865 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_7864 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_7863 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_7862 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_7861 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_7860 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_7859 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_7858 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_7857 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_7856 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_7855 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_7854 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_7853 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_7852 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_7851 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_7850 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_7849 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_7848 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_7847 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_7846 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_7845 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_7844 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_7843 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_7842 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_7841 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_7873 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_7874 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7875 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7876 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7877 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7878 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7879 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7880 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7881 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7882 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7883 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7884 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7885 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7886 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7887 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7888 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7889 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7890 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7891 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7892 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7893 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7894 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7895 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7896 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7897 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7898 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7899 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7900 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7901 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7902 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_7903 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_250 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_7903 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_7902 \FAINST[2].FA_  ( .A(A[2]), .B(B[2]), .CI(1'b0), .S(S[2]), .CO(C[3])
         );
  FA_7901 \FAINST[3].FA_  ( .A(A[3]), .B(B[3]), .CI(C[3]), .S(S[3]), .CO(C[4])
         );
  FA_7900 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_7899 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_7898 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_7897 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_7896 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_7895 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_7894 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_7893 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_7892 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_7891 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_7890 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_7889 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_7888 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_7887 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_7886 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_7885 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_7884 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_7883 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_7882 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_7881 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_7880 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_7879 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_7878 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_7877 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_7876 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_7875 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_7874 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_7873 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_7905 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_7906 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_7907 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_7908 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_7909 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_7910 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_7911 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_7912 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_7913 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_7914 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_7915 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_7916 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_7917 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_7918 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_7919 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_7920 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_7921 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_7922 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_7923 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_7924 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_7925 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_7926 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_7927 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_7928 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_7929 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_7930 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_7931 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_7932 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_7933 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_7934 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_7935 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module ADD_N32_251 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;


  FA_7935 \FAINST[1].FA_  ( .A(A[1]), .B(1'b0), .CI(1'b0), .S(S[1]) );
  FA_7934 \FAINST[2].FA_  ( .A(A[2]), .B(1'b0), .CI(1'b0), .S(S[2]) );
  FA_7933 \FAINST[3].FA_  ( .A(A[3]), .B(1'b0), .CI(1'b0), .S(S[3]) );
  FA_7932 \FAINST[4].FA_  ( .A(A[4]), .B(1'b0), .CI(1'b0), .S(S[4]) );
  FA_7931 \FAINST[5].FA_  ( .A(A[5]), .B(1'b0), .CI(1'b0), .S(S[5]) );
  FA_7930 \FAINST[6].FA_  ( .A(A[6]), .B(1'b0), .CI(1'b0), .S(S[6]) );
  FA_7929 \FAINST[7].FA_  ( .A(A[7]), .B(1'b0), .CI(1'b0), .S(S[7]) );
  FA_7928 \FAINST[8].FA_  ( .A(A[8]), .B(1'b0), .CI(1'b0), .S(S[8]) );
  FA_7927 \FAINST[9].FA_  ( .A(A[9]), .B(1'b0), .CI(1'b0), .S(S[9]) );
  FA_7926 \FAINST[10].FA_  ( .A(A[10]), .B(1'b0), .CI(1'b0), .S(S[10]) );
  FA_7925 \FAINST[11].FA_  ( .A(A[11]), .B(1'b0), .CI(1'b0), .S(S[11]) );
  FA_7924 \FAINST[12].FA_  ( .A(A[12]), .B(1'b0), .CI(1'b0), .S(S[12]) );
  FA_7923 \FAINST[13].FA_  ( .A(A[13]), .B(1'b0), .CI(1'b0), .S(S[13]) );
  FA_7922 \FAINST[14].FA_  ( .A(A[14]), .B(1'b0), .CI(1'b0), .S(S[14]) );
  FA_7921 \FAINST[15].FA_  ( .A(A[15]), .B(1'b0), .CI(1'b0), .S(S[15]) );
  FA_7920 \FAINST[16].FA_  ( .A(A[16]), .B(1'b0), .CI(1'b0), .S(S[16]) );
  FA_7919 \FAINST[17].FA_  ( .A(A[17]), .B(1'b0), .CI(1'b0), .S(S[17]) );
  FA_7918 \FAINST[18].FA_  ( .A(A[18]), .B(1'b0), .CI(1'b0), .S(S[18]) );
  FA_7917 \FAINST[19].FA_  ( .A(A[19]), .B(1'b0), .CI(1'b0), .S(S[19]) );
  FA_7916 \FAINST[20].FA_  ( .A(A[20]), .B(1'b0), .CI(1'b0), .S(S[20]) );
  FA_7915 \FAINST[21].FA_  ( .A(A[21]), .B(1'b0), .CI(1'b0), .S(S[21]) );
  FA_7914 \FAINST[22].FA_  ( .A(A[22]), .B(1'b0), .CI(1'b0), .S(S[22]) );
  FA_7913 \FAINST[23].FA_  ( .A(A[23]), .B(1'b0), .CI(1'b0), .S(S[23]) );
  FA_7912 \FAINST[24].FA_  ( .A(A[24]), .B(1'b0), .CI(1'b0), .S(S[24]) );
  FA_7911 \FAINST[25].FA_  ( .A(A[25]), .B(1'b0), .CI(1'b0), .S(S[25]) );
  FA_7910 \FAINST[26].FA_  ( .A(A[26]), .B(1'b0), .CI(1'b0), .S(S[26]) );
  FA_7909 \FAINST[27].FA_  ( .A(A[27]), .B(1'b0), .CI(1'b0), .S(S[27]) );
  FA_7908 \FAINST[28].FA_  ( .A(A[28]), .B(1'b0), .CI(1'b0), .S(S[28]) );
  FA_7907 \FAINST[29].FA_  ( .A(A[29]), .B(1'b0), .CI(1'b0), .S(S[29]) );
  FA_7906 \FAINST[30].FA_  ( .A(A[30]), .B(1'b0), .CI(1'b0), .S(S[30]) );
  FA_7905 \FAINST[31].FA_  ( .A(A[31]), .B(1'b0), .CI(1'b0), .S(S[31]) );
endmodule


module MULT_N32_3 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   \w[31][31] , \w[31][30] , \w[31][29] , \w[31][28] , \w[31][27] ,
         \w[31][26] , \w[31][25] , \w[31][24] , \w[31][23] , \w[31][22] ,
         \w[31][21] , \w[31][20] , \w[31][19] , \w[31][18] , \w[31][17] ,
         \w[31][16] , \w[31][15] , \w[31][14] , \w[31][13] , \w[31][12] ,
         \w[31][11] , \w[31][10] , \w[31][9] , \w[31][8] , \w[31][7] ,
         \w[31][6] , \w[31][5] , \w[31][4] , \w[31][3] , \w[31][2] ,
         \w[31][1] , \w[30][31] , \w[30][30] , \w[30][29] , \w[30][28] ,
         \w[30][27] , \w[30][26] , \w[30][25] , \w[30][24] , \w[30][23] ,
         \w[30][22] , \w[30][21] , \w[30][20] , \w[30][19] , \w[30][18] ,
         \w[30][17] , \w[30][16] , \w[30][15] , \w[30][14] , \w[30][13] ,
         \w[30][12] , \w[30][11] , \w[30][10] , \w[30][9] , \w[30][8] ,
         \w[30][7] , \w[30][6] , \w[30][5] , \w[30][4] , \w[30][3] ,
         \w[30][2] , \w[30][1] , \w[29][31] , \w[29][30] , \w[29][29] ,
         \w[29][28] , \w[29][27] , \w[29][26] , \w[29][25] , \w[29][24] ,
         \w[29][23] , \w[29][22] , \w[29][21] , \w[29][20] , \w[29][19] ,
         \w[29][18] , \w[29][17] , \w[29][16] , \w[29][15] , \w[29][14] ,
         \w[29][13] , \w[29][12] , \w[29][11] , \w[29][10] , \w[29][9] ,
         \w[29][8] , \w[29][7] , \w[29][6] , \w[29][5] , \w[29][4] ,
         \w[29][3] , \w[29][2] , \w[29][1] , \w[28][31] , \w[28][30] ,
         \w[28][29] , \w[28][28] , \w[28][27] , \w[28][26] , \w[28][25] ,
         \w[28][24] , \w[28][23] , \w[28][22] , \w[28][21] , \w[28][20] ,
         \w[28][19] , \w[28][18] , \w[28][17] , \w[28][16] , \w[28][15] ,
         \w[28][14] , \w[28][13] , \w[28][12] , \w[28][11] , \w[28][10] ,
         \w[28][9] , \w[28][8] , \w[28][7] , \w[28][6] , \w[28][5] ,
         \w[28][4] , \w[28][3] , \w[28][2] , \w[28][1] , \w[27][31] ,
         \w[27][30] , \w[27][29] , \w[27][28] , \w[27][27] , \w[27][26] ,
         \w[27][25] , \w[27][24] , \w[27][23] , \w[27][22] , \w[27][21] ,
         \w[27][20] , \w[27][19] , \w[27][18] , \w[27][17] , \w[27][16] ,
         \w[27][15] , \w[27][14] , \w[27][13] , \w[27][12] , \w[27][11] ,
         \w[27][10] , \w[27][9] , \w[27][8] , \w[27][7] , \w[27][6] ,
         \w[27][5] , \w[27][4] , \w[27][3] , \w[27][2] , \w[27][1] ,
         \w[26][31] , \w[26][30] , \w[26][29] , \w[26][28] , \w[26][27] ,
         \w[26][26] , \w[26][25] , \w[26][24] , \w[26][23] , \w[26][22] ,
         \w[26][21] , \w[26][20] , \w[26][19] , \w[26][18] , \w[26][17] ,
         \w[26][16] , \w[26][15] , \w[26][14] , \w[26][13] , \w[26][12] ,
         \w[26][11] , \w[26][10] , \w[26][9] , \w[26][8] , \w[26][7] ,
         \w[26][6] , \w[26][5] , \w[26][4] , \w[26][3] , \w[26][2] ,
         \w[26][1] , \w[25][31] , \w[25][30] , \w[25][29] , \w[25][28] ,
         \w[25][27] , \w[25][26] , \w[25][25] , \w[25][24] , \w[25][23] ,
         \w[25][22] , \w[25][21] , \w[25][20] , \w[25][19] , \w[25][18] ,
         \w[25][17] , \w[25][16] , \w[25][15] , \w[25][14] , \w[25][13] ,
         \w[25][12] , \w[25][11] , \w[25][10] , \w[25][9] , \w[25][8] ,
         \w[25][7] , \w[25][6] , \w[25][5] , \w[25][4] , \w[25][3] ,
         \w[25][2] , \w[25][1] , \w[24][31] , \w[24][30] , \w[24][29] ,
         \w[24][28] , \w[24][27] , \w[24][26] , \w[24][25] , \w[24][24] ,
         \w[24][23] , \w[24][22] , \w[24][21] , \w[24][20] , \w[24][19] ,
         \w[24][18] , \w[24][17] , \w[24][16] , \w[24][15] , \w[24][14] ,
         \w[24][13] , \w[24][12] , \w[24][11] , \w[24][10] , \w[24][9] ,
         \w[24][8] , \w[24][7] , \w[24][6] , \w[24][5] , \w[24][4] ,
         \w[24][3] , \w[24][2] , \w[24][1] , \w[23][31] , \w[23][30] ,
         \w[23][29] , \w[23][28] , \w[23][27] , \w[23][26] , \w[23][25] ,
         \w[23][24] , \w[23][23] , \w[23][22] , \w[23][21] , \w[23][20] ,
         \w[23][19] , \w[23][18] , \w[23][17] , \w[23][16] , \w[23][15] ,
         \w[23][14] , \w[23][13] , \w[23][12] , \w[23][11] , \w[23][10] ,
         \w[23][9] , \w[23][8] , \w[23][7] , \w[23][6] , \w[23][5] ,
         \w[23][4] , \w[23][3] , \w[23][2] , \w[23][1] , \w[22][31] ,
         \w[22][30] , \w[22][29] , \w[22][28] , \w[22][27] , \w[22][26] ,
         \w[22][25] , \w[22][24] , \w[22][23] , \w[22][22] , \w[22][21] ,
         \w[22][20] , \w[22][19] , \w[22][18] , \w[22][17] , \w[22][16] ,
         \w[22][15] , \w[22][14] , \w[22][13] , \w[22][12] , \w[22][11] ,
         \w[22][10] , \w[22][9] , \w[22][8] , \w[22][7] , \w[22][6] ,
         \w[22][5] , \w[22][4] , \w[22][3] , \w[22][2] , \w[22][1] ,
         \w[21][31] , \w[21][30] , \w[21][29] , \w[21][28] , \w[21][27] ,
         \w[21][26] , \w[21][25] , \w[21][24] , \w[21][23] , \w[21][22] ,
         \w[21][21] , \w[21][20] , \w[21][19] , \w[21][18] , \w[21][17] ,
         \w[21][16] , \w[21][15] , \w[21][14] , \w[21][13] , \w[21][12] ,
         \w[21][11] , \w[21][10] , \w[21][9] , \w[21][8] , \w[21][7] ,
         \w[21][6] , \w[21][5] , \w[21][4] , \w[21][3] , \w[21][2] ,
         \w[21][1] , \w[20][31] , \w[20][30] , \w[20][29] , \w[20][28] ,
         \w[20][27] , \w[20][26] , \w[20][25] , \w[20][24] , \w[20][23] ,
         \w[20][22] , \w[20][21] , \w[20][20] , \w[20][19] , \w[20][18] ,
         \w[20][17] , \w[20][16] , \w[20][15] , \w[20][14] , \w[20][13] ,
         \w[20][12] , \w[20][11] , \w[20][10] , \w[20][9] , \w[20][8] ,
         \w[20][7] , \w[20][6] , \w[20][5] , \w[20][4] , \w[20][3] ,
         \w[20][2] , \w[20][1] , \w[19][31] , \w[19][30] , \w[19][29] ,
         \w[19][28] , \w[19][27] , \w[19][26] , \w[19][25] , \w[19][24] ,
         \w[19][23] , \w[19][22] , \w[19][21] , \w[19][20] , \w[19][19] ,
         \w[19][18] , \w[19][17] , \w[19][16] , \w[19][15] , \w[19][14] ,
         \w[19][13] , \w[19][12] , \w[19][11] , \w[19][10] , \w[19][9] ,
         \w[19][8] , \w[19][7] , \w[19][6] , \w[19][5] , \w[19][4] ,
         \w[19][3] , \w[19][2] , \w[19][1] , \w[18][31] , \w[18][30] ,
         \w[18][29] , \w[18][28] , \w[18][27] , \w[18][26] , \w[18][25] ,
         \w[18][24] , \w[18][23] , \w[18][22] , \w[18][21] , \w[18][20] ,
         \w[18][19] , \w[18][18] , \w[18][17] , \w[18][16] , \w[18][15] ,
         \w[18][14] , \w[18][13] , \w[18][12] , \w[18][11] , \w[18][10] ,
         \w[18][9] , \w[18][8] , \w[18][7] , \w[18][6] , \w[18][5] ,
         \w[18][4] , \w[18][3] , \w[18][2] , \w[18][1] , \w[17][31] ,
         \w[17][30] , \w[17][29] , \w[17][28] , \w[17][27] , \w[17][26] ,
         \w[17][25] , \w[17][24] , \w[17][23] , \w[17][22] , \w[17][21] ,
         \w[17][20] , \w[17][19] , \w[17][18] , \w[17][17] , \w[17][16] ,
         \w[17][15] , \w[17][14] , \w[17][13] , \w[17][12] , \w[17][11] ,
         \w[17][10] , \w[17][9] , \w[17][8] , \w[17][7] , \w[17][6] ,
         \w[17][5] , \w[17][4] , \w[17][3] , \w[17][2] , \w[17][1] ,
         \w[16][31] , \w[16][30] , \w[16][29] , \w[16][28] , \w[16][27] ,
         \w[16][26] , \w[16][25] , \w[16][24] , \w[16][23] , \w[16][22] ,
         \w[16][21] , \w[16][20] , \w[16][19] , \w[16][18] , \w[16][17] ,
         \w[16][16] , \w[16][15] , \w[16][14] , \w[16][13] , \w[16][12] ,
         \w[16][11] , \w[16][10] , \w[16][9] , \w[16][8] , \w[16][7] ,
         \w[16][6] , \w[16][5] , \w[16][4] , \w[16][3] , \w[16][2] ,
         \w[16][1] , \w[15][31] , \w[15][30] , \w[15][29] , \w[15][28] ,
         \w[15][27] , \w[15][26] , \w[15][25] , \w[15][24] , \w[15][23] ,
         \w[15][22] , \w[15][21] , \w[15][20] , \w[15][19] , \w[15][18] ,
         \w[15][17] , \w[15][16] , \w[15][15] , \w[15][14] , \w[15][13] ,
         \w[15][12] , \w[15][11] , \w[15][10] , \w[15][9] , \w[15][8] ,
         \w[15][7] , \w[15][6] , \w[15][5] , \w[15][4] , \w[15][3] ,
         \w[15][2] , \w[15][1] , \w[14][31] , \w[14][30] , \w[14][29] ,
         \w[14][28] , \w[14][27] , \w[14][26] , \w[14][25] , \w[14][24] ,
         \w[14][23] , \w[14][22] , \w[14][21] , \w[14][20] , \w[14][19] ,
         \w[14][18] , \w[14][17] , \w[14][16] , \w[14][15] , \w[14][14] ,
         \w[14][13] , \w[14][12] , \w[14][11] , \w[14][10] , \w[14][9] ,
         \w[14][8] , \w[14][7] , \w[14][6] , \w[14][5] , \w[14][4] ,
         \w[14][3] , \w[14][2] , \w[14][1] , \w[13][31] , \w[13][30] ,
         \w[13][29] , \w[13][28] , \w[13][27] , \w[13][26] , \w[13][25] ,
         \w[13][24] , \w[13][23] , \w[13][22] , \w[13][21] , \w[13][20] ,
         \w[13][19] , \w[13][18] , \w[13][17] , \w[13][16] , \w[13][15] ,
         \w[13][14] , \w[13][13] , \w[13][12] , \w[13][11] , \w[13][10] ,
         \w[13][9] , \w[13][8] , \w[13][7] , \w[13][6] , \w[13][5] ,
         \w[13][4] , \w[13][3] , \w[13][2] , \w[13][1] , \w[12][31] ,
         \w[12][30] , \w[12][29] , \w[12][28] , \w[12][27] , \w[12][26] ,
         \w[12][25] , \w[12][24] , \w[12][23] , \w[12][22] , \w[12][21] ,
         \w[12][20] , \w[12][19] , \w[12][18] , \w[12][17] , \w[12][16] ,
         \w[12][15] , \w[12][14] , \w[12][13] , \w[12][12] , \w[12][11] ,
         \w[12][10] , \w[12][9] , \w[12][8] , \w[12][7] , \w[12][6] ,
         \w[12][5] , \w[12][4] , \w[12][3] , \w[12][2] , \w[12][1] ,
         \w[11][31] , \w[11][30] , \w[11][29] , \w[11][28] , \w[11][27] ,
         \w[11][26] , \w[11][25] , \w[11][24] , \w[11][23] , \w[11][22] ,
         \w[11][21] , \w[11][20] , \w[11][19] , \w[11][18] , \w[11][17] ,
         \w[11][16] , \w[11][15] , \w[11][14] , \w[11][13] , \w[11][12] ,
         \w[11][11] , \w[11][10] , \w[11][9] , \w[11][8] , \w[11][7] ,
         \w[11][6] , \w[11][5] , \w[11][4] , \w[11][3] , \w[11][2] ,
         \w[11][1] , \w[10][31] , \w[10][30] , \w[10][29] , \w[10][28] ,
         \w[10][27] , \w[10][26] , \w[10][25] , \w[10][24] , \w[10][23] ,
         \w[10][22] , \w[10][21] , \w[10][20] , \w[10][19] , \w[10][18] ,
         \w[10][17] , \w[10][16] , \w[10][15] , \w[10][14] , \w[10][13] ,
         \w[10][12] , \w[10][11] , \w[10][10] , \w[10][9] , \w[10][8] ,
         \w[10][7] , \w[10][6] , \w[10][5] , \w[10][4] , \w[10][3] ,
         \w[10][2] , \w[10][1] , \w[9][31] , \w[9][30] , \w[9][29] ,
         \w[9][28] , \w[9][27] , \w[9][26] , \w[9][25] , \w[9][24] ,
         \w[9][23] , \w[9][22] , \w[9][21] , \w[9][20] , \w[9][19] ,
         \w[9][18] , \w[9][17] , \w[9][16] , \w[9][15] , \w[9][14] ,
         \w[9][13] , \w[9][12] , \w[9][11] , \w[9][10] , \w[9][9] , \w[9][8] ,
         \w[9][7] , \w[9][6] , \w[9][5] , \w[9][4] , \w[9][3] , \w[9][2] ,
         \w[9][1] , \w[8][31] , \w[8][30] , \w[8][29] , \w[8][28] , \w[8][27] ,
         \w[8][26] , \w[8][25] , \w[8][24] , \w[8][23] , \w[8][22] ,
         \w[8][21] , \w[8][20] , \w[8][19] , \w[8][18] , \w[8][17] ,
         \w[8][16] , \w[8][15] , \w[8][14] , \w[8][13] , \w[8][12] ,
         \w[8][11] , \w[8][10] , \w[8][9] , \w[8][8] , \w[8][7] , \w[8][6] ,
         \w[8][5] , \w[8][4] , \w[8][3] , \w[8][2] , \w[8][1] , \w[7][31] ,
         \w[7][30] , \w[7][29] , \w[7][28] , \w[7][27] , \w[7][26] ,
         \w[7][25] , \w[7][24] , \w[7][23] , \w[7][22] , \w[7][21] ,
         \w[7][20] , \w[7][19] , \w[7][18] , \w[7][17] , \w[7][16] ,
         \w[7][15] , \w[7][14] , \w[7][13] , \w[7][12] , \w[7][11] ,
         \w[7][10] , \w[7][9] , \w[7][8] , \w[7][7] , \w[7][6] , \w[7][5] ,
         \w[7][4] , \w[7][3] , \w[7][2] , \w[7][1] , \w[6][31] , \w[6][30] ,
         \w[6][29] , \w[6][28] , \w[6][27] , \w[6][26] , \w[6][25] ,
         \w[6][24] , \w[6][23] , \w[6][22] , \w[6][21] , \w[6][20] ,
         \w[6][19] , \w[6][18] , \w[6][17] , \w[6][16] , \w[6][15] ,
         \w[6][14] , \w[6][13] , \w[6][12] , \w[6][11] , \w[6][10] , \w[6][9] ,
         \w[6][8] , \w[6][7] , \w[6][6] , \w[6][5] , \w[6][4] , \w[6][3] ,
         \w[6][2] , \w[6][1] , \w[5][31] , \w[5][30] , \w[5][29] , \w[5][28] ,
         \w[5][27] , \w[5][26] , \w[5][25] , \w[5][24] , \w[5][23] ,
         \w[5][22] , \w[5][21] , \w[5][20] , \w[5][19] , \w[5][18] ,
         \w[5][17] , \w[5][16] , \w[5][15] , \w[5][14] , \w[5][13] ,
         \w[5][12] , \w[5][11] , \w[5][10] , \w[5][9] , \w[5][8] , \w[5][7] ,
         \w[5][6] , \w[5][5] , \w[5][4] , \w[5][3] , \w[5][2] , \w[5][1] ,
         \w[4][31] , \w[4][30] , \w[4][29] , \w[4][28] , \w[4][27] ,
         \w[4][26] , \w[4][25] , \w[4][24] , \w[4][23] , \w[4][22] ,
         \w[4][21] , \w[4][20] , \w[4][19] , \w[4][18] , \w[4][17] ,
         \w[4][16] , \w[4][15] , \w[4][14] , \w[4][13] , \w[4][12] ,
         \w[4][11] , \w[4][10] , \w[4][9] , \w[4][8] , \w[4][7] , \w[4][6] ,
         \w[4][5] , \w[4][4] , \w[4][3] , \w[4][2] , \w[4][1] , \w[3][31] ,
         \w[3][30] , \w[3][29] , \w[3][28] , \w[3][27] , \w[3][26] ,
         \w[3][25] , \w[3][24] , \w[3][23] , \w[3][22] , \w[3][21] ,
         \w[3][20] , \w[3][19] , \w[3][18] , \w[3][17] , \w[3][16] ,
         \w[3][15] , \w[3][14] , \w[3][13] , \w[3][12] , \w[3][11] ,
         \w[3][10] , \w[3][9] , \w[3][8] , \w[3][7] , \w[3][6] , \w[3][5] ,
         \w[3][4] , \w[3][3] , \w[3][2] , \w[3][1] , \w[2][31] , \w[2][30] ,
         \w[2][29] , \w[2][28] , \w[2][27] , \w[2][26] , \w[2][25] ,
         \w[2][24] , \w[2][23] , \w[2][22] , \w[2][21] , \w[2][20] ,
         \w[2][19] , \w[2][18] , \w[2][17] , \w[2][16] , \w[2][15] ,
         \w[2][14] , \w[2][13] , \w[2][12] , \w[2][11] , \w[2][10] , \w[2][9] ,
         \w[2][8] , \w[2][7] , \w[2][6] , \w[2][5] , \w[2][4] , \w[2][3] ,
         \w[2][2] , \w[2][1] , \_0_net_[31] , \_0_net_[30] , \_0_net_[29] ,
         \_0_net_[28] , \_0_net_[27] , \_0_net_[26] , \_0_net_[25] ,
         \_0_net_[24] , \_0_net_[23] , \_0_net_[22] , \_0_net_[21] ,
         \_0_net_[20] , \_0_net_[19] , \_0_net_[18] , \_0_net_[17] ,
         \_0_net_[16] , \_0_net_[15] , \_0_net_[14] , \_0_net_[13] ,
         \_0_net_[12] , \_0_net_[11] , \_0_net_[10] , \_0_net_[9] ,
         \_0_net_[8] , \_0_net_[7] , \_0_net_[6] , \_0_net_[5] , \_0_net_[4] ,
         \_0_net_[3] , \_0_net_[2] , \_0_net_[1] , \_2_net_[31] ,
         \_2_net_[30] , \_2_net_[29] , \_2_net_[28] , \_2_net_[27] ,
         \_2_net_[26] , \_2_net_[25] , \_2_net_[24] , \_2_net_[23] ,
         \_2_net_[22] , \_2_net_[21] , \_2_net_[20] , \_2_net_[19] ,
         \_2_net_[18] , \_2_net_[17] , \_2_net_[16] , \_2_net_[15] ,
         \_2_net_[14] , \_2_net_[13] , \_2_net_[12] , \_2_net_[11] ,
         \_2_net_[10] , \_2_net_[9] , \_2_net_[8] , \_2_net_[7] , \_2_net_[6] ,
         \_2_net_[5] , \_2_net_[4] , \_2_net_[3] , \_2_net_[2] , \_4_net_[31] ,
         \_4_net_[30] , \_4_net_[29] , \_4_net_[28] , \_4_net_[27] ,
         \_4_net_[26] , \_4_net_[25] , \_4_net_[24] , \_4_net_[23] ,
         \_4_net_[22] , \_4_net_[21] , \_4_net_[20] , \_4_net_[19] ,
         \_4_net_[18] , \_4_net_[17] , \_4_net_[16] , \_4_net_[15] ,
         \_4_net_[14] , \_4_net_[13] , \_4_net_[12] , \_4_net_[11] ,
         \_4_net_[10] , \_4_net_[9] , \_4_net_[8] , \_4_net_[7] , \_4_net_[6] ,
         \_4_net_[5] , \_4_net_[4] , \_4_net_[3] , \_6_net_[31] ,
         \_6_net_[30] , \_6_net_[29] , \_6_net_[28] , \_6_net_[27] ,
         \_6_net_[26] , \_6_net_[25] , \_6_net_[24] , \_6_net_[23] ,
         \_6_net_[22] , \_6_net_[21] , \_6_net_[20] , \_6_net_[19] ,
         \_6_net_[18] , \_6_net_[17] , \_6_net_[16] , \_6_net_[15] ,
         \_6_net_[14] , \_6_net_[13] , \_6_net_[12] , \_6_net_[11] ,
         \_6_net_[10] , \_6_net_[9] , \_6_net_[8] , \_6_net_[7] , \_6_net_[6] ,
         \_6_net_[5] , \_6_net_[4] , \_8_net_[31] , \_8_net_[30] ,
         \_8_net_[29] , \_8_net_[28] , \_8_net_[27] , \_8_net_[26] ,
         \_8_net_[25] , \_8_net_[24] , \_8_net_[23] , \_8_net_[22] ,
         \_8_net_[21] , \_8_net_[20] , \_8_net_[19] , \_8_net_[18] ,
         \_8_net_[17] , \_8_net_[16] , \_8_net_[15] , \_8_net_[14] ,
         \_8_net_[13] , \_8_net_[12] , \_8_net_[11] , \_8_net_[10] ,
         \_8_net_[9] , \_8_net_[8] , \_8_net_[7] , \_8_net_[6] , \_8_net_[5] ,
         \_10_net_[31] , \_10_net_[30] , \_10_net_[29] , \_10_net_[28] ,
         \_10_net_[27] , \_10_net_[26] , \_10_net_[25] , \_10_net_[24] ,
         \_10_net_[23] , \_10_net_[22] , \_10_net_[21] , \_10_net_[20] ,
         \_10_net_[19] , \_10_net_[18] , \_10_net_[17] , \_10_net_[16] ,
         \_10_net_[15] , \_10_net_[14] , \_10_net_[13] , \_10_net_[12] ,
         \_10_net_[11] , \_10_net_[10] , \_10_net_[9] , \_10_net_[8] ,
         \_10_net_[7] , \_10_net_[6] , \_12_net_[31] , \_12_net_[30] ,
         \_12_net_[29] , \_12_net_[28] , \_12_net_[27] , \_12_net_[26] ,
         \_12_net_[25] , \_12_net_[24] , \_12_net_[23] , \_12_net_[22] ,
         \_12_net_[21] , \_12_net_[20] , \_12_net_[19] , \_12_net_[18] ,
         \_12_net_[17] , \_12_net_[16] , \_12_net_[15] , \_12_net_[14] ,
         \_12_net_[13] , \_12_net_[12] , \_12_net_[11] , \_12_net_[10] ,
         \_12_net_[9] , \_12_net_[8] , \_12_net_[7] , \_14_net_[31] ,
         \_14_net_[30] , \_14_net_[29] , \_14_net_[28] , \_14_net_[27] ,
         \_14_net_[26] , \_14_net_[25] , \_14_net_[24] , \_14_net_[23] ,
         \_14_net_[22] , \_14_net_[21] , \_14_net_[20] , \_14_net_[19] ,
         \_14_net_[18] , \_14_net_[17] , \_14_net_[16] , \_14_net_[15] ,
         \_14_net_[14] , \_14_net_[13] , \_14_net_[12] , \_14_net_[11] ,
         \_14_net_[10] , \_14_net_[9] , \_14_net_[8] , \_16_net_[31] ,
         \_16_net_[30] , \_16_net_[29] , \_16_net_[28] , \_16_net_[27] ,
         \_16_net_[26] , \_16_net_[25] , \_16_net_[24] , \_16_net_[23] ,
         \_16_net_[22] , \_16_net_[21] , \_16_net_[20] , \_16_net_[19] ,
         \_16_net_[18] , \_16_net_[17] , \_16_net_[16] , \_16_net_[15] ,
         \_16_net_[14] , \_16_net_[13] , \_16_net_[12] , \_16_net_[11] ,
         \_16_net_[10] , \_16_net_[9] , \_18_net_[31] , \_18_net_[30] ,
         \_18_net_[29] , \_18_net_[28] , \_18_net_[27] , \_18_net_[26] ,
         \_18_net_[25] , \_18_net_[24] , \_18_net_[23] , \_18_net_[22] ,
         \_18_net_[21] , \_18_net_[20] , \_18_net_[19] , \_18_net_[18] ,
         \_18_net_[17] , \_18_net_[16] , \_18_net_[15] , \_18_net_[14] ,
         \_18_net_[13] , \_18_net_[12] , \_18_net_[11] , \_18_net_[10] ,
         \_20_net_[31] , \_20_net_[30] , \_20_net_[29] , \_20_net_[28] ,
         \_20_net_[27] , \_20_net_[26] , \_20_net_[25] , \_20_net_[24] ,
         \_20_net_[23] , \_20_net_[22] , \_20_net_[21] , \_20_net_[20] ,
         \_20_net_[19] , \_20_net_[18] , \_20_net_[17] , \_20_net_[16] ,
         \_20_net_[15] , \_20_net_[14] , \_20_net_[13] , \_20_net_[12] ,
         \_20_net_[11] , \_22_net_[31] , \_22_net_[30] , \_22_net_[29] ,
         \_22_net_[28] , \_22_net_[27] , \_22_net_[26] , \_22_net_[25] ,
         \_22_net_[24] , \_22_net_[23] , \_22_net_[22] , \_22_net_[21] ,
         \_22_net_[20] , \_22_net_[19] , \_22_net_[18] , \_22_net_[17] ,
         \_22_net_[16] , \_22_net_[15] , \_22_net_[14] , \_22_net_[13] ,
         \_22_net_[12] , \_24_net_[31] , \_24_net_[30] , \_24_net_[29] ,
         \_24_net_[28] , \_24_net_[27] , \_24_net_[26] , \_24_net_[25] ,
         \_24_net_[24] , \_24_net_[23] , \_24_net_[22] , \_24_net_[21] ,
         \_24_net_[20] , \_24_net_[19] , \_24_net_[18] , \_24_net_[17] ,
         \_24_net_[16] , \_24_net_[15] , \_24_net_[14] , \_24_net_[13] ,
         \_26_net_[31] , \_26_net_[30] , \_26_net_[29] , \_26_net_[28] ,
         \_26_net_[27] , \_26_net_[26] , \_26_net_[25] , \_26_net_[24] ,
         \_26_net_[23] , \_26_net_[22] , \_26_net_[21] , \_26_net_[20] ,
         \_26_net_[19] , \_26_net_[18] , \_26_net_[17] , \_26_net_[16] ,
         \_26_net_[15] , \_26_net_[14] , \_28_net_[31] , \_28_net_[30] ,
         \_28_net_[29] , \_28_net_[28] , \_28_net_[27] , \_28_net_[26] ,
         \_28_net_[25] , \_28_net_[24] , \_28_net_[23] , \_28_net_[22] ,
         \_28_net_[21] , \_28_net_[20] , \_28_net_[19] , \_28_net_[18] ,
         \_28_net_[17] , \_28_net_[16] , \_28_net_[15] , \_30_net_[31] ,
         \_30_net_[30] , \_30_net_[29] , \_30_net_[28] , \_30_net_[27] ,
         \_30_net_[26] , \_30_net_[25] , \_30_net_[24] , \_30_net_[23] ,
         \_30_net_[22] , \_30_net_[21] , \_30_net_[20] , \_30_net_[19] ,
         \_30_net_[18] , \_30_net_[17] , \_30_net_[16] , \_32_net_[31] ,
         \_32_net_[30] , \_32_net_[29] , \_32_net_[28] , \_32_net_[27] ,
         \_32_net_[26] , \_32_net_[25] , \_32_net_[24] , \_32_net_[23] ,
         \_32_net_[22] , \_32_net_[21] , \_32_net_[20] , \_32_net_[19] ,
         \_32_net_[18] , \_32_net_[17] , \_34_net_[31] , \_34_net_[30] ,
         \_34_net_[29] , \_34_net_[28] , \_34_net_[27] , \_34_net_[26] ,
         \_34_net_[25] , \_34_net_[24] , \_34_net_[23] , \_34_net_[22] ,
         \_34_net_[21] , \_34_net_[20] , \_34_net_[19] , \_34_net_[18] ,
         \_36_net_[31] , \_36_net_[30] , \_36_net_[29] , \_36_net_[28] ,
         \_36_net_[27] , \_36_net_[26] , \_36_net_[25] , \_36_net_[24] ,
         \_36_net_[23] , \_36_net_[22] , \_36_net_[21] , \_36_net_[20] ,
         \_36_net_[19] , \_38_net_[31] , \_38_net_[30] , \_38_net_[29] ,
         \_38_net_[28] , \_38_net_[27] , \_38_net_[26] , \_38_net_[25] ,
         \_38_net_[24] , \_38_net_[23] , \_38_net_[22] , \_38_net_[21] ,
         \_38_net_[20] , \_40_net_[31] , \_40_net_[30] , \_40_net_[29] ,
         \_40_net_[28] , \_40_net_[27] , \_40_net_[26] , \_40_net_[25] ,
         \_40_net_[24] , \_40_net_[23] , \_40_net_[22] , \_40_net_[21] ,
         \_42_net_[31] , \_42_net_[30] , \_42_net_[29] , \_42_net_[28] ,
         \_42_net_[27] , \_42_net_[26] , \_42_net_[25] , \_42_net_[24] ,
         \_42_net_[23] , \_42_net_[22] , \_44_net_[31] , \_44_net_[30] ,
         \_44_net_[29] , \_44_net_[28] , \_44_net_[27] , \_44_net_[26] ,
         \_44_net_[25] , \_44_net_[24] , \_44_net_[23] , \_46_net_[31] ,
         \_46_net_[30] , \_46_net_[29] , \_46_net_[28] , \_46_net_[27] ,
         \_46_net_[26] , \_46_net_[25] , \_46_net_[24] , \_48_net_[31] ,
         \_48_net_[30] , \_48_net_[29] , \_48_net_[28] , \_48_net_[27] ,
         \_48_net_[26] , \_48_net_[25] , \_50_net_[31] , \_50_net_[30] ,
         \_50_net_[29] , \_50_net_[28] , \_50_net_[27] , \_50_net_[26] ,
         \_52_net_[31] , \_52_net_[30] , \_52_net_[29] , \_52_net_[28] ,
         \_52_net_[27] , \_54_net_[31] , \_54_net_[30] , \_54_net_[29] ,
         \_54_net_[28] , \_56_net_[31] , \_56_net_[30] , \_56_net_[29] ,
         \_58_net_[31] , \_58_net_[30] , \_60_net_[31] ;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30;

  ADD_N32_251 \FAINST[1].ADD_  ( .A({\_0_net_[31] , \_0_net_[30] , 
        \_0_net_[29] , \_0_net_[28] , \_0_net_[27] , \_0_net_[26] , 
        \_0_net_[25] , \_0_net_[24] , \_0_net_[23] , \_0_net_[22] , 
        \_0_net_[21] , \_0_net_[20] , \_0_net_[19] , \_0_net_[18] , 
        \_0_net_[17] , \_0_net_[16] , \_0_net_[15] , \_0_net_[14] , 
        \_0_net_[13] , \_0_net_[12] , \_0_net_[11] , \_0_net_[10] , 
        \_0_net_[9] , \_0_net_[8] , \_0_net_[7] , \_0_net_[6] , \_0_net_[5] , 
        \_0_net_[4] , \_0_net_[3] , \_0_net_[2] , \_0_net_[1] , 1'b0}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .S({
        \w[2][31] , \w[2][30] , \w[2][29] , \w[2][28] , \w[2][27] , \w[2][26] , 
        \w[2][25] , \w[2][24] , \w[2][23] , \w[2][22] , \w[2][21] , \w[2][20] , 
        \w[2][19] , \w[2][18] , \w[2][17] , \w[2][16] , \w[2][15] , \w[2][14] , 
        \w[2][13] , \w[2][12] , \w[2][11] , \w[2][10] , \w[2][9] , \w[2][8] , 
        \w[2][7] , \w[2][6] , \w[2][5] , \w[2][4] , \w[2][3] , \w[2][2] , 
        \w[2][1] , SYNOPSYS_UNCONNECTED__0}) );
  ADD_N32_250 \FAINST[2].ADD_  ( .A({\_2_net_[31] , \_2_net_[30] , 
        \_2_net_[29] , \_2_net_[28] , \_2_net_[27] , \_2_net_[26] , 
        \_2_net_[25] , \_2_net_[24] , \_2_net_[23] , \_2_net_[22] , 
        \_2_net_[21] , \_2_net_[20] , \_2_net_[19] , \_2_net_[18] , 
        \_2_net_[17] , \_2_net_[16] , \_2_net_[15] , \_2_net_[14] , 
        \_2_net_[13] , \_2_net_[12] , \_2_net_[11] , \_2_net_[10] , 
        \_2_net_[9] , \_2_net_[8] , \_2_net_[7] , \_2_net_[6] , \_2_net_[5] , 
        \_2_net_[4] , \_2_net_[3] , \_2_net_[2] , 1'b0, 1'b0}), .B({\w[2][31] , 
        \w[2][30] , \w[2][29] , \w[2][28] , \w[2][27] , \w[2][26] , \w[2][25] , 
        \w[2][24] , \w[2][23] , \w[2][22] , \w[2][21] , \w[2][20] , \w[2][19] , 
        \w[2][18] , \w[2][17] , \w[2][16] , \w[2][15] , \w[2][14] , \w[2][13] , 
        \w[2][12] , \w[2][11] , \w[2][10] , \w[2][9] , \w[2][8] , \w[2][7] , 
        \w[2][6] , \w[2][5] , \w[2][4] , \w[2][3] , \w[2][2] , \w[2][1] , 1'b0}), .CI(1'b0), .S({\w[3][31] , \w[3][30] , \w[3][29] , \w[3][28] , \w[3][27] , 
        \w[3][26] , \w[3][25] , \w[3][24] , \w[3][23] , \w[3][22] , \w[3][21] , 
        \w[3][20] , \w[3][19] , \w[3][18] , \w[3][17] , \w[3][16] , \w[3][15] , 
        \w[3][14] , \w[3][13] , \w[3][12] , \w[3][11] , \w[3][10] , \w[3][9] , 
        \w[3][8] , \w[3][7] , \w[3][6] , \w[3][5] , \w[3][4] , \w[3][3] , 
        \w[3][2] , \w[3][1] , SYNOPSYS_UNCONNECTED__1}) );
  ADD_N32_249 \FAINST[3].ADD_  ( .A({\_4_net_[31] , \_4_net_[30] , 
        \_4_net_[29] , \_4_net_[28] , \_4_net_[27] , \_4_net_[26] , 
        \_4_net_[25] , \_4_net_[24] , \_4_net_[23] , \_4_net_[22] , 
        \_4_net_[21] , \_4_net_[20] , \_4_net_[19] , \_4_net_[18] , 
        \_4_net_[17] , \_4_net_[16] , \_4_net_[15] , \_4_net_[14] , 
        \_4_net_[13] , \_4_net_[12] , \_4_net_[11] , \_4_net_[10] , 
        \_4_net_[9] , \_4_net_[8] , \_4_net_[7] , \_4_net_[6] , \_4_net_[5] , 
        \_4_net_[4] , \_4_net_[3] , 1'b0, 1'b0, 1'b0}), .B({\w[3][31] , 
        \w[3][30] , \w[3][29] , \w[3][28] , \w[3][27] , \w[3][26] , \w[3][25] , 
        \w[3][24] , \w[3][23] , \w[3][22] , \w[3][21] , \w[3][20] , \w[3][19] , 
        \w[3][18] , \w[3][17] , \w[3][16] , \w[3][15] , \w[3][14] , \w[3][13] , 
        \w[3][12] , \w[3][11] , \w[3][10] , \w[3][9] , \w[3][8] , \w[3][7] , 
        \w[3][6] , \w[3][5] , \w[3][4] , \w[3][3] , \w[3][2] , \w[3][1] , 1'b0}), .CI(1'b0), .S({\w[4][31] , \w[4][30] , \w[4][29] , \w[4][28] , \w[4][27] , 
        \w[4][26] , \w[4][25] , \w[4][24] , \w[4][23] , \w[4][22] , \w[4][21] , 
        \w[4][20] , \w[4][19] , \w[4][18] , \w[4][17] , \w[4][16] , \w[4][15] , 
        \w[4][14] , \w[4][13] , \w[4][12] , \w[4][11] , \w[4][10] , \w[4][9] , 
        \w[4][8] , \w[4][7] , \w[4][6] , \w[4][5] , \w[4][4] , \w[4][3] , 
        \w[4][2] , \w[4][1] , SYNOPSYS_UNCONNECTED__2}) );
  ADD_N32_248 \FAINST[4].ADD_  ( .A({\_6_net_[31] , \_6_net_[30] , 
        \_6_net_[29] , \_6_net_[28] , \_6_net_[27] , \_6_net_[26] , 
        \_6_net_[25] , \_6_net_[24] , \_6_net_[23] , \_6_net_[22] , 
        \_6_net_[21] , \_6_net_[20] , \_6_net_[19] , \_6_net_[18] , 
        \_6_net_[17] , \_6_net_[16] , \_6_net_[15] , \_6_net_[14] , 
        \_6_net_[13] , \_6_net_[12] , \_6_net_[11] , \_6_net_[10] , 
        \_6_net_[9] , \_6_net_[8] , \_6_net_[7] , \_6_net_[6] , \_6_net_[5] , 
        \_6_net_[4] , 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[4][31] , \w[4][30] , 
        \w[4][29] , \w[4][28] , \w[4][27] , \w[4][26] , \w[4][25] , \w[4][24] , 
        \w[4][23] , \w[4][22] , \w[4][21] , \w[4][20] , \w[4][19] , \w[4][18] , 
        \w[4][17] , \w[4][16] , \w[4][15] , \w[4][14] , \w[4][13] , \w[4][12] , 
        \w[4][11] , \w[4][10] , \w[4][9] , \w[4][8] , \w[4][7] , \w[4][6] , 
        \w[4][5] , \w[4][4] , \w[4][3] , \w[4][2] , \w[4][1] , 1'b0}), .CI(
        1'b0), .S({\w[5][31] , \w[5][30] , \w[5][29] , \w[5][28] , \w[5][27] , 
        \w[5][26] , \w[5][25] , \w[5][24] , \w[5][23] , \w[5][22] , \w[5][21] , 
        \w[5][20] , \w[5][19] , \w[5][18] , \w[5][17] , \w[5][16] , \w[5][15] , 
        \w[5][14] , \w[5][13] , \w[5][12] , \w[5][11] , \w[5][10] , \w[5][9] , 
        \w[5][8] , \w[5][7] , \w[5][6] , \w[5][5] , \w[5][4] , \w[5][3] , 
        \w[5][2] , \w[5][1] , SYNOPSYS_UNCONNECTED__3}) );
  ADD_N32_247 \FAINST[5].ADD_  ( .A({\_8_net_[31] , \_8_net_[30] , 
        \_8_net_[29] , \_8_net_[28] , \_8_net_[27] , \_8_net_[26] , 
        \_8_net_[25] , \_8_net_[24] , \_8_net_[23] , \_8_net_[22] , 
        \_8_net_[21] , \_8_net_[20] , \_8_net_[19] , \_8_net_[18] , 
        \_8_net_[17] , \_8_net_[16] , \_8_net_[15] , \_8_net_[14] , 
        \_8_net_[13] , \_8_net_[12] , \_8_net_[11] , \_8_net_[10] , 
        \_8_net_[9] , \_8_net_[8] , \_8_net_[7] , \_8_net_[6] , \_8_net_[5] , 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[5][31] , \w[5][30] , \w[5][29] , 
        \w[5][28] , \w[5][27] , \w[5][26] , \w[5][25] , \w[5][24] , \w[5][23] , 
        \w[5][22] , \w[5][21] , \w[5][20] , \w[5][19] , \w[5][18] , \w[5][17] , 
        \w[5][16] , \w[5][15] , \w[5][14] , \w[5][13] , \w[5][12] , \w[5][11] , 
        \w[5][10] , \w[5][9] , \w[5][8] , \w[5][7] , \w[5][6] , \w[5][5] , 
        \w[5][4] , \w[5][3] , \w[5][2] , \w[5][1] , 1'b0}), .CI(1'b0), .S({
        \w[6][31] , \w[6][30] , \w[6][29] , \w[6][28] , \w[6][27] , \w[6][26] , 
        \w[6][25] , \w[6][24] , \w[6][23] , \w[6][22] , \w[6][21] , \w[6][20] , 
        \w[6][19] , \w[6][18] , \w[6][17] , \w[6][16] , \w[6][15] , \w[6][14] , 
        \w[6][13] , \w[6][12] , \w[6][11] , \w[6][10] , \w[6][9] , \w[6][8] , 
        \w[6][7] , \w[6][6] , \w[6][5] , \w[6][4] , \w[6][3] , \w[6][2] , 
        \w[6][1] , SYNOPSYS_UNCONNECTED__4}) );
  ADD_N32_246 \FAINST[6].ADD_  ( .A({\_10_net_[31] , \_10_net_[30] , 
        \_10_net_[29] , \_10_net_[28] , \_10_net_[27] , \_10_net_[26] , 
        \_10_net_[25] , \_10_net_[24] , \_10_net_[23] , \_10_net_[22] , 
        \_10_net_[21] , \_10_net_[20] , \_10_net_[19] , \_10_net_[18] , 
        \_10_net_[17] , \_10_net_[16] , \_10_net_[15] , \_10_net_[14] , 
        \_10_net_[13] , \_10_net_[12] , \_10_net_[11] , \_10_net_[10] , 
        \_10_net_[9] , \_10_net_[8] , \_10_net_[7] , \_10_net_[6] , 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[6][31] , \w[6][30] , \w[6][29] , 
        \w[6][28] , \w[6][27] , \w[6][26] , \w[6][25] , \w[6][24] , \w[6][23] , 
        \w[6][22] , \w[6][21] , \w[6][20] , \w[6][19] , \w[6][18] , \w[6][17] , 
        \w[6][16] , \w[6][15] , \w[6][14] , \w[6][13] , \w[6][12] , \w[6][11] , 
        \w[6][10] , \w[6][9] , \w[6][8] , \w[6][7] , \w[6][6] , \w[6][5] , 
        \w[6][4] , \w[6][3] , \w[6][2] , \w[6][1] , 1'b0}), .CI(1'b0), .S({
        \w[7][31] , \w[7][30] , \w[7][29] , \w[7][28] , \w[7][27] , \w[7][26] , 
        \w[7][25] , \w[7][24] , \w[7][23] , \w[7][22] , \w[7][21] , \w[7][20] , 
        \w[7][19] , \w[7][18] , \w[7][17] , \w[7][16] , \w[7][15] , \w[7][14] , 
        \w[7][13] , \w[7][12] , \w[7][11] , \w[7][10] , \w[7][9] , \w[7][8] , 
        \w[7][7] , \w[7][6] , \w[7][5] , \w[7][4] , \w[7][3] , \w[7][2] , 
        \w[7][1] , SYNOPSYS_UNCONNECTED__5}) );
  ADD_N32_245 \FAINST[7].ADD_  ( .A({\_12_net_[31] , \_12_net_[30] , 
        \_12_net_[29] , \_12_net_[28] , \_12_net_[27] , \_12_net_[26] , 
        \_12_net_[25] , \_12_net_[24] , \_12_net_[23] , \_12_net_[22] , 
        \_12_net_[21] , \_12_net_[20] , \_12_net_[19] , \_12_net_[18] , 
        \_12_net_[17] , \_12_net_[16] , \_12_net_[15] , \_12_net_[14] , 
        \_12_net_[13] , \_12_net_[12] , \_12_net_[11] , \_12_net_[10] , 
        \_12_net_[9] , \_12_net_[8] , \_12_net_[7] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({\w[7][31] , \w[7][30] , \w[7][29] , \w[7][28] , 
        \w[7][27] , \w[7][26] , \w[7][25] , \w[7][24] , \w[7][23] , \w[7][22] , 
        \w[7][21] , \w[7][20] , \w[7][19] , \w[7][18] , \w[7][17] , \w[7][16] , 
        \w[7][15] , \w[7][14] , \w[7][13] , \w[7][12] , \w[7][11] , \w[7][10] , 
        \w[7][9] , \w[7][8] , \w[7][7] , \w[7][6] , \w[7][5] , \w[7][4] , 
        \w[7][3] , \w[7][2] , \w[7][1] , 1'b0}), .CI(1'b0), .S({\w[8][31] , 
        \w[8][30] , \w[8][29] , \w[8][28] , \w[8][27] , \w[8][26] , \w[8][25] , 
        \w[8][24] , \w[8][23] , \w[8][22] , \w[8][21] , \w[8][20] , \w[8][19] , 
        \w[8][18] , \w[8][17] , \w[8][16] , \w[8][15] , \w[8][14] , \w[8][13] , 
        \w[8][12] , \w[8][11] , \w[8][10] , \w[8][9] , \w[8][8] , \w[8][7] , 
        \w[8][6] , \w[8][5] , \w[8][4] , \w[8][3] , \w[8][2] , \w[8][1] , 
        SYNOPSYS_UNCONNECTED__6}) );
  ADD_N32_244 \FAINST[8].ADD_  ( .A({\_14_net_[31] , \_14_net_[30] , 
        \_14_net_[29] , \_14_net_[28] , \_14_net_[27] , \_14_net_[26] , 
        \_14_net_[25] , \_14_net_[24] , \_14_net_[23] , \_14_net_[22] , 
        \_14_net_[21] , \_14_net_[20] , \_14_net_[19] , \_14_net_[18] , 
        \_14_net_[17] , \_14_net_[16] , \_14_net_[15] , \_14_net_[14] , 
        \_14_net_[13] , \_14_net_[12] , \_14_net_[11] , \_14_net_[10] , 
        \_14_net_[9] , \_14_net_[8] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({\w[8][31] , \w[8][30] , \w[8][29] , \w[8][28] , \w[8][27] , 
        \w[8][26] , \w[8][25] , \w[8][24] , \w[8][23] , \w[8][22] , \w[8][21] , 
        \w[8][20] , \w[8][19] , \w[8][18] , \w[8][17] , \w[8][16] , \w[8][15] , 
        \w[8][14] , \w[8][13] , \w[8][12] , \w[8][11] , \w[8][10] , \w[8][9] , 
        \w[8][8] , \w[8][7] , \w[8][6] , \w[8][5] , \w[8][4] , \w[8][3] , 
        \w[8][2] , \w[8][1] , 1'b0}), .CI(1'b0), .S({\w[9][31] , \w[9][30] , 
        \w[9][29] , \w[9][28] , \w[9][27] , \w[9][26] , \w[9][25] , \w[9][24] , 
        \w[9][23] , \w[9][22] , \w[9][21] , \w[9][20] , \w[9][19] , \w[9][18] , 
        \w[9][17] , \w[9][16] , \w[9][15] , \w[9][14] , \w[9][13] , \w[9][12] , 
        \w[9][11] , \w[9][10] , \w[9][9] , \w[9][8] , \w[9][7] , \w[9][6] , 
        \w[9][5] , \w[9][4] , \w[9][3] , \w[9][2] , \w[9][1] , 
        SYNOPSYS_UNCONNECTED__7}) );
  ADD_N32_243 \FAINST[9].ADD_  ( .A({\_16_net_[31] , \_16_net_[30] , 
        \_16_net_[29] , \_16_net_[28] , \_16_net_[27] , \_16_net_[26] , 
        \_16_net_[25] , \_16_net_[24] , \_16_net_[23] , \_16_net_[22] , 
        \_16_net_[21] , \_16_net_[20] , \_16_net_[19] , \_16_net_[18] , 
        \_16_net_[17] , \_16_net_[16] , \_16_net_[15] , \_16_net_[14] , 
        \_16_net_[13] , \_16_net_[12] , \_16_net_[11] , \_16_net_[10] , 
        \_16_net_[9] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({\w[9][31] , \w[9][30] , \w[9][29] , \w[9][28] , \w[9][27] , 
        \w[9][26] , \w[9][25] , \w[9][24] , \w[9][23] , \w[9][22] , \w[9][21] , 
        \w[9][20] , \w[9][19] , \w[9][18] , \w[9][17] , \w[9][16] , \w[9][15] , 
        \w[9][14] , \w[9][13] , \w[9][12] , \w[9][11] , \w[9][10] , \w[9][9] , 
        \w[9][8] , \w[9][7] , \w[9][6] , \w[9][5] , \w[9][4] , \w[9][3] , 
        \w[9][2] , \w[9][1] , 1'b0}), .CI(1'b0), .S({\w[10][31] , \w[10][30] , 
        \w[10][29] , \w[10][28] , \w[10][27] , \w[10][26] , \w[10][25] , 
        \w[10][24] , \w[10][23] , \w[10][22] , \w[10][21] , \w[10][20] , 
        \w[10][19] , \w[10][18] , \w[10][17] , \w[10][16] , \w[10][15] , 
        \w[10][14] , \w[10][13] , \w[10][12] , \w[10][11] , \w[10][10] , 
        \w[10][9] , \w[10][8] , \w[10][7] , \w[10][6] , \w[10][5] , \w[10][4] , 
        \w[10][3] , \w[10][2] , \w[10][1] , SYNOPSYS_UNCONNECTED__8}) );
  ADD_N32_242 \FAINST[10].ADD_  ( .A({\_18_net_[31] , \_18_net_[30] , 
        \_18_net_[29] , \_18_net_[28] , \_18_net_[27] , \_18_net_[26] , 
        \_18_net_[25] , \_18_net_[24] , \_18_net_[23] , \_18_net_[22] , 
        \_18_net_[21] , \_18_net_[20] , \_18_net_[19] , \_18_net_[18] , 
        \_18_net_[17] , \_18_net_[16] , \_18_net_[15] , \_18_net_[14] , 
        \_18_net_[13] , \_18_net_[12] , \_18_net_[11] , \_18_net_[10] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[10][31] , \w[10][30] , \w[10][29] , \w[10][28] , \w[10][27] , 
        \w[10][26] , \w[10][25] , \w[10][24] , \w[10][23] , \w[10][22] , 
        \w[10][21] , \w[10][20] , \w[10][19] , \w[10][18] , \w[10][17] , 
        \w[10][16] , \w[10][15] , \w[10][14] , \w[10][13] , \w[10][12] , 
        \w[10][11] , \w[10][10] , \w[10][9] , \w[10][8] , \w[10][7] , 
        \w[10][6] , \w[10][5] , \w[10][4] , \w[10][3] , \w[10][2] , \w[10][1] , 
        1'b0}), .CI(1'b0), .S({\w[11][31] , \w[11][30] , \w[11][29] , 
        \w[11][28] , \w[11][27] , \w[11][26] , \w[11][25] , \w[11][24] , 
        \w[11][23] , \w[11][22] , \w[11][21] , \w[11][20] , \w[11][19] , 
        \w[11][18] , \w[11][17] , \w[11][16] , \w[11][15] , \w[11][14] , 
        \w[11][13] , \w[11][12] , \w[11][11] , \w[11][10] , \w[11][9] , 
        \w[11][8] , \w[11][7] , \w[11][6] , \w[11][5] , \w[11][4] , \w[11][3] , 
        \w[11][2] , \w[11][1] , SYNOPSYS_UNCONNECTED__9}) );
  ADD_N32_241 \FAINST[11].ADD_  ( .A({\_20_net_[31] , \_20_net_[30] , 
        \_20_net_[29] , \_20_net_[28] , \_20_net_[27] , \_20_net_[26] , 
        \_20_net_[25] , \_20_net_[24] , \_20_net_[23] , \_20_net_[22] , 
        \_20_net_[21] , \_20_net_[20] , \_20_net_[19] , \_20_net_[18] , 
        \_20_net_[17] , \_20_net_[16] , \_20_net_[15] , \_20_net_[14] , 
        \_20_net_[13] , \_20_net_[12] , \_20_net_[11] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[11][31] , 
        \w[11][30] , \w[11][29] , \w[11][28] , \w[11][27] , \w[11][26] , 
        \w[11][25] , \w[11][24] , \w[11][23] , \w[11][22] , \w[11][21] , 
        \w[11][20] , \w[11][19] , \w[11][18] , \w[11][17] , \w[11][16] , 
        \w[11][15] , \w[11][14] , \w[11][13] , \w[11][12] , \w[11][11] , 
        \w[11][10] , \w[11][9] , \w[11][8] , \w[11][7] , \w[11][6] , 
        \w[11][5] , \w[11][4] , \w[11][3] , \w[11][2] , \w[11][1] , 1'b0}), 
        .CI(1'b0), .S({\w[12][31] , \w[12][30] , \w[12][29] , \w[12][28] , 
        \w[12][27] , \w[12][26] , \w[12][25] , \w[12][24] , \w[12][23] , 
        \w[12][22] , \w[12][21] , \w[12][20] , \w[12][19] , \w[12][18] , 
        \w[12][17] , \w[12][16] , \w[12][15] , \w[12][14] , \w[12][13] , 
        \w[12][12] , \w[12][11] , \w[12][10] , \w[12][9] , \w[12][8] , 
        \w[12][7] , \w[12][6] , \w[12][5] , \w[12][4] , \w[12][3] , \w[12][2] , 
        \w[12][1] , SYNOPSYS_UNCONNECTED__10}) );
  ADD_N32_240 \FAINST[12].ADD_  ( .A({\_22_net_[31] , \_22_net_[30] , 
        \_22_net_[29] , \_22_net_[28] , \_22_net_[27] , \_22_net_[26] , 
        \_22_net_[25] , \_22_net_[24] , \_22_net_[23] , \_22_net_[22] , 
        \_22_net_[21] , \_22_net_[20] , \_22_net_[19] , \_22_net_[18] , 
        \_22_net_[17] , \_22_net_[16] , \_22_net_[15] , \_22_net_[14] , 
        \_22_net_[13] , \_22_net_[12] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[12][31] , \w[12][30] , 
        \w[12][29] , \w[12][28] , \w[12][27] , \w[12][26] , \w[12][25] , 
        \w[12][24] , \w[12][23] , \w[12][22] , \w[12][21] , \w[12][20] , 
        \w[12][19] , \w[12][18] , \w[12][17] , \w[12][16] , \w[12][15] , 
        \w[12][14] , \w[12][13] , \w[12][12] , \w[12][11] , \w[12][10] , 
        \w[12][9] , \w[12][8] , \w[12][7] , \w[12][6] , \w[12][5] , \w[12][4] , 
        \w[12][3] , \w[12][2] , \w[12][1] , 1'b0}), .CI(1'b0), .S({\w[13][31] , 
        \w[13][30] , \w[13][29] , \w[13][28] , \w[13][27] , \w[13][26] , 
        \w[13][25] , \w[13][24] , \w[13][23] , \w[13][22] , \w[13][21] , 
        \w[13][20] , \w[13][19] , \w[13][18] , \w[13][17] , \w[13][16] , 
        \w[13][15] , \w[13][14] , \w[13][13] , \w[13][12] , \w[13][11] , 
        \w[13][10] , \w[13][9] , \w[13][8] , \w[13][7] , \w[13][6] , 
        \w[13][5] , \w[13][4] , \w[13][3] , \w[13][2] , \w[13][1] , 
        SYNOPSYS_UNCONNECTED__11}) );
  ADD_N32_239 \FAINST[13].ADD_  ( .A({\_24_net_[31] , \_24_net_[30] , 
        \_24_net_[29] , \_24_net_[28] , \_24_net_[27] , \_24_net_[26] , 
        \_24_net_[25] , \_24_net_[24] , \_24_net_[23] , \_24_net_[22] , 
        \_24_net_[21] , \_24_net_[20] , \_24_net_[19] , \_24_net_[18] , 
        \_24_net_[17] , \_24_net_[16] , \_24_net_[15] , \_24_net_[14] , 
        \_24_net_[13] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[13][31] , \w[13][30] , \w[13][29] , 
        \w[13][28] , \w[13][27] , \w[13][26] , \w[13][25] , \w[13][24] , 
        \w[13][23] , \w[13][22] , \w[13][21] , \w[13][20] , \w[13][19] , 
        \w[13][18] , \w[13][17] , \w[13][16] , \w[13][15] , \w[13][14] , 
        \w[13][13] , \w[13][12] , \w[13][11] , \w[13][10] , \w[13][9] , 
        \w[13][8] , \w[13][7] , \w[13][6] , \w[13][5] , \w[13][4] , \w[13][3] , 
        \w[13][2] , \w[13][1] , 1'b0}), .CI(1'b0), .S({\w[14][31] , 
        \w[14][30] , \w[14][29] , \w[14][28] , \w[14][27] , \w[14][26] , 
        \w[14][25] , \w[14][24] , \w[14][23] , \w[14][22] , \w[14][21] , 
        \w[14][20] , \w[14][19] , \w[14][18] , \w[14][17] , \w[14][16] , 
        \w[14][15] , \w[14][14] , \w[14][13] , \w[14][12] , \w[14][11] , 
        \w[14][10] , \w[14][9] , \w[14][8] , \w[14][7] , \w[14][6] , 
        \w[14][5] , \w[14][4] , \w[14][3] , \w[14][2] , \w[14][1] , 
        SYNOPSYS_UNCONNECTED__12}) );
  ADD_N32_238 \FAINST[14].ADD_  ( .A({\_26_net_[31] , \_26_net_[30] , 
        \_26_net_[29] , \_26_net_[28] , \_26_net_[27] , \_26_net_[26] , 
        \_26_net_[25] , \_26_net_[24] , \_26_net_[23] , \_26_net_[22] , 
        \_26_net_[21] , \_26_net_[20] , \_26_net_[19] , \_26_net_[18] , 
        \_26_net_[17] , \_26_net_[16] , \_26_net_[15] , \_26_net_[14] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({\w[14][31] , \w[14][30] , \w[14][29] , \w[14][28] , 
        \w[14][27] , \w[14][26] , \w[14][25] , \w[14][24] , \w[14][23] , 
        \w[14][22] , \w[14][21] , \w[14][20] , \w[14][19] , \w[14][18] , 
        \w[14][17] , \w[14][16] , \w[14][15] , \w[14][14] , \w[14][13] , 
        \w[14][12] , \w[14][11] , \w[14][10] , \w[14][9] , \w[14][8] , 
        \w[14][7] , \w[14][6] , \w[14][5] , \w[14][4] , \w[14][3] , \w[14][2] , 
        \w[14][1] , 1'b0}), .CI(1'b0), .S({\w[15][31] , \w[15][30] , 
        \w[15][29] , \w[15][28] , \w[15][27] , \w[15][26] , \w[15][25] , 
        \w[15][24] , \w[15][23] , \w[15][22] , \w[15][21] , \w[15][20] , 
        \w[15][19] , \w[15][18] , \w[15][17] , \w[15][16] , \w[15][15] , 
        \w[15][14] , \w[15][13] , \w[15][12] , \w[15][11] , \w[15][10] , 
        \w[15][9] , \w[15][8] , \w[15][7] , \w[15][6] , \w[15][5] , \w[15][4] , 
        \w[15][3] , \w[15][2] , \w[15][1] , SYNOPSYS_UNCONNECTED__13}) );
  ADD_N32_237 \FAINST[15].ADD_  ( .A({\_28_net_[31] , \_28_net_[30] , 
        \_28_net_[29] , \_28_net_[28] , \_28_net_[27] , \_28_net_[26] , 
        \_28_net_[25] , \_28_net_[24] , \_28_net_[23] , \_28_net_[22] , 
        \_28_net_[21] , \_28_net_[20] , \_28_net_[19] , \_28_net_[18] , 
        \_28_net_[17] , \_28_net_[16] , \_28_net_[15] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({\w[15][31] , \w[15][30] , \w[15][29] , \w[15][28] , \w[15][27] , 
        \w[15][26] , \w[15][25] , \w[15][24] , \w[15][23] , \w[15][22] , 
        \w[15][21] , \w[15][20] , \w[15][19] , \w[15][18] , \w[15][17] , 
        \w[15][16] , \w[15][15] , \w[15][14] , \w[15][13] , \w[15][12] , 
        \w[15][11] , \w[15][10] , \w[15][9] , \w[15][8] , \w[15][7] , 
        \w[15][6] , \w[15][5] , \w[15][4] , \w[15][3] , \w[15][2] , \w[15][1] , 
        1'b0}), .CI(1'b0), .S({\w[16][31] , \w[16][30] , \w[16][29] , 
        \w[16][28] , \w[16][27] , \w[16][26] , \w[16][25] , \w[16][24] , 
        \w[16][23] , \w[16][22] , \w[16][21] , \w[16][20] , \w[16][19] , 
        \w[16][18] , \w[16][17] , \w[16][16] , \w[16][15] , \w[16][14] , 
        \w[16][13] , \w[16][12] , \w[16][11] , \w[16][10] , \w[16][9] , 
        \w[16][8] , \w[16][7] , \w[16][6] , \w[16][5] , \w[16][4] , \w[16][3] , 
        \w[16][2] , \w[16][1] , SYNOPSYS_UNCONNECTED__14}) );
  ADD_N32_236 \FAINST[16].ADD_  ( .A({\_30_net_[31] , \_30_net_[30] , 
        \_30_net_[29] , \_30_net_[28] , \_30_net_[27] , \_30_net_[26] , 
        \_30_net_[25] , \_30_net_[24] , \_30_net_[23] , \_30_net_[22] , 
        \_30_net_[21] , \_30_net_[20] , \_30_net_[19] , \_30_net_[18] , 
        \_30_net_[17] , \_30_net_[16] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[16][31] , \w[16][30] , \w[16][29] , \w[16][28] , \w[16][27] , 
        \w[16][26] , \w[16][25] , \w[16][24] , \w[16][23] , \w[16][22] , 
        \w[16][21] , \w[16][20] , \w[16][19] , \w[16][18] , \w[16][17] , 
        \w[16][16] , \w[16][15] , \w[16][14] , \w[16][13] , \w[16][12] , 
        \w[16][11] , \w[16][10] , \w[16][9] , \w[16][8] , \w[16][7] , 
        \w[16][6] , \w[16][5] , \w[16][4] , \w[16][3] , \w[16][2] , \w[16][1] , 
        1'b0}), .CI(1'b0), .S({\w[17][31] , \w[17][30] , \w[17][29] , 
        \w[17][28] , \w[17][27] , \w[17][26] , \w[17][25] , \w[17][24] , 
        \w[17][23] , \w[17][22] , \w[17][21] , \w[17][20] , \w[17][19] , 
        \w[17][18] , \w[17][17] , \w[17][16] , \w[17][15] , \w[17][14] , 
        \w[17][13] , \w[17][12] , \w[17][11] , \w[17][10] , \w[17][9] , 
        \w[17][8] , \w[17][7] , \w[17][6] , \w[17][5] , \w[17][4] , \w[17][3] , 
        \w[17][2] , \w[17][1] , SYNOPSYS_UNCONNECTED__15}) );
  ADD_N32_235 \FAINST[17].ADD_  ( .A({\_32_net_[31] , \_32_net_[30] , 
        \_32_net_[29] , \_32_net_[28] , \_32_net_[27] , \_32_net_[26] , 
        \_32_net_[25] , \_32_net_[24] , \_32_net_[23] , \_32_net_[22] , 
        \_32_net_[21] , \_32_net_[20] , \_32_net_[19] , \_32_net_[18] , 
        \_32_net_[17] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[17][31] , 
        \w[17][30] , \w[17][29] , \w[17][28] , \w[17][27] , \w[17][26] , 
        \w[17][25] , \w[17][24] , \w[17][23] , \w[17][22] , \w[17][21] , 
        \w[17][20] , \w[17][19] , \w[17][18] , \w[17][17] , \w[17][16] , 
        \w[17][15] , \w[17][14] , \w[17][13] , \w[17][12] , \w[17][11] , 
        \w[17][10] , \w[17][9] , \w[17][8] , \w[17][7] , \w[17][6] , 
        \w[17][5] , \w[17][4] , \w[17][3] , \w[17][2] , \w[17][1] , 1'b0}), 
        .CI(1'b0), .S({\w[18][31] , \w[18][30] , \w[18][29] , \w[18][28] , 
        \w[18][27] , \w[18][26] , \w[18][25] , \w[18][24] , \w[18][23] , 
        \w[18][22] , \w[18][21] , \w[18][20] , \w[18][19] , \w[18][18] , 
        \w[18][17] , \w[18][16] , \w[18][15] , \w[18][14] , \w[18][13] , 
        \w[18][12] , \w[18][11] , \w[18][10] , \w[18][9] , \w[18][8] , 
        \w[18][7] , \w[18][6] , \w[18][5] , \w[18][4] , \w[18][3] , \w[18][2] , 
        \w[18][1] , SYNOPSYS_UNCONNECTED__16}) );
  ADD_N32_234 \FAINST[18].ADD_  ( .A({\_34_net_[31] , \_34_net_[30] , 
        \_34_net_[29] , \_34_net_[28] , \_34_net_[27] , \_34_net_[26] , 
        \_34_net_[25] , \_34_net_[24] , \_34_net_[23] , \_34_net_[22] , 
        \_34_net_[21] , \_34_net_[20] , \_34_net_[19] , \_34_net_[18] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[18][31] , \w[18][30] , 
        \w[18][29] , \w[18][28] , \w[18][27] , \w[18][26] , \w[18][25] , 
        \w[18][24] , \w[18][23] , \w[18][22] , \w[18][21] , \w[18][20] , 
        \w[18][19] , \w[18][18] , \w[18][17] , \w[18][16] , \w[18][15] , 
        \w[18][14] , \w[18][13] , \w[18][12] , \w[18][11] , \w[18][10] , 
        \w[18][9] , \w[18][8] , \w[18][7] , \w[18][6] , \w[18][5] , \w[18][4] , 
        \w[18][3] , \w[18][2] , \w[18][1] , 1'b0}), .CI(1'b0), .S({\w[19][31] , 
        \w[19][30] , \w[19][29] , \w[19][28] , \w[19][27] , \w[19][26] , 
        \w[19][25] , \w[19][24] , \w[19][23] , \w[19][22] , \w[19][21] , 
        \w[19][20] , \w[19][19] , \w[19][18] , \w[19][17] , \w[19][16] , 
        \w[19][15] , \w[19][14] , \w[19][13] , \w[19][12] , \w[19][11] , 
        \w[19][10] , \w[19][9] , \w[19][8] , \w[19][7] , \w[19][6] , 
        \w[19][5] , \w[19][4] , \w[19][3] , \w[19][2] , \w[19][1] , 
        SYNOPSYS_UNCONNECTED__17}) );
  ADD_N32_233 \FAINST[19].ADD_  ( .A({\_36_net_[31] , \_36_net_[30] , 
        \_36_net_[29] , \_36_net_[28] , \_36_net_[27] , \_36_net_[26] , 
        \_36_net_[25] , \_36_net_[24] , \_36_net_[23] , \_36_net_[22] , 
        \_36_net_[21] , \_36_net_[20] , \_36_net_[19] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({\w[19][31] , \w[19][30] , \w[19][29] , 
        \w[19][28] , \w[19][27] , \w[19][26] , \w[19][25] , \w[19][24] , 
        \w[19][23] , \w[19][22] , \w[19][21] , \w[19][20] , \w[19][19] , 
        \w[19][18] , \w[19][17] , \w[19][16] , \w[19][15] , \w[19][14] , 
        \w[19][13] , \w[19][12] , \w[19][11] , \w[19][10] , \w[19][9] , 
        \w[19][8] , \w[19][7] , \w[19][6] , \w[19][5] , \w[19][4] , \w[19][3] , 
        \w[19][2] , \w[19][1] , 1'b0}), .CI(1'b0), .S({\w[20][31] , 
        \w[20][30] , \w[20][29] , \w[20][28] , \w[20][27] , \w[20][26] , 
        \w[20][25] , \w[20][24] , \w[20][23] , \w[20][22] , \w[20][21] , 
        \w[20][20] , \w[20][19] , \w[20][18] , \w[20][17] , \w[20][16] , 
        \w[20][15] , \w[20][14] , \w[20][13] , \w[20][12] , \w[20][11] , 
        \w[20][10] , \w[20][9] , \w[20][8] , \w[20][7] , \w[20][6] , 
        \w[20][5] , \w[20][4] , \w[20][3] , \w[20][2] , \w[20][1] , 
        SYNOPSYS_UNCONNECTED__18}) );
  ADD_N32_232 \FAINST[20].ADD_  ( .A({\_38_net_[31] , \_38_net_[30] , 
        \_38_net_[29] , \_38_net_[28] , \_38_net_[27] , \_38_net_[26] , 
        \_38_net_[25] , \_38_net_[24] , \_38_net_[23] , \_38_net_[22] , 
        \_38_net_[21] , \_38_net_[20] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .B({\w[20][31] , \w[20][30] , \w[20][29] , \w[20][28] , 
        \w[20][27] , \w[20][26] , \w[20][25] , \w[20][24] , \w[20][23] , 
        \w[20][22] , \w[20][21] , \w[20][20] , \w[20][19] , \w[20][18] , 
        \w[20][17] , \w[20][16] , \w[20][15] , \w[20][14] , \w[20][13] , 
        \w[20][12] , \w[20][11] , \w[20][10] , \w[20][9] , \w[20][8] , 
        \w[20][7] , \w[20][6] , \w[20][5] , \w[20][4] , \w[20][3] , \w[20][2] , 
        \w[20][1] , 1'b0}), .CI(1'b0), .S({\w[21][31] , \w[21][30] , 
        \w[21][29] , \w[21][28] , \w[21][27] , \w[21][26] , \w[21][25] , 
        \w[21][24] , \w[21][23] , \w[21][22] , \w[21][21] , \w[21][20] , 
        \w[21][19] , \w[21][18] , \w[21][17] , \w[21][16] , \w[21][15] , 
        \w[21][14] , \w[21][13] , \w[21][12] , \w[21][11] , \w[21][10] , 
        \w[21][9] , \w[21][8] , \w[21][7] , \w[21][6] , \w[21][5] , \w[21][4] , 
        \w[21][3] , \w[21][2] , \w[21][1] , SYNOPSYS_UNCONNECTED__19}) );
  ADD_N32_231 \FAINST[21].ADD_  ( .A({\_40_net_[31] , \_40_net_[30] , 
        \_40_net_[29] , \_40_net_[28] , \_40_net_[27] , \_40_net_[26] , 
        \_40_net_[25] , \_40_net_[24] , \_40_net_[23] , \_40_net_[22] , 
        \_40_net_[21] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[21][31] , \w[21][30] , \w[21][29] , \w[21][28] , \w[21][27] , 
        \w[21][26] , \w[21][25] , \w[21][24] , \w[21][23] , \w[21][22] , 
        \w[21][21] , \w[21][20] , \w[21][19] , \w[21][18] , \w[21][17] , 
        \w[21][16] , \w[21][15] , \w[21][14] , \w[21][13] , \w[21][12] , 
        \w[21][11] , \w[21][10] , \w[21][9] , \w[21][8] , \w[21][7] , 
        \w[21][6] , \w[21][5] , \w[21][4] , \w[21][3] , \w[21][2] , \w[21][1] , 
        1'b0}), .CI(1'b0), .S({\w[22][31] , \w[22][30] , \w[22][29] , 
        \w[22][28] , \w[22][27] , \w[22][26] , \w[22][25] , \w[22][24] , 
        \w[22][23] , \w[22][22] , \w[22][21] , \w[22][20] , \w[22][19] , 
        \w[22][18] , \w[22][17] , \w[22][16] , \w[22][15] , \w[22][14] , 
        \w[22][13] , \w[22][12] , \w[22][11] , \w[22][10] , \w[22][9] , 
        \w[22][8] , \w[22][7] , \w[22][6] , \w[22][5] , \w[22][4] , \w[22][3] , 
        \w[22][2] , \w[22][1] , SYNOPSYS_UNCONNECTED__20}) );
  ADD_N32_230 \FAINST[22].ADD_  ( .A({\_42_net_[31] , \_42_net_[30] , 
        \_42_net_[29] , \_42_net_[28] , \_42_net_[27] , \_42_net_[26] , 
        \_42_net_[25] , \_42_net_[24] , \_42_net_[23] , \_42_net_[22] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[22][31] , \w[22][30] , \w[22][29] , \w[22][28] , \w[22][27] , 
        \w[22][26] , \w[22][25] , \w[22][24] , \w[22][23] , \w[22][22] , 
        \w[22][21] , \w[22][20] , \w[22][19] , \w[22][18] , \w[22][17] , 
        \w[22][16] , \w[22][15] , \w[22][14] , \w[22][13] , \w[22][12] , 
        \w[22][11] , \w[22][10] , \w[22][9] , \w[22][8] , \w[22][7] , 
        \w[22][6] , \w[22][5] , \w[22][4] , \w[22][3] , \w[22][2] , \w[22][1] , 
        1'b0}), .CI(1'b0), .S({\w[23][31] , \w[23][30] , \w[23][29] , 
        \w[23][28] , \w[23][27] , \w[23][26] , \w[23][25] , \w[23][24] , 
        \w[23][23] , \w[23][22] , \w[23][21] , \w[23][20] , \w[23][19] , 
        \w[23][18] , \w[23][17] , \w[23][16] , \w[23][15] , \w[23][14] , 
        \w[23][13] , \w[23][12] , \w[23][11] , \w[23][10] , \w[23][9] , 
        \w[23][8] , \w[23][7] , \w[23][6] , \w[23][5] , \w[23][4] , \w[23][3] , 
        \w[23][2] , \w[23][1] , SYNOPSYS_UNCONNECTED__21}) );
  ADD_N32_229 \FAINST[23].ADD_  ( .A({\_44_net_[31] , \_44_net_[30] , 
        \_44_net_[29] , \_44_net_[28] , \_44_net_[27] , \_44_net_[26] , 
        \_44_net_[25] , \_44_net_[24] , \_44_net_[23] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[23][31] , 
        \w[23][30] , \w[23][29] , \w[23][28] , \w[23][27] , \w[23][26] , 
        \w[23][25] , \w[23][24] , \w[23][23] , \w[23][22] , \w[23][21] , 
        \w[23][20] , \w[23][19] , \w[23][18] , \w[23][17] , \w[23][16] , 
        \w[23][15] , \w[23][14] , \w[23][13] , \w[23][12] , \w[23][11] , 
        \w[23][10] , \w[23][9] , \w[23][8] , \w[23][7] , \w[23][6] , 
        \w[23][5] , \w[23][4] , \w[23][3] , \w[23][2] , \w[23][1] , 1'b0}), 
        .CI(1'b0), .S({\w[24][31] , \w[24][30] , \w[24][29] , \w[24][28] , 
        \w[24][27] , \w[24][26] , \w[24][25] , \w[24][24] , \w[24][23] , 
        \w[24][22] , \w[24][21] , \w[24][20] , \w[24][19] , \w[24][18] , 
        \w[24][17] , \w[24][16] , \w[24][15] , \w[24][14] , \w[24][13] , 
        \w[24][12] , \w[24][11] , \w[24][10] , \w[24][9] , \w[24][8] , 
        \w[24][7] , \w[24][6] , \w[24][5] , \w[24][4] , \w[24][3] , \w[24][2] , 
        \w[24][1] , SYNOPSYS_UNCONNECTED__22}) );
  ADD_N32_228 \FAINST[24].ADD_  ( .A({\_46_net_[31] , \_46_net_[30] , 
        \_46_net_[29] , \_46_net_[28] , \_46_net_[27] , \_46_net_[26] , 
        \_46_net_[25] , \_46_net_[24] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[24][31] , \w[24][30] , 
        \w[24][29] , \w[24][28] , \w[24][27] , \w[24][26] , \w[24][25] , 
        \w[24][24] , \w[24][23] , \w[24][22] , \w[24][21] , \w[24][20] , 
        \w[24][19] , \w[24][18] , \w[24][17] , \w[24][16] , \w[24][15] , 
        \w[24][14] , \w[24][13] , \w[24][12] , \w[24][11] , \w[24][10] , 
        \w[24][9] , \w[24][8] , \w[24][7] , \w[24][6] , \w[24][5] , \w[24][4] , 
        \w[24][3] , \w[24][2] , \w[24][1] , 1'b0}), .CI(1'b0), .S({\w[25][31] , 
        \w[25][30] , \w[25][29] , \w[25][28] , \w[25][27] , \w[25][26] , 
        \w[25][25] , \w[25][24] , \w[25][23] , \w[25][22] , \w[25][21] , 
        \w[25][20] , \w[25][19] , \w[25][18] , \w[25][17] , \w[25][16] , 
        \w[25][15] , \w[25][14] , \w[25][13] , \w[25][12] , \w[25][11] , 
        \w[25][10] , \w[25][9] , \w[25][8] , \w[25][7] , \w[25][6] , 
        \w[25][5] , \w[25][4] , \w[25][3] , \w[25][2] , \w[25][1] , 
        SYNOPSYS_UNCONNECTED__23}) );
  ADD_N32_227 \FAINST[25].ADD_  ( .A({\_48_net_[31] , \_48_net_[30] , 
        \_48_net_[29] , \_48_net_[28] , \_48_net_[27] , \_48_net_[26] , 
        \_48_net_[25] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[25][31] , \w[25][30] , \w[25][29] , 
        \w[25][28] , \w[25][27] , \w[25][26] , \w[25][25] , \w[25][24] , 
        \w[25][23] , \w[25][22] , \w[25][21] , \w[25][20] , \w[25][19] , 
        \w[25][18] , \w[25][17] , \w[25][16] , \w[25][15] , \w[25][14] , 
        \w[25][13] , \w[25][12] , \w[25][11] , \w[25][10] , \w[25][9] , 
        \w[25][8] , \w[25][7] , \w[25][6] , \w[25][5] , \w[25][4] , \w[25][3] , 
        \w[25][2] , \w[25][1] , 1'b0}), .CI(1'b0), .S({\w[26][31] , 
        \w[26][30] , \w[26][29] , \w[26][28] , \w[26][27] , \w[26][26] , 
        \w[26][25] , \w[26][24] , \w[26][23] , \w[26][22] , \w[26][21] , 
        \w[26][20] , \w[26][19] , \w[26][18] , \w[26][17] , \w[26][16] , 
        \w[26][15] , \w[26][14] , \w[26][13] , \w[26][12] , \w[26][11] , 
        \w[26][10] , \w[26][9] , \w[26][8] , \w[26][7] , \w[26][6] , 
        \w[26][5] , \w[26][4] , \w[26][3] , \w[26][2] , \w[26][1] , 
        SYNOPSYS_UNCONNECTED__24}) );
  ADD_N32_226 \FAINST[26].ADD_  ( .A({\_50_net_[31] , \_50_net_[30] , 
        \_50_net_[29] , \_50_net_[28] , \_50_net_[27] , \_50_net_[26] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({\w[26][31] , \w[26][30] , \w[26][29] , \w[26][28] , 
        \w[26][27] , \w[26][26] , \w[26][25] , \w[26][24] , \w[26][23] , 
        \w[26][22] , \w[26][21] , \w[26][20] , \w[26][19] , \w[26][18] , 
        \w[26][17] , \w[26][16] , \w[26][15] , \w[26][14] , \w[26][13] , 
        \w[26][12] , \w[26][11] , \w[26][10] , \w[26][9] , \w[26][8] , 
        \w[26][7] , \w[26][6] , \w[26][5] , \w[26][4] , \w[26][3] , \w[26][2] , 
        \w[26][1] , 1'b0}), .CI(1'b0), .S({\w[27][31] , \w[27][30] , 
        \w[27][29] , \w[27][28] , \w[27][27] , \w[27][26] , \w[27][25] , 
        \w[27][24] , \w[27][23] , \w[27][22] , \w[27][21] , \w[27][20] , 
        \w[27][19] , \w[27][18] , \w[27][17] , \w[27][16] , \w[27][15] , 
        \w[27][14] , \w[27][13] , \w[27][12] , \w[27][11] , \w[27][10] , 
        \w[27][9] , \w[27][8] , \w[27][7] , \w[27][6] , \w[27][5] , \w[27][4] , 
        \w[27][3] , \w[27][2] , \w[27][1] , SYNOPSYS_UNCONNECTED__25}) );
  ADD_N32_225 \FAINST[27].ADD_  ( .A({\_52_net_[31] , \_52_net_[30] , 
        \_52_net_[29] , \_52_net_[28] , \_52_net_[27] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({\w[27][31] , \w[27][30] , \w[27][29] , \w[27][28] , \w[27][27] , 
        \w[27][26] , \w[27][25] , \w[27][24] , \w[27][23] , \w[27][22] , 
        \w[27][21] , \w[27][20] , \w[27][19] , \w[27][18] , \w[27][17] , 
        \w[27][16] , \w[27][15] , \w[27][14] , \w[27][13] , \w[27][12] , 
        \w[27][11] , \w[27][10] , \w[27][9] , \w[27][8] , \w[27][7] , 
        \w[27][6] , \w[27][5] , \w[27][4] , \w[27][3] , \w[27][2] , \w[27][1] , 
        1'b0}), .CI(1'b0), .S({\w[28][31] , \w[28][30] , \w[28][29] , 
        \w[28][28] , \w[28][27] , \w[28][26] , \w[28][25] , \w[28][24] , 
        \w[28][23] , \w[28][22] , \w[28][21] , \w[28][20] , \w[28][19] , 
        \w[28][18] , \w[28][17] , \w[28][16] , \w[28][15] , \w[28][14] , 
        \w[28][13] , \w[28][12] , \w[28][11] , \w[28][10] , \w[28][9] , 
        \w[28][8] , \w[28][7] , \w[28][6] , \w[28][5] , \w[28][4] , \w[28][3] , 
        \w[28][2] , \w[28][1] , SYNOPSYS_UNCONNECTED__26}) );
  ADD_N32_224 \FAINST[28].ADD_  ( .A({\_54_net_[31] , \_54_net_[30] , 
        \_54_net_[29] , \_54_net_[28] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[28][31] , \w[28][30] , \w[28][29] , \w[28][28] , \w[28][27] , 
        \w[28][26] , \w[28][25] , \w[28][24] , \w[28][23] , \w[28][22] , 
        \w[28][21] , \w[28][20] , \w[28][19] , \w[28][18] , \w[28][17] , 
        \w[28][16] , \w[28][15] , \w[28][14] , \w[28][13] , \w[28][12] , 
        \w[28][11] , \w[28][10] , \w[28][9] , \w[28][8] , \w[28][7] , 
        \w[28][6] , \w[28][5] , \w[28][4] , \w[28][3] , \w[28][2] , \w[28][1] , 
        1'b0}), .CI(1'b0), .S({\w[29][31] , \w[29][30] , \w[29][29] , 
        \w[29][28] , \w[29][27] , \w[29][26] , \w[29][25] , \w[29][24] , 
        \w[29][23] , \w[29][22] , \w[29][21] , \w[29][20] , \w[29][19] , 
        \w[29][18] , \w[29][17] , \w[29][16] , \w[29][15] , \w[29][14] , 
        \w[29][13] , \w[29][12] , \w[29][11] , \w[29][10] , \w[29][9] , 
        \w[29][8] , \w[29][7] , \w[29][6] , \w[29][5] , \w[29][4] , \w[29][3] , 
        \w[29][2] , \w[29][1] , SYNOPSYS_UNCONNECTED__27}) );
  ADD_N32_223 \FAINST[29].ADD_  ( .A({\_56_net_[31] , \_56_net_[30] , 
        \_56_net_[29] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[29][31] , 
        \w[29][30] , \w[29][29] , \w[29][28] , \w[29][27] , \w[29][26] , 
        \w[29][25] , \w[29][24] , \w[29][23] , \w[29][22] , \w[29][21] , 
        \w[29][20] , \w[29][19] , \w[29][18] , \w[29][17] , \w[29][16] , 
        \w[29][15] , \w[29][14] , \w[29][13] , \w[29][12] , \w[29][11] , 
        \w[29][10] , \w[29][9] , \w[29][8] , \w[29][7] , \w[29][6] , 
        \w[29][5] , \w[29][4] , \w[29][3] , \w[29][2] , \w[29][1] , 1'b0}), 
        .CI(1'b0), .S({\w[30][31] , \w[30][30] , \w[30][29] , \w[30][28] , 
        \w[30][27] , \w[30][26] , \w[30][25] , \w[30][24] , \w[30][23] , 
        \w[30][22] , \w[30][21] , \w[30][20] , \w[30][19] , \w[30][18] , 
        \w[30][17] , \w[30][16] , \w[30][15] , \w[30][14] , \w[30][13] , 
        \w[30][12] , \w[30][11] , \w[30][10] , \w[30][9] , \w[30][8] , 
        \w[30][7] , \w[30][6] , \w[30][5] , \w[30][4] , \w[30][3] , \w[30][2] , 
        \w[30][1] , SYNOPSYS_UNCONNECTED__28}) );
  ADD_N32_222 \FAINST[30].ADD_  ( .A({\_58_net_[31] , \_58_net_[30] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[30][31] , \w[30][30] , 
        \w[30][29] , \w[30][28] , \w[30][27] , \w[30][26] , \w[30][25] , 
        \w[30][24] , \w[30][23] , \w[30][22] , \w[30][21] , \w[30][20] , 
        \w[30][19] , \w[30][18] , \w[30][17] , \w[30][16] , \w[30][15] , 
        \w[30][14] , \w[30][13] , \w[30][12] , \w[30][11] , \w[30][10] , 
        \w[30][9] , \w[30][8] , \w[30][7] , \w[30][6] , \w[30][5] , \w[30][4] , 
        \w[30][3] , \w[30][2] , \w[30][1] , 1'b0}), .CI(1'b0), .S({\w[31][31] , 
        \w[31][30] , \w[31][29] , \w[31][28] , \w[31][27] , \w[31][26] , 
        \w[31][25] , \w[31][24] , \w[31][23] , \w[31][22] , \w[31][21] , 
        \w[31][20] , \w[31][19] , \w[31][18] , \w[31][17] , \w[31][16] , 
        \w[31][15] , \w[31][14] , \w[31][13] , \w[31][12] , \w[31][11] , 
        \w[31][10] , \w[31][9] , \w[31][8] , \w[31][7] , \w[31][6] , 
        \w[31][5] , \w[31][4] , \w[31][3] , \w[31][2] , \w[31][1] , 
        SYNOPSYS_UNCONNECTED__29}) );
  ADD_N32_221 \FAINST[31].ADD_  ( .A({\_60_net_[31] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({\w[31][31] , \w[31][30] , \w[31][29] , 
        \w[31][28] , \w[31][27] , \w[31][26] , \w[31][25] , \w[31][24] , 
        \w[31][23] , \w[31][22] , \w[31][21] , \w[31][20] , \w[31][19] , 
        \w[31][18] , \w[31][17] , \w[31][16] , \w[31][15] , \w[31][14] , 
        \w[31][13] , \w[31][12] , \w[31][11] , \w[31][10] , \w[31][9] , 
        \w[31][8] , \w[31][7] , \w[31][6] , \w[31][5] , \w[31][4] , \w[31][3] , 
        \w[31][2] , \w[31][1] , 1'b0}), .CI(1'b0), .S({O[31:1], 
        SYNOPSYS_UNCONNECTED__30}) );
  AND U2 ( .A(A[5]), .B(B[4]), .Z(\_8_net_[9] ) );
  AND U3 ( .A(A[5]), .B(B[3]), .Z(\_8_net_[8] ) );
  AND U4 ( .A(A[5]), .B(B[2]), .Z(\_8_net_[7] ) );
  AND U5 ( .A(A[5]), .B(B[1]), .Z(\_8_net_[6] ) );
  AND U6 ( .A(A[5]), .B(B[0]), .Z(\_8_net_[5] ) );
  AND U7 ( .A(A[5]), .B(B[26]), .Z(\_8_net_[31] ) );
  AND U8 ( .A(A[5]), .B(B[25]), .Z(\_8_net_[30] ) );
  AND U9 ( .A(A[5]), .B(B[24]), .Z(\_8_net_[29] ) );
  AND U10 ( .A(A[5]), .B(B[23]), .Z(\_8_net_[28] ) );
  AND U11 ( .A(A[5]), .B(B[22]), .Z(\_8_net_[27] ) );
  AND U12 ( .A(A[5]), .B(B[21]), .Z(\_8_net_[26] ) );
  AND U13 ( .A(A[5]), .B(B[20]), .Z(\_8_net_[25] ) );
  AND U14 ( .A(A[5]), .B(B[19]), .Z(\_8_net_[24] ) );
  AND U15 ( .A(A[5]), .B(B[18]), .Z(\_8_net_[23] ) );
  AND U16 ( .A(A[5]), .B(B[17]), .Z(\_8_net_[22] ) );
  AND U17 ( .A(A[5]), .B(B[16]), .Z(\_8_net_[21] ) );
  AND U18 ( .A(A[5]), .B(B[15]), .Z(\_8_net_[20] ) );
  AND U19 ( .A(A[5]), .B(B[14]), .Z(\_8_net_[19] ) );
  AND U20 ( .A(A[5]), .B(B[13]), .Z(\_8_net_[18] ) );
  AND U21 ( .A(A[5]), .B(B[12]), .Z(\_8_net_[17] ) );
  AND U22 ( .A(A[5]), .B(B[11]), .Z(\_8_net_[16] ) );
  AND U23 ( .A(A[5]), .B(B[10]), .Z(\_8_net_[15] ) );
  AND U24 ( .A(A[5]), .B(B[9]), .Z(\_8_net_[14] ) );
  AND U25 ( .A(A[5]), .B(B[8]), .Z(\_8_net_[13] ) );
  AND U26 ( .A(A[5]), .B(B[7]), .Z(\_8_net_[12] ) );
  AND U27 ( .A(A[5]), .B(B[6]), .Z(\_8_net_[11] ) );
  AND U28 ( .A(A[5]), .B(B[5]), .Z(\_8_net_[10] ) );
  AND U29 ( .A(B[5]), .B(A[4]), .Z(\_6_net_[9] ) );
  AND U30 ( .A(B[4]), .B(A[4]), .Z(\_6_net_[8] ) );
  AND U31 ( .A(B[3]), .B(A[4]), .Z(\_6_net_[7] ) );
  AND U32 ( .A(B[2]), .B(A[4]), .Z(\_6_net_[6] ) );
  AND U33 ( .A(B[1]), .B(A[4]), .Z(\_6_net_[5] ) );
  AND U34 ( .A(B[0]), .B(A[4]), .Z(\_6_net_[4] ) );
  AND U35 ( .A(A[4]), .B(B[27]), .Z(\_6_net_[31] ) );
  AND U36 ( .A(B[26]), .B(A[4]), .Z(\_6_net_[30] ) );
  AND U37 ( .A(B[25]), .B(A[4]), .Z(\_6_net_[29] ) );
  AND U38 ( .A(B[24]), .B(A[4]), .Z(\_6_net_[28] ) );
  AND U39 ( .A(B[23]), .B(A[4]), .Z(\_6_net_[27] ) );
  AND U40 ( .A(B[22]), .B(A[4]), .Z(\_6_net_[26] ) );
  AND U41 ( .A(B[21]), .B(A[4]), .Z(\_6_net_[25] ) );
  AND U42 ( .A(B[20]), .B(A[4]), .Z(\_6_net_[24] ) );
  AND U43 ( .A(B[19]), .B(A[4]), .Z(\_6_net_[23] ) );
  AND U44 ( .A(B[18]), .B(A[4]), .Z(\_6_net_[22] ) );
  AND U45 ( .A(B[17]), .B(A[4]), .Z(\_6_net_[21] ) );
  AND U46 ( .A(B[16]), .B(A[4]), .Z(\_6_net_[20] ) );
  AND U47 ( .A(B[15]), .B(A[4]), .Z(\_6_net_[19] ) );
  AND U48 ( .A(B[14]), .B(A[4]), .Z(\_6_net_[18] ) );
  AND U49 ( .A(B[13]), .B(A[4]), .Z(\_6_net_[17] ) );
  AND U50 ( .A(B[12]), .B(A[4]), .Z(\_6_net_[16] ) );
  AND U51 ( .A(B[11]), .B(A[4]), .Z(\_6_net_[15] ) );
  AND U52 ( .A(B[10]), .B(A[4]), .Z(\_6_net_[14] ) );
  AND U53 ( .A(B[9]), .B(A[4]), .Z(\_6_net_[13] ) );
  AND U54 ( .A(B[8]), .B(A[4]), .Z(\_6_net_[12] ) );
  AND U55 ( .A(B[7]), .B(A[4]), .Z(\_6_net_[11] ) );
  AND U56 ( .A(B[6]), .B(A[4]), .Z(\_6_net_[10] ) );
  AND U57 ( .A(A[31]), .B(B[0]), .Z(\_60_net_[31] ) );
  AND U58 ( .A(B[1]), .B(A[30]), .Z(\_58_net_[31] ) );
  AND U59 ( .A(A[30]), .B(B[0]), .Z(\_58_net_[30] ) );
  AND U60 ( .A(B[2]), .B(A[29]), .Z(\_56_net_[31] ) );
  AND U61 ( .A(B[1]), .B(A[29]), .Z(\_56_net_[30] ) );
  AND U62 ( .A(A[29]), .B(B[0]), .Z(\_56_net_[29] ) );
  AND U63 ( .A(B[3]), .B(A[28]), .Z(\_54_net_[31] ) );
  AND U64 ( .A(B[2]), .B(A[28]), .Z(\_54_net_[30] ) );
  AND U65 ( .A(B[1]), .B(A[28]), .Z(\_54_net_[29] ) );
  AND U66 ( .A(A[28]), .B(B[0]), .Z(\_54_net_[28] ) );
  AND U67 ( .A(B[4]), .B(A[27]), .Z(\_52_net_[31] ) );
  AND U68 ( .A(B[3]), .B(A[27]), .Z(\_52_net_[30] ) );
  AND U69 ( .A(B[2]), .B(A[27]), .Z(\_52_net_[29] ) );
  AND U70 ( .A(B[1]), .B(A[27]), .Z(\_52_net_[28] ) );
  AND U71 ( .A(A[27]), .B(B[0]), .Z(\_52_net_[27] ) );
  AND U72 ( .A(B[5]), .B(A[26]), .Z(\_50_net_[31] ) );
  AND U73 ( .A(B[4]), .B(A[26]), .Z(\_50_net_[30] ) );
  AND U74 ( .A(B[3]), .B(A[26]), .Z(\_50_net_[29] ) );
  AND U75 ( .A(B[2]), .B(A[26]), .Z(\_50_net_[28] ) );
  AND U76 ( .A(B[1]), .B(A[26]), .Z(\_50_net_[27] ) );
  AND U77 ( .A(A[26]), .B(B[0]), .Z(\_50_net_[26] ) );
  AND U78 ( .A(B[6]), .B(A[3]), .Z(\_4_net_[9] ) );
  AND U79 ( .A(B[5]), .B(A[3]), .Z(\_4_net_[8] ) );
  AND U80 ( .A(B[4]), .B(A[3]), .Z(\_4_net_[7] ) );
  AND U81 ( .A(B[3]), .B(A[3]), .Z(\_4_net_[6] ) );
  AND U82 ( .A(B[2]), .B(A[3]), .Z(\_4_net_[5] ) );
  AND U83 ( .A(B[1]), .B(A[3]), .Z(\_4_net_[4] ) );
  AND U84 ( .A(B[0]), .B(A[3]), .Z(\_4_net_[3] ) );
  AND U85 ( .A(A[3]), .B(B[28]), .Z(\_4_net_[31] ) );
  AND U86 ( .A(B[27]), .B(A[3]), .Z(\_4_net_[30] ) );
  AND U87 ( .A(B[26]), .B(A[3]), .Z(\_4_net_[29] ) );
  AND U88 ( .A(B[25]), .B(A[3]), .Z(\_4_net_[28] ) );
  AND U89 ( .A(B[24]), .B(A[3]), .Z(\_4_net_[27] ) );
  AND U90 ( .A(B[23]), .B(A[3]), .Z(\_4_net_[26] ) );
  AND U91 ( .A(B[22]), .B(A[3]), .Z(\_4_net_[25] ) );
  AND U92 ( .A(B[21]), .B(A[3]), .Z(\_4_net_[24] ) );
  AND U93 ( .A(B[20]), .B(A[3]), .Z(\_4_net_[23] ) );
  AND U94 ( .A(B[19]), .B(A[3]), .Z(\_4_net_[22] ) );
  AND U95 ( .A(B[18]), .B(A[3]), .Z(\_4_net_[21] ) );
  AND U96 ( .A(B[17]), .B(A[3]), .Z(\_4_net_[20] ) );
  AND U97 ( .A(B[16]), .B(A[3]), .Z(\_4_net_[19] ) );
  AND U98 ( .A(B[15]), .B(A[3]), .Z(\_4_net_[18] ) );
  AND U99 ( .A(B[14]), .B(A[3]), .Z(\_4_net_[17] ) );
  AND U100 ( .A(B[13]), .B(A[3]), .Z(\_4_net_[16] ) );
  AND U101 ( .A(B[12]), .B(A[3]), .Z(\_4_net_[15] ) );
  AND U102 ( .A(B[11]), .B(A[3]), .Z(\_4_net_[14] ) );
  AND U103 ( .A(B[10]), .B(A[3]), .Z(\_4_net_[13] ) );
  AND U104 ( .A(B[9]), .B(A[3]), .Z(\_4_net_[12] ) );
  AND U105 ( .A(B[8]), .B(A[3]), .Z(\_4_net_[11] ) );
  AND U106 ( .A(B[7]), .B(A[3]), .Z(\_4_net_[10] ) );
  AND U107 ( .A(B[6]), .B(A[25]), .Z(\_48_net_[31] ) );
  AND U108 ( .A(B[5]), .B(A[25]), .Z(\_48_net_[30] ) );
  AND U109 ( .A(B[4]), .B(A[25]), .Z(\_48_net_[29] ) );
  AND U110 ( .A(B[3]), .B(A[25]), .Z(\_48_net_[28] ) );
  AND U111 ( .A(B[2]), .B(A[25]), .Z(\_48_net_[27] ) );
  AND U112 ( .A(B[1]), .B(A[25]), .Z(\_48_net_[26] ) );
  AND U113 ( .A(A[25]), .B(B[0]), .Z(\_48_net_[25] ) );
  AND U114 ( .A(B[7]), .B(A[24]), .Z(\_46_net_[31] ) );
  AND U115 ( .A(B[6]), .B(A[24]), .Z(\_46_net_[30] ) );
  AND U116 ( .A(B[5]), .B(A[24]), .Z(\_46_net_[29] ) );
  AND U117 ( .A(B[4]), .B(A[24]), .Z(\_46_net_[28] ) );
  AND U118 ( .A(B[3]), .B(A[24]), .Z(\_46_net_[27] ) );
  AND U119 ( .A(B[2]), .B(A[24]), .Z(\_46_net_[26] ) );
  AND U120 ( .A(B[1]), .B(A[24]), .Z(\_46_net_[25] ) );
  AND U121 ( .A(A[24]), .B(B[0]), .Z(\_46_net_[24] ) );
  AND U122 ( .A(B[8]), .B(A[23]), .Z(\_44_net_[31] ) );
  AND U123 ( .A(B[7]), .B(A[23]), .Z(\_44_net_[30] ) );
  AND U124 ( .A(B[6]), .B(A[23]), .Z(\_44_net_[29] ) );
  AND U125 ( .A(B[5]), .B(A[23]), .Z(\_44_net_[28] ) );
  AND U126 ( .A(B[4]), .B(A[23]), .Z(\_44_net_[27] ) );
  AND U127 ( .A(B[3]), .B(A[23]), .Z(\_44_net_[26] ) );
  AND U128 ( .A(B[2]), .B(A[23]), .Z(\_44_net_[25] ) );
  AND U129 ( .A(B[1]), .B(A[23]), .Z(\_44_net_[24] ) );
  AND U130 ( .A(A[23]), .B(B[0]), .Z(\_44_net_[23] ) );
  AND U131 ( .A(B[9]), .B(A[22]), .Z(\_42_net_[31] ) );
  AND U132 ( .A(B[8]), .B(A[22]), .Z(\_42_net_[30] ) );
  AND U133 ( .A(B[7]), .B(A[22]), .Z(\_42_net_[29] ) );
  AND U134 ( .A(B[6]), .B(A[22]), .Z(\_42_net_[28] ) );
  AND U135 ( .A(B[5]), .B(A[22]), .Z(\_42_net_[27] ) );
  AND U136 ( .A(B[4]), .B(A[22]), .Z(\_42_net_[26] ) );
  AND U137 ( .A(B[3]), .B(A[22]), .Z(\_42_net_[25] ) );
  AND U138 ( .A(B[2]), .B(A[22]), .Z(\_42_net_[24] ) );
  AND U139 ( .A(B[1]), .B(A[22]), .Z(\_42_net_[23] ) );
  AND U140 ( .A(A[22]), .B(B[0]), .Z(\_42_net_[22] ) );
  AND U141 ( .A(B[10]), .B(A[21]), .Z(\_40_net_[31] ) );
  AND U142 ( .A(B[9]), .B(A[21]), .Z(\_40_net_[30] ) );
  AND U143 ( .A(B[8]), .B(A[21]), .Z(\_40_net_[29] ) );
  AND U144 ( .A(B[7]), .B(A[21]), .Z(\_40_net_[28] ) );
  AND U145 ( .A(B[6]), .B(A[21]), .Z(\_40_net_[27] ) );
  AND U146 ( .A(B[5]), .B(A[21]), .Z(\_40_net_[26] ) );
  AND U147 ( .A(B[4]), .B(A[21]), .Z(\_40_net_[25] ) );
  AND U148 ( .A(B[3]), .B(A[21]), .Z(\_40_net_[24] ) );
  AND U149 ( .A(B[2]), .B(A[21]), .Z(\_40_net_[23] ) );
  AND U150 ( .A(B[1]), .B(A[21]), .Z(\_40_net_[22] ) );
  AND U151 ( .A(A[21]), .B(B[0]), .Z(\_40_net_[21] ) );
  AND U152 ( .A(B[11]), .B(A[20]), .Z(\_38_net_[31] ) );
  AND U153 ( .A(B[10]), .B(A[20]), .Z(\_38_net_[30] ) );
  AND U154 ( .A(B[9]), .B(A[20]), .Z(\_38_net_[29] ) );
  AND U155 ( .A(B[8]), .B(A[20]), .Z(\_38_net_[28] ) );
  AND U156 ( .A(B[7]), .B(A[20]), .Z(\_38_net_[27] ) );
  AND U157 ( .A(B[6]), .B(A[20]), .Z(\_38_net_[26] ) );
  AND U158 ( .A(B[5]), .B(A[20]), .Z(\_38_net_[25] ) );
  AND U159 ( .A(B[4]), .B(A[20]), .Z(\_38_net_[24] ) );
  AND U160 ( .A(B[3]), .B(A[20]), .Z(\_38_net_[23] ) );
  AND U161 ( .A(B[2]), .B(A[20]), .Z(\_38_net_[22] ) );
  AND U162 ( .A(B[1]), .B(A[20]), .Z(\_38_net_[21] ) );
  AND U163 ( .A(A[20]), .B(B[0]), .Z(\_38_net_[20] ) );
  AND U164 ( .A(B[12]), .B(A[19]), .Z(\_36_net_[31] ) );
  AND U165 ( .A(B[11]), .B(A[19]), .Z(\_36_net_[30] ) );
  AND U166 ( .A(B[10]), .B(A[19]), .Z(\_36_net_[29] ) );
  AND U167 ( .A(B[9]), .B(A[19]), .Z(\_36_net_[28] ) );
  AND U168 ( .A(B[8]), .B(A[19]), .Z(\_36_net_[27] ) );
  AND U169 ( .A(B[7]), .B(A[19]), .Z(\_36_net_[26] ) );
  AND U170 ( .A(B[6]), .B(A[19]), .Z(\_36_net_[25] ) );
  AND U171 ( .A(B[5]), .B(A[19]), .Z(\_36_net_[24] ) );
  AND U172 ( .A(B[4]), .B(A[19]), .Z(\_36_net_[23] ) );
  AND U173 ( .A(B[3]), .B(A[19]), .Z(\_36_net_[22] ) );
  AND U174 ( .A(B[2]), .B(A[19]), .Z(\_36_net_[21] ) );
  AND U175 ( .A(B[1]), .B(A[19]), .Z(\_36_net_[20] ) );
  AND U176 ( .A(A[19]), .B(B[0]), .Z(\_36_net_[19] ) );
  AND U177 ( .A(B[13]), .B(A[18]), .Z(\_34_net_[31] ) );
  AND U178 ( .A(B[12]), .B(A[18]), .Z(\_34_net_[30] ) );
  AND U179 ( .A(B[11]), .B(A[18]), .Z(\_34_net_[29] ) );
  AND U180 ( .A(B[10]), .B(A[18]), .Z(\_34_net_[28] ) );
  AND U181 ( .A(B[9]), .B(A[18]), .Z(\_34_net_[27] ) );
  AND U182 ( .A(B[8]), .B(A[18]), .Z(\_34_net_[26] ) );
  AND U183 ( .A(B[7]), .B(A[18]), .Z(\_34_net_[25] ) );
  AND U184 ( .A(B[6]), .B(A[18]), .Z(\_34_net_[24] ) );
  AND U185 ( .A(B[5]), .B(A[18]), .Z(\_34_net_[23] ) );
  AND U186 ( .A(B[4]), .B(A[18]), .Z(\_34_net_[22] ) );
  AND U187 ( .A(B[3]), .B(A[18]), .Z(\_34_net_[21] ) );
  AND U188 ( .A(B[2]), .B(A[18]), .Z(\_34_net_[20] ) );
  AND U189 ( .A(B[1]), .B(A[18]), .Z(\_34_net_[19] ) );
  AND U190 ( .A(A[18]), .B(B[0]), .Z(\_34_net_[18] ) );
  AND U191 ( .A(B[14]), .B(A[17]), .Z(\_32_net_[31] ) );
  AND U192 ( .A(B[13]), .B(A[17]), .Z(\_32_net_[30] ) );
  AND U193 ( .A(B[12]), .B(A[17]), .Z(\_32_net_[29] ) );
  AND U194 ( .A(B[11]), .B(A[17]), .Z(\_32_net_[28] ) );
  AND U195 ( .A(B[10]), .B(A[17]), .Z(\_32_net_[27] ) );
  AND U196 ( .A(B[9]), .B(A[17]), .Z(\_32_net_[26] ) );
  AND U197 ( .A(B[8]), .B(A[17]), .Z(\_32_net_[25] ) );
  AND U198 ( .A(B[7]), .B(A[17]), .Z(\_32_net_[24] ) );
  AND U199 ( .A(B[6]), .B(A[17]), .Z(\_32_net_[23] ) );
  AND U200 ( .A(B[5]), .B(A[17]), .Z(\_32_net_[22] ) );
  AND U201 ( .A(B[4]), .B(A[17]), .Z(\_32_net_[21] ) );
  AND U202 ( .A(B[3]), .B(A[17]), .Z(\_32_net_[20] ) );
  AND U203 ( .A(B[2]), .B(A[17]), .Z(\_32_net_[19] ) );
  AND U204 ( .A(B[1]), .B(A[17]), .Z(\_32_net_[18] ) );
  AND U205 ( .A(A[17]), .B(B[0]), .Z(\_32_net_[17] ) );
  AND U206 ( .A(B[15]), .B(A[16]), .Z(\_30_net_[31] ) );
  AND U207 ( .A(B[14]), .B(A[16]), .Z(\_30_net_[30] ) );
  AND U208 ( .A(B[13]), .B(A[16]), .Z(\_30_net_[29] ) );
  AND U209 ( .A(B[12]), .B(A[16]), .Z(\_30_net_[28] ) );
  AND U210 ( .A(B[11]), .B(A[16]), .Z(\_30_net_[27] ) );
  AND U211 ( .A(B[10]), .B(A[16]), .Z(\_30_net_[26] ) );
  AND U212 ( .A(B[9]), .B(A[16]), .Z(\_30_net_[25] ) );
  AND U213 ( .A(B[8]), .B(A[16]), .Z(\_30_net_[24] ) );
  AND U214 ( .A(B[7]), .B(A[16]), .Z(\_30_net_[23] ) );
  AND U215 ( .A(B[6]), .B(A[16]), .Z(\_30_net_[22] ) );
  AND U216 ( .A(B[5]), .B(A[16]), .Z(\_30_net_[21] ) );
  AND U217 ( .A(B[4]), .B(A[16]), .Z(\_30_net_[20] ) );
  AND U218 ( .A(B[3]), .B(A[16]), .Z(\_30_net_[19] ) );
  AND U219 ( .A(B[2]), .B(A[16]), .Z(\_30_net_[18] ) );
  AND U220 ( .A(B[1]), .B(A[16]), .Z(\_30_net_[17] ) );
  AND U221 ( .A(A[16]), .B(B[0]), .Z(\_30_net_[16] ) );
  AND U222 ( .A(B[7]), .B(A[2]), .Z(\_2_net_[9] ) );
  AND U223 ( .A(B[6]), .B(A[2]), .Z(\_2_net_[8] ) );
  AND U224 ( .A(B[5]), .B(A[2]), .Z(\_2_net_[7] ) );
  AND U225 ( .A(B[4]), .B(A[2]), .Z(\_2_net_[6] ) );
  AND U226 ( .A(B[3]), .B(A[2]), .Z(\_2_net_[5] ) );
  AND U227 ( .A(B[2]), .B(A[2]), .Z(\_2_net_[4] ) );
  AND U228 ( .A(B[1]), .B(A[2]), .Z(\_2_net_[3] ) );
  AND U229 ( .A(A[2]), .B(B[29]), .Z(\_2_net_[31] ) );
  AND U230 ( .A(B[28]), .B(A[2]), .Z(\_2_net_[30] ) );
  AND U231 ( .A(B[0]), .B(A[2]), .Z(\_2_net_[2] ) );
  AND U232 ( .A(B[27]), .B(A[2]), .Z(\_2_net_[29] ) );
  AND U233 ( .A(B[26]), .B(A[2]), .Z(\_2_net_[28] ) );
  AND U234 ( .A(B[25]), .B(A[2]), .Z(\_2_net_[27] ) );
  AND U235 ( .A(B[24]), .B(A[2]), .Z(\_2_net_[26] ) );
  AND U236 ( .A(B[23]), .B(A[2]), .Z(\_2_net_[25] ) );
  AND U237 ( .A(B[22]), .B(A[2]), .Z(\_2_net_[24] ) );
  AND U238 ( .A(B[21]), .B(A[2]), .Z(\_2_net_[23] ) );
  AND U239 ( .A(B[20]), .B(A[2]), .Z(\_2_net_[22] ) );
  AND U240 ( .A(B[19]), .B(A[2]), .Z(\_2_net_[21] ) );
  AND U241 ( .A(B[18]), .B(A[2]), .Z(\_2_net_[20] ) );
  AND U242 ( .A(B[17]), .B(A[2]), .Z(\_2_net_[19] ) );
  AND U243 ( .A(B[16]), .B(A[2]), .Z(\_2_net_[18] ) );
  AND U244 ( .A(B[15]), .B(A[2]), .Z(\_2_net_[17] ) );
  AND U245 ( .A(B[14]), .B(A[2]), .Z(\_2_net_[16] ) );
  AND U246 ( .A(B[13]), .B(A[2]), .Z(\_2_net_[15] ) );
  AND U247 ( .A(B[12]), .B(A[2]), .Z(\_2_net_[14] ) );
  AND U248 ( .A(B[11]), .B(A[2]), .Z(\_2_net_[13] ) );
  AND U249 ( .A(B[10]), .B(A[2]), .Z(\_2_net_[12] ) );
  AND U250 ( .A(B[9]), .B(A[2]), .Z(\_2_net_[11] ) );
  AND U251 ( .A(B[8]), .B(A[2]), .Z(\_2_net_[10] ) );
  AND U252 ( .A(B[16]), .B(A[15]), .Z(\_28_net_[31] ) );
  AND U253 ( .A(B[15]), .B(A[15]), .Z(\_28_net_[30] ) );
  AND U254 ( .A(B[14]), .B(A[15]), .Z(\_28_net_[29] ) );
  AND U255 ( .A(B[13]), .B(A[15]), .Z(\_28_net_[28] ) );
  AND U256 ( .A(B[12]), .B(A[15]), .Z(\_28_net_[27] ) );
  AND U257 ( .A(B[11]), .B(A[15]), .Z(\_28_net_[26] ) );
  AND U258 ( .A(B[10]), .B(A[15]), .Z(\_28_net_[25] ) );
  AND U259 ( .A(B[9]), .B(A[15]), .Z(\_28_net_[24] ) );
  AND U260 ( .A(B[8]), .B(A[15]), .Z(\_28_net_[23] ) );
  AND U261 ( .A(B[7]), .B(A[15]), .Z(\_28_net_[22] ) );
  AND U262 ( .A(B[6]), .B(A[15]), .Z(\_28_net_[21] ) );
  AND U263 ( .A(B[5]), .B(A[15]), .Z(\_28_net_[20] ) );
  AND U264 ( .A(B[4]), .B(A[15]), .Z(\_28_net_[19] ) );
  AND U265 ( .A(B[3]), .B(A[15]), .Z(\_28_net_[18] ) );
  AND U266 ( .A(B[2]), .B(A[15]), .Z(\_28_net_[17] ) );
  AND U267 ( .A(B[1]), .B(A[15]), .Z(\_28_net_[16] ) );
  AND U268 ( .A(A[15]), .B(B[0]), .Z(\_28_net_[15] ) );
  AND U269 ( .A(B[17]), .B(A[14]), .Z(\_26_net_[31] ) );
  AND U270 ( .A(B[16]), .B(A[14]), .Z(\_26_net_[30] ) );
  AND U271 ( .A(B[15]), .B(A[14]), .Z(\_26_net_[29] ) );
  AND U272 ( .A(B[14]), .B(A[14]), .Z(\_26_net_[28] ) );
  AND U273 ( .A(B[13]), .B(A[14]), .Z(\_26_net_[27] ) );
  AND U274 ( .A(B[12]), .B(A[14]), .Z(\_26_net_[26] ) );
  AND U275 ( .A(B[11]), .B(A[14]), .Z(\_26_net_[25] ) );
  AND U276 ( .A(B[10]), .B(A[14]), .Z(\_26_net_[24] ) );
  AND U277 ( .A(B[9]), .B(A[14]), .Z(\_26_net_[23] ) );
  AND U278 ( .A(B[8]), .B(A[14]), .Z(\_26_net_[22] ) );
  AND U279 ( .A(B[7]), .B(A[14]), .Z(\_26_net_[21] ) );
  AND U280 ( .A(B[6]), .B(A[14]), .Z(\_26_net_[20] ) );
  AND U281 ( .A(B[5]), .B(A[14]), .Z(\_26_net_[19] ) );
  AND U282 ( .A(B[4]), .B(A[14]), .Z(\_26_net_[18] ) );
  AND U283 ( .A(B[3]), .B(A[14]), .Z(\_26_net_[17] ) );
  AND U284 ( .A(B[2]), .B(A[14]), .Z(\_26_net_[16] ) );
  AND U285 ( .A(B[1]), .B(A[14]), .Z(\_26_net_[15] ) );
  AND U286 ( .A(A[14]), .B(B[0]), .Z(\_26_net_[14] ) );
  AND U287 ( .A(B[18]), .B(A[13]), .Z(\_24_net_[31] ) );
  AND U288 ( .A(B[17]), .B(A[13]), .Z(\_24_net_[30] ) );
  AND U289 ( .A(B[16]), .B(A[13]), .Z(\_24_net_[29] ) );
  AND U290 ( .A(B[15]), .B(A[13]), .Z(\_24_net_[28] ) );
  AND U291 ( .A(B[14]), .B(A[13]), .Z(\_24_net_[27] ) );
  AND U292 ( .A(B[13]), .B(A[13]), .Z(\_24_net_[26] ) );
  AND U293 ( .A(B[12]), .B(A[13]), .Z(\_24_net_[25] ) );
  AND U294 ( .A(B[11]), .B(A[13]), .Z(\_24_net_[24] ) );
  AND U295 ( .A(B[10]), .B(A[13]), .Z(\_24_net_[23] ) );
  AND U296 ( .A(B[9]), .B(A[13]), .Z(\_24_net_[22] ) );
  AND U297 ( .A(B[8]), .B(A[13]), .Z(\_24_net_[21] ) );
  AND U298 ( .A(B[7]), .B(A[13]), .Z(\_24_net_[20] ) );
  AND U299 ( .A(B[6]), .B(A[13]), .Z(\_24_net_[19] ) );
  AND U300 ( .A(B[5]), .B(A[13]), .Z(\_24_net_[18] ) );
  AND U301 ( .A(B[4]), .B(A[13]), .Z(\_24_net_[17] ) );
  AND U302 ( .A(B[3]), .B(A[13]), .Z(\_24_net_[16] ) );
  AND U303 ( .A(B[2]), .B(A[13]), .Z(\_24_net_[15] ) );
  AND U304 ( .A(B[1]), .B(A[13]), .Z(\_24_net_[14] ) );
  AND U305 ( .A(A[13]), .B(B[0]), .Z(\_24_net_[13] ) );
  AND U306 ( .A(B[19]), .B(A[12]), .Z(\_22_net_[31] ) );
  AND U307 ( .A(B[18]), .B(A[12]), .Z(\_22_net_[30] ) );
  AND U308 ( .A(B[17]), .B(A[12]), .Z(\_22_net_[29] ) );
  AND U309 ( .A(B[16]), .B(A[12]), .Z(\_22_net_[28] ) );
  AND U310 ( .A(B[15]), .B(A[12]), .Z(\_22_net_[27] ) );
  AND U311 ( .A(B[14]), .B(A[12]), .Z(\_22_net_[26] ) );
  AND U312 ( .A(B[13]), .B(A[12]), .Z(\_22_net_[25] ) );
  AND U313 ( .A(B[12]), .B(A[12]), .Z(\_22_net_[24] ) );
  AND U314 ( .A(B[11]), .B(A[12]), .Z(\_22_net_[23] ) );
  AND U315 ( .A(B[10]), .B(A[12]), .Z(\_22_net_[22] ) );
  AND U316 ( .A(B[9]), .B(A[12]), .Z(\_22_net_[21] ) );
  AND U317 ( .A(B[8]), .B(A[12]), .Z(\_22_net_[20] ) );
  AND U318 ( .A(B[7]), .B(A[12]), .Z(\_22_net_[19] ) );
  AND U319 ( .A(B[6]), .B(A[12]), .Z(\_22_net_[18] ) );
  AND U320 ( .A(B[5]), .B(A[12]), .Z(\_22_net_[17] ) );
  AND U321 ( .A(B[4]), .B(A[12]), .Z(\_22_net_[16] ) );
  AND U322 ( .A(B[3]), .B(A[12]), .Z(\_22_net_[15] ) );
  AND U323 ( .A(B[2]), .B(A[12]), .Z(\_22_net_[14] ) );
  AND U324 ( .A(B[1]), .B(A[12]), .Z(\_22_net_[13] ) );
  AND U325 ( .A(A[12]), .B(B[0]), .Z(\_22_net_[12] ) );
  AND U326 ( .A(B[20]), .B(A[11]), .Z(\_20_net_[31] ) );
  AND U327 ( .A(B[19]), .B(A[11]), .Z(\_20_net_[30] ) );
  AND U328 ( .A(B[18]), .B(A[11]), .Z(\_20_net_[29] ) );
  AND U329 ( .A(B[17]), .B(A[11]), .Z(\_20_net_[28] ) );
  AND U330 ( .A(B[16]), .B(A[11]), .Z(\_20_net_[27] ) );
  AND U331 ( .A(B[15]), .B(A[11]), .Z(\_20_net_[26] ) );
  AND U332 ( .A(B[14]), .B(A[11]), .Z(\_20_net_[25] ) );
  AND U333 ( .A(B[13]), .B(A[11]), .Z(\_20_net_[24] ) );
  AND U334 ( .A(B[12]), .B(A[11]), .Z(\_20_net_[23] ) );
  AND U335 ( .A(B[11]), .B(A[11]), .Z(\_20_net_[22] ) );
  AND U336 ( .A(B[10]), .B(A[11]), .Z(\_20_net_[21] ) );
  AND U337 ( .A(B[9]), .B(A[11]), .Z(\_20_net_[20] ) );
  AND U338 ( .A(B[8]), .B(A[11]), .Z(\_20_net_[19] ) );
  AND U339 ( .A(B[7]), .B(A[11]), .Z(\_20_net_[18] ) );
  AND U340 ( .A(B[6]), .B(A[11]), .Z(\_20_net_[17] ) );
  AND U341 ( .A(B[5]), .B(A[11]), .Z(\_20_net_[16] ) );
  AND U342 ( .A(B[4]), .B(A[11]), .Z(\_20_net_[15] ) );
  AND U343 ( .A(B[3]), .B(A[11]), .Z(\_20_net_[14] ) );
  AND U344 ( .A(B[2]), .B(A[11]), .Z(\_20_net_[13] ) );
  AND U345 ( .A(B[1]), .B(A[11]), .Z(\_20_net_[12] ) );
  AND U346 ( .A(A[11]), .B(B[0]), .Z(\_20_net_[11] ) );
  AND U347 ( .A(B[21]), .B(A[10]), .Z(\_18_net_[31] ) );
  AND U348 ( .A(B[20]), .B(A[10]), .Z(\_18_net_[30] ) );
  AND U349 ( .A(B[19]), .B(A[10]), .Z(\_18_net_[29] ) );
  AND U350 ( .A(B[18]), .B(A[10]), .Z(\_18_net_[28] ) );
  AND U351 ( .A(B[17]), .B(A[10]), .Z(\_18_net_[27] ) );
  AND U352 ( .A(B[16]), .B(A[10]), .Z(\_18_net_[26] ) );
  AND U353 ( .A(B[15]), .B(A[10]), .Z(\_18_net_[25] ) );
  AND U354 ( .A(B[14]), .B(A[10]), .Z(\_18_net_[24] ) );
  AND U355 ( .A(B[13]), .B(A[10]), .Z(\_18_net_[23] ) );
  AND U356 ( .A(B[12]), .B(A[10]), .Z(\_18_net_[22] ) );
  AND U357 ( .A(B[11]), .B(A[10]), .Z(\_18_net_[21] ) );
  AND U358 ( .A(B[10]), .B(A[10]), .Z(\_18_net_[20] ) );
  AND U359 ( .A(B[9]), .B(A[10]), .Z(\_18_net_[19] ) );
  AND U360 ( .A(B[8]), .B(A[10]), .Z(\_18_net_[18] ) );
  AND U361 ( .A(B[7]), .B(A[10]), .Z(\_18_net_[17] ) );
  AND U362 ( .A(B[6]), .B(A[10]), .Z(\_18_net_[16] ) );
  AND U363 ( .A(B[5]), .B(A[10]), .Z(\_18_net_[15] ) );
  AND U364 ( .A(B[4]), .B(A[10]), .Z(\_18_net_[14] ) );
  AND U365 ( .A(B[3]), .B(A[10]), .Z(\_18_net_[13] ) );
  AND U366 ( .A(B[2]), .B(A[10]), .Z(\_18_net_[12] ) );
  AND U367 ( .A(B[1]), .B(A[10]), .Z(\_18_net_[11] ) );
  AND U368 ( .A(A[10]), .B(B[0]), .Z(\_18_net_[10] ) );
  AND U369 ( .A(B[0]), .B(A[9]), .Z(\_16_net_[9] ) );
  AND U370 ( .A(B[22]), .B(A[9]), .Z(\_16_net_[31] ) );
  AND U371 ( .A(B[21]), .B(A[9]), .Z(\_16_net_[30] ) );
  AND U372 ( .A(B[20]), .B(A[9]), .Z(\_16_net_[29] ) );
  AND U373 ( .A(B[19]), .B(A[9]), .Z(\_16_net_[28] ) );
  AND U374 ( .A(B[18]), .B(A[9]), .Z(\_16_net_[27] ) );
  AND U375 ( .A(B[17]), .B(A[9]), .Z(\_16_net_[26] ) );
  AND U376 ( .A(B[16]), .B(A[9]), .Z(\_16_net_[25] ) );
  AND U377 ( .A(B[15]), .B(A[9]), .Z(\_16_net_[24] ) );
  AND U378 ( .A(B[14]), .B(A[9]), .Z(\_16_net_[23] ) );
  AND U379 ( .A(B[13]), .B(A[9]), .Z(\_16_net_[22] ) );
  AND U380 ( .A(B[12]), .B(A[9]), .Z(\_16_net_[21] ) );
  AND U381 ( .A(B[11]), .B(A[9]), .Z(\_16_net_[20] ) );
  AND U382 ( .A(B[10]), .B(A[9]), .Z(\_16_net_[19] ) );
  AND U383 ( .A(B[9]), .B(A[9]), .Z(\_16_net_[18] ) );
  AND U384 ( .A(B[8]), .B(A[9]), .Z(\_16_net_[17] ) );
  AND U385 ( .A(B[7]), .B(A[9]), .Z(\_16_net_[16] ) );
  AND U386 ( .A(B[6]), .B(A[9]), .Z(\_16_net_[15] ) );
  AND U387 ( .A(B[5]), .B(A[9]), .Z(\_16_net_[14] ) );
  AND U388 ( .A(B[4]), .B(A[9]), .Z(\_16_net_[13] ) );
  AND U389 ( .A(B[3]), .B(A[9]), .Z(\_16_net_[12] ) );
  AND U390 ( .A(B[2]), .B(A[9]), .Z(\_16_net_[11] ) );
  AND U391 ( .A(A[9]), .B(B[1]), .Z(\_16_net_[10] ) );
  AND U392 ( .A(B[1]), .B(A[8]), .Z(\_14_net_[9] ) );
  AND U393 ( .A(B[0]), .B(A[8]), .Z(\_14_net_[8] ) );
  AND U394 ( .A(B[23]), .B(A[8]), .Z(\_14_net_[31] ) );
  AND U395 ( .A(B[22]), .B(A[8]), .Z(\_14_net_[30] ) );
  AND U396 ( .A(B[21]), .B(A[8]), .Z(\_14_net_[29] ) );
  AND U397 ( .A(B[20]), .B(A[8]), .Z(\_14_net_[28] ) );
  AND U398 ( .A(B[19]), .B(A[8]), .Z(\_14_net_[27] ) );
  AND U399 ( .A(B[18]), .B(A[8]), .Z(\_14_net_[26] ) );
  AND U400 ( .A(B[17]), .B(A[8]), .Z(\_14_net_[25] ) );
  AND U401 ( .A(B[16]), .B(A[8]), .Z(\_14_net_[24] ) );
  AND U402 ( .A(B[15]), .B(A[8]), .Z(\_14_net_[23] ) );
  AND U403 ( .A(B[14]), .B(A[8]), .Z(\_14_net_[22] ) );
  AND U404 ( .A(B[13]), .B(A[8]), .Z(\_14_net_[21] ) );
  AND U405 ( .A(B[12]), .B(A[8]), .Z(\_14_net_[20] ) );
  AND U406 ( .A(B[11]), .B(A[8]), .Z(\_14_net_[19] ) );
  AND U407 ( .A(B[10]), .B(A[8]), .Z(\_14_net_[18] ) );
  AND U408 ( .A(B[9]), .B(A[8]), .Z(\_14_net_[17] ) );
  AND U409 ( .A(B[8]), .B(A[8]), .Z(\_14_net_[16] ) );
  AND U410 ( .A(B[7]), .B(A[8]), .Z(\_14_net_[15] ) );
  AND U411 ( .A(B[6]), .B(A[8]), .Z(\_14_net_[14] ) );
  AND U412 ( .A(B[5]), .B(A[8]), .Z(\_14_net_[13] ) );
  AND U413 ( .A(B[4]), .B(A[8]), .Z(\_14_net_[12] ) );
  AND U414 ( .A(B[3]), .B(A[8]), .Z(\_14_net_[11] ) );
  AND U415 ( .A(A[8]), .B(B[2]), .Z(\_14_net_[10] ) );
  AND U416 ( .A(B[2]), .B(A[7]), .Z(\_12_net_[9] ) );
  AND U417 ( .A(B[1]), .B(A[7]), .Z(\_12_net_[8] ) );
  AND U418 ( .A(B[0]), .B(A[7]), .Z(\_12_net_[7] ) );
  AND U419 ( .A(B[24]), .B(A[7]), .Z(\_12_net_[31] ) );
  AND U420 ( .A(B[23]), .B(A[7]), .Z(\_12_net_[30] ) );
  AND U421 ( .A(B[22]), .B(A[7]), .Z(\_12_net_[29] ) );
  AND U422 ( .A(B[21]), .B(A[7]), .Z(\_12_net_[28] ) );
  AND U423 ( .A(B[20]), .B(A[7]), .Z(\_12_net_[27] ) );
  AND U424 ( .A(B[19]), .B(A[7]), .Z(\_12_net_[26] ) );
  AND U425 ( .A(B[18]), .B(A[7]), .Z(\_12_net_[25] ) );
  AND U426 ( .A(B[17]), .B(A[7]), .Z(\_12_net_[24] ) );
  AND U427 ( .A(B[16]), .B(A[7]), .Z(\_12_net_[23] ) );
  AND U428 ( .A(B[15]), .B(A[7]), .Z(\_12_net_[22] ) );
  AND U429 ( .A(B[14]), .B(A[7]), .Z(\_12_net_[21] ) );
  AND U430 ( .A(B[13]), .B(A[7]), .Z(\_12_net_[20] ) );
  AND U431 ( .A(B[12]), .B(A[7]), .Z(\_12_net_[19] ) );
  AND U432 ( .A(B[11]), .B(A[7]), .Z(\_12_net_[18] ) );
  AND U433 ( .A(B[10]), .B(A[7]), .Z(\_12_net_[17] ) );
  AND U434 ( .A(B[9]), .B(A[7]), .Z(\_12_net_[16] ) );
  AND U435 ( .A(B[8]), .B(A[7]), .Z(\_12_net_[15] ) );
  AND U436 ( .A(B[7]), .B(A[7]), .Z(\_12_net_[14] ) );
  AND U437 ( .A(B[6]), .B(A[7]), .Z(\_12_net_[13] ) );
  AND U438 ( .A(B[5]), .B(A[7]), .Z(\_12_net_[12] ) );
  AND U439 ( .A(B[4]), .B(A[7]), .Z(\_12_net_[11] ) );
  AND U440 ( .A(A[7]), .B(B[3]), .Z(\_12_net_[10] ) );
  AND U441 ( .A(B[3]), .B(A[6]), .Z(\_10_net_[9] ) );
  AND U442 ( .A(B[2]), .B(A[6]), .Z(\_10_net_[8] ) );
  AND U443 ( .A(B[1]), .B(A[6]), .Z(\_10_net_[7] ) );
  AND U444 ( .A(B[0]), .B(A[6]), .Z(\_10_net_[6] ) );
  AND U445 ( .A(B[25]), .B(A[6]), .Z(\_10_net_[31] ) );
  AND U446 ( .A(B[24]), .B(A[6]), .Z(\_10_net_[30] ) );
  AND U447 ( .A(B[23]), .B(A[6]), .Z(\_10_net_[29] ) );
  AND U448 ( .A(B[22]), .B(A[6]), .Z(\_10_net_[28] ) );
  AND U449 ( .A(B[21]), .B(A[6]), .Z(\_10_net_[27] ) );
  AND U450 ( .A(B[20]), .B(A[6]), .Z(\_10_net_[26] ) );
  AND U451 ( .A(B[19]), .B(A[6]), .Z(\_10_net_[25] ) );
  AND U452 ( .A(B[18]), .B(A[6]), .Z(\_10_net_[24] ) );
  AND U453 ( .A(B[17]), .B(A[6]), .Z(\_10_net_[23] ) );
  AND U454 ( .A(B[16]), .B(A[6]), .Z(\_10_net_[22] ) );
  AND U455 ( .A(B[15]), .B(A[6]), .Z(\_10_net_[21] ) );
  AND U456 ( .A(B[14]), .B(A[6]), .Z(\_10_net_[20] ) );
  AND U457 ( .A(B[13]), .B(A[6]), .Z(\_10_net_[19] ) );
  AND U458 ( .A(B[12]), .B(A[6]), .Z(\_10_net_[18] ) );
  AND U459 ( .A(B[11]), .B(A[6]), .Z(\_10_net_[17] ) );
  AND U460 ( .A(B[10]), .B(A[6]), .Z(\_10_net_[16] ) );
  AND U461 ( .A(B[9]), .B(A[6]), .Z(\_10_net_[15] ) );
  AND U462 ( .A(B[8]), .B(A[6]), .Z(\_10_net_[14] ) );
  AND U463 ( .A(B[7]), .B(A[6]), .Z(\_10_net_[13] ) );
  AND U464 ( .A(B[6]), .B(A[6]), .Z(\_10_net_[12] ) );
  AND U465 ( .A(B[5]), .B(A[6]), .Z(\_10_net_[11] ) );
  AND U466 ( .A(A[6]), .B(B[4]), .Z(\_10_net_[10] ) );
  AND U467 ( .A(B[8]), .B(A[1]), .Z(\_0_net_[9] ) );
  AND U468 ( .A(B[7]), .B(A[1]), .Z(\_0_net_[8] ) );
  AND U469 ( .A(B[6]), .B(A[1]), .Z(\_0_net_[7] ) );
  AND U470 ( .A(B[5]), .B(A[1]), .Z(\_0_net_[6] ) );
  AND U471 ( .A(B[4]), .B(A[1]), .Z(\_0_net_[5] ) );
  AND U472 ( .A(B[3]), .B(A[1]), .Z(\_0_net_[4] ) );
  AND U473 ( .A(B[2]), .B(A[1]), .Z(\_0_net_[3] ) );
  AND U474 ( .A(B[30]), .B(A[1]), .Z(\_0_net_[31] ) );
  AND U475 ( .A(B[29]), .B(A[1]), .Z(\_0_net_[30] ) );
  AND U476 ( .A(B[1]), .B(A[1]), .Z(\_0_net_[2] ) );
  AND U477 ( .A(B[28]), .B(A[1]), .Z(\_0_net_[29] ) );
  AND U478 ( .A(B[27]), .B(A[1]), .Z(\_0_net_[28] ) );
  AND U479 ( .A(B[26]), .B(A[1]), .Z(\_0_net_[27] ) );
  AND U480 ( .A(B[25]), .B(A[1]), .Z(\_0_net_[26] ) );
  AND U481 ( .A(B[24]), .B(A[1]), .Z(\_0_net_[25] ) );
  AND U482 ( .A(B[23]), .B(A[1]), .Z(\_0_net_[24] ) );
  AND U483 ( .A(B[22]), .B(A[1]), .Z(\_0_net_[23] ) );
  AND U484 ( .A(B[21]), .B(A[1]), .Z(\_0_net_[22] ) );
  AND U485 ( .A(B[20]), .B(A[1]), .Z(\_0_net_[21] ) );
  AND U486 ( .A(B[19]), .B(A[1]), .Z(\_0_net_[20] ) );
  AND U487 ( .A(B[0]), .B(A[1]), .Z(\_0_net_[1] ) );
  AND U488 ( .A(B[18]), .B(A[1]), .Z(\_0_net_[19] ) );
  AND U489 ( .A(B[17]), .B(A[1]), .Z(\_0_net_[18] ) );
  AND U490 ( .A(B[16]), .B(A[1]), .Z(\_0_net_[17] ) );
  AND U491 ( .A(B[15]), .B(A[1]), .Z(\_0_net_[16] ) );
  AND U492 ( .A(B[14]), .B(A[1]), .Z(\_0_net_[15] ) );
  AND U493 ( .A(B[13]), .B(A[1]), .Z(\_0_net_[14] ) );
  AND U494 ( .A(B[12]), .B(A[1]), .Z(\_0_net_[13] ) );
  AND U495 ( .A(B[11]), .B(A[1]), .Z(\_0_net_[12] ) );
  AND U496 ( .A(B[10]), .B(A[1]), .Z(\_0_net_[11] ) );
  AND U497 ( .A(A[1]), .B(B[9]), .Z(\_0_net_[10] ) );
endmodule


module FA_8065 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_8066 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8067 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8068 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8069 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8070 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8071 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8072 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8073 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8074 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8075 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8076 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8077 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8078 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8079 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8080 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8081 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8082 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8083 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8084 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8085 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8086 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8087 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8088 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8089 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8090 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8091 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8092 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8093 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8094 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8095 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module ADD_N32_96 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_8095 \FAINST[1].FA_  ( .A(A[1]), .B(B[1]), .CI(1'b0), .S(S[1]), .CO(C[2])
         );
  FA_8094 \FAINST[2].FA_  ( .A(A[2]), .B(B[2]), .CI(C[2]), .S(S[2]), .CO(C[3])
         );
  FA_8093 \FAINST[3].FA_  ( .A(A[3]), .B(B[3]), .CI(C[3]), .S(S[3]), .CO(C[4])
         );
  FA_8092 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_8091 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_8090 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_8089 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_8088 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_8087 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_8086 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_8085 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_8084 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_8083 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_8082 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_8081 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_8080 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_8079 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_8078 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_8077 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_8076 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_8075 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_8074 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_8073 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_8072 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_8071 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_8070 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_8069 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_8068 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_8067 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_8066 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_8065 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_32 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_64 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_96 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_512 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_544 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_576 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_608 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_640 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_672 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_704 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_736 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_768 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_800 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_832 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_864 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_896 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_928 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_960 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_992 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_97 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;


  FA_992 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_960 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_928 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_896 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_864 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_832 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_800 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_768 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_736 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_704 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_672 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_640 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_608 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_576 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_544 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_512 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_480 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_448 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_416 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_384 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_352 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_320 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_288 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_256 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_224 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_192 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_160 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_128 \FAINST[28].FA_  ( .A(1'b0), .B(B[28]), .CI(1'b0), .S(S[28]) );
  FA_96 \FAINST[29].FA_  ( .A(1'b0), .B(B[29]), .CI(1'b0), .S(S[29]) );
  FA_64 \FAINST[30].FA_  ( .A(1'b0), .B(B[30]), .CI(1'b0), .S(S[30]) );
  FA_32 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(1'b0), .S(S[31]) );
endmodule


module FA_1056 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1088 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1120 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1152 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1184 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1216 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1248 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1280 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1312 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1344 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1376 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1408 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1440 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1472 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1504 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1536 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1568 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1600 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1632 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1664 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1696 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1728 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1760 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1792 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1824 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1856 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1888 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1920 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1952 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1984 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2016 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_98 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;
  wire   \C[31] ;

  FA_2016 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1984 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1952 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1920 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1888 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1856 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1824 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1792 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1760 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1728 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1696 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1664 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1632 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1600 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_1568 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_1536 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_1504 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_1472 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_1440 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_1408 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_1376 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_1344 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_1312 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_1280 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_1248 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_1216 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_1184 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_1152 \FAINST[28].FA_  ( .A(1'b0), .B(B[28]), .CI(1'b0), .S(S[28]) );
  FA_1120 \FAINST[29].FA_  ( .A(1'b0), .B(B[29]), .CI(1'b0), .S(S[29]) );
  FA_1088 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(1'b0), .S(S[30]), .CO(
        \C[31] ) );
  FA_1056 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(\C[31] ), .S(S[31]) );
endmodule


module FA_2080 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_2112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_2176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2528 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2560 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2592 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2624 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2656 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2688 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2720 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2752 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2784 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2816 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2848 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2880 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2912 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2944 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2976 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3008 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3040 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_99 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3040 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3008 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_2976 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_2944 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_2912 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_2880 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_2848 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_2816 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_2784 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_2752 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_2720 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_2688 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_2656 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_2624 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_2592 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_2560 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_2528 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_2496 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_2464 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_2432 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_2400 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_2368 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_2336 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_2304 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_2272 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_2240 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_2208 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_2176 \FAINST[28].FA_  ( .A(1'b0), .B(B[28]), .CI(1'b0), .S(S[28]) );
  FA_2144 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(1'b0), .S(S[29]), .CO(
        C[30]) );
  FA_2112 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_2080 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3073 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3074 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3075 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3076 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3077 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3078 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3079 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3080 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3081 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3082 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3083 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3084 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3085 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3086 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3087 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3088 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3089 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3090 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3091 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3092 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3093 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3094 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3095 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3096 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3097 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3098 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3099 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_100 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3103 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3102 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3101 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3100 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3099 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3098 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3097 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3096 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3095 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3094 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3093 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3092 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_3091 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_3090 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_3089 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_3088 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_3087 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_3086 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_3085 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_3084 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_3083 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_3082 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_3081 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_3080 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_3079 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_3078 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_3077 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_3076 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(1'b0), .S(S[28]), .CO(
        C[29]) );
  FA_3075 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3074 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3073 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3120 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_101 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3135 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3134 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3133 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3132 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3131 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3130 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3129 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3128 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3127 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3126 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3125 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3124 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_3123 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_3122 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_3121 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_3120 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_3119 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_3118 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_3117 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_3116 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_3115 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_3114 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_3113 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_3112 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_3111 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_3110 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_3109 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(1'b0), .S(S[27]), .CO(
        C[28]) );
  FA_3108 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3107 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3106 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3105 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3152 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_102 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3167 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3166 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3165 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3164 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3163 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3162 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3161 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3160 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3159 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3158 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3157 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3156 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_3155 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_3154 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_3153 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_3152 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_3151 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_3150 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_3149 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_3148 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_3147 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_3146 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_3145 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_3144 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_3143 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_3142 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(1'b0), .S(S[26]), .CO(
        C[27]) );
  FA_3141 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3140 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3139 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3138 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3137 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3184 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_103 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3199 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3198 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3197 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3196 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3195 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3194 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3193 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3192 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3191 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3190 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3189 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3188 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_3187 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_3186 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_3185 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_3184 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_3183 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_3182 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_3181 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_3180 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_3179 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_3178 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_3177 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_3176 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_3175 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(1'b0), .S(S[25]), .CO(
        C[26]) );
  FA_3174 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3173 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3172 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3171 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3170 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3169 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3216 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_104 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3231 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3230 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3229 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3228 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3227 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3226 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3225 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3224 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3223 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3222 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3221 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3220 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_3219 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_3218 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_3217 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_3216 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_3215 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_3214 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_3213 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_3212 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_3211 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_3210 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_3209 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_3208 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(1'b0), .S(S[24]), .CO(
        C[25]) );
  FA_3207 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3206 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3205 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3204 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3203 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3202 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3201 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3248 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_105 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3263 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3262 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3261 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3260 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3259 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3258 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3257 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3256 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3255 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3254 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3253 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3252 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_3251 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_3250 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_3249 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_3248 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_3247 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_3246 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_3245 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_3244 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_3243 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_3242 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_3241 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(1'b0), .S(S[23]), .CO(
        C[24]) );
  FA_3240 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3239 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3238 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3237 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3236 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3235 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3234 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3233 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3280 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_106 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3295 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3294 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3293 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3292 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3291 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3290 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3289 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3288 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3287 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3286 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3285 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3284 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_3283 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_3282 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_3281 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_3280 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_3279 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_3278 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_3277 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_3276 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_3275 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_3274 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(1'b0), .S(S[22]), .CO(
        C[23]) );
  FA_3273 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3272 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3271 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3270 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3269 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3268 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3267 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3266 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3265 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3312 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_107 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3327 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3326 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3325 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3324 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3323 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3322 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3321 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3320 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3319 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3318 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3317 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3316 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_3315 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_3314 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_3313 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_3312 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_3311 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_3310 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_3309 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_3308 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_3307 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(1'b0), .S(S[21]), .CO(
        C[22]) );
  FA_3306 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3305 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3304 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3303 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3302 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3301 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3300 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3299 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3298 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3297 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3344 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_108 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3359 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3358 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3357 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3356 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3355 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3354 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3353 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3352 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3351 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3350 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3349 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3348 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_3347 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_3346 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_3345 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_3344 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_3343 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_3342 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_3341 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_3340 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(1'b0), .S(S[20]), .CO(
        C[21]) );
  FA_3339 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3338 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3337 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3336 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3335 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3334 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3333 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3332 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3331 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3330 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3329 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3376 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_109 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3391 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3390 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3389 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3388 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3387 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3386 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3385 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3384 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3383 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3382 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3381 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3380 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_3379 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_3378 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_3377 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_3376 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_3375 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_3374 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_3373 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(1'b0), .S(S[19]), .CO(
        C[20]) );
  FA_3372 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3371 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3370 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3369 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3368 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3367 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3366 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3365 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3364 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3363 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3362 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3361 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3408 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_110 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3423 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3422 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3421 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3420 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3419 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3418 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3417 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3416 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3415 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3414 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3413 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3412 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_3411 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_3410 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_3409 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_3408 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_3407 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_3406 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(1'b0), .S(S[18]), .CO(
        C[19]) );
  FA_3405 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3404 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3403 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3402 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3401 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3400 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3399 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3398 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3397 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3396 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3395 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3394 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3393 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3440 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_111 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3455 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3454 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3453 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3452 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3451 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3450 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3449 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3448 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3447 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3446 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3445 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3444 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_3443 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_3442 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_3441 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_3440 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_3439 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(1'b0), .S(S[17]), .CO(
        C[18]) );
  FA_3438 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3437 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3436 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3435 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3434 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3433 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3432 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3431 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3430 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3429 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3428 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3427 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3426 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3425 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3472 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_112 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3487 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3486 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3485 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3484 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3483 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3482 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3481 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3480 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3479 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3478 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3477 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3476 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_3475 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_3474 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_3473 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_3472 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(1'b0), .S(S[16]), .CO(
        C[17]) );
  FA_3471 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_3470 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3469 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3468 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3467 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3466 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3465 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3464 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3463 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3462 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3461 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3460 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3459 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3458 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3457 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3504 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3512 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3513 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3514 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3515 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3516 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3517 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3518 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3519 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_113 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3519 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3518 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3517 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3516 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3515 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3514 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3513 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3512 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3511 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3510 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3509 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3508 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_3507 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_3506 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_3505 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(1'b0), .S(S[15]), .CO(
        C[16]) );
  FA_3504 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_3503 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_3502 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3501 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3500 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3499 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3498 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3497 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3496 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3495 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3494 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3493 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3492 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3491 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3490 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3489 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3521 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3522 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3523 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3524 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3525 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3526 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3527 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3528 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3529 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3530 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3531 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3532 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3533 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3534 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3535 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3536 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3537 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3538 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3539 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3540 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3541 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3542 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3543 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3544 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3545 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3546 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3547 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3548 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3549 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3550 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3551 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_114 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3551 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3550 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3549 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3548 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3547 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3546 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3545 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3544 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3543 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3542 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3541 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3540 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_3539 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_3538 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(1'b0), .S(S[14]), .CO(
        C[15]) );
  FA_3537 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_3536 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_3535 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_3534 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3533 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3532 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3531 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3530 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3529 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3528 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3527 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3526 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3525 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3524 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3523 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3522 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3521 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3553 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3554 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3555 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3556 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3557 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3558 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3559 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3560 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3561 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3562 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3563 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3564 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3565 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3566 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3567 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3568 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3569 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3570 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3571 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3572 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3573 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3574 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3575 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3576 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3577 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3578 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3579 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3580 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3581 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3582 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3583 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_115 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3583 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3582 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3581 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3580 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3579 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3578 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3577 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3576 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3575 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3574 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3573 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3572 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_3571 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(1'b0), .S(S[13]), .CO(
        C[14]) );
  FA_3570 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_3569 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_3568 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_3567 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_3566 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3565 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3564 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3563 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3562 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3561 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3560 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3559 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3558 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3557 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3556 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3555 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3554 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3553 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3585 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3586 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3587 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3588 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3589 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3590 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3591 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3592 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3593 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3594 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3595 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3596 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3597 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3598 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3599 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3600 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3601 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3602 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3603 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3604 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3605 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3606 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3607 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3608 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3609 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3610 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3611 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3612 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3613 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3614 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3615 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_116 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3615 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3614 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3613 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3612 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3611 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3610 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3609 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3608 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3607 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3606 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3605 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3604 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(1'b0), .S(S[12]), .CO(
        C[13]) );
  FA_3603 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_3602 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_3601 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_3600 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_3599 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_3598 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3597 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3596 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3595 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3594 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3593 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3592 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3591 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3590 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3589 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3588 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3587 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3586 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3585 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3617 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3618 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3619 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3620 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3621 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3622 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3623 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3624 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3625 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3626 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3627 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3628 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3629 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3630 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3631 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3632 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3633 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3634 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3635 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3636 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3637 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3638 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3639 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3640 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3641 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3642 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3643 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3644 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3645 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3646 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3647 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_117 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3647 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3646 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3645 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3644 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3643 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3642 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3641 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3640 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3639 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3638 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3637 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(1'b0), .S(S[11]), .CO(
        C[12]) );
  FA_3636 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_3635 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_3634 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_3633 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_3632 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_3631 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_3630 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3629 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3628 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3627 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3626 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3625 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3624 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3623 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3622 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3621 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3620 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3619 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3618 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3617 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3649 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3650 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3651 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3652 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3653 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3654 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3655 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3656 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3657 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3658 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3659 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3660 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3661 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3662 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3663 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3664 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3665 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3666 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3667 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3668 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3669 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3670 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3671 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3672 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3673 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3674 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3675 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3676 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3677 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3678 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3679 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_118 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3679 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3678 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3677 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3676 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3675 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3674 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3673 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3672 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3671 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3670 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(1'b0), .S(S[10]), .CO(
        C[11]) );
  FA_3669 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_3668 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_3667 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_3666 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_3665 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_3664 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_3663 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_3662 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3661 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3660 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3659 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3658 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3657 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3656 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3655 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3654 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3653 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3652 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3651 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3650 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3649 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3681 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3682 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3683 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3684 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3685 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3686 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3687 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3688 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3689 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3690 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3691 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3692 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3693 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3694 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3695 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3696 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3697 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3698 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3699 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3700 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3701 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3702 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3703 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3704 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3705 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3706 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3707 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3708 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3709 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3710 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3711 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_119 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3711 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3710 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3709 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3708 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3707 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3706 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3705 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3704 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3703 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(1'b0), .S(S[9]), .CO(C[10]) );
  FA_3702 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_3701 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_3700 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_3699 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_3698 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_3697 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_3696 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_3695 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_3694 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3693 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3692 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3691 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3690 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3689 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3688 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3687 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3686 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3685 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3684 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3683 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3682 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3681 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3713 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3714 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3715 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3716 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3717 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3718 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3719 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3720 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3721 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3722 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3723 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3724 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3725 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3726 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3727 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3728 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3729 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3730 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3731 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3732 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3733 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3734 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3735 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3736 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3737 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3738 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3739 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3740 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3741 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3742 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3743 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_120 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3743 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3742 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3741 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3740 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3739 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3738 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3737 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3736 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(1'b0), .S(S[8]), .CO(C[9])
         );
  FA_3735 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_3734 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_3733 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_3732 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_3731 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_3730 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_3729 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_3728 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_3727 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_3726 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3725 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3724 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3723 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3722 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3721 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3720 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3719 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3718 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3717 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3716 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3715 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3714 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3713 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3745 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3746 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3747 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3748 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3749 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3750 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3751 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3752 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3753 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3754 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3755 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3756 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3757 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3758 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3759 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3760 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3761 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3762 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3763 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3764 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3765 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3766 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3767 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3768 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3769 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3770 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3771 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3772 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3773 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3774 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3775 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_121 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3775 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3774 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3773 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3772 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3771 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3770 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3769 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(1'b0), .S(S[7]), .CO(C[8])
         );
  FA_3768 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_3767 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_3766 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_3765 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_3764 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_3763 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_3762 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_3761 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_3760 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_3759 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_3758 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3757 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3756 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3755 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3754 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3753 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3752 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3751 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3750 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3749 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3748 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3747 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3746 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3745 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3777 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3778 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3779 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3780 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3781 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3782 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3783 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3784 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3785 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3786 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3787 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3788 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3789 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3790 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3791 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3792 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3793 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3794 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3795 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3796 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3797 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3798 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3799 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3800 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3801 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3802 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3803 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3804 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3805 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3806 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3807 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_122 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3807 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3806 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3805 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3804 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3803 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3802 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(1'b0), .S(S[6]), .CO(C[7])
         );
  FA_3801 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_3800 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_3799 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_3798 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_3797 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_3796 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_3795 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_3794 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_3793 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_3792 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_3791 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_3790 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3789 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3788 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3787 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3786 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3785 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3784 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3783 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3782 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3781 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3780 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3779 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3778 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3777 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3809 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3810 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3811 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3812 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3813 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3814 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3815 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3816 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3817 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3818 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3819 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3820 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3821 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3822 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3823 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3824 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3825 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3826 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3827 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3828 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3829 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3830 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3831 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3832 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3833 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3834 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3835 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3836 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3837 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3838 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3839 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_123 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3839 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3838 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3837 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3836 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3835 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(1'b0), .S(S[5]), .CO(C[6])
         );
  FA_3834 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_3833 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_3832 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_3831 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_3830 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_3829 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_3828 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_3827 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_3826 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_3825 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_3824 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_3823 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_3822 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3821 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3820 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3819 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3818 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3817 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3816 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3815 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3814 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3813 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3812 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3811 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3810 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3809 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3841 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3842 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3843 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3844 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3845 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3846 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3847 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3848 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3849 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3850 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3851 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3852 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3853 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3854 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3855 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3856 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3857 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3858 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3859 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3860 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3861 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3862 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3863 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3864 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3865 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3866 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3867 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3868 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3869 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3870 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3871 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_124 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3871 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3870 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3869 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3868 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(1'b0), .S(S[4]), .CO(C[5])
         );
  FA_3867 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_3866 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_3865 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_3864 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_3863 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_3862 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_3861 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_3860 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_3859 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_3858 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_3857 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_3856 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_3855 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_3854 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3853 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3852 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3851 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3850 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3849 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3848 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3847 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3846 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3845 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3844 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3843 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3842 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3841 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3873 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3874 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3875 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3876 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3877 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3878 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3879 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3880 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3881 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3882 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3883 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3884 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3885 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3886 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3887 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3888 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3889 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3890 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3891 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3892 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3893 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3894 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3895 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3896 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3897 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3898 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3899 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3900 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3901 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3902 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3903 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_125 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3903 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3902 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3901 \FAINST[3].FA_  ( .A(A[3]), .B(B[3]), .CI(1'b0), .S(S[3]), .CO(C[4])
         );
  FA_3900 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_3899 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_3898 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_3897 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_3896 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_3895 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_3894 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_3893 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_3892 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_3891 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_3890 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_3889 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_3888 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_3887 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_3886 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3885 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3884 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3883 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3882 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3881 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3880 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3879 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3878 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3877 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3876 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3875 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3874 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3873 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3905 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3906 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3907 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3908 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3909 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3910 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3911 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3912 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3913 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3914 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3915 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3916 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3917 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3918 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3919 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3920 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3921 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3922 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3923 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3924 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3925 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3926 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3927 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3928 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3929 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3930 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3931 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3932 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3933 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3934 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3935 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_126 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3935 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3934 \FAINST[2].FA_  ( .A(A[2]), .B(B[2]), .CI(1'b0), .S(S[2]), .CO(C[3])
         );
  FA_3933 \FAINST[3].FA_  ( .A(A[3]), .B(B[3]), .CI(C[3]), .S(S[3]), .CO(C[4])
         );
  FA_3932 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_3931 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_3930 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_3929 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_3928 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_3927 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_3926 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_3925 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_3924 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_3923 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_3922 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_3921 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_3920 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_3919 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_3918 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3917 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3916 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3915 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3914 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3913 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3912 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3911 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3910 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3909 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3908 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3907 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3906 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3905 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3937 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3938 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3939 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3940 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3941 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3942 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3943 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3944 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3945 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3946 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3947 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3948 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3949 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3950 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3951 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3952 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3953 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3954 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3955 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3956 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3957 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3958 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3959 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3960 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3961 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3962 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3963 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3964 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3965 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3966 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3967 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module ADD_N32_127 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;


  FA_3967 \FAINST[1].FA_  ( .A(A[1]), .B(1'b0), .CI(1'b0), .S(S[1]) );
  FA_3966 \FAINST[2].FA_  ( .A(A[2]), .B(1'b0), .CI(1'b0), .S(S[2]) );
  FA_3965 \FAINST[3].FA_  ( .A(A[3]), .B(1'b0), .CI(1'b0), .S(S[3]) );
  FA_3964 \FAINST[4].FA_  ( .A(A[4]), .B(1'b0), .CI(1'b0), .S(S[4]) );
  FA_3963 \FAINST[5].FA_  ( .A(A[5]), .B(1'b0), .CI(1'b0), .S(S[5]) );
  FA_3962 \FAINST[6].FA_  ( .A(A[6]), .B(1'b0), .CI(1'b0), .S(S[6]) );
  FA_3961 \FAINST[7].FA_  ( .A(A[7]), .B(1'b0), .CI(1'b0), .S(S[7]) );
  FA_3960 \FAINST[8].FA_  ( .A(A[8]), .B(1'b0), .CI(1'b0), .S(S[8]) );
  FA_3959 \FAINST[9].FA_  ( .A(A[9]), .B(1'b0), .CI(1'b0), .S(S[9]) );
  FA_3958 \FAINST[10].FA_  ( .A(A[10]), .B(1'b0), .CI(1'b0), .S(S[10]) );
  FA_3957 \FAINST[11].FA_  ( .A(A[11]), .B(1'b0), .CI(1'b0), .S(S[11]) );
  FA_3956 \FAINST[12].FA_  ( .A(A[12]), .B(1'b0), .CI(1'b0), .S(S[12]) );
  FA_3955 \FAINST[13].FA_  ( .A(A[13]), .B(1'b0), .CI(1'b0), .S(S[13]) );
  FA_3954 \FAINST[14].FA_  ( .A(A[14]), .B(1'b0), .CI(1'b0), .S(S[14]) );
  FA_3953 \FAINST[15].FA_  ( .A(A[15]), .B(1'b0), .CI(1'b0), .S(S[15]) );
  FA_3952 \FAINST[16].FA_  ( .A(A[16]), .B(1'b0), .CI(1'b0), .S(S[16]) );
  FA_3951 \FAINST[17].FA_  ( .A(A[17]), .B(1'b0), .CI(1'b0), .S(S[17]) );
  FA_3950 \FAINST[18].FA_  ( .A(A[18]), .B(1'b0), .CI(1'b0), .S(S[18]) );
  FA_3949 \FAINST[19].FA_  ( .A(A[19]), .B(1'b0), .CI(1'b0), .S(S[19]) );
  FA_3948 \FAINST[20].FA_  ( .A(A[20]), .B(1'b0), .CI(1'b0), .S(S[20]) );
  FA_3947 \FAINST[21].FA_  ( .A(A[21]), .B(1'b0), .CI(1'b0), .S(S[21]) );
  FA_3946 \FAINST[22].FA_  ( .A(A[22]), .B(1'b0), .CI(1'b0), .S(S[22]) );
  FA_3945 \FAINST[23].FA_  ( .A(A[23]), .B(1'b0), .CI(1'b0), .S(S[23]) );
  FA_3944 \FAINST[24].FA_  ( .A(A[24]), .B(1'b0), .CI(1'b0), .S(S[24]) );
  FA_3943 \FAINST[25].FA_  ( .A(A[25]), .B(1'b0), .CI(1'b0), .S(S[25]) );
  FA_3942 \FAINST[26].FA_  ( .A(A[26]), .B(1'b0), .CI(1'b0), .S(S[26]) );
  FA_3941 \FAINST[27].FA_  ( .A(A[27]), .B(1'b0), .CI(1'b0), .S(S[27]) );
  FA_3940 \FAINST[28].FA_  ( .A(A[28]), .B(1'b0), .CI(1'b0), .S(S[28]) );
  FA_3939 \FAINST[29].FA_  ( .A(A[29]), .B(1'b0), .CI(1'b0), .S(S[29]) );
  FA_3938 \FAINST[30].FA_  ( .A(A[30]), .B(1'b0), .CI(1'b0), .S(S[30]) );
  FA_3937 \FAINST[31].FA_  ( .A(A[31]), .B(1'b0), .CI(1'b0), .S(S[31]) );
endmodule


module MULT_N32_4 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   \w[31][31] , \w[31][30] , \w[31][29] , \w[31][28] , \w[31][27] ,
         \w[31][26] , \w[31][25] , \w[31][24] , \w[31][23] , \w[31][22] ,
         \w[31][21] , \w[31][20] , \w[31][19] , \w[31][18] , \w[31][17] ,
         \w[31][16] , \w[31][15] , \w[31][14] , \w[31][13] , \w[31][12] ,
         \w[31][11] , \w[31][10] , \w[31][9] , \w[31][8] , \w[31][7] ,
         \w[31][6] , \w[31][5] , \w[31][4] , \w[31][3] , \w[31][2] ,
         \w[31][1] , \w[30][31] , \w[30][30] , \w[30][29] , \w[30][28] ,
         \w[30][27] , \w[30][26] , \w[30][25] , \w[30][24] , \w[30][23] ,
         \w[30][22] , \w[30][21] , \w[30][20] , \w[30][19] , \w[30][18] ,
         \w[30][17] , \w[30][16] , \w[30][15] , \w[30][14] , \w[30][13] ,
         \w[30][12] , \w[30][11] , \w[30][10] , \w[30][9] , \w[30][8] ,
         \w[30][7] , \w[30][6] , \w[30][5] , \w[30][4] , \w[30][3] ,
         \w[30][2] , \w[30][1] , \w[29][31] , \w[29][30] , \w[29][29] ,
         \w[29][28] , \w[29][27] , \w[29][26] , \w[29][25] , \w[29][24] ,
         \w[29][23] , \w[29][22] , \w[29][21] , \w[29][20] , \w[29][19] ,
         \w[29][18] , \w[29][17] , \w[29][16] , \w[29][15] , \w[29][14] ,
         \w[29][13] , \w[29][12] , \w[29][11] , \w[29][10] , \w[29][9] ,
         \w[29][8] , \w[29][7] , \w[29][6] , \w[29][5] , \w[29][4] ,
         \w[29][3] , \w[29][2] , \w[29][1] , \w[28][31] , \w[28][30] ,
         \w[28][29] , \w[28][28] , \w[28][27] , \w[28][26] , \w[28][25] ,
         \w[28][24] , \w[28][23] , \w[28][22] , \w[28][21] , \w[28][20] ,
         \w[28][19] , \w[28][18] , \w[28][17] , \w[28][16] , \w[28][15] ,
         \w[28][14] , \w[28][13] , \w[28][12] , \w[28][11] , \w[28][10] ,
         \w[28][9] , \w[28][8] , \w[28][7] , \w[28][6] , \w[28][5] ,
         \w[28][4] , \w[28][3] , \w[28][2] , \w[28][1] , \w[27][31] ,
         \w[27][30] , \w[27][29] , \w[27][28] , \w[27][27] , \w[27][26] ,
         \w[27][25] , \w[27][24] , \w[27][23] , \w[27][22] , \w[27][21] ,
         \w[27][20] , \w[27][19] , \w[27][18] , \w[27][17] , \w[27][16] ,
         \w[27][15] , \w[27][14] , \w[27][13] , \w[27][12] , \w[27][11] ,
         \w[27][10] , \w[27][9] , \w[27][8] , \w[27][7] , \w[27][6] ,
         \w[27][5] , \w[27][4] , \w[27][3] , \w[27][2] , \w[27][1] ,
         \w[26][31] , \w[26][30] , \w[26][29] , \w[26][28] , \w[26][27] ,
         \w[26][26] , \w[26][25] , \w[26][24] , \w[26][23] , \w[26][22] ,
         \w[26][21] , \w[26][20] , \w[26][19] , \w[26][18] , \w[26][17] ,
         \w[26][16] , \w[26][15] , \w[26][14] , \w[26][13] , \w[26][12] ,
         \w[26][11] , \w[26][10] , \w[26][9] , \w[26][8] , \w[26][7] ,
         \w[26][6] , \w[26][5] , \w[26][4] , \w[26][3] , \w[26][2] ,
         \w[26][1] , \w[25][31] , \w[25][30] , \w[25][29] , \w[25][28] ,
         \w[25][27] , \w[25][26] , \w[25][25] , \w[25][24] , \w[25][23] ,
         \w[25][22] , \w[25][21] , \w[25][20] , \w[25][19] , \w[25][18] ,
         \w[25][17] , \w[25][16] , \w[25][15] , \w[25][14] , \w[25][13] ,
         \w[25][12] , \w[25][11] , \w[25][10] , \w[25][9] , \w[25][8] ,
         \w[25][7] , \w[25][6] , \w[25][5] , \w[25][4] , \w[25][3] ,
         \w[25][2] , \w[25][1] , \w[24][31] , \w[24][30] , \w[24][29] ,
         \w[24][28] , \w[24][27] , \w[24][26] , \w[24][25] , \w[24][24] ,
         \w[24][23] , \w[24][22] , \w[24][21] , \w[24][20] , \w[24][19] ,
         \w[24][18] , \w[24][17] , \w[24][16] , \w[24][15] , \w[24][14] ,
         \w[24][13] , \w[24][12] , \w[24][11] , \w[24][10] , \w[24][9] ,
         \w[24][8] , \w[24][7] , \w[24][6] , \w[24][5] , \w[24][4] ,
         \w[24][3] , \w[24][2] , \w[24][1] , \w[23][31] , \w[23][30] ,
         \w[23][29] , \w[23][28] , \w[23][27] , \w[23][26] , \w[23][25] ,
         \w[23][24] , \w[23][23] , \w[23][22] , \w[23][21] , \w[23][20] ,
         \w[23][19] , \w[23][18] , \w[23][17] , \w[23][16] , \w[23][15] ,
         \w[23][14] , \w[23][13] , \w[23][12] , \w[23][11] , \w[23][10] ,
         \w[23][9] , \w[23][8] , \w[23][7] , \w[23][6] , \w[23][5] ,
         \w[23][4] , \w[23][3] , \w[23][2] , \w[23][1] , \w[22][31] ,
         \w[22][30] , \w[22][29] , \w[22][28] , \w[22][27] , \w[22][26] ,
         \w[22][25] , \w[22][24] , \w[22][23] , \w[22][22] , \w[22][21] ,
         \w[22][20] , \w[22][19] , \w[22][18] , \w[22][17] , \w[22][16] ,
         \w[22][15] , \w[22][14] , \w[22][13] , \w[22][12] , \w[22][11] ,
         \w[22][10] , \w[22][9] , \w[22][8] , \w[22][7] , \w[22][6] ,
         \w[22][5] , \w[22][4] , \w[22][3] , \w[22][2] , \w[22][1] ,
         \w[21][31] , \w[21][30] , \w[21][29] , \w[21][28] , \w[21][27] ,
         \w[21][26] , \w[21][25] , \w[21][24] , \w[21][23] , \w[21][22] ,
         \w[21][21] , \w[21][20] , \w[21][19] , \w[21][18] , \w[21][17] ,
         \w[21][16] , \w[21][15] , \w[21][14] , \w[21][13] , \w[21][12] ,
         \w[21][11] , \w[21][10] , \w[21][9] , \w[21][8] , \w[21][7] ,
         \w[21][6] , \w[21][5] , \w[21][4] , \w[21][3] , \w[21][2] ,
         \w[21][1] , \w[20][31] , \w[20][30] , \w[20][29] , \w[20][28] ,
         \w[20][27] , \w[20][26] , \w[20][25] , \w[20][24] , \w[20][23] ,
         \w[20][22] , \w[20][21] , \w[20][20] , \w[20][19] , \w[20][18] ,
         \w[20][17] , \w[20][16] , \w[20][15] , \w[20][14] , \w[20][13] ,
         \w[20][12] , \w[20][11] , \w[20][10] , \w[20][9] , \w[20][8] ,
         \w[20][7] , \w[20][6] , \w[20][5] , \w[20][4] , \w[20][3] ,
         \w[20][2] , \w[20][1] , \w[19][31] , \w[19][30] , \w[19][29] ,
         \w[19][28] , \w[19][27] , \w[19][26] , \w[19][25] , \w[19][24] ,
         \w[19][23] , \w[19][22] , \w[19][21] , \w[19][20] , \w[19][19] ,
         \w[19][18] , \w[19][17] , \w[19][16] , \w[19][15] , \w[19][14] ,
         \w[19][13] , \w[19][12] , \w[19][11] , \w[19][10] , \w[19][9] ,
         \w[19][8] , \w[19][7] , \w[19][6] , \w[19][5] , \w[19][4] ,
         \w[19][3] , \w[19][2] , \w[19][1] , \w[18][31] , \w[18][30] ,
         \w[18][29] , \w[18][28] , \w[18][27] , \w[18][26] , \w[18][25] ,
         \w[18][24] , \w[18][23] , \w[18][22] , \w[18][21] , \w[18][20] ,
         \w[18][19] , \w[18][18] , \w[18][17] , \w[18][16] , \w[18][15] ,
         \w[18][14] , \w[18][13] , \w[18][12] , \w[18][11] , \w[18][10] ,
         \w[18][9] , \w[18][8] , \w[18][7] , \w[18][6] , \w[18][5] ,
         \w[18][4] , \w[18][3] , \w[18][2] , \w[18][1] , \w[17][31] ,
         \w[17][30] , \w[17][29] , \w[17][28] , \w[17][27] , \w[17][26] ,
         \w[17][25] , \w[17][24] , \w[17][23] , \w[17][22] , \w[17][21] ,
         \w[17][20] , \w[17][19] , \w[17][18] , \w[17][17] , \w[17][16] ,
         \w[17][15] , \w[17][14] , \w[17][13] , \w[17][12] , \w[17][11] ,
         \w[17][10] , \w[17][9] , \w[17][8] , \w[17][7] , \w[17][6] ,
         \w[17][5] , \w[17][4] , \w[17][3] , \w[17][2] , \w[17][1] ,
         \w[16][31] , \w[16][30] , \w[16][29] , \w[16][28] , \w[16][27] ,
         \w[16][26] , \w[16][25] , \w[16][24] , \w[16][23] , \w[16][22] ,
         \w[16][21] , \w[16][20] , \w[16][19] , \w[16][18] , \w[16][17] ,
         \w[16][16] , \w[16][15] , \w[16][14] , \w[16][13] , \w[16][12] ,
         \w[16][11] , \w[16][10] , \w[16][9] , \w[16][8] , \w[16][7] ,
         \w[16][6] , \w[16][5] , \w[16][4] , \w[16][3] , \w[16][2] ,
         \w[16][1] , \w[15][31] , \w[15][30] , \w[15][29] , \w[15][28] ,
         \w[15][27] , \w[15][26] , \w[15][25] , \w[15][24] , \w[15][23] ,
         \w[15][22] , \w[15][21] , \w[15][20] , \w[15][19] , \w[15][18] ,
         \w[15][17] , \w[15][16] , \w[15][15] , \w[15][14] , \w[15][13] ,
         \w[15][12] , \w[15][11] , \w[15][10] , \w[15][9] , \w[15][8] ,
         \w[15][7] , \w[15][6] , \w[15][5] , \w[15][4] , \w[15][3] ,
         \w[15][2] , \w[15][1] , \w[14][31] , \w[14][30] , \w[14][29] ,
         \w[14][28] , \w[14][27] , \w[14][26] , \w[14][25] , \w[14][24] ,
         \w[14][23] , \w[14][22] , \w[14][21] , \w[14][20] , \w[14][19] ,
         \w[14][18] , \w[14][17] , \w[14][16] , \w[14][15] , \w[14][14] ,
         \w[14][13] , \w[14][12] , \w[14][11] , \w[14][10] , \w[14][9] ,
         \w[14][8] , \w[14][7] , \w[14][6] , \w[14][5] , \w[14][4] ,
         \w[14][3] , \w[14][2] , \w[14][1] , \w[13][31] , \w[13][30] ,
         \w[13][29] , \w[13][28] , \w[13][27] , \w[13][26] , \w[13][25] ,
         \w[13][24] , \w[13][23] , \w[13][22] , \w[13][21] , \w[13][20] ,
         \w[13][19] , \w[13][18] , \w[13][17] , \w[13][16] , \w[13][15] ,
         \w[13][14] , \w[13][13] , \w[13][12] , \w[13][11] , \w[13][10] ,
         \w[13][9] , \w[13][8] , \w[13][7] , \w[13][6] , \w[13][5] ,
         \w[13][4] , \w[13][3] , \w[13][2] , \w[13][1] , \w[12][31] ,
         \w[12][30] , \w[12][29] , \w[12][28] , \w[12][27] , \w[12][26] ,
         \w[12][25] , \w[12][24] , \w[12][23] , \w[12][22] , \w[12][21] ,
         \w[12][20] , \w[12][19] , \w[12][18] , \w[12][17] , \w[12][16] ,
         \w[12][15] , \w[12][14] , \w[12][13] , \w[12][12] , \w[12][11] ,
         \w[12][10] , \w[12][9] , \w[12][8] , \w[12][7] , \w[12][6] ,
         \w[12][5] , \w[12][4] , \w[12][3] , \w[12][2] , \w[12][1] ,
         \w[11][31] , \w[11][30] , \w[11][29] , \w[11][28] , \w[11][27] ,
         \w[11][26] , \w[11][25] , \w[11][24] , \w[11][23] , \w[11][22] ,
         \w[11][21] , \w[11][20] , \w[11][19] , \w[11][18] , \w[11][17] ,
         \w[11][16] , \w[11][15] , \w[11][14] , \w[11][13] , \w[11][12] ,
         \w[11][11] , \w[11][10] , \w[11][9] , \w[11][8] , \w[11][7] ,
         \w[11][6] , \w[11][5] , \w[11][4] , \w[11][3] , \w[11][2] ,
         \w[11][1] , \w[10][31] , \w[10][30] , \w[10][29] , \w[10][28] ,
         \w[10][27] , \w[10][26] , \w[10][25] , \w[10][24] , \w[10][23] ,
         \w[10][22] , \w[10][21] , \w[10][20] , \w[10][19] , \w[10][18] ,
         \w[10][17] , \w[10][16] , \w[10][15] , \w[10][14] , \w[10][13] ,
         \w[10][12] , \w[10][11] , \w[10][10] , \w[10][9] , \w[10][8] ,
         \w[10][7] , \w[10][6] , \w[10][5] , \w[10][4] , \w[10][3] ,
         \w[10][2] , \w[10][1] , \w[9][31] , \w[9][30] , \w[9][29] ,
         \w[9][28] , \w[9][27] , \w[9][26] , \w[9][25] , \w[9][24] ,
         \w[9][23] , \w[9][22] , \w[9][21] , \w[9][20] , \w[9][19] ,
         \w[9][18] , \w[9][17] , \w[9][16] , \w[9][15] , \w[9][14] ,
         \w[9][13] , \w[9][12] , \w[9][11] , \w[9][10] , \w[9][9] , \w[9][8] ,
         \w[9][7] , \w[9][6] , \w[9][5] , \w[9][4] , \w[9][3] , \w[9][2] ,
         \w[9][1] , \w[8][31] , \w[8][30] , \w[8][29] , \w[8][28] , \w[8][27] ,
         \w[8][26] , \w[8][25] , \w[8][24] , \w[8][23] , \w[8][22] ,
         \w[8][21] , \w[8][20] , \w[8][19] , \w[8][18] , \w[8][17] ,
         \w[8][16] , \w[8][15] , \w[8][14] , \w[8][13] , \w[8][12] ,
         \w[8][11] , \w[8][10] , \w[8][9] , \w[8][8] , \w[8][7] , \w[8][6] ,
         \w[8][5] , \w[8][4] , \w[8][3] , \w[8][2] , \w[8][1] , \w[7][31] ,
         \w[7][30] , \w[7][29] , \w[7][28] , \w[7][27] , \w[7][26] ,
         \w[7][25] , \w[7][24] , \w[7][23] , \w[7][22] , \w[7][21] ,
         \w[7][20] , \w[7][19] , \w[7][18] , \w[7][17] , \w[7][16] ,
         \w[7][15] , \w[7][14] , \w[7][13] , \w[7][12] , \w[7][11] ,
         \w[7][10] , \w[7][9] , \w[7][8] , \w[7][7] , \w[7][6] , \w[7][5] ,
         \w[7][4] , \w[7][3] , \w[7][2] , \w[7][1] , \w[6][31] , \w[6][30] ,
         \w[6][29] , \w[6][28] , \w[6][27] , \w[6][26] , \w[6][25] ,
         \w[6][24] , \w[6][23] , \w[6][22] , \w[6][21] , \w[6][20] ,
         \w[6][19] , \w[6][18] , \w[6][17] , \w[6][16] , \w[6][15] ,
         \w[6][14] , \w[6][13] , \w[6][12] , \w[6][11] , \w[6][10] , \w[6][9] ,
         \w[6][8] , \w[6][7] , \w[6][6] , \w[6][5] , \w[6][4] , \w[6][3] ,
         \w[6][2] , \w[6][1] , \w[5][31] , \w[5][30] , \w[5][29] , \w[5][28] ,
         \w[5][27] , \w[5][26] , \w[5][25] , \w[5][24] , \w[5][23] ,
         \w[5][22] , \w[5][21] , \w[5][20] , \w[5][19] , \w[5][18] ,
         \w[5][17] , \w[5][16] , \w[5][15] , \w[5][14] , \w[5][13] ,
         \w[5][12] , \w[5][11] , \w[5][10] , \w[5][9] , \w[5][8] , \w[5][7] ,
         \w[5][6] , \w[5][5] , \w[5][4] , \w[5][3] , \w[5][2] , \w[5][1] ,
         \w[4][31] , \w[4][30] , \w[4][29] , \w[4][28] , \w[4][27] ,
         \w[4][26] , \w[4][25] , \w[4][24] , \w[4][23] , \w[4][22] ,
         \w[4][21] , \w[4][20] , \w[4][19] , \w[4][18] , \w[4][17] ,
         \w[4][16] , \w[4][15] , \w[4][14] , \w[4][13] , \w[4][12] ,
         \w[4][11] , \w[4][10] , \w[4][9] , \w[4][8] , \w[4][7] , \w[4][6] ,
         \w[4][5] , \w[4][4] , \w[4][3] , \w[4][2] , \w[4][1] , \w[3][31] ,
         \w[3][30] , \w[3][29] , \w[3][28] , \w[3][27] , \w[3][26] ,
         \w[3][25] , \w[3][24] , \w[3][23] , \w[3][22] , \w[3][21] ,
         \w[3][20] , \w[3][19] , \w[3][18] , \w[3][17] , \w[3][16] ,
         \w[3][15] , \w[3][14] , \w[3][13] , \w[3][12] , \w[3][11] ,
         \w[3][10] , \w[3][9] , \w[3][8] , \w[3][7] , \w[3][6] , \w[3][5] ,
         \w[3][4] , \w[3][3] , \w[3][2] , \w[3][1] , \w[2][31] , \w[2][30] ,
         \w[2][29] , \w[2][28] , \w[2][27] , \w[2][26] , \w[2][25] ,
         \w[2][24] , \w[2][23] , \w[2][22] , \w[2][21] , \w[2][20] ,
         \w[2][19] , \w[2][18] , \w[2][17] , \w[2][16] , \w[2][15] ,
         \w[2][14] , \w[2][13] , \w[2][12] , \w[2][11] , \w[2][10] , \w[2][9] ,
         \w[2][8] , \w[2][7] , \w[2][6] , \w[2][5] , \w[2][4] , \w[2][3] ,
         \w[2][2] , \w[2][1] , \_0_net_[31] , \_0_net_[30] , \_0_net_[29] ,
         \_0_net_[28] , \_0_net_[27] , \_0_net_[26] , \_0_net_[25] ,
         \_0_net_[24] , \_0_net_[23] , \_0_net_[22] , \_0_net_[21] ,
         \_0_net_[20] , \_0_net_[19] , \_0_net_[18] , \_0_net_[17] ,
         \_0_net_[16] , \_0_net_[15] , \_0_net_[14] , \_0_net_[13] ,
         \_0_net_[12] , \_0_net_[11] , \_0_net_[10] , \_0_net_[9] ,
         \_0_net_[8] , \_0_net_[7] , \_0_net_[6] , \_0_net_[5] , \_0_net_[4] ,
         \_0_net_[3] , \_0_net_[2] , \_0_net_[1] , \_2_net_[31] ,
         \_2_net_[30] , \_2_net_[29] , \_2_net_[28] , \_2_net_[27] ,
         \_2_net_[26] , \_2_net_[25] , \_2_net_[24] , \_2_net_[23] ,
         \_2_net_[22] , \_2_net_[21] , \_2_net_[20] , \_2_net_[19] ,
         \_2_net_[18] , \_2_net_[17] , \_2_net_[16] , \_2_net_[15] ,
         \_2_net_[14] , \_2_net_[13] , \_2_net_[12] , \_2_net_[11] ,
         \_2_net_[10] , \_2_net_[9] , \_2_net_[8] , \_2_net_[7] , \_2_net_[6] ,
         \_2_net_[5] , \_2_net_[4] , \_2_net_[3] , \_2_net_[2] , \_4_net_[31] ,
         \_4_net_[30] , \_4_net_[29] , \_4_net_[28] , \_4_net_[27] ,
         \_4_net_[26] , \_4_net_[25] , \_4_net_[24] , \_4_net_[23] ,
         \_4_net_[22] , \_4_net_[21] , \_4_net_[20] , \_4_net_[19] ,
         \_4_net_[18] , \_4_net_[17] , \_4_net_[16] , \_4_net_[15] ,
         \_4_net_[14] , \_4_net_[13] , \_4_net_[12] , \_4_net_[11] ,
         \_4_net_[10] , \_4_net_[9] , \_4_net_[8] , \_4_net_[7] , \_4_net_[6] ,
         \_4_net_[5] , \_4_net_[4] , \_4_net_[3] , \_6_net_[31] ,
         \_6_net_[30] , \_6_net_[29] , \_6_net_[28] , \_6_net_[27] ,
         \_6_net_[26] , \_6_net_[25] , \_6_net_[24] , \_6_net_[23] ,
         \_6_net_[22] , \_6_net_[21] , \_6_net_[20] , \_6_net_[19] ,
         \_6_net_[18] , \_6_net_[17] , \_6_net_[16] , \_6_net_[15] ,
         \_6_net_[14] , \_6_net_[13] , \_6_net_[12] , \_6_net_[11] ,
         \_6_net_[10] , \_6_net_[9] , \_6_net_[8] , \_6_net_[7] , \_6_net_[6] ,
         \_6_net_[5] , \_6_net_[4] , \_8_net_[31] , \_8_net_[30] ,
         \_8_net_[29] , \_8_net_[28] , \_8_net_[27] , \_8_net_[26] ,
         \_8_net_[25] , \_8_net_[24] , \_8_net_[23] , \_8_net_[22] ,
         \_8_net_[21] , \_8_net_[20] , \_8_net_[19] , \_8_net_[18] ,
         \_8_net_[17] , \_8_net_[16] , \_8_net_[15] , \_8_net_[14] ,
         \_8_net_[13] , \_8_net_[12] , \_8_net_[11] , \_8_net_[10] ,
         \_8_net_[9] , \_8_net_[8] , \_8_net_[7] , \_8_net_[6] , \_8_net_[5] ,
         \_10_net_[31] , \_10_net_[30] , \_10_net_[29] , \_10_net_[28] ,
         \_10_net_[27] , \_10_net_[26] , \_10_net_[25] , \_10_net_[24] ,
         \_10_net_[23] , \_10_net_[22] , \_10_net_[21] , \_10_net_[20] ,
         \_10_net_[19] , \_10_net_[18] , \_10_net_[17] , \_10_net_[16] ,
         \_10_net_[15] , \_10_net_[14] , \_10_net_[13] , \_10_net_[12] ,
         \_10_net_[11] , \_10_net_[10] , \_10_net_[9] , \_10_net_[8] ,
         \_10_net_[7] , \_10_net_[6] , \_12_net_[31] , \_12_net_[30] ,
         \_12_net_[29] , \_12_net_[28] , \_12_net_[27] , \_12_net_[26] ,
         \_12_net_[25] , \_12_net_[24] , \_12_net_[23] , \_12_net_[22] ,
         \_12_net_[21] , \_12_net_[20] , \_12_net_[19] , \_12_net_[18] ,
         \_12_net_[17] , \_12_net_[16] , \_12_net_[15] , \_12_net_[14] ,
         \_12_net_[13] , \_12_net_[12] , \_12_net_[11] , \_12_net_[10] ,
         \_12_net_[9] , \_12_net_[8] , \_12_net_[7] , \_14_net_[31] ,
         \_14_net_[30] , \_14_net_[29] , \_14_net_[28] , \_14_net_[27] ,
         \_14_net_[26] , \_14_net_[25] , \_14_net_[24] , \_14_net_[23] ,
         \_14_net_[22] , \_14_net_[21] , \_14_net_[20] , \_14_net_[19] ,
         \_14_net_[18] , \_14_net_[17] , \_14_net_[16] , \_14_net_[15] ,
         \_14_net_[14] , \_14_net_[13] , \_14_net_[12] , \_14_net_[11] ,
         \_14_net_[10] , \_14_net_[9] , \_14_net_[8] , \_16_net_[31] ,
         \_16_net_[30] , \_16_net_[29] , \_16_net_[28] , \_16_net_[27] ,
         \_16_net_[26] , \_16_net_[25] , \_16_net_[24] , \_16_net_[23] ,
         \_16_net_[22] , \_16_net_[21] , \_16_net_[20] , \_16_net_[19] ,
         \_16_net_[18] , \_16_net_[17] , \_16_net_[16] , \_16_net_[15] ,
         \_16_net_[14] , \_16_net_[13] , \_16_net_[12] , \_16_net_[11] ,
         \_16_net_[10] , \_16_net_[9] , \_18_net_[31] , \_18_net_[30] ,
         \_18_net_[29] , \_18_net_[28] , \_18_net_[27] , \_18_net_[26] ,
         \_18_net_[25] , \_18_net_[24] , \_18_net_[23] , \_18_net_[22] ,
         \_18_net_[21] , \_18_net_[20] , \_18_net_[19] , \_18_net_[18] ,
         \_18_net_[17] , \_18_net_[16] , \_18_net_[15] , \_18_net_[14] ,
         \_18_net_[13] , \_18_net_[12] , \_18_net_[11] , \_18_net_[10] ,
         \_20_net_[31] , \_20_net_[30] , \_20_net_[29] , \_20_net_[28] ,
         \_20_net_[27] , \_20_net_[26] , \_20_net_[25] , \_20_net_[24] ,
         \_20_net_[23] , \_20_net_[22] , \_20_net_[21] , \_20_net_[20] ,
         \_20_net_[19] , \_20_net_[18] , \_20_net_[17] , \_20_net_[16] ,
         \_20_net_[15] , \_20_net_[14] , \_20_net_[13] , \_20_net_[12] ,
         \_20_net_[11] , \_22_net_[31] , \_22_net_[30] , \_22_net_[29] ,
         \_22_net_[28] , \_22_net_[27] , \_22_net_[26] , \_22_net_[25] ,
         \_22_net_[24] , \_22_net_[23] , \_22_net_[22] , \_22_net_[21] ,
         \_22_net_[20] , \_22_net_[19] , \_22_net_[18] , \_22_net_[17] ,
         \_22_net_[16] , \_22_net_[15] , \_22_net_[14] , \_22_net_[13] ,
         \_22_net_[12] , \_24_net_[31] , \_24_net_[30] , \_24_net_[29] ,
         \_24_net_[28] , \_24_net_[27] , \_24_net_[26] , \_24_net_[25] ,
         \_24_net_[24] , \_24_net_[23] , \_24_net_[22] , \_24_net_[21] ,
         \_24_net_[20] , \_24_net_[19] , \_24_net_[18] , \_24_net_[17] ,
         \_24_net_[16] , \_24_net_[15] , \_24_net_[14] , \_24_net_[13] ,
         \_26_net_[31] , \_26_net_[30] , \_26_net_[29] , \_26_net_[28] ,
         \_26_net_[27] , \_26_net_[26] , \_26_net_[25] , \_26_net_[24] ,
         \_26_net_[23] , \_26_net_[22] , \_26_net_[21] , \_26_net_[20] ,
         \_26_net_[19] , \_26_net_[18] , \_26_net_[17] , \_26_net_[16] ,
         \_26_net_[15] , \_26_net_[14] , \_28_net_[31] , \_28_net_[30] ,
         \_28_net_[29] , \_28_net_[28] , \_28_net_[27] , \_28_net_[26] ,
         \_28_net_[25] , \_28_net_[24] , \_28_net_[23] , \_28_net_[22] ,
         \_28_net_[21] , \_28_net_[20] , \_28_net_[19] , \_28_net_[18] ,
         \_28_net_[17] , \_28_net_[16] , \_28_net_[15] , \_30_net_[31] ,
         \_30_net_[30] , \_30_net_[29] , \_30_net_[28] , \_30_net_[27] ,
         \_30_net_[26] , \_30_net_[25] , \_30_net_[24] , \_30_net_[23] ,
         \_30_net_[22] , \_30_net_[21] , \_30_net_[20] , \_30_net_[19] ,
         \_30_net_[18] , \_30_net_[17] , \_30_net_[16] , \_32_net_[31] ,
         \_32_net_[30] , \_32_net_[29] , \_32_net_[28] , \_32_net_[27] ,
         \_32_net_[26] , \_32_net_[25] , \_32_net_[24] , \_32_net_[23] ,
         \_32_net_[22] , \_32_net_[21] , \_32_net_[20] , \_32_net_[19] ,
         \_32_net_[18] , \_32_net_[17] , \_34_net_[31] , \_34_net_[30] ,
         \_34_net_[29] , \_34_net_[28] , \_34_net_[27] , \_34_net_[26] ,
         \_34_net_[25] , \_34_net_[24] , \_34_net_[23] , \_34_net_[22] ,
         \_34_net_[21] , \_34_net_[20] , \_34_net_[19] , \_34_net_[18] ,
         \_36_net_[31] , \_36_net_[30] , \_36_net_[29] , \_36_net_[28] ,
         \_36_net_[27] , \_36_net_[26] , \_36_net_[25] , \_36_net_[24] ,
         \_36_net_[23] , \_36_net_[22] , \_36_net_[21] , \_36_net_[20] ,
         \_36_net_[19] , \_38_net_[31] , \_38_net_[30] , \_38_net_[29] ,
         \_38_net_[28] , \_38_net_[27] , \_38_net_[26] , \_38_net_[25] ,
         \_38_net_[24] , \_38_net_[23] , \_38_net_[22] , \_38_net_[21] ,
         \_38_net_[20] , \_40_net_[31] , \_40_net_[30] , \_40_net_[29] ,
         \_40_net_[28] , \_40_net_[27] , \_40_net_[26] , \_40_net_[25] ,
         \_40_net_[24] , \_40_net_[23] , \_40_net_[22] , \_40_net_[21] ,
         \_42_net_[31] , \_42_net_[30] , \_42_net_[29] , \_42_net_[28] ,
         \_42_net_[27] , \_42_net_[26] , \_42_net_[25] , \_42_net_[24] ,
         \_42_net_[23] , \_42_net_[22] , \_44_net_[31] , \_44_net_[30] ,
         \_44_net_[29] , \_44_net_[28] , \_44_net_[27] , \_44_net_[26] ,
         \_44_net_[25] , \_44_net_[24] , \_44_net_[23] , \_46_net_[31] ,
         \_46_net_[30] , \_46_net_[29] , \_46_net_[28] , \_46_net_[27] ,
         \_46_net_[26] , \_46_net_[25] , \_46_net_[24] , \_48_net_[31] ,
         \_48_net_[30] , \_48_net_[29] , \_48_net_[28] , \_48_net_[27] ,
         \_48_net_[26] , \_48_net_[25] , \_50_net_[31] , \_50_net_[30] ,
         \_50_net_[29] , \_50_net_[28] , \_50_net_[27] , \_50_net_[26] ,
         \_52_net_[31] , \_52_net_[30] , \_52_net_[29] , \_52_net_[28] ,
         \_52_net_[27] , \_54_net_[31] , \_54_net_[30] , \_54_net_[29] ,
         \_54_net_[28] , \_56_net_[31] , \_56_net_[30] , \_56_net_[29] ,
         \_58_net_[31] , \_58_net_[30] , \_60_net_[31] ;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30;

  ADD_N32_127 \FAINST[1].ADD_  ( .A({\_0_net_[31] , \_0_net_[30] , 
        \_0_net_[29] , \_0_net_[28] , \_0_net_[27] , \_0_net_[26] , 
        \_0_net_[25] , \_0_net_[24] , \_0_net_[23] , \_0_net_[22] , 
        \_0_net_[21] , \_0_net_[20] , \_0_net_[19] , \_0_net_[18] , 
        \_0_net_[17] , \_0_net_[16] , \_0_net_[15] , \_0_net_[14] , 
        \_0_net_[13] , \_0_net_[12] , \_0_net_[11] , \_0_net_[10] , 
        \_0_net_[9] , \_0_net_[8] , \_0_net_[7] , \_0_net_[6] , \_0_net_[5] , 
        \_0_net_[4] , \_0_net_[3] , \_0_net_[2] , \_0_net_[1] , 1'b0}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .S({
        \w[2][31] , \w[2][30] , \w[2][29] , \w[2][28] , \w[2][27] , \w[2][26] , 
        \w[2][25] , \w[2][24] , \w[2][23] , \w[2][22] , \w[2][21] , \w[2][20] , 
        \w[2][19] , \w[2][18] , \w[2][17] , \w[2][16] , \w[2][15] , \w[2][14] , 
        \w[2][13] , \w[2][12] , \w[2][11] , \w[2][10] , \w[2][9] , \w[2][8] , 
        \w[2][7] , \w[2][6] , \w[2][5] , \w[2][4] , \w[2][3] , \w[2][2] , 
        \w[2][1] , SYNOPSYS_UNCONNECTED__0}) );
  ADD_N32_126 \FAINST[2].ADD_  ( .A({\_2_net_[31] , \_2_net_[30] , 
        \_2_net_[29] , \_2_net_[28] , \_2_net_[27] , \_2_net_[26] , 
        \_2_net_[25] , \_2_net_[24] , \_2_net_[23] , \_2_net_[22] , 
        \_2_net_[21] , \_2_net_[20] , \_2_net_[19] , \_2_net_[18] , 
        \_2_net_[17] , \_2_net_[16] , \_2_net_[15] , \_2_net_[14] , 
        \_2_net_[13] , \_2_net_[12] , \_2_net_[11] , \_2_net_[10] , 
        \_2_net_[9] , \_2_net_[8] , \_2_net_[7] , \_2_net_[6] , \_2_net_[5] , 
        \_2_net_[4] , \_2_net_[3] , \_2_net_[2] , 1'b0, 1'b0}), .B({\w[2][31] , 
        \w[2][30] , \w[2][29] , \w[2][28] , \w[2][27] , \w[2][26] , \w[2][25] , 
        \w[2][24] , \w[2][23] , \w[2][22] , \w[2][21] , \w[2][20] , \w[2][19] , 
        \w[2][18] , \w[2][17] , \w[2][16] , \w[2][15] , \w[2][14] , \w[2][13] , 
        \w[2][12] , \w[2][11] , \w[2][10] , \w[2][9] , \w[2][8] , \w[2][7] , 
        \w[2][6] , \w[2][5] , \w[2][4] , \w[2][3] , \w[2][2] , \w[2][1] , 1'b0}), .CI(1'b0), .S({\w[3][31] , \w[3][30] , \w[3][29] , \w[3][28] , \w[3][27] , 
        \w[3][26] , \w[3][25] , \w[3][24] , \w[3][23] , \w[3][22] , \w[3][21] , 
        \w[3][20] , \w[3][19] , \w[3][18] , \w[3][17] , \w[3][16] , \w[3][15] , 
        \w[3][14] , \w[3][13] , \w[3][12] , \w[3][11] , \w[3][10] , \w[3][9] , 
        \w[3][8] , \w[3][7] , \w[3][6] , \w[3][5] , \w[3][4] , \w[3][3] , 
        \w[3][2] , \w[3][1] , SYNOPSYS_UNCONNECTED__1}) );
  ADD_N32_125 \FAINST[3].ADD_  ( .A({\_4_net_[31] , \_4_net_[30] , 
        \_4_net_[29] , \_4_net_[28] , \_4_net_[27] , \_4_net_[26] , 
        \_4_net_[25] , \_4_net_[24] , \_4_net_[23] , \_4_net_[22] , 
        \_4_net_[21] , \_4_net_[20] , \_4_net_[19] , \_4_net_[18] , 
        \_4_net_[17] , \_4_net_[16] , \_4_net_[15] , \_4_net_[14] , 
        \_4_net_[13] , \_4_net_[12] , \_4_net_[11] , \_4_net_[10] , 
        \_4_net_[9] , \_4_net_[8] , \_4_net_[7] , \_4_net_[6] , \_4_net_[5] , 
        \_4_net_[4] , \_4_net_[3] , 1'b0, 1'b0, 1'b0}), .B({\w[3][31] , 
        \w[3][30] , \w[3][29] , \w[3][28] , \w[3][27] , \w[3][26] , \w[3][25] , 
        \w[3][24] , \w[3][23] , \w[3][22] , \w[3][21] , \w[3][20] , \w[3][19] , 
        \w[3][18] , \w[3][17] , \w[3][16] , \w[3][15] , \w[3][14] , \w[3][13] , 
        \w[3][12] , \w[3][11] , \w[3][10] , \w[3][9] , \w[3][8] , \w[3][7] , 
        \w[3][6] , \w[3][5] , \w[3][4] , \w[3][3] , \w[3][2] , \w[3][1] , 1'b0}), .CI(1'b0), .S({\w[4][31] , \w[4][30] , \w[4][29] , \w[4][28] , \w[4][27] , 
        \w[4][26] , \w[4][25] , \w[4][24] , \w[4][23] , \w[4][22] , \w[4][21] , 
        \w[4][20] , \w[4][19] , \w[4][18] , \w[4][17] , \w[4][16] , \w[4][15] , 
        \w[4][14] , \w[4][13] , \w[4][12] , \w[4][11] , \w[4][10] , \w[4][9] , 
        \w[4][8] , \w[4][7] , \w[4][6] , \w[4][5] , \w[4][4] , \w[4][3] , 
        \w[4][2] , \w[4][1] , SYNOPSYS_UNCONNECTED__2}) );
  ADD_N32_124 \FAINST[4].ADD_  ( .A({\_6_net_[31] , \_6_net_[30] , 
        \_6_net_[29] , \_6_net_[28] , \_6_net_[27] , \_6_net_[26] , 
        \_6_net_[25] , \_6_net_[24] , \_6_net_[23] , \_6_net_[22] , 
        \_6_net_[21] , \_6_net_[20] , \_6_net_[19] , \_6_net_[18] , 
        \_6_net_[17] , \_6_net_[16] , \_6_net_[15] , \_6_net_[14] , 
        \_6_net_[13] , \_6_net_[12] , \_6_net_[11] , \_6_net_[10] , 
        \_6_net_[9] , \_6_net_[8] , \_6_net_[7] , \_6_net_[6] , \_6_net_[5] , 
        \_6_net_[4] , 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[4][31] , \w[4][30] , 
        \w[4][29] , \w[4][28] , \w[4][27] , \w[4][26] , \w[4][25] , \w[4][24] , 
        \w[4][23] , \w[4][22] , \w[4][21] , \w[4][20] , \w[4][19] , \w[4][18] , 
        \w[4][17] , \w[4][16] , \w[4][15] , \w[4][14] , \w[4][13] , \w[4][12] , 
        \w[4][11] , \w[4][10] , \w[4][9] , \w[4][8] , \w[4][7] , \w[4][6] , 
        \w[4][5] , \w[4][4] , \w[4][3] , \w[4][2] , \w[4][1] , 1'b0}), .CI(
        1'b0), .S({\w[5][31] , \w[5][30] , \w[5][29] , \w[5][28] , \w[5][27] , 
        \w[5][26] , \w[5][25] , \w[5][24] , \w[5][23] , \w[5][22] , \w[5][21] , 
        \w[5][20] , \w[5][19] , \w[5][18] , \w[5][17] , \w[5][16] , \w[5][15] , 
        \w[5][14] , \w[5][13] , \w[5][12] , \w[5][11] , \w[5][10] , \w[5][9] , 
        \w[5][8] , \w[5][7] , \w[5][6] , \w[5][5] , \w[5][4] , \w[5][3] , 
        \w[5][2] , \w[5][1] , SYNOPSYS_UNCONNECTED__3}) );
  ADD_N32_123 \FAINST[5].ADD_  ( .A({\_8_net_[31] , \_8_net_[30] , 
        \_8_net_[29] , \_8_net_[28] , \_8_net_[27] , \_8_net_[26] , 
        \_8_net_[25] , \_8_net_[24] , \_8_net_[23] , \_8_net_[22] , 
        \_8_net_[21] , \_8_net_[20] , \_8_net_[19] , \_8_net_[18] , 
        \_8_net_[17] , \_8_net_[16] , \_8_net_[15] , \_8_net_[14] , 
        \_8_net_[13] , \_8_net_[12] , \_8_net_[11] , \_8_net_[10] , 
        \_8_net_[9] , \_8_net_[8] , \_8_net_[7] , \_8_net_[6] , \_8_net_[5] , 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[5][31] , \w[5][30] , \w[5][29] , 
        \w[5][28] , \w[5][27] , \w[5][26] , \w[5][25] , \w[5][24] , \w[5][23] , 
        \w[5][22] , \w[5][21] , \w[5][20] , \w[5][19] , \w[5][18] , \w[5][17] , 
        \w[5][16] , \w[5][15] , \w[5][14] , \w[5][13] , \w[5][12] , \w[5][11] , 
        \w[5][10] , \w[5][9] , \w[5][8] , \w[5][7] , \w[5][6] , \w[5][5] , 
        \w[5][4] , \w[5][3] , \w[5][2] , \w[5][1] , 1'b0}), .CI(1'b0), .S({
        \w[6][31] , \w[6][30] , \w[6][29] , \w[6][28] , \w[6][27] , \w[6][26] , 
        \w[6][25] , \w[6][24] , \w[6][23] , \w[6][22] , \w[6][21] , \w[6][20] , 
        \w[6][19] , \w[6][18] , \w[6][17] , \w[6][16] , \w[6][15] , \w[6][14] , 
        \w[6][13] , \w[6][12] , \w[6][11] , \w[6][10] , \w[6][9] , \w[6][8] , 
        \w[6][7] , \w[6][6] , \w[6][5] , \w[6][4] , \w[6][3] , \w[6][2] , 
        \w[6][1] , SYNOPSYS_UNCONNECTED__4}) );
  ADD_N32_122 \FAINST[6].ADD_  ( .A({\_10_net_[31] , \_10_net_[30] , 
        \_10_net_[29] , \_10_net_[28] , \_10_net_[27] , \_10_net_[26] , 
        \_10_net_[25] , \_10_net_[24] , \_10_net_[23] , \_10_net_[22] , 
        \_10_net_[21] , \_10_net_[20] , \_10_net_[19] , \_10_net_[18] , 
        \_10_net_[17] , \_10_net_[16] , \_10_net_[15] , \_10_net_[14] , 
        \_10_net_[13] , \_10_net_[12] , \_10_net_[11] , \_10_net_[10] , 
        \_10_net_[9] , \_10_net_[8] , \_10_net_[7] , \_10_net_[6] , 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[6][31] , \w[6][30] , \w[6][29] , 
        \w[6][28] , \w[6][27] , \w[6][26] , \w[6][25] , \w[6][24] , \w[6][23] , 
        \w[6][22] , \w[6][21] , \w[6][20] , \w[6][19] , \w[6][18] , \w[6][17] , 
        \w[6][16] , \w[6][15] , \w[6][14] , \w[6][13] , \w[6][12] , \w[6][11] , 
        \w[6][10] , \w[6][9] , \w[6][8] , \w[6][7] , \w[6][6] , \w[6][5] , 
        \w[6][4] , \w[6][3] , \w[6][2] , \w[6][1] , 1'b0}), .CI(1'b0), .S({
        \w[7][31] , \w[7][30] , \w[7][29] , \w[7][28] , \w[7][27] , \w[7][26] , 
        \w[7][25] , \w[7][24] , \w[7][23] , \w[7][22] , \w[7][21] , \w[7][20] , 
        \w[7][19] , \w[7][18] , \w[7][17] , \w[7][16] , \w[7][15] , \w[7][14] , 
        \w[7][13] , \w[7][12] , \w[7][11] , \w[7][10] , \w[7][9] , \w[7][8] , 
        \w[7][7] , \w[7][6] , \w[7][5] , \w[7][4] , \w[7][3] , \w[7][2] , 
        \w[7][1] , SYNOPSYS_UNCONNECTED__5}) );
  ADD_N32_121 \FAINST[7].ADD_  ( .A({\_12_net_[31] , \_12_net_[30] , 
        \_12_net_[29] , \_12_net_[28] , \_12_net_[27] , \_12_net_[26] , 
        \_12_net_[25] , \_12_net_[24] , \_12_net_[23] , \_12_net_[22] , 
        \_12_net_[21] , \_12_net_[20] , \_12_net_[19] , \_12_net_[18] , 
        \_12_net_[17] , \_12_net_[16] , \_12_net_[15] , \_12_net_[14] , 
        \_12_net_[13] , \_12_net_[12] , \_12_net_[11] , \_12_net_[10] , 
        \_12_net_[9] , \_12_net_[8] , \_12_net_[7] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({\w[7][31] , \w[7][30] , \w[7][29] , \w[7][28] , 
        \w[7][27] , \w[7][26] , \w[7][25] , \w[7][24] , \w[7][23] , \w[7][22] , 
        \w[7][21] , \w[7][20] , \w[7][19] , \w[7][18] , \w[7][17] , \w[7][16] , 
        \w[7][15] , \w[7][14] , \w[7][13] , \w[7][12] , \w[7][11] , \w[7][10] , 
        \w[7][9] , \w[7][8] , \w[7][7] , \w[7][6] , \w[7][5] , \w[7][4] , 
        \w[7][3] , \w[7][2] , \w[7][1] , 1'b0}), .CI(1'b0), .S({\w[8][31] , 
        \w[8][30] , \w[8][29] , \w[8][28] , \w[8][27] , \w[8][26] , \w[8][25] , 
        \w[8][24] , \w[8][23] , \w[8][22] , \w[8][21] , \w[8][20] , \w[8][19] , 
        \w[8][18] , \w[8][17] , \w[8][16] , \w[8][15] , \w[8][14] , \w[8][13] , 
        \w[8][12] , \w[8][11] , \w[8][10] , \w[8][9] , \w[8][8] , \w[8][7] , 
        \w[8][6] , \w[8][5] , \w[8][4] , \w[8][3] , \w[8][2] , \w[8][1] , 
        SYNOPSYS_UNCONNECTED__6}) );
  ADD_N32_120 \FAINST[8].ADD_  ( .A({\_14_net_[31] , \_14_net_[30] , 
        \_14_net_[29] , \_14_net_[28] , \_14_net_[27] , \_14_net_[26] , 
        \_14_net_[25] , \_14_net_[24] , \_14_net_[23] , \_14_net_[22] , 
        \_14_net_[21] , \_14_net_[20] , \_14_net_[19] , \_14_net_[18] , 
        \_14_net_[17] , \_14_net_[16] , \_14_net_[15] , \_14_net_[14] , 
        \_14_net_[13] , \_14_net_[12] , \_14_net_[11] , \_14_net_[10] , 
        \_14_net_[9] , \_14_net_[8] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({\w[8][31] , \w[8][30] , \w[8][29] , \w[8][28] , \w[8][27] , 
        \w[8][26] , \w[8][25] , \w[8][24] , \w[8][23] , \w[8][22] , \w[8][21] , 
        \w[8][20] , \w[8][19] , \w[8][18] , \w[8][17] , \w[8][16] , \w[8][15] , 
        \w[8][14] , \w[8][13] , \w[8][12] , \w[8][11] , \w[8][10] , \w[8][9] , 
        \w[8][8] , \w[8][7] , \w[8][6] , \w[8][5] , \w[8][4] , \w[8][3] , 
        \w[8][2] , \w[8][1] , 1'b0}), .CI(1'b0), .S({\w[9][31] , \w[9][30] , 
        \w[9][29] , \w[9][28] , \w[9][27] , \w[9][26] , \w[9][25] , \w[9][24] , 
        \w[9][23] , \w[9][22] , \w[9][21] , \w[9][20] , \w[9][19] , \w[9][18] , 
        \w[9][17] , \w[9][16] , \w[9][15] , \w[9][14] , \w[9][13] , \w[9][12] , 
        \w[9][11] , \w[9][10] , \w[9][9] , \w[9][8] , \w[9][7] , \w[9][6] , 
        \w[9][5] , \w[9][4] , \w[9][3] , \w[9][2] , \w[9][1] , 
        SYNOPSYS_UNCONNECTED__7}) );
  ADD_N32_119 \FAINST[9].ADD_  ( .A({\_16_net_[31] , \_16_net_[30] , 
        \_16_net_[29] , \_16_net_[28] , \_16_net_[27] , \_16_net_[26] , 
        \_16_net_[25] , \_16_net_[24] , \_16_net_[23] , \_16_net_[22] , 
        \_16_net_[21] , \_16_net_[20] , \_16_net_[19] , \_16_net_[18] , 
        \_16_net_[17] , \_16_net_[16] , \_16_net_[15] , \_16_net_[14] , 
        \_16_net_[13] , \_16_net_[12] , \_16_net_[11] , \_16_net_[10] , 
        \_16_net_[9] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({\w[9][31] , \w[9][30] , \w[9][29] , \w[9][28] , \w[9][27] , 
        \w[9][26] , \w[9][25] , \w[9][24] , \w[9][23] , \w[9][22] , \w[9][21] , 
        \w[9][20] , \w[9][19] , \w[9][18] , \w[9][17] , \w[9][16] , \w[9][15] , 
        \w[9][14] , \w[9][13] , \w[9][12] , \w[9][11] , \w[9][10] , \w[9][9] , 
        \w[9][8] , \w[9][7] , \w[9][6] , \w[9][5] , \w[9][4] , \w[9][3] , 
        \w[9][2] , \w[9][1] , 1'b0}), .CI(1'b0), .S({\w[10][31] , \w[10][30] , 
        \w[10][29] , \w[10][28] , \w[10][27] , \w[10][26] , \w[10][25] , 
        \w[10][24] , \w[10][23] , \w[10][22] , \w[10][21] , \w[10][20] , 
        \w[10][19] , \w[10][18] , \w[10][17] , \w[10][16] , \w[10][15] , 
        \w[10][14] , \w[10][13] , \w[10][12] , \w[10][11] , \w[10][10] , 
        \w[10][9] , \w[10][8] , \w[10][7] , \w[10][6] , \w[10][5] , \w[10][4] , 
        \w[10][3] , \w[10][2] , \w[10][1] , SYNOPSYS_UNCONNECTED__8}) );
  ADD_N32_118 \FAINST[10].ADD_  ( .A({\_18_net_[31] , \_18_net_[30] , 
        \_18_net_[29] , \_18_net_[28] , \_18_net_[27] , \_18_net_[26] , 
        \_18_net_[25] , \_18_net_[24] , \_18_net_[23] , \_18_net_[22] , 
        \_18_net_[21] , \_18_net_[20] , \_18_net_[19] , \_18_net_[18] , 
        \_18_net_[17] , \_18_net_[16] , \_18_net_[15] , \_18_net_[14] , 
        \_18_net_[13] , \_18_net_[12] , \_18_net_[11] , \_18_net_[10] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[10][31] , \w[10][30] , \w[10][29] , \w[10][28] , \w[10][27] , 
        \w[10][26] , \w[10][25] , \w[10][24] , \w[10][23] , \w[10][22] , 
        \w[10][21] , \w[10][20] , \w[10][19] , \w[10][18] , \w[10][17] , 
        \w[10][16] , \w[10][15] , \w[10][14] , \w[10][13] , \w[10][12] , 
        \w[10][11] , \w[10][10] , \w[10][9] , \w[10][8] , \w[10][7] , 
        \w[10][6] , \w[10][5] , \w[10][4] , \w[10][3] , \w[10][2] , \w[10][1] , 
        1'b0}), .CI(1'b0), .S({\w[11][31] , \w[11][30] , \w[11][29] , 
        \w[11][28] , \w[11][27] , \w[11][26] , \w[11][25] , \w[11][24] , 
        \w[11][23] , \w[11][22] , \w[11][21] , \w[11][20] , \w[11][19] , 
        \w[11][18] , \w[11][17] , \w[11][16] , \w[11][15] , \w[11][14] , 
        \w[11][13] , \w[11][12] , \w[11][11] , \w[11][10] , \w[11][9] , 
        \w[11][8] , \w[11][7] , \w[11][6] , \w[11][5] , \w[11][4] , \w[11][3] , 
        \w[11][2] , \w[11][1] , SYNOPSYS_UNCONNECTED__9}) );
  ADD_N32_117 \FAINST[11].ADD_  ( .A({\_20_net_[31] , \_20_net_[30] , 
        \_20_net_[29] , \_20_net_[28] , \_20_net_[27] , \_20_net_[26] , 
        \_20_net_[25] , \_20_net_[24] , \_20_net_[23] , \_20_net_[22] , 
        \_20_net_[21] , \_20_net_[20] , \_20_net_[19] , \_20_net_[18] , 
        \_20_net_[17] , \_20_net_[16] , \_20_net_[15] , \_20_net_[14] , 
        \_20_net_[13] , \_20_net_[12] , \_20_net_[11] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[11][31] , 
        \w[11][30] , \w[11][29] , \w[11][28] , \w[11][27] , \w[11][26] , 
        \w[11][25] , \w[11][24] , \w[11][23] , \w[11][22] , \w[11][21] , 
        \w[11][20] , \w[11][19] , \w[11][18] , \w[11][17] , \w[11][16] , 
        \w[11][15] , \w[11][14] , \w[11][13] , \w[11][12] , \w[11][11] , 
        \w[11][10] , \w[11][9] , \w[11][8] , \w[11][7] , \w[11][6] , 
        \w[11][5] , \w[11][4] , \w[11][3] , \w[11][2] , \w[11][1] , 1'b0}), 
        .CI(1'b0), .S({\w[12][31] , \w[12][30] , \w[12][29] , \w[12][28] , 
        \w[12][27] , \w[12][26] , \w[12][25] , \w[12][24] , \w[12][23] , 
        \w[12][22] , \w[12][21] , \w[12][20] , \w[12][19] , \w[12][18] , 
        \w[12][17] , \w[12][16] , \w[12][15] , \w[12][14] , \w[12][13] , 
        \w[12][12] , \w[12][11] , \w[12][10] , \w[12][9] , \w[12][8] , 
        \w[12][7] , \w[12][6] , \w[12][5] , \w[12][4] , \w[12][3] , \w[12][2] , 
        \w[12][1] , SYNOPSYS_UNCONNECTED__10}) );
  ADD_N32_116 \FAINST[12].ADD_  ( .A({\_22_net_[31] , \_22_net_[30] , 
        \_22_net_[29] , \_22_net_[28] , \_22_net_[27] , \_22_net_[26] , 
        \_22_net_[25] , \_22_net_[24] , \_22_net_[23] , \_22_net_[22] , 
        \_22_net_[21] , \_22_net_[20] , \_22_net_[19] , \_22_net_[18] , 
        \_22_net_[17] , \_22_net_[16] , \_22_net_[15] , \_22_net_[14] , 
        \_22_net_[13] , \_22_net_[12] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[12][31] , \w[12][30] , 
        \w[12][29] , \w[12][28] , \w[12][27] , \w[12][26] , \w[12][25] , 
        \w[12][24] , \w[12][23] , \w[12][22] , \w[12][21] , \w[12][20] , 
        \w[12][19] , \w[12][18] , \w[12][17] , \w[12][16] , \w[12][15] , 
        \w[12][14] , \w[12][13] , \w[12][12] , \w[12][11] , \w[12][10] , 
        \w[12][9] , \w[12][8] , \w[12][7] , \w[12][6] , \w[12][5] , \w[12][4] , 
        \w[12][3] , \w[12][2] , \w[12][1] , 1'b0}), .CI(1'b0), .S({\w[13][31] , 
        \w[13][30] , \w[13][29] , \w[13][28] , \w[13][27] , \w[13][26] , 
        \w[13][25] , \w[13][24] , \w[13][23] , \w[13][22] , \w[13][21] , 
        \w[13][20] , \w[13][19] , \w[13][18] , \w[13][17] , \w[13][16] , 
        \w[13][15] , \w[13][14] , \w[13][13] , \w[13][12] , \w[13][11] , 
        \w[13][10] , \w[13][9] , \w[13][8] , \w[13][7] , \w[13][6] , 
        \w[13][5] , \w[13][4] , \w[13][3] , \w[13][2] , \w[13][1] , 
        SYNOPSYS_UNCONNECTED__11}) );
  ADD_N32_115 \FAINST[13].ADD_  ( .A({\_24_net_[31] , \_24_net_[30] , 
        \_24_net_[29] , \_24_net_[28] , \_24_net_[27] , \_24_net_[26] , 
        \_24_net_[25] , \_24_net_[24] , \_24_net_[23] , \_24_net_[22] , 
        \_24_net_[21] , \_24_net_[20] , \_24_net_[19] , \_24_net_[18] , 
        \_24_net_[17] , \_24_net_[16] , \_24_net_[15] , \_24_net_[14] , 
        \_24_net_[13] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[13][31] , \w[13][30] , \w[13][29] , 
        \w[13][28] , \w[13][27] , \w[13][26] , \w[13][25] , \w[13][24] , 
        \w[13][23] , \w[13][22] , \w[13][21] , \w[13][20] , \w[13][19] , 
        \w[13][18] , \w[13][17] , \w[13][16] , \w[13][15] , \w[13][14] , 
        \w[13][13] , \w[13][12] , \w[13][11] , \w[13][10] , \w[13][9] , 
        \w[13][8] , \w[13][7] , \w[13][6] , \w[13][5] , \w[13][4] , \w[13][3] , 
        \w[13][2] , \w[13][1] , 1'b0}), .CI(1'b0), .S({\w[14][31] , 
        \w[14][30] , \w[14][29] , \w[14][28] , \w[14][27] , \w[14][26] , 
        \w[14][25] , \w[14][24] , \w[14][23] , \w[14][22] , \w[14][21] , 
        \w[14][20] , \w[14][19] , \w[14][18] , \w[14][17] , \w[14][16] , 
        \w[14][15] , \w[14][14] , \w[14][13] , \w[14][12] , \w[14][11] , 
        \w[14][10] , \w[14][9] , \w[14][8] , \w[14][7] , \w[14][6] , 
        \w[14][5] , \w[14][4] , \w[14][3] , \w[14][2] , \w[14][1] , 
        SYNOPSYS_UNCONNECTED__12}) );
  ADD_N32_114 \FAINST[14].ADD_  ( .A({\_26_net_[31] , \_26_net_[30] , 
        \_26_net_[29] , \_26_net_[28] , \_26_net_[27] , \_26_net_[26] , 
        \_26_net_[25] , \_26_net_[24] , \_26_net_[23] , \_26_net_[22] , 
        \_26_net_[21] , \_26_net_[20] , \_26_net_[19] , \_26_net_[18] , 
        \_26_net_[17] , \_26_net_[16] , \_26_net_[15] , \_26_net_[14] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({\w[14][31] , \w[14][30] , \w[14][29] , \w[14][28] , 
        \w[14][27] , \w[14][26] , \w[14][25] , \w[14][24] , \w[14][23] , 
        \w[14][22] , \w[14][21] , \w[14][20] , \w[14][19] , \w[14][18] , 
        \w[14][17] , \w[14][16] , \w[14][15] , \w[14][14] , \w[14][13] , 
        \w[14][12] , \w[14][11] , \w[14][10] , \w[14][9] , \w[14][8] , 
        \w[14][7] , \w[14][6] , \w[14][5] , \w[14][4] , \w[14][3] , \w[14][2] , 
        \w[14][1] , 1'b0}), .CI(1'b0), .S({\w[15][31] , \w[15][30] , 
        \w[15][29] , \w[15][28] , \w[15][27] , \w[15][26] , \w[15][25] , 
        \w[15][24] , \w[15][23] , \w[15][22] , \w[15][21] , \w[15][20] , 
        \w[15][19] , \w[15][18] , \w[15][17] , \w[15][16] , \w[15][15] , 
        \w[15][14] , \w[15][13] , \w[15][12] , \w[15][11] , \w[15][10] , 
        \w[15][9] , \w[15][8] , \w[15][7] , \w[15][6] , \w[15][5] , \w[15][4] , 
        \w[15][3] , \w[15][2] , \w[15][1] , SYNOPSYS_UNCONNECTED__13}) );
  ADD_N32_113 \FAINST[15].ADD_  ( .A({\_28_net_[31] , \_28_net_[30] , 
        \_28_net_[29] , \_28_net_[28] , \_28_net_[27] , \_28_net_[26] , 
        \_28_net_[25] , \_28_net_[24] , \_28_net_[23] , \_28_net_[22] , 
        \_28_net_[21] , \_28_net_[20] , \_28_net_[19] , \_28_net_[18] , 
        \_28_net_[17] , \_28_net_[16] , \_28_net_[15] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({\w[15][31] , \w[15][30] , \w[15][29] , \w[15][28] , \w[15][27] , 
        \w[15][26] , \w[15][25] , \w[15][24] , \w[15][23] , \w[15][22] , 
        \w[15][21] , \w[15][20] , \w[15][19] , \w[15][18] , \w[15][17] , 
        \w[15][16] , \w[15][15] , \w[15][14] , \w[15][13] , \w[15][12] , 
        \w[15][11] , \w[15][10] , \w[15][9] , \w[15][8] , \w[15][7] , 
        \w[15][6] , \w[15][5] , \w[15][4] , \w[15][3] , \w[15][2] , \w[15][1] , 
        1'b0}), .CI(1'b0), .S({\w[16][31] , \w[16][30] , \w[16][29] , 
        \w[16][28] , \w[16][27] , \w[16][26] , \w[16][25] , \w[16][24] , 
        \w[16][23] , \w[16][22] , \w[16][21] , \w[16][20] , \w[16][19] , 
        \w[16][18] , \w[16][17] , \w[16][16] , \w[16][15] , \w[16][14] , 
        \w[16][13] , \w[16][12] , \w[16][11] , \w[16][10] , \w[16][9] , 
        \w[16][8] , \w[16][7] , \w[16][6] , \w[16][5] , \w[16][4] , \w[16][3] , 
        \w[16][2] , \w[16][1] , SYNOPSYS_UNCONNECTED__14}) );
  ADD_N32_112 \FAINST[16].ADD_  ( .A({\_30_net_[31] , \_30_net_[30] , 
        \_30_net_[29] , \_30_net_[28] , \_30_net_[27] , \_30_net_[26] , 
        \_30_net_[25] , \_30_net_[24] , \_30_net_[23] , \_30_net_[22] , 
        \_30_net_[21] , \_30_net_[20] , \_30_net_[19] , \_30_net_[18] , 
        \_30_net_[17] , \_30_net_[16] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[16][31] , \w[16][30] , \w[16][29] , \w[16][28] , \w[16][27] , 
        \w[16][26] , \w[16][25] , \w[16][24] , \w[16][23] , \w[16][22] , 
        \w[16][21] , \w[16][20] , \w[16][19] , \w[16][18] , \w[16][17] , 
        \w[16][16] , \w[16][15] , \w[16][14] , \w[16][13] , \w[16][12] , 
        \w[16][11] , \w[16][10] , \w[16][9] , \w[16][8] , \w[16][7] , 
        \w[16][6] , \w[16][5] , \w[16][4] , \w[16][3] , \w[16][2] , \w[16][1] , 
        1'b0}), .CI(1'b0), .S({\w[17][31] , \w[17][30] , \w[17][29] , 
        \w[17][28] , \w[17][27] , \w[17][26] , \w[17][25] , \w[17][24] , 
        \w[17][23] , \w[17][22] , \w[17][21] , \w[17][20] , \w[17][19] , 
        \w[17][18] , \w[17][17] , \w[17][16] , \w[17][15] , \w[17][14] , 
        \w[17][13] , \w[17][12] , \w[17][11] , \w[17][10] , \w[17][9] , 
        \w[17][8] , \w[17][7] , \w[17][6] , \w[17][5] , \w[17][4] , \w[17][3] , 
        \w[17][2] , \w[17][1] , SYNOPSYS_UNCONNECTED__15}) );
  ADD_N32_111 \FAINST[17].ADD_  ( .A({\_32_net_[31] , \_32_net_[30] , 
        \_32_net_[29] , \_32_net_[28] , \_32_net_[27] , \_32_net_[26] , 
        \_32_net_[25] , \_32_net_[24] , \_32_net_[23] , \_32_net_[22] , 
        \_32_net_[21] , \_32_net_[20] , \_32_net_[19] , \_32_net_[18] , 
        \_32_net_[17] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[17][31] , 
        \w[17][30] , \w[17][29] , \w[17][28] , \w[17][27] , \w[17][26] , 
        \w[17][25] , \w[17][24] , \w[17][23] , \w[17][22] , \w[17][21] , 
        \w[17][20] , \w[17][19] , \w[17][18] , \w[17][17] , \w[17][16] , 
        \w[17][15] , \w[17][14] , \w[17][13] , \w[17][12] , \w[17][11] , 
        \w[17][10] , \w[17][9] , \w[17][8] , \w[17][7] , \w[17][6] , 
        \w[17][5] , \w[17][4] , \w[17][3] , \w[17][2] , \w[17][1] , 1'b0}), 
        .CI(1'b0), .S({\w[18][31] , \w[18][30] , \w[18][29] , \w[18][28] , 
        \w[18][27] , \w[18][26] , \w[18][25] , \w[18][24] , \w[18][23] , 
        \w[18][22] , \w[18][21] , \w[18][20] , \w[18][19] , \w[18][18] , 
        \w[18][17] , \w[18][16] , \w[18][15] , \w[18][14] , \w[18][13] , 
        \w[18][12] , \w[18][11] , \w[18][10] , \w[18][9] , \w[18][8] , 
        \w[18][7] , \w[18][6] , \w[18][5] , \w[18][4] , \w[18][3] , \w[18][2] , 
        \w[18][1] , SYNOPSYS_UNCONNECTED__16}) );
  ADD_N32_110 \FAINST[18].ADD_  ( .A({\_34_net_[31] , \_34_net_[30] , 
        \_34_net_[29] , \_34_net_[28] , \_34_net_[27] , \_34_net_[26] , 
        \_34_net_[25] , \_34_net_[24] , \_34_net_[23] , \_34_net_[22] , 
        \_34_net_[21] , \_34_net_[20] , \_34_net_[19] , \_34_net_[18] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[18][31] , \w[18][30] , 
        \w[18][29] , \w[18][28] , \w[18][27] , \w[18][26] , \w[18][25] , 
        \w[18][24] , \w[18][23] , \w[18][22] , \w[18][21] , \w[18][20] , 
        \w[18][19] , \w[18][18] , \w[18][17] , \w[18][16] , \w[18][15] , 
        \w[18][14] , \w[18][13] , \w[18][12] , \w[18][11] , \w[18][10] , 
        \w[18][9] , \w[18][8] , \w[18][7] , \w[18][6] , \w[18][5] , \w[18][4] , 
        \w[18][3] , \w[18][2] , \w[18][1] , 1'b0}), .CI(1'b0), .S({\w[19][31] , 
        \w[19][30] , \w[19][29] , \w[19][28] , \w[19][27] , \w[19][26] , 
        \w[19][25] , \w[19][24] , \w[19][23] , \w[19][22] , \w[19][21] , 
        \w[19][20] , \w[19][19] , \w[19][18] , \w[19][17] , \w[19][16] , 
        \w[19][15] , \w[19][14] , \w[19][13] , \w[19][12] , \w[19][11] , 
        \w[19][10] , \w[19][9] , \w[19][8] , \w[19][7] , \w[19][6] , 
        \w[19][5] , \w[19][4] , \w[19][3] , \w[19][2] , \w[19][1] , 
        SYNOPSYS_UNCONNECTED__17}) );
  ADD_N32_109 \FAINST[19].ADD_  ( .A({\_36_net_[31] , \_36_net_[30] , 
        \_36_net_[29] , \_36_net_[28] , \_36_net_[27] , \_36_net_[26] , 
        \_36_net_[25] , \_36_net_[24] , \_36_net_[23] , \_36_net_[22] , 
        \_36_net_[21] , \_36_net_[20] , \_36_net_[19] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({\w[19][31] , \w[19][30] , \w[19][29] , 
        \w[19][28] , \w[19][27] , \w[19][26] , \w[19][25] , \w[19][24] , 
        \w[19][23] , \w[19][22] , \w[19][21] , \w[19][20] , \w[19][19] , 
        \w[19][18] , \w[19][17] , \w[19][16] , \w[19][15] , \w[19][14] , 
        \w[19][13] , \w[19][12] , \w[19][11] , \w[19][10] , \w[19][9] , 
        \w[19][8] , \w[19][7] , \w[19][6] , \w[19][5] , \w[19][4] , \w[19][3] , 
        \w[19][2] , \w[19][1] , 1'b0}), .CI(1'b0), .S({\w[20][31] , 
        \w[20][30] , \w[20][29] , \w[20][28] , \w[20][27] , \w[20][26] , 
        \w[20][25] , \w[20][24] , \w[20][23] , \w[20][22] , \w[20][21] , 
        \w[20][20] , \w[20][19] , \w[20][18] , \w[20][17] , \w[20][16] , 
        \w[20][15] , \w[20][14] , \w[20][13] , \w[20][12] , \w[20][11] , 
        \w[20][10] , \w[20][9] , \w[20][8] , \w[20][7] , \w[20][6] , 
        \w[20][5] , \w[20][4] , \w[20][3] , \w[20][2] , \w[20][1] , 
        SYNOPSYS_UNCONNECTED__18}) );
  ADD_N32_108 \FAINST[20].ADD_  ( .A({\_38_net_[31] , \_38_net_[30] , 
        \_38_net_[29] , \_38_net_[28] , \_38_net_[27] , \_38_net_[26] , 
        \_38_net_[25] , \_38_net_[24] , \_38_net_[23] , \_38_net_[22] , 
        \_38_net_[21] , \_38_net_[20] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .B({\w[20][31] , \w[20][30] , \w[20][29] , \w[20][28] , 
        \w[20][27] , \w[20][26] , \w[20][25] , \w[20][24] , \w[20][23] , 
        \w[20][22] , \w[20][21] , \w[20][20] , \w[20][19] , \w[20][18] , 
        \w[20][17] , \w[20][16] , \w[20][15] , \w[20][14] , \w[20][13] , 
        \w[20][12] , \w[20][11] , \w[20][10] , \w[20][9] , \w[20][8] , 
        \w[20][7] , \w[20][6] , \w[20][5] , \w[20][4] , \w[20][3] , \w[20][2] , 
        \w[20][1] , 1'b0}), .CI(1'b0), .S({\w[21][31] , \w[21][30] , 
        \w[21][29] , \w[21][28] , \w[21][27] , \w[21][26] , \w[21][25] , 
        \w[21][24] , \w[21][23] , \w[21][22] , \w[21][21] , \w[21][20] , 
        \w[21][19] , \w[21][18] , \w[21][17] , \w[21][16] , \w[21][15] , 
        \w[21][14] , \w[21][13] , \w[21][12] , \w[21][11] , \w[21][10] , 
        \w[21][9] , \w[21][8] , \w[21][7] , \w[21][6] , \w[21][5] , \w[21][4] , 
        \w[21][3] , \w[21][2] , \w[21][1] , SYNOPSYS_UNCONNECTED__19}) );
  ADD_N32_107 \FAINST[21].ADD_  ( .A({\_40_net_[31] , \_40_net_[30] , 
        \_40_net_[29] , \_40_net_[28] , \_40_net_[27] , \_40_net_[26] , 
        \_40_net_[25] , \_40_net_[24] , \_40_net_[23] , \_40_net_[22] , 
        \_40_net_[21] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[21][31] , \w[21][30] , \w[21][29] , \w[21][28] , \w[21][27] , 
        \w[21][26] , \w[21][25] , \w[21][24] , \w[21][23] , \w[21][22] , 
        \w[21][21] , \w[21][20] , \w[21][19] , \w[21][18] , \w[21][17] , 
        \w[21][16] , \w[21][15] , \w[21][14] , \w[21][13] , \w[21][12] , 
        \w[21][11] , \w[21][10] , \w[21][9] , \w[21][8] , \w[21][7] , 
        \w[21][6] , \w[21][5] , \w[21][4] , \w[21][3] , \w[21][2] , \w[21][1] , 
        1'b0}), .CI(1'b0), .S({\w[22][31] , \w[22][30] , \w[22][29] , 
        \w[22][28] , \w[22][27] , \w[22][26] , \w[22][25] , \w[22][24] , 
        \w[22][23] , \w[22][22] , \w[22][21] , \w[22][20] , \w[22][19] , 
        \w[22][18] , \w[22][17] , \w[22][16] , \w[22][15] , \w[22][14] , 
        \w[22][13] , \w[22][12] , \w[22][11] , \w[22][10] , \w[22][9] , 
        \w[22][8] , \w[22][7] , \w[22][6] , \w[22][5] , \w[22][4] , \w[22][3] , 
        \w[22][2] , \w[22][1] , SYNOPSYS_UNCONNECTED__20}) );
  ADD_N32_106 \FAINST[22].ADD_  ( .A({\_42_net_[31] , \_42_net_[30] , 
        \_42_net_[29] , \_42_net_[28] , \_42_net_[27] , \_42_net_[26] , 
        \_42_net_[25] , \_42_net_[24] , \_42_net_[23] , \_42_net_[22] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[22][31] , \w[22][30] , \w[22][29] , \w[22][28] , \w[22][27] , 
        \w[22][26] , \w[22][25] , \w[22][24] , \w[22][23] , \w[22][22] , 
        \w[22][21] , \w[22][20] , \w[22][19] , \w[22][18] , \w[22][17] , 
        \w[22][16] , \w[22][15] , \w[22][14] , \w[22][13] , \w[22][12] , 
        \w[22][11] , \w[22][10] , \w[22][9] , \w[22][8] , \w[22][7] , 
        \w[22][6] , \w[22][5] , \w[22][4] , \w[22][3] , \w[22][2] , \w[22][1] , 
        1'b0}), .CI(1'b0), .S({\w[23][31] , \w[23][30] , \w[23][29] , 
        \w[23][28] , \w[23][27] , \w[23][26] , \w[23][25] , \w[23][24] , 
        \w[23][23] , \w[23][22] , \w[23][21] , \w[23][20] , \w[23][19] , 
        \w[23][18] , \w[23][17] , \w[23][16] , \w[23][15] , \w[23][14] , 
        \w[23][13] , \w[23][12] , \w[23][11] , \w[23][10] , \w[23][9] , 
        \w[23][8] , \w[23][7] , \w[23][6] , \w[23][5] , \w[23][4] , \w[23][3] , 
        \w[23][2] , \w[23][1] , SYNOPSYS_UNCONNECTED__21}) );
  ADD_N32_105 \FAINST[23].ADD_  ( .A({\_44_net_[31] , \_44_net_[30] , 
        \_44_net_[29] , \_44_net_[28] , \_44_net_[27] , \_44_net_[26] , 
        \_44_net_[25] , \_44_net_[24] , \_44_net_[23] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[23][31] , 
        \w[23][30] , \w[23][29] , \w[23][28] , \w[23][27] , \w[23][26] , 
        \w[23][25] , \w[23][24] , \w[23][23] , \w[23][22] , \w[23][21] , 
        \w[23][20] , \w[23][19] , \w[23][18] , \w[23][17] , \w[23][16] , 
        \w[23][15] , \w[23][14] , \w[23][13] , \w[23][12] , \w[23][11] , 
        \w[23][10] , \w[23][9] , \w[23][8] , \w[23][7] , \w[23][6] , 
        \w[23][5] , \w[23][4] , \w[23][3] , \w[23][2] , \w[23][1] , 1'b0}), 
        .CI(1'b0), .S({\w[24][31] , \w[24][30] , \w[24][29] , \w[24][28] , 
        \w[24][27] , \w[24][26] , \w[24][25] , \w[24][24] , \w[24][23] , 
        \w[24][22] , \w[24][21] , \w[24][20] , \w[24][19] , \w[24][18] , 
        \w[24][17] , \w[24][16] , \w[24][15] , \w[24][14] , \w[24][13] , 
        \w[24][12] , \w[24][11] , \w[24][10] , \w[24][9] , \w[24][8] , 
        \w[24][7] , \w[24][6] , \w[24][5] , \w[24][4] , \w[24][3] , \w[24][2] , 
        \w[24][1] , SYNOPSYS_UNCONNECTED__22}) );
  ADD_N32_104 \FAINST[24].ADD_  ( .A({\_46_net_[31] , \_46_net_[30] , 
        \_46_net_[29] , \_46_net_[28] , \_46_net_[27] , \_46_net_[26] , 
        \_46_net_[25] , \_46_net_[24] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[24][31] , \w[24][30] , 
        \w[24][29] , \w[24][28] , \w[24][27] , \w[24][26] , \w[24][25] , 
        \w[24][24] , \w[24][23] , \w[24][22] , \w[24][21] , \w[24][20] , 
        \w[24][19] , \w[24][18] , \w[24][17] , \w[24][16] , \w[24][15] , 
        \w[24][14] , \w[24][13] , \w[24][12] , \w[24][11] , \w[24][10] , 
        \w[24][9] , \w[24][8] , \w[24][7] , \w[24][6] , \w[24][5] , \w[24][4] , 
        \w[24][3] , \w[24][2] , \w[24][1] , 1'b0}), .CI(1'b0), .S({\w[25][31] , 
        \w[25][30] , \w[25][29] , \w[25][28] , \w[25][27] , \w[25][26] , 
        \w[25][25] , \w[25][24] , \w[25][23] , \w[25][22] , \w[25][21] , 
        \w[25][20] , \w[25][19] , \w[25][18] , \w[25][17] , \w[25][16] , 
        \w[25][15] , \w[25][14] , \w[25][13] , \w[25][12] , \w[25][11] , 
        \w[25][10] , \w[25][9] , \w[25][8] , \w[25][7] , \w[25][6] , 
        \w[25][5] , \w[25][4] , \w[25][3] , \w[25][2] , \w[25][1] , 
        SYNOPSYS_UNCONNECTED__23}) );
  ADD_N32_103 \FAINST[25].ADD_  ( .A({\_48_net_[31] , \_48_net_[30] , 
        \_48_net_[29] , \_48_net_[28] , \_48_net_[27] , \_48_net_[26] , 
        \_48_net_[25] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[25][31] , \w[25][30] , \w[25][29] , 
        \w[25][28] , \w[25][27] , \w[25][26] , \w[25][25] , \w[25][24] , 
        \w[25][23] , \w[25][22] , \w[25][21] , \w[25][20] , \w[25][19] , 
        \w[25][18] , \w[25][17] , \w[25][16] , \w[25][15] , \w[25][14] , 
        \w[25][13] , \w[25][12] , \w[25][11] , \w[25][10] , \w[25][9] , 
        \w[25][8] , \w[25][7] , \w[25][6] , \w[25][5] , \w[25][4] , \w[25][3] , 
        \w[25][2] , \w[25][1] , 1'b0}), .CI(1'b0), .S({\w[26][31] , 
        \w[26][30] , \w[26][29] , \w[26][28] , \w[26][27] , \w[26][26] , 
        \w[26][25] , \w[26][24] , \w[26][23] , \w[26][22] , \w[26][21] , 
        \w[26][20] , \w[26][19] , \w[26][18] , \w[26][17] , \w[26][16] , 
        \w[26][15] , \w[26][14] , \w[26][13] , \w[26][12] , \w[26][11] , 
        \w[26][10] , \w[26][9] , \w[26][8] , \w[26][7] , \w[26][6] , 
        \w[26][5] , \w[26][4] , \w[26][3] , \w[26][2] , \w[26][1] , 
        SYNOPSYS_UNCONNECTED__24}) );
  ADD_N32_102 \FAINST[26].ADD_  ( .A({\_50_net_[31] , \_50_net_[30] , 
        \_50_net_[29] , \_50_net_[28] , \_50_net_[27] , \_50_net_[26] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({\w[26][31] , \w[26][30] , \w[26][29] , \w[26][28] , 
        \w[26][27] , \w[26][26] , \w[26][25] , \w[26][24] , \w[26][23] , 
        \w[26][22] , \w[26][21] , \w[26][20] , \w[26][19] , \w[26][18] , 
        \w[26][17] , \w[26][16] , \w[26][15] , \w[26][14] , \w[26][13] , 
        \w[26][12] , \w[26][11] , \w[26][10] , \w[26][9] , \w[26][8] , 
        \w[26][7] , \w[26][6] , \w[26][5] , \w[26][4] , \w[26][3] , \w[26][2] , 
        \w[26][1] , 1'b0}), .CI(1'b0), .S({\w[27][31] , \w[27][30] , 
        \w[27][29] , \w[27][28] , \w[27][27] , \w[27][26] , \w[27][25] , 
        \w[27][24] , \w[27][23] , \w[27][22] , \w[27][21] , \w[27][20] , 
        \w[27][19] , \w[27][18] , \w[27][17] , \w[27][16] , \w[27][15] , 
        \w[27][14] , \w[27][13] , \w[27][12] , \w[27][11] , \w[27][10] , 
        \w[27][9] , \w[27][8] , \w[27][7] , \w[27][6] , \w[27][5] , \w[27][4] , 
        \w[27][3] , \w[27][2] , \w[27][1] , SYNOPSYS_UNCONNECTED__25}) );
  ADD_N32_101 \FAINST[27].ADD_  ( .A({\_52_net_[31] , \_52_net_[30] , 
        \_52_net_[29] , \_52_net_[28] , \_52_net_[27] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({\w[27][31] , \w[27][30] , \w[27][29] , \w[27][28] , \w[27][27] , 
        \w[27][26] , \w[27][25] , \w[27][24] , \w[27][23] , \w[27][22] , 
        \w[27][21] , \w[27][20] , \w[27][19] , \w[27][18] , \w[27][17] , 
        \w[27][16] , \w[27][15] , \w[27][14] , \w[27][13] , \w[27][12] , 
        \w[27][11] , \w[27][10] , \w[27][9] , \w[27][8] , \w[27][7] , 
        \w[27][6] , \w[27][5] , \w[27][4] , \w[27][3] , \w[27][2] , \w[27][1] , 
        1'b0}), .CI(1'b0), .S({\w[28][31] , \w[28][30] , \w[28][29] , 
        \w[28][28] , \w[28][27] , \w[28][26] , \w[28][25] , \w[28][24] , 
        \w[28][23] , \w[28][22] , \w[28][21] , \w[28][20] , \w[28][19] , 
        \w[28][18] , \w[28][17] , \w[28][16] , \w[28][15] , \w[28][14] , 
        \w[28][13] , \w[28][12] , \w[28][11] , \w[28][10] , \w[28][9] , 
        \w[28][8] , \w[28][7] , \w[28][6] , \w[28][5] , \w[28][4] , \w[28][3] , 
        \w[28][2] , \w[28][1] , SYNOPSYS_UNCONNECTED__26}) );
  ADD_N32_100 \FAINST[28].ADD_  ( .A({\_54_net_[31] , \_54_net_[30] , 
        \_54_net_[29] , \_54_net_[28] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[28][31] , \w[28][30] , \w[28][29] , \w[28][28] , \w[28][27] , 
        \w[28][26] , \w[28][25] , \w[28][24] , \w[28][23] , \w[28][22] , 
        \w[28][21] , \w[28][20] , \w[28][19] , \w[28][18] , \w[28][17] , 
        \w[28][16] , \w[28][15] , \w[28][14] , \w[28][13] , \w[28][12] , 
        \w[28][11] , \w[28][10] , \w[28][9] , \w[28][8] , \w[28][7] , 
        \w[28][6] , \w[28][5] , \w[28][4] , \w[28][3] , \w[28][2] , \w[28][1] , 
        1'b0}), .CI(1'b0), .S({\w[29][31] , \w[29][30] , \w[29][29] , 
        \w[29][28] , \w[29][27] , \w[29][26] , \w[29][25] , \w[29][24] , 
        \w[29][23] , \w[29][22] , \w[29][21] , \w[29][20] , \w[29][19] , 
        \w[29][18] , \w[29][17] , \w[29][16] , \w[29][15] , \w[29][14] , 
        \w[29][13] , \w[29][12] , \w[29][11] , \w[29][10] , \w[29][9] , 
        \w[29][8] , \w[29][7] , \w[29][6] , \w[29][5] , \w[29][4] , \w[29][3] , 
        \w[29][2] , \w[29][1] , SYNOPSYS_UNCONNECTED__27}) );
  ADD_N32_99 \FAINST[29].ADD_  ( .A({\_56_net_[31] , \_56_net_[30] , 
        \_56_net_[29] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[29][31] , 
        \w[29][30] , \w[29][29] , \w[29][28] , \w[29][27] , \w[29][26] , 
        \w[29][25] , \w[29][24] , \w[29][23] , \w[29][22] , \w[29][21] , 
        \w[29][20] , \w[29][19] , \w[29][18] , \w[29][17] , \w[29][16] , 
        \w[29][15] , \w[29][14] , \w[29][13] , \w[29][12] , \w[29][11] , 
        \w[29][10] , \w[29][9] , \w[29][8] , \w[29][7] , \w[29][6] , 
        \w[29][5] , \w[29][4] , \w[29][3] , \w[29][2] , \w[29][1] , 1'b0}), 
        .CI(1'b0), .S({\w[30][31] , \w[30][30] , \w[30][29] , \w[30][28] , 
        \w[30][27] , \w[30][26] , \w[30][25] , \w[30][24] , \w[30][23] , 
        \w[30][22] , \w[30][21] , \w[30][20] , \w[30][19] , \w[30][18] , 
        \w[30][17] , \w[30][16] , \w[30][15] , \w[30][14] , \w[30][13] , 
        \w[30][12] , \w[30][11] , \w[30][10] , \w[30][9] , \w[30][8] , 
        \w[30][7] , \w[30][6] , \w[30][5] , \w[30][4] , \w[30][3] , \w[30][2] , 
        \w[30][1] , SYNOPSYS_UNCONNECTED__28}) );
  ADD_N32_98 \FAINST[30].ADD_  ( .A({\_58_net_[31] , \_58_net_[30] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[30][31] , \w[30][30] , 
        \w[30][29] , \w[30][28] , \w[30][27] , \w[30][26] , \w[30][25] , 
        \w[30][24] , \w[30][23] , \w[30][22] , \w[30][21] , \w[30][20] , 
        \w[30][19] , \w[30][18] , \w[30][17] , \w[30][16] , \w[30][15] , 
        \w[30][14] , \w[30][13] , \w[30][12] , \w[30][11] , \w[30][10] , 
        \w[30][9] , \w[30][8] , \w[30][7] , \w[30][6] , \w[30][5] , \w[30][4] , 
        \w[30][3] , \w[30][2] , \w[30][1] , 1'b0}), .CI(1'b0), .S({\w[31][31] , 
        \w[31][30] , \w[31][29] , \w[31][28] , \w[31][27] , \w[31][26] , 
        \w[31][25] , \w[31][24] , \w[31][23] , \w[31][22] , \w[31][21] , 
        \w[31][20] , \w[31][19] , \w[31][18] , \w[31][17] , \w[31][16] , 
        \w[31][15] , \w[31][14] , \w[31][13] , \w[31][12] , \w[31][11] , 
        \w[31][10] , \w[31][9] , \w[31][8] , \w[31][7] , \w[31][6] , 
        \w[31][5] , \w[31][4] , \w[31][3] , \w[31][2] , \w[31][1] , 
        SYNOPSYS_UNCONNECTED__29}) );
  ADD_N32_97 \FAINST[31].ADD_  ( .A({\_60_net_[31] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({\w[31][31] , \w[31][30] , \w[31][29] , 
        \w[31][28] , \w[31][27] , \w[31][26] , \w[31][25] , \w[31][24] , 
        \w[31][23] , \w[31][22] , \w[31][21] , \w[31][20] , \w[31][19] , 
        \w[31][18] , \w[31][17] , \w[31][16] , \w[31][15] , \w[31][14] , 
        \w[31][13] , \w[31][12] , \w[31][11] , \w[31][10] , \w[31][9] , 
        \w[31][8] , \w[31][7] , \w[31][6] , \w[31][5] , \w[31][4] , \w[31][3] , 
        \w[31][2] , \w[31][1] , 1'b0}), .CI(1'b0), .S({O[31:1], 
        SYNOPSYS_UNCONNECTED__30}) );
  AND U2 ( .A(A[5]), .B(B[4]), .Z(\_8_net_[9] ) );
  AND U3 ( .A(A[5]), .B(B[3]), .Z(\_8_net_[8] ) );
  AND U4 ( .A(A[5]), .B(B[2]), .Z(\_8_net_[7] ) );
  AND U5 ( .A(A[5]), .B(B[1]), .Z(\_8_net_[6] ) );
  AND U6 ( .A(A[5]), .B(B[0]), .Z(\_8_net_[5] ) );
  AND U7 ( .A(A[5]), .B(B[26]), .Z(\_8_net_[31] ) );
  AND U8 ( .A(A[5]), .B(B[25]), .Z(\_8_net_[30] ) );
  AND U9 ( .A(A[5]), .B(B[24]), .Z(\_8_net_[29] ) );
  AND U10 ( .A(A[5]), .B(B[23]), .Z(\_8_net_[28] ) );
  AND U11 ( .A(A[5]), .B(B[22]), .Z(\_8_net_[27] ) );
  AND U12 ( .A(A[5]), .B(B[21]), .Z(\_8_net_[26] ) );
  AND U13 ( .A(A[5]), .B(B[20]), .Z(\_8_net_[25] ) );
  AND U14 ( .A(A[5]), .B(B[19]), .Z(\_8_net_[24] ) );
  AND U15 ( .A(A[5]), .B(B[18]), .Z(\_8_net_[23] ) );
  AND U16 ( .A(A[5]), .B(B[17]), .Z(\_8_net_[22] ) );
  AND U17 ( .A(A[5]), .B(B[16]), .Z(\_8_net_[21] ) );
  AND U18 ( .A(A[5]), .B(B[15]), .Z(\_8_net_[20] ) );
  AND U19 ( .A(A[5]), .B(B[14]), .Z(\_8_net_[19] ) );
  AND U20 ( .A(A[5]), .B(B[13]), .Z(\_8_net_[18] ) );
  AND U21 ( .A(A[5]), .B(B[12]), .Z(\_8_net_[17] ) );
  AND U22 ( .A(A[5]), .B(B[11]), .Z(\_8_net_[16] ) );
  AND U23 ( .A(A[5]), .B(B[10]), .Z(\_8_net_[15] ) );
  AND U24 ( .A(A[5]), .B(B[9]), .Z(\_8_net_[14] ) );
  AND U25 ( .A(A[5]), .B(B[8]), .Z(\_8_net_[13] ) );
  AND U26 ( .A(A[5]), .B(B[7]), .Z(\_8_net_[12] ) );
  AND U27 ( .A(A[5]), .B(B[6]), .Z(\_8_net_[11] ) );
  AND U28 ( .A(A[5]), .B(B[5]), .Z(\_8_net_[10] ) );
  AND U29 ( .A(B[5]), .B(A[4]), .Z(\_6_net_[9] ) );
  AND U30 ( .A(B[4]), .B(A[4]), .Z(\_6_net_[8] ) );
  AND U31 ( .A(B[3]), .B(A[4]), .Z(\_6_net_[7] ) );
  AND U32 ( .A(B[2]), .B(A[4]), .Z(\_6_net_[6] ) );
  AND U33 ( .A(B[1]), .B(A[4]), .Z(\_6_net_[5] ) );
  AND U34 ( .A(B[0]), .B(A[4]), .Z(\_6_net_[4] ) );
  AND U35 ( .A(A[4]), .B(B[27]), .Z(\_6_net_[31] ) );
  AND U36 ( .A(B[26]), .B(A[4]), .Z(\_6_net_[30] ) );
  AND U37 ( .A(B[25]), .B(A[4]), .Z(\_6_net_[29] ) );
  AND U38 ( .A(B[24]), .B(A[4]), .Z(\_6_net_[28] ) );
  AND U39 ( .A(B[23]), .B(A[4]), .Z(\_6_net_[27] ) );
  AND U40 ( .A(B[22]), .B(A[4]), .Z(\_6_net_[26] ) );
  AND U41 ( .A(B[21]), .B(A[4]), .Z(\_6_net_[25] ) );
  AND U42 ( .A(B[20]), .B(A[4]), .Z(\_6_net_[24] ) );
  AND U43 ( .A(B[19]), .B(A[4]), .Z(\_6_net_[23] ) );
  AND U44 ( .A(B[18]), .B(A[4]), .Z(\_6_net_[22] ) );
  AND U45 ( .A(B[17]), .B(A[4]), .Z(\_6_net_[21] ) );
  AND U46 ( .A(B[16]), .B(A[4]), .Z(\_6_net_[20] ) );
  AND U47 ( .A(B[15]), .B(A[4]), .Z(\_6_net_[19] ) );
  AND U48 ( .A(B[14]), .B(A[4]), .Z(\_6_net_[18] ) );
  AND U49 ( .A(B[13]), .B(A[4]), .Z(\_6_net_[17] ) );
  AND U50 ( .A(B[12]), .B(A[4]), .Z(\_6_net_[16] ) );
  AND U51 ( .A(B[11]), .B(A[4]), .Z(\_6_net_[15] ) );
  AND U52 ( .A(B[10]), .B(A[4]), .Z(\_6_net_[14] ) );
  AND U53 ( .A(B[9]), .B(A[4]), .Z(\_6_net_[13] ) );
  AND U54 ( .A(B[8]), .B(A[4]), .Z(\_6_net_[12] ) );
  AND U55 ( .A(B[7]), .B(A[4]), .Z(\_6_net_[11] ) );
  AND U56 ( .A(B[6]), .B(A[4]), .Z(\_6_net_[10] ) );
  AND U57 ( .A(A[31]), .B(B[0]), .Z(\_60_net_[31] ) );
  AND U58 ( .A(B[1]), .B(A[30]), .Z(\_58_net_[31] ) );
  AND U59 ( .A(A[30]), .B(B[0]), .Z(\_58_net_[30] ) );
  AND U60 ( .A(B[2]), .B(A[29]), .Z(\_56_net_[31] ) );
  AND U61 ( .A(B[1]), .B(A[29]), .Z(\_56_net_[30] ) );
  AND U62 ( .A(A[29]), .B(B[0]), .Z(\_56_net_[29] ) );
  AND U63 ( .A(B[3]), .B(A[28]), .Z(\_54_net_[31] ) );
  AND U64 ( .A(B[2]), .B(A[28]), .Z(\_54_net_[30] ) );
  AND U65 ( .A(B[1]), .B(A[28]), .Z(\_54_net_[29] ) );
  AND U66 ( .A(A[28]), .B(B[0]), .Z(\_54_net_[28] ) );
  AND U67 ( .A(B[4]), .B(A[27]), .Z(\_52_net_[31] ) );
  AND U68 ( .A(B[3]), .B(A[27]), .Z(\_52_net_[30] ) );
  AND U69 ( .A(B[2]), .B(A[27]), .Z(\_52_net_[29] ) );
  AND U70 ( .A(B[1]), .B(A[27]), .Z(\_52_net_[28] ) );
  AND U71 ( .A(A[27]), .B(B[0]), .Z(\_52_net_[27] ) );
  AND U72 ( .A(B[5]), .B(A[26]), .Z(\_50_net_[31] ) );
  AND U73 ( .A(B[4]), .B(A[26]), .Z(\_50_net_[30] ) );
  AND U74 ( .A(B[3]), .B(A[26]), .Z(\_50_net_[29] ) );
  AND U75 ( .A(B[2]), .B(A[26]), .Z(\_50_net_[28] ) );
  AND U76 ( .A(B[1]), .B(A[26]), .Z(\_50_net_[27] ) );
  AND U77 ( .A(A[26]), .B(B[0]), .Z(\_50_net_[26] ) );
  AND U78 ( .A(B[6]), .B(A[3]), .Z(\_4_net_[9] ) );
  AND U79 ( .A(B[5]), .B(A[3]), .Z(\_4_net_[8] ) );
  AND U80 ( .A(B[4]), .B(A[3]), .Z(\_4_net_[7] ) );
  AND U81 ( .A(B[3]), .B(A[3]), .Z(\_4_net_[6] ) );
  AND U82 ( .A(B[2]), .B(A[3]), .Z(\_4_net_[5] ) );
  AND U83 ( .A(B[1]), .B(A[3]), .Z(\_4_net_[4] ) );
  AND U84 ( .A(B[0]), .B(A[3]), .Z(\_4_net_[3] ) );
  AND U85 ( .A(A[3]), .B(B[28]), .Z(\_4_net_[31] ) );
  AND U86 ( .A(B[27]), .B(A[3]), .Z(\_4_net_[30] ) );
  AND U87 ( .A(B[26]), .B(A[3]), .Z(\_4_net_[29] ) );
  AND U88 ( .A(B[25]), .B(A[3]), .Z(\_4_net_[28] ) );
  AND U89 ( .A(B[24]), .B(A[3]), .Z(\_4_net_[27] ) );
  AND U90 ( .A(B[23]), .B(A[3]), .Z(\_4_net_[26] ) );
  AND U91 ( .A(B[22]), .B(A[3]), .Z(\_4_net_[25] ) );
  AND U92 ( .A(B[21]), .B(A[3]), .Z(\_4_net_[24] ) );
  AND U93 ( .A(B[20]), .B(A[3]), .Z(\_4_net_[23] ) );
  AND U94 ( .A(B[19]), .B(A[3]), .Z(\_4_net_[22] ) );
  AND U95 ( .A(B[18]), .B(A[3]), .Z(\_4_net_[21] ) );
  AND U96 ( .A(B[17]), .B(A[3]), .Z(\_4_net_[20] ) );
  AND U97 ( .A(B[16]), .B(A[3]), .Z(\_4_net_[19] ) );
  AND U98 ( .A(B[15]), .B(A[3]), .Z(\_4_net_[18] ) );
  AND U99 ( .A(B[14]), .B(A[3]), .Z(\_4_net_[17] ) );
  AND U100 ( .A(B[13]), .B(A[3]), .Z(\_4_net_[16] ) );
  AND U101 ( .A(B[12]), .B(A[3]), .Z(\_4_net_[15] ) );
  AND U102 ( .A(B[11]), .B(A[3]), .Z(\_4_net_[14] ) );
  AND U103 ( .A(B[10]), .B(A[3]), .Z(\_4_net_[13] ) );
  AND U104 ( .A(B[9]), .B(A[3]), .Z(\_4_net_[12] ) );
  AND U105 ( .A(B[8]), .B(A[3]), .Z(\_4_net_[11] ) );
  AND U106 ( .A(B[7]), .B(A[3]), .Z(\_4_net_[10] ) );
  AND U107 ( .A(B[6]), .B(A[25]), .Z(\_48_net_[31] ) );
  AND U108 ( .A(B[5]), .B(A[25]), .Z(\_48_net_[30] ) );
  AND U109 ( .A(B[4]), .B(A[25]), .Z(\_48_net_[29] ) );
  AND U110 ( .A(B[3]), .B(A[25]), .Z(\_48_net_[28] ) );
  AND U111 ( .A(B[2]), .B(A[25]), .Z(\_48_net_[27] ) );
  AND U112 ( .A(B[1]), .B(A[25]), .Z(\_48_net_[26] ) );
  AND U113 ( .A(A[25]), .B(B[0]), .Z(\_48_net_[25] ) );
  AND U114 ( .A(B[7]), .B(A[24]), .Z(\_46_net_[31] ) );
  AND U115 ( .A(B[6]), .B(A[24]), .Z(\_46_net_[30] ) );
  AND U116 ( .A(B[5]), .B(A[24]), .Z(\_46_net_[29] ) );
  AND U117 ( .A(B[4]), .B(A[24]), .Z(\_46_net_[28] ) );
  AND U118 ( .A(B[3]), .B(A[24]), .Z(\_46_net_[27] ) );
  AND U119 ( .A(B[2]), .B(A[24]), .Z(\_46_net_[26] ) );
  AND U120 ( .A(B[1]), .B(A[24]), .Z(\_46_net_[25] ) );
  AND U121 ( .A(A[24]), .B(B[0]), .Z(\_46_net_[24] ) );
  AND U122 ( .A(B[8]), .B(A[23]), .Z(\_44_net_[31] ) );
  AND U123 ( .A(B[7]), .B(A[23]), .Z(\_44_net_[30] ) );
  AND U124 ( .A(B[6]), .B(A[23]), .Z(\_44_net_[29] ) );
  AND U125 ( .A(B[5]), .B(A[23]), .Z(\_44_net_[28] ) );
  AND U126 ( .A(B[4]), .B(A[23]), .Z(\_44_net_[27] ) );
  AND U127 ( .A(B[3]), .B(A[23]), .Z(\_44_net_[26] ) );
  AND U128 ( .A(B[2]), .B(A[23]), .Z(\_44_net_[25] ) );
  AND U129 ( .A(B[1]), .B(A[23]), .Z(\_44_net_[24] ) );
  AND U130 ( .A(A[23]), .B(B[0]), .Z(\_44_net_[23] ) );
  AND U131 ( .A(B[9]), .B(A[22]), .Z(\_42_net_[31] ) );
  AND U132 ( .A(B[8]), .B(A[22]), .Z(\_42_net_[30] ) );
  AND U133 ( .A(B[7]), .B(A[22]), .Z(\_42_net_[29] ) );
  AND U134 ( .A(B[6]), .B(A[22]), .Z(\_42_net_[28] ) );
  AND U135 ( .A(B[5]), .B(A[22]), .Z(\_42_net_[27] ) );
  AND U136 ( .A(B[4]), .B(A[22]), .Z(\_42_net_[26] ) );
  AND U137 ( .A(B[3]), .B(A[22]), .Z(\_42_net_[25] ) );
  AND U138 ( .A(B[2]), .B(A[22]), .Z(\_42_net_[24] ) );
  AND U139 ( .A(B[1]), .B(A[22]), .Z(\_42_net_[23] ) );
  AND U140 ( .A(A[22]), .B(B[0]), .Z(\_42_net_[22] ) );
  AND U141 ( .A(B[10]), .B(A[21]), .Z(\_40_net_[31] ) );
  AND U142 ( .A(B[9]), .B(A[21]), .Z(\_40_net_[30] ) );
  AND U143 ( .A(B[8]), .B(A[21]), .Z(\_40_net_[29] ) );
  AND U144 ( .A(B[7]), .B(A[21]), .Z(\_40_net_[28] ) );
  AND U145 ( .A(B[6]), .B(A[21]), .Z(\_40_net_[27] ) );
  AND U146 ( .A(B[5]), .B(A[21]), .Z(\_40_net_[26] ) );
  AND U147 ( .A(B[4]), .B(A[21]), .Z(\_40_net_[25] ) );
  AND U148 ( .A(B[3]), .B(A[21]), .Z(\_40_net_[24] ) );
  AND U149 ( .A(B[2]), .B(A[21]), .Z(\_40_net_[23] ) );
  AND U150 ( .A(B[1]), .B(A[21]), .Z(\_40_net_[22] ) );
  AND U151 ( .A(A[21]), .B(B[0]), .Z(\_40_net_[21] ) );
  AND U152 ( .A(B[11]), .B(A[20]), .Z(\_38_net_[31] ) );
  AND U153 ( .A(B[10]), .B(A[20]), .Z(\_38_net_[30] ) );
  AND U154 ( .A(B[9]), .B(A[20]), .Z(\_38_net_[29] ) );
  AND U155 ( .A(B[8]), .B(A[20]), .Z(\_38_net_[28] ) );
  AND U156 ( .A(B[7]), .B(A[20]), .Z(\_38_net_[27] ) );
  AND U157 ( .A(B[6]), .B(A[20]), .Z(\_38_net_[26] ) );
  AND U158 ( .A(B[5]), .B(A[20]), .Z(\_38_net_[25] ) );
  AND U159 ( .A(B[4]), .B(A[20]), .Z(\_38_net_[24] ) );
  AND U160 ( .A(B[3]), .B(A[20]), .Z(\_38_net_[23] ) );
  AND U161 ( .A(B[2]), .B(A[20]), .Z(\_38_net_[22] ) );
  AND U162 ( .A(B[1]), .B(A[20]), .Z(\_38_net_[21] ) );
  AND U163 ( .A(A[20]), .B(B[0]), .Z(\_38_net_[20] ) );
  AND U164 ( .A(B[12]), .B(A[19]), .Z(\_36_net_[31] ) );
  AND U165 ( .A(B[11]), .B(A[19]), .Z(\_36_net_[30] ) );
  AND U166 ( .A(B[10]), .B(A[19]), .Z(\_36_net_[29] ) );
  AND U167 ( .A(B[9]), .B(A[19]), .Z(\_36_net_[28] ) );
  AND U168 ( .A(B[8]), .B(A[19]), .Z(\_36_net_[27] ) );
  AND U169 ( .A(B[7]), .B(A[19]), .Z(\_36_net_[26] ) );
  AND U170 ( .A(B[6]), .B(A[19]), .Z(\_36_net_[25] ) );
  AND U171 ( .A(B[5]), .B(A[19]), .Z(\_36_net_[24] ) );
  AND U172 ( .A(B[4]), .B(A[19]), .Z(\_36_net_[23] ) );
  AND U173 ( .A(B[3]), .B(A[19]), .Z(\_36_net_[22] ) );
  AND U174 ( .A(B[2]), .B(A[19]), .Z(\_36_net_[21] ) );
  AND U175 ( .A(B[1]), .B(A[19]), .Z(\_36_net_[20] ) );
  AND U176 ( .A(A[19]), .B(B[0]), .Z(\_36_net_[19] ) );
  AND U177 ( .A(B[13]), .B(A[18]), .Z(\_34_net_[31] ) );
  AND U178 ( .A(B[12]), .B(A[18]), .Z(\_34_net_[30] ) );
  AND U179 ( .A(B[11]), .B(A[18]), .Z(\_34_net_[29] ) );
  AND U180 ( .A(B[10]), .B(A[18]), .Z(\_34_net_[28] ) );
  AND U181 ( .A(B[9]), .B(A[18]), .Z(\_34_net_[27] ) );
  AND U182 ( .A(B[8]), .B(A[18]), .Z(\_34_net_[26] ) );
  AND U183 ( .A(B[7]), .B(A[18]), .Z(\_34_net_[25] ) );
  AND U184 ( .A(B[6]), .B(A[18]), .Z(\_34_net_[24] ) );
  AND U185 ( .A(B[5]), .B(A[18]), .Z(\_34_net_[23] ) );
  AND U186 ( .A(B[4]), .B(A[18]), .Z(\_34_net_[22] ) );
  AND U187 ( .A(B[3]), .B(A[18]), .Z(\_34_net_[21] ) );
  AND U188 ( .A(B[2]), .B(A[18]), .Z(\_34_net_[20] ) );
  AND U189 ( .A(B[1]), .B(A[18]), .Z(\_34_net_[19] ) );
  AND U190 ( .A(A[18]), .B(B[0]), .Z(\_34_net_[18] ) );
  AND U191 ( .A(B[14]), .B(A[17]), .Z(\_32_net_[31] ) );
  AND U192 ( .A(B[13]), .B(A[17]), .Z(\_32_net_[30] ) );
  AND U193 ( .A(B[12]), .B(A[17]), .Z(\_32_net_[29] ) );
  AND U194 ( .A(B[11]), .B(A[17]), .Z(\_32_net_[28] ) );
  AND U195 ( .A(B[10]), .B(A[17]), .Z(\_32_net_[27] ) );
  AND U196 ( .A(B[9]), .B(A[17]), .Z(\_32_net_[26] ) );
  AND U197 ( .A(B[8]), .B(A[17]), .Z(\_32_net_[25] ) );
  AND U198 ( .A(B[7]), .B(A[17]), .Z(\_32_net_[24] ) );
  AND U199 ( .A(B[6]), .B(A[17]), .Z(\_32_net_[23] ) );
  AND U200 ( .A(B[5]), .B(A[17]), .Z(\_32_net_[22] ) );
  AND U201 ( .A(B[4]), .B(A[17]), .Z(\_32_net_[21] ) );
  AND U202 ( .A(B[3]), .B(A[17]), .Z(\_32_net_[20] ) );
  AND U203 ( .A(B[2]), .B(A[17]), .Z(\_32_net_[19] ) );
  AND U204 ( .A(B[1]), .B(A[17]), .Z(\_32_net_[18] ) );
  AND U205 ( .A(A[17]), .B(B[0]), .Z(\_32_net_[17] ) );
  AND U206 ( .A(B[15]), .B(A[16]), .Z(\_30_net_[31] ) );
  AND U207 ( .A(B[14]), .B(A[16]), .Z(\_30_net_[30] ) );
  AND U208 ( .A(B[13]), .B(A[16]), .Z(\_30_net_[29] ) );
  AND U209 ( .A(B[12]), .B(A[16]), .Z(\_30_net_[28] ) );
  AND U210 ( .A(B[11]), .B(A[16]), .Z(\_30_net_[27] ) );
  AND U211 ( .A(B[10]), .B(A[16]), .Z(\_30_net_[26] ) );
  AND U212 ( .A(B[9]), .B(A[16]), .Z(\_30_net_[25] ) );
  AND U213 ( .A(B[8]), .B(A[16]), .Z(\_30_net_[24] ) );
  AND U214 ( .A(B[7]), .B(A[16]), .Z(\_30_net_[23] ) );
  AND U215 ( .A(B[6]), .B(A[16]), .Z(\_30_net_[22] ) );
  AND U216 ( .A(B[5]), .B(A[16]), .Z(\_30_net_[21] ) );
  AND U217 ( .A(B[4]), .B(A[16]), .Z(\_30_net_[20] ) );
  AND U218 ( .A(B[3]), .B(A[16]), .Z(\_30_net_[19] ) );
  AND U219 ( .A(B[2]), .B(A[16]), .Z(\_30_net_[18] ) );
  AND U220 ( .A(B[1]), .B(A[16]), .Z(\_30_net_[17] ) );
  AND U221 ( .A(A[16]), .B(B[0]), .Z(\_30_net_[16] ) );
  AND U222 ( .A(B[7]), .B(A[2]), .Z(\_2_net_[9] ) );
  AND U223 ( .A(B[6]), .B(A[2]), .Z(\_2_net_[8] ) );
  AND U224 ( .A(B[5]), .B(A[2]), .Z(\_2_net_[7] ) );
  AND U225 ( .A(B[4]), .B(A[2]), .Z(\_2_net_[6] ) );
  AND U226 ( .A(B[3]), .B(A[2]), .Z(\_2_net_[5] ) );
  AND U227 ( .A(B[2]), .B(A[2]), .Z(\_2_net_[4] ) );
  AND U228 ( .A(B[1]), .B(A[2]), .Z(\_2_net_[3] ) );
  AND U229 ( .A(A[2]), .B(B[29]), .Z(\_2_net_[31] ) );
  AND U230 ( .A(B[28]), .B(A[2]), .Z(\_2_net_[30] ) );
  AND U231 ( .A(B[0]), .B(A[2]), .Z(\_2_net_[2] ) );
  AND U232 ( .A(B[27]), .B(A[2]), .Z(\_2_net_[29] ) );
  AND U233 ( .A(B[26]), .B(A[2]), .Z(\_2_net_[28] ) );
  AND U234 ( .A(B[25]), .B(A[2]), .Z(\_2_net_[27] ) );
  AND U235 ( .A(B[24]), .B(A[2]), .Z(\_2_net_[26] ) );
  AND U236 ( .A(B[23]), .B(A[2]), .Z(\_2_net_[25] ) );
  AND U237 ( .A(B[22]), .B(A[2]), .Z(\_2_net_[24] ) );
  AND U238 ( .A(B[21]), .B(A[2]), .Z(\_2_net_[23] ) );
  AND U239 ( .A(B[20]), .B(A[2]), .Z(\_2_net_[22] ) );
  AND U240 ( .A(B[19]), .B(A[2]), .Z(\_2_net_[21] ) );
  AND U241 ( .A(B[18]), .B(A[2]), .Z(\_2_net_[20] ) );
  AND U242 ( .A(B[17]), .B(A[2]), .Z(\_2_net_[19] ) );
  AND U243 ( .A(B[16]), .B(A[2]), .Z(\_2_net_[18] ) );
  AND U244 ( .A(B[15]), .B(A[2]), .Z(\_2_net_[17] ) );
  AND U245 ( .A(B[14]), .B(A[2]), .Z(\_2_net_[16] ) );
  AND U246 ( .A(B[13]), .B(A[2]), .Z(\_2_net_[15] ) );
  AND U247 ( .A(B[12]), .B(A[2]), .Z(\_2_net_[14] ) );
  AND U248 ( .A(B[11]), .B(A[2]), .Z(\_2_net_[13] ) );
  AND U249 ( .A(B[10]), .B(A[2]), .Z(\_2_net_[12] ) );
  AND U250 ( .A(B[9]), .B(A[2]), .Z(\_2_net_[11] ) );
  AND U251 ( .A(B[8]), .B(A[2]), .Z(\_2_net_[10] ) );
  AND U252 ( .A(B[16]), .B(A[15]), .Z(\_28_net_[31] ) );
  AND U253 ( .A(B[15]), .B(A[15]), .Z(\_28_net_[30] ) );
  AND U254 ( .A(B[14]), .B(A[15]), .Z(\_28_net_[29] ) );
  AND U255 ( .A(B[13]), .B(A[15]), .Z(\_28_net_[28] ) );
  AND U256 ( .A(B[12]), .B(A[15]), .Z(\_28_net_[27] ) );
  AND U257 ( .A(B[11]), .B(A[15]), .Z(\_28_net_[26] ) );
  AND U258 ( .A(B[10]), .B(A[15]), .Z(\_28_net_[25] ) );
  AND U259 ( .A(B[9]), .B(A[15]), .Z(\_28_net_[24] ) );
  AND U260 ( .A(B[8]), .B(A[15]), .Z(\_28_net_[23] ) );
  AND U261 ( .A(B[7]), .B(A[15]), .Z(\_28_net_[22] ) );
  AND U262 ( .A(B[6]), .B(A[15]), .Z(\_28_net_[21] ) );
  AND U263 ( .A(B[5]), .B(A[15]), .Z(\_28_net_[20] ) );
  AND U264 ( .A(B[4]), .B(A[15]), .Z(\_28_net_[19] ) );
  AND U265 ( .A(B[3]), .B(A[15]), .Z(\_28_net_[18] ) );
  AND U266 ( .A(B[2]), .B(A[15]), .Z(\_28_net_[17] ) );
  AND U267 ( .A(B[1]), .B(A[15]), .Z(\_28_net_[16] ) );
  AND U268 ( .A(A[15]), .B(B[0]), .Z(\_28_net_[15] ) );
  AND U269 ( .A(B[17]), .B(A[14]), .Z(\_26_net_[31] ) );
  AND U270 ( .A(B[16]), .B(A[14]), .Z(\_26_net_[30] ) );
  AND U271 ( .A(B[15]), .B(A[14]), .Z(\_26_net_[29] ) );
  AND U272 ( .A(B[14]), .B(A[14]), .Z(\_26_net_[28] ) );
  AND U273 ( .A(B[13]), .B(A[14]), .Z(\_26_net_[27] ) );
  AND U274 ( .A(B[12]), .B(A[14]), .Z(\_26_net_[26] ) );
  AND U275 ( .A(B[11]), .B(A[14]), .Z(\_26_net_[25] ) );
  AND U276 ( .A(B[10]), .B(A[14]), .Z(\_26_net_[24] ) );
  AND U277 ( .A(B[9]), .B(A[14]), .Z(\_26_net_[23] ) );
  AND U278 ( .A(B[8]), .B(A[14]), .Z(\_26_net_[22] ) );
  AND U279 ( .A(B[7]), .B(A[14]), .Z(\_26_net_[21] ) );
  AND U280 ( .A(B[6]), .B(A[14]), .Z(\_26_net_[20] ) );
  AND U281 ( .A(B[5]), .B(A[14]), .Z(\_26_net_[19] ) );
  AND U282 ( .A(B[4]), .B(A[14]), .Z(\_26_net_[18] ) );
  AND U283 ( .A(B[3]), .B(A[14]), .Z(\_26_net_[17] ) );
  AND U284 ( .A(B[2]), .B(A[14]), .Z(\_26_net_[16] ) );
  AND U285 ( .A(B[1]), .B(A[14]), .Z(\_26_net_[15] ) );
  AND U286 ( .A(A[14]), .B(B[0]), .Z(\_26_net_[14] ) );
  AND U287 ( .A(B[18]), .B(A[13]), .Z(\_24_net_[31] ) );
  AND U288 ( .A(B[17]), .B(A[13]), .Z(\_24_net_[30] ) );
  AND U289 ( .A(B[16]), .B(A[13]), .Z(\_24_net_[29] ) );
  AND U290 ( .A(B[15]), .B(A[13]), .Z(\_24_net_[28] ) );
  AND U291 ( .A(B[14]), .B(A[13]), .Z(\_24_net_[27] ) );
  AND U292 ( .A(B[13]), .B(A[13]), .Z(\_24_net_[26] ) );
  AND U293 ( .A(B[12]), .B(A[13]), .Z(\_24_net_[25] ) );
  AND U294 ( .A(B[11]), .B(A[13]), .Z(\_24_net_[24] ) );
  AND U295 ( .A(B[10]), .B(A[13]), .Z(\_24_net_[23] ) );
  AND U296 ( .A(B[9]), .B(A[13]), .Z(\_24_net_[22] ) );
  AND U297 ( .A(B[8]), .B(A[13]), .Z(\_24_net_[21] ) );
  AND U298 ( .A(B[7]), .B(A[13]), .Z(\_24_net_[20] ) );
  AND U299 ( .A(B[6]), .B(A[13]), .Z(\_24_net_[19] ) );
  AND U300 ( .A(B[5]), .B(A[13]), .Z(\_24_net_[18] ) );
  AND U301 ( .A(B[4]), .B(A[13]), .Z(\_24_net_[17] ) );
  AND U302 ( .A(B[3]), .B(A[13]), .Z(\_24_net_[16] ) );
  AND U303 ( .A(B[2]), .B(A[13]), .Z(\_24_net_[15] ) );
  AND U304 ( .A(B[1]), .B(A[13]), .Z(\_24_net_[14] ) );
  AND U305 ( .A(A[13]), .B(B[0]), .Z(\_24_net_[13] ) );
  AND U306 ( .A(B[19]), .B(A[12]), .Z(\_22_net_[31] ) );
  AND U307 ( .A(B[18]), .B(A[12]), .Z(\_22_net_[30] ) );
  AND U308 ( .A(B[17]), .B(A[12]), .Z(\_22_net_[29] ) );
  AND U309 ( .A(B[16]), .B(A[12]), .Z(\_22_net_[28] ) );
  AND U310 ( .A(B[15]), .B(A[12]), .Z(\_22_net_[27] ) );
  AND U311 ( .A(B[14]), .B(A[12]), .Z(\_22_net_[26] ) );
  AND U312 ( .A(B[13]), .B(A[12]), .Z(\_22_net_[25] ) );
  AND U313 ( .A(B[12]), .B(A[12]), .Z(\_22_net_[24] ) );
  AND U314 ( .A(B[11]), .B(A[12]), .Z(\_22_net_[23] ) );
  AND U315 ( .A(B[10]), .B(A[12]), .Z(\_22_net_[22] ) );
  AND U316 ( .A(B[9]), .B(A[12]), .Z(\_22_net_[21] ) );
  AND U317 ( .A(B[8]), .B(A[12]), .Z(\_22_net_[20] ) );
  AND U318 ( .A(B[7]), .B(A[12]), .Z(\_22_net_[19] ) );
  AND U319 ( .A(B[6]), .B(A[12]), .Z(\_22_net_[18] ) );
  AND U320 ( .A(B[5]), .B(A[12]), .Z(\_22_net_[17] ) );
  AND U321 ( .A(B[4]), .B(A[12]), .Z(\_22_net_[16] ) );
  AND U322 ( .A(B[3]), .B(A[12]), .Z(\_22_net_[15] ) );
  AND U323 ( .A(B[2]), .B(A[12]), .Z(\_22_net_[14] ) );
  AND U324 ( .A(B[1]), .B(A[12]), .Z(\_22_net_[13] ) );
  AND U325 ( .A(A[12]), .B(B[0]), .Z(\_22_net_[12] ) );
  AND U326 ( .A(B[20]), .B(A[11]), .Z(\_20_net_[31] ) );
  AND U327 ( .A(B[19]), .B(A[11]), .Z(\_20_net_[30] ) );
  AND U328 ( .A(B[18]), .B(A[11]), .Z(\_20_net_[29] ) );
  AND U329 ( .A(B[17]), .B(A[11]), .Z(\_20_net_[28] ) );
  AND U330 ( .A(B[16]), .B(A[11]), .Z(\_20_net_[27] ) );
  AND U331 ( .A(B[15]), .B(A[11]), .Z(\_20_net_[26] ) );
  AND U332 ( .A(B[14]), .B(A[11]), .Z(\_20_net_[25] ) );
  AND U333 ( .A(B[13]), .B(A[11]), .Z(\_20_net_[24] ) );
  AND U334 ( .A(B[12]), .B(A[11]), .Z(\_20_net_[23] ) );
  AND U335 ( .A(B[11]), .B(A[11]), .Z(\_20_net_[22] ) );
  AND U336 ( .A(B[10]), .B(A[11]), .Z(\_20_net_[21] ) );
  AND U337 ( .A(B[9]), .B(A[11]), .Z(\_20_net_[20] ) );
  AND U338 ( .A(B[8]), .B(A[11]), .Z(\_20_net_[19] ) );
  AND U339 ( .A(B[7]), .B(A[11]), .Z(\_20_net_[18] ) );
  AND U340 ( .A(B[6]), .B(A[11]), .Z(\_20_net_[17] ) );
  AND U341 ( .A(B[5]), .B(A[11]), .Z(\_20_net_[16] ) );
  AND U342 ( .A(B[4]), .B(A[11]), .Z(\_20_net_[15] ) );
  AND U343 ( .A(B[3]), .B(A[11]), .Z(\_20_net_[14] ) );
  AND U344 ( .A(B[2]), .B(A[11]), .Z(\_20_net_[13] ) );
  AND U345 ( .A(B[1]), .B(A[11]), .Z(\_20_net_[12] ) );
  AND U346 ( .A(A[11]), .B(B[0]), .Z(\_20_net_[11] ) );
  AND U347 ( .A(B[21]), .B(A[10]), .Z(\_18_net_[31] ) );
  AND U348 ( .A(B[20]), .B(A[10]), .Z(\_18_net_[30] ) );
  AND U349 ( .A(B[19]), .B(A[10]), .Z(\_18_net_[29] ) );
  AND U350 ( .A(B[18]), .B(A[10]), .Z(\_18_net_[28] ) );
  AND U351 ( .A(B[17]), .B(A[10]), .Z(\_18_net_[27] ) );
  AND U352 ( .A(B[16]), .B(A[10]), .Z(\_18_net_[26] ) );
  AND U353 ( .A(B[15]), .B(A[10]), .Z(\_18_net_[25] ) );
  AND U354 ( .A(B[14]), .B(A[10]), .Z(\_18_net_[24] ) );
  AND U355 ( .A(B[13]), .B(A[10]), .Z(\_18_net_[23] ) );
  AND U356 ( .A(B[12]), .B(A[10]), .Z(\_18_net_[22] ) );
  AND U357 ( .A(B[11]), .B(A[10]), .Z(\_18_net_[21] ) );
  AND U358 ( .A(B[10]), .B(A[10]), .Z(\_18_net_[20] ) );
  AND U359 ( .A(B[9]), .B(A[10]), .Z(\_18_net_[19] ) );
  AND U360 ( .A(B[8]), .B(A[10]), .Z(\_18_net_[18] ) );
  AND U361 ( .A(B[7]), .B(A[10]), .Z(\_18_net_[17] ) );
  AND U362 ( .A(B[6]), .B(A[10]), .Z(\_18_net_[16] ) );
  AND U363 ( .A(B[5]), .B(A[10]), .Z(\_18_net_[15] ) );
  AND U364 ( .A(B[4]), .B(A[10]), .Z(\_18_net_[14] ) );
  AND U365 ( .A(B[3]), .B(A[10]), .Z(\_18_net_[13] ) );
  AND U366 ( .A(B[2]), .B(A[10]), .Z(\_18_net_[12] ) );
  AND U367 ( .A(B[1]), .B(A[10]), .Z(\_18_net_[11] ) );
  AND U368 ( .A(A[10]), .B(B[0]), .Z(\_18_net_[10] ) );
  AND U369 ( .A(B[0]), .B(A[9]), .Z(\_16_net_[9] ) );
  AND U370 ( .A(B[22]), .B(A[9]), .Z(\_16_net_[31] ) );
  AND U371 ( .A(B[21]), .B(A[9]), .Z(\_16_net_[30] ) );
  AND U372 ( .A(B[20]), .B(A[9]), .Z(\_16_net_[29] ) );
  AND U373 ( .A(B[19]), .B(A[9]), .Z(\_16_net_[28] ) );
  AND U374 ( .A(B[18]), .B(A[9]), .Z(\_16_net_[27] ) );
  AND U375 ( .A(B[17]), .B(A[9]), .Z(\_16_net_[26] ) );
  AND U376 ( .A(B[16]), .B(A[9]), .Z(\_16_net_[25] ) );
  AND U377 ( .A(B[15]), .B(A[9]), .Z(\_16_net_[24] ) );
  AND U378 ( .A(B[14]), .B(A[9]), .Z(\_16_net_[23] ) );
  AND U379 ( .A(B[13]), .B(A[9]), .Z(\_16_net_[22] ) );
  AND U380 ( .A(B[12]), .B(A[9]), .Z(\_16_net_[21] ) );
  AND U381 ( .A(B[11]), .B(A[9]), .Z(\_16_net_[20] ) );
  AND U382 ( .A(B[10]), .B(A[9]), .Z(\_16_net_[19] ) );
  AND U383 ( .A(B[9]), .B(A[9]), .Z(\_16_net_[18] ) );
  AND U384 ( .A(B[8]), .B(A[9]), .Z(\_16_net_[17] ) );
  AND U385 ( .A(B[7]), .B(A[9]), .Z(\_16_net_[16] ) );
  AND U386 ( .A(B[6]), .B(A[9]), .Z(\_16_net_[15] ) );
  AND U387 ( .A(B[5]), .B(A[9]), .Z(\_16_net_[14] ) );
  AND U388 ( .A(B[4]), .B(A[9]), .Z(\_16_net_[13] ) );
  AND U389 ( .A(B[3]), .B(A[9]), .Z(\_16_net_[12] ) );
  AND U390 ( .A(B[2]), .B(A[9]), .Z(\_16_net_[11] ) );
  AND U391 ( .A(A[9]), .B(B[1]), .Z(\_16_net_[10] ) );
  AND U392 ( .A(B[1]), .B(A[8]), .Z(\_14_net_[9] ) );
  AND U393 ( .A(B[0]), .B(A[8]), .Z(\_14_net_[8] ) );
  AND U394 ( .A(B[23]), .B(A[8]), .Z(\_14_net_[31] ) );
  AND U395 ( .A(B[22]), .B(A[8]), .Z(\_14_net_[30] ) );
  AND U396 ( .A(B[21]), .B(A[8]), .Z(\_14_net_[29] ) );
  AND U397 ( .A(B[20]), .B(A[8]), .Z(\_14_net_[28] ) );
  AND U398 ( .A(B[19]), .B(A[8]), .Z(\_14_net_[27] ) );
  AND U399 ( .A(B[18]), .B(A[8]), .Z(\_14_net_[26] ) );
  AND U400 ( .A(B[17]), .B(A[8]), .Z(\_14_net_[25] ) );
  AND U401 ( .A(B[16]), .B(A[8]), .Z(\_14_net_[24] ) );
  AND U402 ( .A(B[15]), .B(A[8]), .Z(\_14_net_[23] ) );
  AND U403 ( .A(B[14]), .B(A[8]), .Z(\_14_net_[22] ) );
  AND U404 ( .A(B[13]), .B(A[8]), .Z(\_14_net_[21] ) );
  AND U405 ( .A(B[12]), .B(A[8]), .Z(\_14_net_[20] ) );
  AND U406 ( .A(B[11]), .B(A[8]), .Z(\_14_net_[19] ) );
  AND U407 ( .A(B[10]), .B(A[8]), .Z(\_14_net_[18] ) );
  AND U408 ( .A(B[9]), .B(A[8]), .Z(\_14_net_[17] ) );
  AND U409 ( .A(B[8]), .B(A[8]), .Z(\_14_net_[16] ) );
  AND U410 ( .A(B[7]), .B(A[8]), .Z(\_14_net_[15] ) );
  AND U411 ( .A(B[6]), .B(A[8]), .Z(\_14_net_[14] ) );
  AND U412 ( .A(B[5]), .B(A[8]), .Z(\_14_net_[13] ) );
  AND U413 ( .A(B[4]), .B(A[8]), .Z(\_14_net_[12] ) );
  AND U414 ( .A(B[3]), .B(A[8]), .Z(\_14_net_[11] ) );
  AND U415 ( .A(A[8]), .B(B[2]), .Z(\_14_net_[10] ) );
  AND U416 ( .A(B[2]), .B(A[7]), .Z(\_12_net_[9] ) );
  AND U417 ( .A(B[1]), .B(A[7]), .Z(\_12_net_[8] ) );
  AND U418 ( .A(B[0]), .B(A[7]), .Z(\_12_net_[7] ) );
  AND U419 ( .A(B[24]), .B(A[7]), .Z(\_12_net_[31] ) );
  AND U420 ( .A(B[23]), .B(A[7]), .Z(\_12_net_[30] ) );
  AND U421 ( .A(B[22]), .B(A[7]), .Z(\_12_net_[29] ) );
  AND U422 ( .A(B[21]), .B(A[7]), .Z(\_12_net_[28] ) );
  AND U423 ( .A(B[20]), .B(A[7]), .Z(\_12_net_[27] ) );
  AND U424 ( .A(B[19]), .B(A[7]), .Z(\_12_net_[26] ) );
  AND U425 ( .A(B[18]), .B(A[7]), .Z(\_12_net_[25] ) );
  AND U426 ( .A(B[17]), .B(A[7]), .Z(\_12_net_[24] ) );
  AND U427 ( .A(B[16]), .B(A[7]), .Z(\_12_net_[23] ) );
  AND U428 ( .A(B[15]), .B(A[7]), .Z(\_12_net_[22] ) );
  AND U429 ( .A(B[14]), .B(A[7]), .Z(\_12_net_[21] ) );
  AND U430 ( .A(B[13]), .B(A[7]), .Z(\_12_net_[20] ) );
  AND U431 ( .A(B[12]), .B(A[7]), .Z(\_12_net_[19] ) );
  AND U432 ( .A(B[11]), .B(A[7]), .Z(\_12_net_[18] ) );
  AND U433 ( .A(B[10]), .B(A[7]), .Z(\_12_net_[17] ) );
  AND U434 ( .A(B[9]), .B(A[7]), .Z(\_12_net_[16] ) );
  AND U435 ( .A(B[8]), .B(A[7]), .Z(\_12_net_[15] ) );
  AND U436 ( .A(B[7]), .B(A[7]), .Z(\_12_net_[14] ) );
  AND U437 ( .A(B[6]), .B(A[7]), .Z(\_12_net_[13] ) );
  AND U438 ( .A(B[5]), .B(A[7]), .Z(\_12_net_[12] ) );
  AND U439 ( .A(B[4]), .B(A[7]), .Z(\_12_net_[11] ) );
  AND U440 ( .A(A[7]), .B(B[3]), .Z(\_12_net_[10] ) );
  AND U441 ( .A(B[3]), .B(A[6]), .Z(\_10_net_[9] ) );
  AND U442 ( .A(B[2]), .B(A[6]), .Z(\_10_net_[8] ) );
  AND U443 ( .A(B[1]), .B(A[6]), .Z(\_10_net_[7] ) );
  AND U444 ( .A(B[0]), .B(A[6]), .Z(\_10_net_[6] ) );
  AND U445 ( .A(B[25]), .B(A[6]), .Z(\_10_net_[31] ) );
  AND U446 ( .A(B[24]), .B(A[6]), .Z(\_10_net_[30] ) );
  AND U447 ( .A(B[23]), .B(A[6]), .Z(\_10_net_[29] ) );
  AND U448 ( .A(B[22]), .B(A[6]), .Z(\_10_net_[28] ) );
  AND U449 ( .A(B[21]), .B(A[6]), .Z(\_10_net_[27] ) );
  AND U450 ( .A(B[20]), .B(A[6]), .Z(\_10_net_[26] ) );
  AND U451 ( .A(B[19]), .B(A[6]), .Z(\_10_net_[25] ) );
  AND U452 ( .A(B[18]), .B(A[6]), .Z(\_10_net_[24] ) );
  AND U453 ( .A(B[17]), .B(A[6]), .Z(\_10_net_[23] ) );
  AND U454 ( .A(B[16]), .B(A[6]), .Z(\_10_net_[22] ) );
  AND U455 ( .A(B[15]), .B(A[6]), .Z(\_10_net_[21] ) );
  AND U456 ( .A(B[14]), .B(A[6]), .Z(\_10_net_[20] ) );
  AND U457 ( .A(B[13]), .B(A[6]), .Z(\_10_net_[19] ) );
  AND U458 ( .A(B[12]), .B(A[6]), .Z(\_10_net_[18] ) );
  AND U459 ( .A(B[11]), .B(A[6]), .Z(\_10_net_[17] ) );
  AND U460 ( .A(B[10]), .B(A[6]), .Z(\_10_net_[16] ) );
  AND U461 ( .A(B[9]), .B(A[6]), .Z(\_10_net_[15] ) );
  AND U462 ( .A(B[8]), .B(A[6]), .Z(\_10_net_[14] ) );
  AND U463 ( .A(B[7]), .B(A[6]), .Z(\_10_net_[13] ) );
  AND U464 ( .A(B[6]), .B(A[6]), .Z(\_10_net_[12] ) );
  AND U465 ( .A(B[5]), .B(A[6]), .Z(\_10_net_[11] ) );
  AND U466 ( .A(A[6]), .B(B[4]), .Z(\_10_net_[10] ) );
  AND U467 ( .A(B[8]), .B(A[1]), .Z(\_0_net_[9] ) );
  AND U468 ( .A(B[7]), .B(A[1]), .Z(\_0_net_[8] ) );
  AND U469 ( .A(B[6]), .B(A[1]), .Z(\_0_net_[7] ) );
  AND U470 ( .A(B[5]), .B(A[1]), .Z(\_0_net_[6] ) );
  AND U471 ( .A(B[4]), .B(A[1]), .Z(\_0_net_[5] ) );
  AND U472 ( .A(B[3]), .B(A[1]), .Z(\_0_net_[4] ) );
  AND U473 ( .A(B[2]), .B(A[1]), .Z(\_0_net_[3] ) );
  AND U474 ( .A(B[30]), .B(A[1]), .Z(\_0_net_[31] ) );
  AND U475 ( .A(B[29]), .B(A[1]), .Z(\_0_net_[30] ) );
  AND U476 ( .A(B[1]), .B(A[1]), .Z(\_0_net_[2] ) );
  AND U477 ( .A(B[28]), .B(A[1]), .Z(\_0_net_[29] ) );
  AND U478 ( .A(B[27]), .B(A[1]), .Z(\_0_net_[28] ) );
  AND U479 ( .A(B[26]), .B(A[1]), .Z(\_0_net_[27] ) );
  AND U480 ( .A(B[25]), .B(A[1]), .Z(\_0_net_[26] ) );
  AND U481 ( .A(B[24]), .B(A[1]), .Z(\_0_net_[25] ) );
  AND U482 ( .A(B[23]), .B(A[1]), .Z(\_0_net_[24] ) );
  AND U483 ( .A(B[22]), .B(A[1]), .Z(\_0_net_[23] ) );
  AND U484 ( .A(B[21]), .B(A[1]), .Z(\_0_net_[22] ) );
  AND U485 ( .A(B[20]), .B(A[1]), .Z(\_0_net_[21] ) );
  AND U486 ( .A(B[19]), .B(A[1]), .Z(\_0_net_[20] ) );
  AND U487 ( .A(B[0]), .B(A[1]), .Z(\_0_net_[1] ) );
  AND U488 ( .A(B[18]), .B(A[1]), .Z(\_0_net_[19] ) );
  AND U489 ( .A(B[17]), .B(A[1]), .Z(\_0_net_[18] ) );
  AND U490 ( .A(B[16]), .B(A[1]), .Z(\_0_net_[17] ) );
  AND U491 ( .A(B[15]), .B(A[1]), .Z(\_0_net_[16] ) );
  AND U492 ( .A(B[14]), .B(A[1]), .Z(\_0_net_[15] ) );
  AND U493 ( .A(B[13]), .B(A[1]), .Z(\_0_net_[14] ) );
  AND U494 ( .A(B[12]), .B(A[1]), .Z(\_0_net_[13] ) );
  AND U495 ( .A(B[11]), .B(A[1]), .Z(\_0_net_[12] ) );
  AND U496 ( .A(B[10]), .B(A[1]), .Z(\_0_net_[11] ) );
  AND U497 ( .A(A[1]), .B(B[9]), .Z(\_0_net_[10] ) );
endmodule


module FA_3969 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_3970 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3971 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3972 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3973 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3974 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3975 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3976 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3977 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3978 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3979 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3980 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3981 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3982 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3983 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3984 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3985 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3986 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3987 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3988 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3989 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3990 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3991 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3992 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3993 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3994 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3995 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3996 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3997 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3998 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3999 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_128 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;


  FA_3999 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3998 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3997 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3996 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3995 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3994 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3993 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3992 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3991 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3990 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3989 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3988 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_3987 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_3986 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_3985 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_3984 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_3983 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_3982 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_3981 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_3980 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_3979 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_3978 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_3977 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_3976 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_3975 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_3974 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_3973 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_3972 \FAINST[28].FA_  ( .A(1'b0), .B(B[28]), .CI(1'b0), .S(S[28]) );
  FA_3971 \FAINST[29].FA_  ( .A(1'b0), .B(B[29]), .CI(1'b0), .S(S[29]) );
  FA_3970 \FAINST[30].FA_  ( .A(1'b0), .B(B[30]), .CI(1'b0), .S(S[30]) );
  FA_3969 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(1'b0), .S(S[31]) );
endmodule


module FA_4001 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_4002 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_4003 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4004 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4005 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4006 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4007 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4008 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4009 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4010 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4011 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4012 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4013 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4014 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4015 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4016 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4017 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4018 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4019 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4020 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4021 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4022 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4023 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4024 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4025 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4026 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4027 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4028 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4029 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4030 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4031 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_129 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;
  wire   \C[31] ;

  FA_4031 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_4030 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_4029 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_4028 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_4027 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_4026 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_4025 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_4024 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_4023 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_4022 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_4021 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_4020 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_4019 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_4018 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_4017 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_4016 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_4015 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_4014 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_4013 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_4012 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_4011 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_4010 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_4009 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_4008 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_4007 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_4006 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_4005 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_4004 \FAINST[28].FA_  ( .A(1'b0), .B(B[28]), .CI(1'b0), .S(S[28]) );
  FA_4003 \FAINST[29].FA_  ( .A(1'b0), .B(B[29]), .CI(1'b0), .S(S[29]) );
  FA_4002 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(1'b0), .S(S[30]), .CO(
        \C[31] ) );
  FA_4001 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(\C[31] ), .S(S[31]) );
endmodule


module FA_4033 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_4034 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4035 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_4036 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4037 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4038 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4039 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4040 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4041 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4042 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4043 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4044 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4045 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4046 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4047 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4048 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4049 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4050 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4051 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4052 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4053 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4054 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4055 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4056 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4057 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4058 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4059 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4060 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4061 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4062 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4063 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_130 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_4063 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_4062 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_4061 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_4060 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_4059 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_4058 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_4057 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_4056 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_4055 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_4054 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_4053 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_4052 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_4051 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_4050 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_4049 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_4048 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_4047 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_4046 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_4045 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_4044 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_4043 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_4042 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_4041 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_4040 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_4039 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_4038 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_4037 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_4036 \FAINST[28].FA_  ( .A(1'b0), .B(B[28]), .CI(1'b0), .S(S[28]) );
  FA_4035 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(1'b0), .S(S[29]), .CO(
        C[30]) );
  FA_4034 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_4033 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_4065 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_4066 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4067 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4068 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_4069 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4070 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4071 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4072 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4073 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4074 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4075 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4076 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4077 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4078 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4079 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4080 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4081 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4082 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4083 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4084 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4085 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4086 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4087 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4088 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4089 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4090 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4091 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4092 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4093 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4094 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4095 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_131 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_4095 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_4094 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_4093 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_4092 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_4091 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_4090 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_4089 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_4088 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_4087 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_4086 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_4085 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_4084 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_4083 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_4082 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_4081 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_4080 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_4079 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_4078 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_4077 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_4076 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_4075 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_4074 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_4073 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_4072 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_4071 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_4070 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_4069 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_4068 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(1'b0), .S(S[28]), .CO(
        C[29]) );
  FA_4067 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_4066 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_4065 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_4097 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_4098 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4099 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_4102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4104 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4120 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_132 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_4127 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_4126 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_4125 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_4124 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_4123 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_4122 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_4121 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_4120 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_4119 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_4118 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_4117 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_4116 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_4115 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_4114 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_4113 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_4112 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_4111 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_4110 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_4109 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_4108 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_4107 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_4106 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_4105 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_4104 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_4103 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_4102 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_4101 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(1'b0), .S(S[27]), .CO(
        C[28]) );
  FA_4100 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_4099 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_4098 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_4097 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_4129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_4130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_4135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4136 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4152 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_133 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_4159 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_4158 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_4157 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_4156 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_4155 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_4154 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_4153 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_4152 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_4151 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_4150 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_4149 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_4148 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_4147 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_4146 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_4145 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_4144 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_4143 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_4142 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_4141 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_4140 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_4139 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_4138 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_4137 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_4136 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_4135 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_4134 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(1'b0), .S(S[26]), .CO(
        C[27]) );
  FA_4133 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_4132 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_4131 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_4130 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_4129 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_4161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_4162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_4168 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4184 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_134 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_4191 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_4190 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_4189 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_4188 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_4187 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_4186 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_4185 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_4184 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_4183 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_4182 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_4181 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_4180 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_4179 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_4178 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_4177 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_4176 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_4175 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_4174 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_4173 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_4172 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_4171 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_4170 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_4169 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_4168 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_4167 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(1'b0), .S(S[25]), .CO(
        C[26]) );
  FA_4166 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_4165 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_4164 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_4163 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_4162 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_4161 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_4193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_4194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4200 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_4201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4216 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_135 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_4223 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_4222 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_4221 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_4220 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_4219 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_4218 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_4217 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_4216 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_4215 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_4214 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_4213 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_4212 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_4211 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_4210 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_4209 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_4208 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_4207 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_4206 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_4205 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_4204 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_4203 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_4202 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_4201 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_4200 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(1'b0), .S(S[24]), .CO(
        C[25]) );
  FA_4199 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_4198 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_4197 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_4196 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_4195 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_4194 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_4193 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_4225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_4226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4232 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_4234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4248 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_136 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_4255 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_4254 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_4253 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_4252 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_4251 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_4250 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_4249 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_4248 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_4247 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_4246 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_4245 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_4244 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_4243 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_4242 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_4241 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_4240 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_4239 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_4238 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_4237 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_4236 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_4235 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_4234 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_4233 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(1'b0), .S(S[23]), .CO(
        C[24]) );
  FA_4232 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_4231 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_4230 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_4229 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_4228 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_4227 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_4226 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_4225 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_4257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_4258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4264 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_4267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4280 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_137 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_4287 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_4286 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_4285 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_4284 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_4283 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_4282 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_4281 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_4280 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_4279 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_4278 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_4277 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_4276 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_4275 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_4274 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_4273 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_4272 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_4271 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_4270 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_4269 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_4268 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_4267 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_4266 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(1'b0), .S(S[22]), .CO(
        C[23]) );
  FA_4265 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_4264 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_4263 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_4262 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_4261 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_4260 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_4259 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_4258 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_4257 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_4289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_4290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4296 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_4300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4312 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_138 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_4319 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_4318 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_4317 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_4316 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_4315 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_4314 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_4313 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_4312 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_4311 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_4310 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_4309 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_4308 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_4307 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_4306 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_4305 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_4304 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_4303 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_4302 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_4301 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_4300 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_4299 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(1'b0), .S(S[21]), .CO(
        C[22]) );
  FA_4298 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_4297 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_4296 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_4295 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_4294 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_4293 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_4292 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_4291 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_4290 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_4289 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_4321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_4322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4328 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_4333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4344 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_139 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_4351 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_4350 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_4349 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_4348 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_4347 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_4346 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_4345 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_4344 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_4343 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_4342 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_4341 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_4340 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_4339 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_4338 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_4337 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_4336 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_4335 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_4334 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_4333 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_4332 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(1'b0), .S(S[20]), .CO(
        C[21]) );
  FA_4331 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_4330 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_4329 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_4328 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_4327 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_4326 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_4325 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_4324 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_4323 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_4322 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_4321 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_4353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_4354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4360 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_4366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4376 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_140 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_4383 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_4382 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_4381 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_4380 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_4379 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_4378 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_4377 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_4376 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_4375 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_4374 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_4373 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_4372 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_4371 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_4370 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_4369 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_4368 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_4367 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_4366 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_4365 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(1'b0), .S(S[19]), .CO(
        C[20]) );
  FA_4364 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_4363 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_4362 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_4361 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_4360 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_4359 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_4358 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_4357 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_4356 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_4355 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_4354 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_4353 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_4385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_4386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4392 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_4399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4408 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_141 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_4415 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_4414 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_4413 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_4412 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_4411 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_4410 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_4409 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_4408 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_4407 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_4406 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_4405 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_4404 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_4403 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_4402 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_4401 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_4400 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_4399 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_4398 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(1'b0), .S(S[18]), .CO(
        C[19]) );
  FA_4397 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_4396 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_4395 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_4394 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_4393 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_4392 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_4391 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_4390 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_4389 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_4388 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_4387 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_4386 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_4385 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_4417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_4418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4424 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_4432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4440 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_142 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_4447 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_4446 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_4445 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_4444 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_4443 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_4442 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_4441 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_4440 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_4439 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_4438 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_4437 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_4436 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_4435 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_4434 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_4433 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_4432 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_4431 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(1'b0), .S(S[17]), .CO(
        C[18]) );
  FA_4430 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_4429 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_4428 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_4427 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_4426 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_4425 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_4424 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_4423 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_4422 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_4421 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_4420 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_4419 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_4418 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_4417 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_4449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_4450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4456 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_4465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4472 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_143 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_4479 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_4478 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_4477 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_4476 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_4475 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_4474 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_4473 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_4472 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_4471 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_4470 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_4469 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_4468 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_4467 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_4466 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_4465 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_4464 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(1'b0), .S(S[16]), .CO(
        C[17]) );
  FA_4463 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_4462 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_4461 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_4460 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_4459 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_4458 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_4457 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_4456 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_4455 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_4454 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_4453 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_4452 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_4451 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_4450 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_4449 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_4481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_4482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4488 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_4498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4504 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_144 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_4511 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_4510 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_4509 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_4508 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_4507 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_4506 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_4505 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_4504 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_4503 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_4502 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_4501 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_4500 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_4499 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_4498 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_4497 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(1'b0), .S(S[15]), .CO(
        C[16]) );
  FA_4496 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_4495 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_4494 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_4493 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_4492 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_4491 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_4490 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_4489 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_4488 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_4487 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_4486 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_4485 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_4484 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_4483 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_4482 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_4481 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_4513 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_4514 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4515 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4516 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4517 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4518 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4519 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4520 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4521 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4522 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4523 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4524 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4525 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4526 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4527 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4528 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4529 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4530 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_4531 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4532 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4533 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4534 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4535 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4536 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4537 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4538 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4539 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4540 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4541 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4542 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4543 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_145 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_4543 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_4542 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_4541 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_4540 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_4539 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_4538 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_4537 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_4536 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_4535 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_4534 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_4533 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_4532 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_4531 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_4530 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(1'b0), .S(S[14]), .CO(
        C[15]) );
  FA_4529 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_4528 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_4527 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_4526 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_4525 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_4524 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_4523 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_4522 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_4521 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_4520 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_4519 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_4518 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_4517 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_4516 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_4515 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_4514 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_4513 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_4545 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_4546 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4547 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4548 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4549 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4550 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4551 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4552 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4553 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4554 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4555 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4556 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4557 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4558 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4559 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4560 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4561 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4562 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4563 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_4564 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4565 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4566 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4567 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4568 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4569 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4570 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4571 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4572 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4573 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4574 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4575 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_146 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_4575 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_4574 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_4573 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_4572 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_4571 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_4570 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_4569 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_4568 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_4567 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_4566 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_4565 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_4564 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_4563 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(1'b0), .S(S[13]), .CO(
        C[14]) );
  FA_4562 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_4561 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_4560 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_4559 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_4558 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_4557 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_4556 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_4555 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_4554 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_4553 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_4552 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_4551 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_4550 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_4549 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_4548 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_4547 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_4546 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_4545 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_4577 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_4578 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4579 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4580 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4581 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4582 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4583 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4584 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4585 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4586 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4587 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4588 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4589 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4590 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4591 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4592 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4593 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4594 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4595 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4596 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_4597 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4598 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4599 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4600 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4601 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4602 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4603 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4604 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4605 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4606 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4607 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_147 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_4607 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_4606 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_4605 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_4604 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_4603 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_4602 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_4601 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_4600 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_4599 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_4598 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_4597 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_4596 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(1'b0), .S(S[12]), .CO(
        C[13]) );
  FA_4595 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_4594 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_4593 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_4592 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_4591 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_4590 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_4589 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_4588 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_4587 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_4586 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_4585 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_4584 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_4583 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_4582 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_4581 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_4580 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_4579 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_4578 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_4577 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_4609 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_4610 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4611 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4612 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4613 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4614 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4615 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4616 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4617 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4618 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4619 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4620 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4621 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4622 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4623 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4624 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4625 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4626 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4627 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4628 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4629 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_4630 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4631 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4632 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4633 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4634 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4635 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4636 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4637 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4638 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4639 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_148 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_4639 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_4638 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_4637 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_4636 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_4635 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_4634 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_4633 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_4632 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_4631 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_4630 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_4629 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(1'b0), .S(S[11]), .CO(
        C[12]) );
  FA_4628 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_4627 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_4626 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_4625 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_4624 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_4623 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_4622 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_4621 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_4620 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_4619 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_4618 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_4617 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_4616 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_4615 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_4614 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_4613 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_4612 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_4611 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_4610 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_4609 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_4641 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_4642 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4643 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4644 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4645 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4646 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4647 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4648 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4649 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4650 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4651 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4652 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4653 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4654 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4655 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4656 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4657 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4658 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4659 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4660 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4661 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4662 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_4663 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4664 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4665 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4666 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4667 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4668 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4669 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4670 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4671 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_149 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_4671 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_4670 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_4669 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_4668 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_4667 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_4666 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_4665 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_4664 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_4663 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_4662 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(1'b0), .S(S[10]), .CO(
        C[11]) );
  FA_4661 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_4660 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_4659 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_4658 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_4657 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_4656 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_4655 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_4654 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_4653 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_4652 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_4651 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_4650 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_4649 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_4648 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_4647 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_4646 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_4645 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_4644 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_4643 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_4642 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_4641 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_4673 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_4674 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4675 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4676 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4677 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4678 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4679 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4680 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4681 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4682 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4683 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4684 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4685 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4686 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4687 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4688 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4689 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4690 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4691 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4692 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4693 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4694 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4695 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_4696 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4697 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4698 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4699 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4700 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4701 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4702 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4703 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_150 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_4703 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_4702 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_4701 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_4700 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_4699 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_4698 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_4697 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_4696 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_4695 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(1'b0), .S(S[9]), .CO(C[10]) );
  FA_4694 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_4693 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_4692 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_4691 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_4690 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_4689 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_4688 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_4687 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_4686 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_4685 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_4684 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_4683 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_4682 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_4681 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_4680 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_4679 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_4678 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_4677 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_4676 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_4675 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_4674 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_4673 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_4705 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_4706 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4707 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4708 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4709 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4710 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4711 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4712 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4713 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4714 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4715 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4716 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4717 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4718 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4719 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4720 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4721 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4722 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4723 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4724 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4725 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4726 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4727 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4728 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_4729 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4730 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4731 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4732 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4733 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4734 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4735 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_151 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_4735 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_4734 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_4733 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_4732 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_4731 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_4730 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_4729 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_4728 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(1'b0), .S(S[8]), .CO(C[9])
         );
  FA_4727 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_4726 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_4725 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_4724 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_4723 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_4722 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_4721 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_4720 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_4719 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_4718 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_4717 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_4716 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_4715 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_4714 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_4713 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_4712 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_4711 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_4710 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_4709 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_4708 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_4707 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_4706 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_4705 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_4737 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_4738 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4739 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4740 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4741 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4742 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4743 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4744 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4745 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4746 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4747 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4748 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4749 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4750 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4751 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4752 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4753 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4754 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4755 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4756 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4757 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4758 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4759 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4760 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4761 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_4762 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4763 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4764 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4765 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4766 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4767 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_152 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_4767 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_4766 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_4765 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_4764 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_4763 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_4762 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_4761 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(1'b0), .S(S[7]), .CO(C[8])
         );
  FA_4760 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_4759 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_4758 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_4757 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_4756 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_4755 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_4754 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_4753 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_4752 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_4751 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_4750 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_4749 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_4748 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_4747 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_4746 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_4745 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_4744 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_4743 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_4742 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_4741 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_4740 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_4739 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_4738 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_4737 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_4769 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_4770 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4771 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4772 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4773 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4774 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4775 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4776 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4777 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4778 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4779 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4780 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4781 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4782 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4783 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4784 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4785 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4786 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4787 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4788 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4789 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4790 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4791 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4792 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4793 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4794 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_4795 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4796 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4797 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4798 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4799 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_153 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_4799 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_4798 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_4797 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_4796 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_4795 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_4794 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(1'b0), .S(S[6]), .CO(C[7])
         );
  FA_4793 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_4792 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_4791 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_4790 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_4789 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_4788 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_4787 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_4786 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_4785 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_4784 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_4783 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_4782 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_4781 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_4780 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_4779 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_4778 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_4777 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_4776 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_4775 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_4774 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_4773 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_4772 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_4771 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_4770 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_4769 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_4801 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_4802 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4803 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4804 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4805 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4806 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4807 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4808 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4809 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4810 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4811 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4812 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4813 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4814 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4815 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4816 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4817 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4818 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4819 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4820 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4821 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4822 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4823 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4824 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4825 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4826 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4827 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_4828 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4829 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4830 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4831 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_154 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_4831 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_4830 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_4829 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_4828 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_4827 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(1'b0), .S(S[5]), .CO(C[6])
         );
  FA_4826 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_4825 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_4824 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_4823 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_4822 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_4821 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_4820 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_4819 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_4818 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_4817 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_4816 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_4815 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_4814 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_4813 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_4812 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_4811 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_4810 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_4809 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_4808 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_4807 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_4806 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_4805 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_4804 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_4803 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_4802 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_4801 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_4833 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_4834 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4835 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4836 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4837 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4838 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4839 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4840 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4841 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4842 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4843 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4844 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4845 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4846 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4847 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4848 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4849 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4850 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4851 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4852 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4853 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4854 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4855 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4856 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4857 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4858 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4859 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4860 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_4861 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4862 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4863 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_155 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_4863 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_4862 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_4861 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_4860 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(1'b0), .S(S[4]), .CO(C[5])
         );
  FA_4859 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_4858 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_4857 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_4856 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_4855 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_4854 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_4853 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_4852 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_4851 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_4850 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_4849 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_4848 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_4847 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_4846 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_4845 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_4844 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_4843 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_4842 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_4841 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_4840 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_4839 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_4838 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_4837 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_4836 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_4835 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_4834 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_4833 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_4865 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_4866 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4867 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4868 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4869 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4870 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4871 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4872 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4873 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4874 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4875 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4876 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4877 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4878 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4879 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4880 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4881 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4882 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4883 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4884 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4885 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4886 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4887 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4888 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4889 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4890 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4891 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4892 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4893 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_4894 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4895 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_156 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_4895 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_4894 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_4893 \FAINST[3].FA_  ( .A(A[3]), .B(B[3]), .CI(1'b0), .S(S[3]), .CO(C[4])
         );
  FA_4892 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_4891 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_4890 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_4889 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_4888 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_4887 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_4886 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_4885 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_4884 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_4883 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_4882 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_4881 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_4880 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_4879 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_4878 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_4877 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_4876 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_4875 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_4874 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_4873 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_4872 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_4871 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_4870 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_4869 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_4868 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_4867 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_4866 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_4865 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_4897 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_4898 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4899 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4900 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4901 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4902 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4903 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4904 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4905 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4906 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4907 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4908 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4909 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4910 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4911 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4912 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4913 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4914 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4915 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4916 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4917 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4918 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4919 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4920 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4921 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4922 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4923 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4924 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4925 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4926 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_4927 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_157 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_4927 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_4926 \FAINST[2].FA_  ( .A(A[2]), .B(B[2]), .CI(1'b0), .S(S[2]), .CO(C[3])
         );
  FA_4925 \FAINST[3].FA_  ( .A(A[3]), .B(B[3]), .CI(C[3]), .S(S[3]), .CO(C[4])
         );
  FA_4924 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_4923 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_4922 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_4921 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_4920 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_4919 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_4918 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_4917 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_4916 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_4915 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_4914 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_4913 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_4912 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_4911 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_4910 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_4909 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_4908 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_4907 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_4906 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_4905 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_4904 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_4903 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_4902 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_4901 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_4900 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_4899 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_4898 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_4897 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_4929 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_4930 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_4931 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_4932 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_4933 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_4934 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_4935 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_4936 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_4937 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_4938 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_4939 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_4940 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_4941 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_4942 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_4943 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_4944 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_4945 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_4946 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_4947 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_4948 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_4949 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_4950 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_4951 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_4952 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_4953 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_4954 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_4955 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_4956 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_4957 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_4958 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_4959 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module ADD_N32_158 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;


  FA_4959 \FAINST[1].FA_  ( .A(A[1]), .B(1'b0), .CI(1'b0), .S(S[1]) );
  FA_4958 \FAINST[2].FA_  ( .A(A[2]), .B(1'b0), .CI(1'b0), .S(S[2]) );
  FA_4957 \FAINST[3].FA_  ( .A(A[3]), .B(1'b0), .CI(1'b0), .S(S[3]) );
  FA_4956 \FAINST[4].FA_  ( .A(A[4]), .B(1'b0), .CI(1'b0), .S(S[4]) );
  FA_4955 \FAINST[5].FA_  ( .A(A[5]), .B(1'b0), .CI(1'b0), .S(S[5]) );
  FA_4954 \FAINST[6].FA_  ( .A(A[6]), .B(1'b0), .CI(1'b0), .S(S[6]) );
  FA_4953 \FAINST[7].FA_  ( .A(A[7]), .B(1'b0), .CI(1'b0), .S(S[7]) );
  FA_4952 \FAINST[8].FA_  ( .A(A[8]), .B(1'b0), .CI(1'b0), .S(S[8]) );
  FA_4951 \FAINST[9].FA_  ( .A(A[9]), .B(1'b0), .CI(1'b0), .S(S[9]) );
  FA_4950 \FAINST[10].FA_  ( .A(A[10]), .B(1'b0), .CI(1'b0), .S(S[10]) );
  FA_4949 \FAINST[11].FA_  ( .A(A[11]), .B(1'b0), .CI(1'b0), .S(S[11]) );
  FA_4948 \FAINST[12].FA_  ( .A(A[12]), .B(1'b0), .CI(1'b0), .S(S[12]) );
  FA_4947 \FAINST[13].FA_  ( .A(A[13]), .B(1'b0), .CI(1'b0), .S(S[13]) );
  FA_4946 \FAINST[14].FA_  ( .A(A[14]), .B(1'b0), .CI(1'b0), .S(S[14]) );
  FA_4945 \FAINST[15].FA_  ( .A(A[15]), .B(1'b0), .CI(1'b0), .S(S[15]) );
  FA_4944 \FAINST[16].FA_  ( .A(A[16]), .B(1'b0), .CI(1'b0), .S(S[16]) );
  FA_4943 \FAINST[17].FA_  ( .A(A[17]), .B(1'b0), .CI(1'b0), .S(S[17]) );
  FA_4942 \FAINST[18].FA_  ( .A(A[18]), .B(1'b0), .CI(1'b0), .S(S[18]) );
  FA_4941 \FAINST[19].FA_  ( .A(A[19]), .B(1'b0), .CI(1'b0), .S(S[19]) );
  FA_4940 \FAINST[20].FA_  ( .A(A[20]), .B(1'b0), .CI(1'b0), .S(S[20]) );
  FA_4939 \FAINST[21].FA_  ( .A(A[21]), .B(1'b0), .CI(1'b0), .S(S[21]) );
  FA_4938 \FAINST[22].FA_  ( .A(A[22]), .B(1'b0), .CI(1'b0), .S(S[22]) );
  FA_4937 \FAINST[23].FA_  ( .A(A[23]), .B(1'b0), .CI(1'b0), .S(S[23]) );
  FA_4936 \FAINST[24].FA_  ( .A(A[24]), .B(1'b0), .CI(1'b0), .S(S[24]) );
  FA_4935 \FAINST[25].FA_  ( .A(A[25]), .B(1'b0), .CI(1'b0), .S(S[25]) );
  FA_4934 \FAINST[26].FA_  ( .A(A[26]), .B(1'b0), .CI(1'b0), .S(S[26]) );
  FA_4933 \FAINST[27].FA_  ( .A(A[27]), .B(1'b0), .CI(1'b0), .S(S[27]) );
  FA_4932 \FAINST[28].FA_  ( .A(A[28]), .B(1'b0), .CI(1'b0), .S(S[28]) );
  FA_4931 \FAINST[29].FA_  ( .A(A[29]), .B(1'b0), .CI(1'b0), .S(S[29]) );
  FA_4930 \FAINST[30].FA_  ( .A(A[30]), .B(1'b0), .CI(1'b0), .S(S[30]) );
  FA_4929 \FAINST[31].FA_  ( .A(A[31]), .B(1'b0), .CI(1'b0), .S(S[31]) );
endmodule


module MULT_N32_5 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   \w[31][31] , \w[31][30] , \w[31][29] , \w[31][28] , \w[31][27] ,
         \w[31][26] , \w[31][25] , \w[31][24] , \w[31][23] , \w[31][22] ,
         \w[31][21] , \w[31][20] , \w[31][19] , \w[31][18] , \w[31][17] ,
         \w[31][16] , \w[31][15] , \w[31][14] , \w[31][13] , \w[31][12] ,
         \w[31][11] , \w[31][10] , \w[31][9] , \w[31][8] , \w[31][7] ,
         \w[31][6] , \w[31][5] , \w[31][4] , \w[31][3] , \w[31][2] ,
         \w[31][1] , \w[30][31] , \w[30][30] , \w[30][29] , \w[30][28] ,
         \w[30][27] , \w[30][26] , \w[30][25] , \w[30][24] , \w[30][23] ,
         \w[30][22] , \w[30][21] , \w[30][20] , \w[30][19] , \w[30][18] ,
         \w[30][17] , \w[30][16] , \w[30][15] , \w[30][14] , \w[30][13] ,
         \w[30][12] , \w[30][11] , \w[30][10] , \w[30][9] , \w[30][8] ,
         \w[30][7] , \w[30][6] , \w[30][5] , \w[30][4] , \w[30][3] ,
         \w[30][2] , \w[30][1] , \w[29][31] , \w[29][30] , \w[29][29] ,
         \w[29][28] , \w[29][27] , \w[29][26] , \w[29][25] , \w[29][24] ,
         \w[29][23] , \w[29][22] , \w[29][21] , \w[29][20] , \w[29][19] ,
         \w[29][18] , \w[29][17] , \w[29][16] , \w[29][15] , \w[29][14] ,
         \w[29][13] , \w[29][12] , \w[29][11] , \w[29][10] , \w[29][9] ,
         \w[29][8] , \w[29][7] , \w[29][6] , \w[29][5] , \w[29][4] ,
         \w[29][3] , \w[29][2] , \w[29][1] , \w[28][31] , \w[28][30] ,
         \w[28][29] , \w[28][28] , \w[28][27] , \w[28][26] , \w[28][25] ,
         \w[28][24] , \w[28][23] , \w[28][22] , \w[28][21] , \w[28][20] ,
         \w[28][19] , \w[28][18] , \w[28][17] , \w[28][16] , \w[28][15] ,
         \w[28][14] , \w[28][13] , \w[28][12] , \w[28][11] , \w[28][10] ,
         \w[28][9] , \w[28][8] , \w[28][7] , \w[28][6] , \w[28][5] ,
         \w[28][4] , \w[28][3] , \w[28][2] , \w[28][1] , \w[27][31] ,
         \w[27][30] , \w[27][29] , \w[27][28] , \w[27][27] , \w[27][26] ,
         \w[27][25] , \w[27][24] , \w[27][23] , \w[27][22] , \w[27][21] ,
         \w[27][20] , \w[27][19] , \w[27][18] , \w[27][17] , \w[27][16] ,
         \w[27][15] , \w[27][14] , \w[27][13] , \w[27][12] , \w[27][11] ,
         \w[27][10] , \w[27][9] , \w[27][8] , \w[27][7] , \w[27][6] ,
         \w[27][5] , \w[27][4] , \w[27][3] , \w[27][2] , \w[27][1] ,
         \w[26][31] , \w[26][30] , \w[26][29] , \w[26][28] , \w[26][27] ,
         \w[26][26] , \w[26][25] , \w[26][24] , \w[26][23] , \w[26][22] ,
         \w[26][21] , \w[26][20] , \w[26][19] , \w[26][18] , \w[26][17] ,
         \w[26][16] , \w[26][15] , \w[26][14] , \w[26][13] , \w[26][12] ,
         \w[26][11] , \w[26][10] , \w[26][9] , \w[26][8] , \w[26][7] ,
         \w[26][6] , \w[26][5] , \w[26][4] , \w[26][3] , \w[26][2] ,
         \w[26][1] , \w[25][31] , \w[25][30] , \w[25][29] , \w[25][28] ,
         \w[25][27] , \w[25][26] , \w[25][25] , \w[25][24] , \w[25][23] ,
         \w[25][22] , \w[25][21] , \w[25][20] , \w[25][19] , \w[25][18] ,
         \w[25][17] , \w[25][16] , \w[25][15] , \w[25][14] , \w[25][13] ,
         \w[25][12] , \w[25][11] , \w[25][10] , \w[25][9] , \w[25][8] ,
         \w[25][7] , \w[25][6] , \w[25][5] , \w[25][4] , \w[25][3] ,
         \w[25][2] , \w[25][1] , \w[24][31] , \w[24][30] , \w[24][29] ,
         \w[24][28] , \w[24][27] , \w[24][26] , \w[24][25] , \w[24][24] ,
         \w[24][23] , \w[24][22] , \w[24][21] , \w[24][20] , \w[24][19] ,
         \w[24][18] , \w[24][17] , \w[24][16] , \w[24][15] , \w[24][14] ,
         \w[24][13] , \w[24][12] , \w[24][11] , \w[24][10] , \w[24][9] ,
         \w[24][8] , \w[24][7] , \w[24][6] , \w[24][5] , \w[24][4] ,
         \w[24][3] , \w[24][2] , \w[24][1] , \w[23][31] , \w[23][30] ,
         \w[23][29] , \w[23][28] , \w[23][27] , \w[23][26] , \w[23][25] ,
         \w[23][24] , \w[23][23] , \w[23][22] , \w[23][21] , \w[23][20] ,
         \w[23][19] , \w[23][18] , \w[23][17] , \w[23][16] , \w[23][15] ,
         \w[23][14] , \w[23][13] , \w[23][12] , \w[23][11] , \w[23][10] ,
         \w[23][9] , \w[23][8] , \w[23][7] , \w[23][6] , \w[23][5] ,
         \w[23][4] , \w[23][3] , \w[23][2] , \w[23][1] , \w[22][31] ,
         \w[22][30] , \w[22][29] , \w[22][28] , \w[22][27] , \w[22][26] ,
         \w[22][25] , \w[22][24] , \w[22][23] , \w[22][22] , \w[22][21] ,
         \w[22][20] , \w[22][19] , \w[22][18] , \w[22][17] , \w[22][16] ,
         \w[22][15] , \w[22][14] , \w[22][13] , \w[22][12] , \w[22][11] ,
         \w[22][10] , \w[22][9] , \w[22][8] , \w[22][7] , \w[22][6] ,
         \w[22][5] , \w[22][4] , \w[22][3] , \w[22][2] , \w[22][1] ,
         \w[21][31] , \w[21][30] , \w[21][29] , \w[21][28] , \w[21][27] ,
         \w[21][26] , \w[21][25] , \w[21][24] , \w[21][23] , \w[21][22] ,
         \w[21][21] , \w[21][20] , \w[21][19] , \w[21][18] , \w[21][17] ,
         \w[21][16] , \w[21][15] , \w[21][14] , \w[21][13] , \w[21][12] ,
         \w[21][11] , \w[21][10] , \w[21][9] , \w[21][8] , \w[21][7] ,
         \w[21][6] , \w[21][5] , \w[21][4] , \w[21][3] , \w[21][2] ,
         \w[21][1] , \w[20][31] , \w[20][30] , \w[20][29] , \w[20][28] ,
         \w[20][27] , \w[20][26] , \w[20][25] , \w[20][24] , \w[20][23] ,
         \w[20][22] , \w[20][21] , \w[20][20] , \w[20][19] , \w[20][18] ,
         \w[20][17] , \w[20][16] , \w[20][15] , \w[20][14] , \w[20][13] ,
         \w[20][12] , \w[20][11] , \w[20][10] , \w[20][9] , \w[20][8] ,
         \w[20][7] , \w[20][6] , \w[20][5] , \w[20][4] , \w[20][3] ,
         \w[20][2] , \w[20][1] , \w[19][31] , \w[19][30] , \w[19][29] ,
         \w[19][28] , \w[19][27] , \w[19][26] , \w[19][25] , \w[19][24] ,
         \w[19][23] , \w[19][22] , \w[19][21] , \w[19][20] , \w[19][19] ,
         \w[19][18] , \w[19][17] , \w[19][16] , \w[19][15] , \w[19][14] ,
         \w[19][13] , \w[19][12] , \w[19][11] , \w[19][10] , \w[19][9] ,
         \w[19][8] , \w[19][7] , \w[19][6] , \w[19][5] , \w[19][4] ,
         \w[19][3] , \w[19][2] , \w[19][1] , \w[18][31] , \w[18][30] ,
         \w[18][29] , \w[18][28] , \w[18][27] , \w[18][26] , \w[18][25] ,
         \w[18][24] , \w[18][23] , \w[18][22] , \w[18][21] , \w[18][20] ,
         \w[18][19] , \w[18][18] , \w[18][17] , \w[18][16] , \w[18][15] ,
         \w[18][14] , \w[18][13] , \w[18][12] , \w[18][11] , \w[18][10] ,
         \w[18][9] , \w[18][8] , \w[18][7] , \w[18][6] , \w[18][5] ,
         \w[18][4] , \w[18][3] , \w[18][2] , \w[18][1] , \w[17][31] ,
         \w[17][30] , \w[17][29] , \w[17][28] , \w[17][27] , \w[17][26] ,
         \w[17][25] , \w[17][24] , \w[17][23] , \w[17][22] , \w[17][21] ,
         \w[17][20] , \w[17][19] , \w[17][18] , \w[17][17] , \w[17][16] ,
         \w[17][15] , \w[17][14] , \w[17][13] , \w[17][12] , \w[17][11] ,
         \w[17][10] , \w[17][9] , \w[17][8] , \w[17][7] , \w[17][6] ,
         \w[17][5] , \w[17][4] , \w[17][3] , \w[17][2] , \w[17][1] ,
         \w[16][31] , \w[16][30] , \w[16][29] , \w[16][28] , \w[16][27] ,
         \w[16][26] , \w[16][25] , \w[16][24] , \w[16][23] , \w[16][22] ,
         \w[16][21] , \w[16][20] , \w[16][19] , \w[16][18] , \w[16][17] ,
         \w[16][16] , \w[16][15] , \w[16][14] , \w[16][13] , \w[16][12] ,
         \w[16][11] , \w[16][10] , \w[16][9] , \w[16][8] , \w[16][7] ,
         \w[16][6] , \w[16][5] , \w[16][4] , \w[16][3] , \w[16][2] ,
         \w[16][1] , \w[15][31] , \w[15][30] , \w[15][29] , \w[15][28] ,
         \w[15][27] , \w[15][26] , \w[15][25] , \w[15][24] , \w[15][23] ,
         \w[15][22] , \w[15][21] , \w[15][20] , \w[15][19] , \w[15][18] ,
         \w[15][17] , \w[15][16] , \w[15][15] , \w[15][14] , \w[15][13] ,
         \w[15][12] , \w[15][11] , \w[15][10] , \w[15][9] , \w[15][8] ,
         \w[15][7] , \w[15][6] , \w[15][5] , \w[15][4] , \w[15][3] ,
         \w[15][2] , \w[15][1] , \w[14][31] , \w[14][30] , \w[14][29] ,
         \w[14][28] , \w[14][27] , \w[14][26] , \w[14][25] , \w[14][24] ,
         \w[14][23] , \w[14][22] , \w[14][21] , \w[14][20] , \w[14][19] ,
         \w[14][18] , \w[14][17] , \w[14][16] , \w[14][15] , \w[14][14] ,
         \w[14][13] , \w[14][12] , \w[14][11] , \w[14][10] , \w[14][9] ,
         \w[14][8] , \w[14][7] , \w[14][6] , \w[14][5] , \w[14][4] ,
         \w[14][3] , \w[14][2] , \w[14][1] , \w[13][31] , \w[13][30] ,
         \w[13][29] , \w[13][28] , \w[13][27] , \w[13][26] , \w[13][25] ,
         \w[13][24] , \w[13][23] , \w[13][22] , \w[13][21] , \w[13][20] ,
         \w[13][19] , \w[13][18] , \w[13][17] , \w[13][16] , \w[13][15] ,
         \w[13][14] , \w[13][13] , \w[13][12] , \w[13][11] , \w[13][10] ,
         \w[13][9] , \w[13][8] , \w[13][7] , \w[13][6] , \w[13][5] ,
         \w[13][4] , \w[13][3] , \w[13][2] , \w[13][1] , \w[12][31] ,
         \w[12][30] , \w[12][29] , \w[12][28] , \w[12][27] , \w[12][26] ,
         \w[12][25] , \w[12][24] , \w[12][23] , \w[12][22] , \w[12][21] ,
         \w[12][20] , \w[12][19] , \w[12][18] , \w[12][17] , \w[12][16] ,
         \w[12][15] , \w[12][14] , \w[12][13] , \w[12][12] , \w[12][11] ,
         \w[12][10] , \w[12][9] , \w[12][8] , \w[12][7] , \w[12][6] ,
         \w[12][5] , \w[12][4] , \w[12][3] , \w[12][2] , \w[12][1] ,
         \w[11][31] , \w[11][30] , \w[11][29] , \w[11][28] , \w[11][27] ,
         \w[11][26] , \w[11][25] , \w[11][24] , \w[11][23] , \w[11][22] ,
         \w[11][21] , \w[11][20] , \w[11][19] , \w[11][18] , \w[11][17] ,
         \w[11][16] , \w[11][15] , \w[11][14] , \w[11][13] , \w[11][12] ,
         \w[11][11] , \w[11][10] , \w[11][9] , \w[11][8] , \w[11][7] ,
         \w[11][6] , \w[11][5] , \w[11][4] , \w[11][3] , \w[11][2] ,
         \w[11][1] , \w[10][31] , \w[10][30] , \w[10][29] , \w[10][28] ,
         \w[10][27] , \w[10][26] , \w[10][25] , \w[10][24] , \w[10][23] ,
         \w[10][22] , \w[10][21] , \w[10][20] , \w[10][19] , \w[10][18] ,
         \w[10][17] , \w[10][16] , \w[10][15] , \w[10][14] , \w[10][13] ,
         \w[10][12] , \w[10][11] , \w[10][10] , \w[10][9] , \w[10][8] ,
         \w[10][7] , \w[10][6] , \w[10][5] , \w[10][4] , \w[10][3] ,
         \w[10][2] , \w[10][1] , \w[9][31] , \w[9][30] , \w[9][29] ,
         \w[9][28] , \w[9][27] , \w[9][26] , \w[9][25] , \w[9][24] ,
         \w[9][23] , \w[9][22] , \w[9][21] , \w[9][20] , \w[9][19] ,
         \w[9][18] , \w[9][17] , \w[9][16] , \w[9][15] , \w[9][14] ,
         \w[9][13] , \w[9][12] , \w[9][11] , \w[9][10] , \w[9][9] , \w[9][8] ,
         \w[9][7] , \w[9][6] , \w[9][5] , \w[9][4] , \w[9][3] , \w[9][2] ,
         \w[9][1] , \w[8][31] , \w[8][30] , \w[8][29] , \w[8][28] , \w[8][27] ,
         \w[8][26] , \w[8][25] , \w[8][24] , \w[8][23] , \w[8][22] ,
         \w[8][21] , \w[8][20] , \w[8][19] , \w[8][18] , \w[8][17] ,
         \w[8][16] , \w[8][15] , \w[8][14] , \w[8][13] , \w[8][12] ,
         \w[8][11] , \w[8][10] , \w[8][9] , \w[8][8] , \w[8][7] , \w[8][6] ,
         \w[8][5] , \w[8][4] , \w[8][3] , \w[8][2] , \w[8][1] , \w[7][31] ,
         \w[7][30] , \w[7][29] , \w[7][28] , \w[7][27] , \w[7][26] ,
         \w[7][25] , \w[7][24] , \w[7][23] , \w[7][22] , \w[7][21] ,
         \w[7][20] , \w[7][19] , \w[7][18] , \w[7][17] , \w[7][16] ,
         \w[7][15] , \w[7][14] , \w[7][13] , \w[7][12] , \w[7][11] ,
         \w[7][10] , \w[7][9] , \w[7][8] , \w[7][7] , \w[7][6] , \w[7][5] ,
         \w[7][4] , \w[7][3] , \w[7][2] , \w[7][1] , \w[6][31] , \w[6][30] ,
         \w[6][29] , \w[6][28] , \w[6][27] , \w[6][26] , \w[6][25] ,
         \w[6][24] , \w[6][23] , \w[6][22] , \w[6][21] , \w[6][20] ,
         \w[6][19] , \w[6][18] , \w[6][17] , \w[6][16] , \w[6][15] ,
         \w[6][14] , \w[6][13] , \w[6][12] , \w[6][11] , \w[6][10] , \w[6][9] ,
         \w[6][8] , \w[6][7] , \w[6][6] , \w[6][5] , \w[6][4] , \w[6][3] ,
         \w[6][2] , \w[6][1] , \w[5][31] , \w[5][30] , \w[5][29] , \w[5][28] ,
         \w[5][27] , \w[5][26] , \w[5][25] , \w[5][24] , \w[5][23] ,
         \w[5][22] , \w[5][21] , \w[5][20] , \w[5][19] , \w[5][18] ,
         \w[5][17] , \w[5][16] , \w[5][15] , \w[5][14] , \w[5][13] ,
         \w[5][12] , \w[5][11] , \w[5][10] , \w[5][9] , \w[5][8] , \w[5][7] ,
         \w[5][6] , \w[5][5] , \w[5][4] , \w[5][3] , \w[5][2] , \w[5][1] ,
         \w[4][31] , \w[4][30] , \w[4][29] , \w[4][28] , \w[4][27] ,
         \w[4][26] , \w[4][25] , \w[4][24] , \w[4][23] , \w[4][22] ,
         \w[4][21] , \w[4][20] , \w[4][19] , \w[4][18] , \w[4][17] ,
         \w[4][16] , \w[4][15] , \w[4][14] , \w[4][13] , \w[4][12] ,
         \w[4][11] , \w[4][10] , \w[4][9] , \w[4][8] , \w[4][7] , \w[4][6] ,
         \w[4][5] , \w[4][4] , \w[4][3] , \w[4][2] , \w[4][1] , \w[3][31] ,
         \w[3][30] , \w[3][29] , \w[3][28] , \w[3][27] , \w[3][26] ,
         \w[3][25] , \w[3][24] , \w[3][23] , \w[3][22] , \w[3][21] ,
         \w[3][20] , \w[3][19] , \w[3][18] , \w[3][17] , \w[3][16] ,
         \w[3][15] , \w[3][14] , \w[3][13] , \w[3][12] , \w[3][11] ,
         \w[3][10] , \w[3][9] , \w[3][8] , \w[3][7] , \w[3][6] , \w[3][5] ,
         \w[3][4] , \w[3][3] , \w[3][2] , \w[3][1] , \w[2][31] , \w[2][30] ,
         \w[2][29] , \w[2][28] , \w[2][27] , \w[2][26] , \w[2][25] ,
         \w[2][24] , \w[2][23] , \w[2][22] , \w[2][21] , \w[2][20] ,
         \w[2][19] , \w[2][18] , \w[2][17] , \w[2][16] , \w[2][15] ,
         \w[2][14] , \w[2][13] , \w[2][12] , \w[2][11] , \w[2][10] , \w[2][9] ,
         \w[2][8] , \w[2][7] , \w[2][6] , \w[2][5] , \w[2][4] , \w[2][3] ,
         \w[2][2] , \w[2][1] , \_0_net_[31] , \_0_net_[30] , \_0_net_[29] ,
         \_0_net_[28] , \_0_net_[27] , \_0_net_[26] , \_0_net_[25] ,
         \_0_net_[24] , \_0_net_[23] , \_0_net_[22] , \_0_net_[21] ,
         \_0_net_[20] , \_0_net_[19] , \_0_net_[18] , \_0_net_[17] ,
         \_0_net_[16] , \_0_net_[15] , \_0_net_[14] , \_0_net_[13] ,
         \_0_net_[12] , \_0_net_[11] , \_0_net_[10] , \_0_net_[9] ,
         \_0_net_[8] , \_0_net_[7] , \_0_net_[6] , \_0_net_[5] , \_0_net_[4] ,
         \_0_net_[3] , \_0_net_[2] , \_0_net_[1] , \_2_net_[31] ,
         \_2_net_[30] , \_2_net_[29] , \_2_net_[28] , \_2_net_[27] ,
         \_2_net_[26] , \_2_net_[25] , \_2_net_[24] , \_2_net_[23] ,
         \_2_net_[22] , \_2_net_[21] , \_2_net_[20] , \_2_net_[19] ,
         \_2_net_[18] , \_2_net_[17] , \_2_net_[16] , \_2_net_[15] ,
         \_2_net_[14] , \_2_net_[13] , \_2_net_[12] , \_2_net_[11] ,
         \_2_net_[10] , \_2_net_[9] , \_2_net_[8] , \_2_net_[7] , \_2_net_[6] ,
         \_2_net_[5] , \_2_net_[4] , \_2_net_[3] , \_2_net_[2] , \_4_net_[31] ,
         \_4_net_[30] , \_4_net_[29] , \_4_net_[28] , \_4_net_[27] ,
         \_4_net_[26] , \_4_net_[25] , \_4_net_[24] , \_4_net_[23] ,
         \_4_net_[22] , \_4_net_[21] , \_4_net_[20] , \_4_net_[19] ,
         \_4_net_[18] , \_4_net_[17] , \_4_net_[16] , \_4_net_[15] ,
         \_4_net_[14] , \_4_net_[13] , \_4_net_[12] , \_4_net_[11] ,
         \_4_net_[10] , \_4_net_[9] , \_4_net_[8] , \_4_net_[7] , \_4_net_[6] ,
         \_4_net_[5] , \_4_net_[4] , \_4_net_[3] , \_6_net_[31] ,
         \_6_net_[30] , \_6_net_[29] , \_6_net_[28] , \_6_net_[27] ,
         \_6_net_[26] , \_6_net_[25] , \_6_net_[24] , \_6_net_[23] ,
         \_6_net_[22] , \_6_net_[21] , \_6_net_[20] , \_6_net_[19] ,
         \_6_net_[18] , \_6_net_[17] , \_6_net_[16] , \_6_net_[15] ,
         \_6_net_[14] , \_6_net_[13] , \_6_net_[12] , \_6_net_[11] ,
         \_6_net_[10] , \_6_net_[9] , \_6_net_[8] , \_6_net_[7] , \_6_net_[6] ,
         \_6_net_[5] , \_6_net_[4] , \_8_net_[31] , \_8_net_[30] ,
         \_8_net_[29] , \_8_net_[28] , \_8_net_[27] , \_8_net_[26] ,
         \_8_net_[25] , \_8_net_[24] , \_8_net_[23] , \_8_net_[22] ,
         \_8_net_[21] , \_8_net_[20] , \_8_net_[19] , \_8_net_[18] ,
         \_8_net_[17] , \_8_net_[16] , \_8_net_[15] , \_8_net_[14] ,
         \_8_net_[13] , \_8_net_[12] , \_8_net_[11] , \_8_net_[10] ,
         \_8_net_[9] , \_8_net_[8] , \_8_net_[7] , \_8_net_[6] , \_8_net_[5] ,
         \_10_net_[31] , \_10_net_[30] , \_10_net_[29] , \_10_net_[28] ,
         \_10_net_[27] , \_10_net_[26] , \_10_net_[25] , \_10_net_[24] ,
         \_10_net_[23] , \_10_net_[22] , \_10_net_[21] , \_10_net_[20] ,
         \_10_net_[19] , \_10_net_[18] , \_10_net_[17] , \_10_net_[16] ,
         \_10_net_[15] , \_10_net_[14] , \_10_net_[13] , \_10_net_[12] ,
         \_10_net_[11] , \_10_net_[10] , \_10_net_[9] , \_10_net_[8] ,
         \_10_net_[7] , \_10_net_[6] , \_12_net_[31] , \_12_net_[30] ,
         \_12_net_[29] , \_12_net_[28] , \_12_net_[27] , \_12_net_[26] ,
         \_12_net_[25] , \_12_net_[24] , \_12_net_[23] , \_12_net_[22] ,
         \_12_net_[21] , \_12_net_[20] , \_12_net_[19] , \_12_net_[18] ,
         \_12_net_[17] , \_12_net_[16] , \_12_net_[15] , \_12_net_[14] ,
         \_12_net_[13] , \_12_net_[12] , \_12_net_[11] , \_12_net_[10] ,
         \_12_net_[9] , \_12_net_[8] , \_12_net_[7] , \_14_net_[31] ,
         \_14_net_[30] , \_14_net_[29] , \_14_net_[28] , \_14_net_[27] ,
         \_14_net_[26] , \_14_net_[25] , \_14_net_[24] , \_14_net_[23] ,
         \_14_net_[22] , \_14_net_[21] , \_14_net_[20] , \_14_net_[19] ,
         \_14_net_[18] , \_14_net_[17] , \_14_net_[16] , \_14_net_[15] ,
         \_14_net_[14] , \_14_net_[13] , \_14_net_[12] , \_14_net_[11] ,
         \_14_net_[10] , \_14_net_[9] , \_14_net_[8] , \_16_net_[31] ,
         \_16_net_[30] , \_16_net_[29] , \_16_net_[28] , \_16_net_[27] ,
         \_16_net_[26] , \_16_net_[25] , \_16_net_[24] , \_16_net_[23] ,
         \_16_net_[22] , \_16_net_[21] , \_16_net_[20] , \_16_net_[19] ,
         \_16_net_[18] , \_16_net_[17] , \_16_net_[16] , \_16_net_[15] ,
         \_16_net_[14] , \_16_net_[13] , \_16_net_[12] , \_16_net_[11] ,
         \_16_net_[10] , \_16_net_[9] , \_18_net_[31] , \_18_net_[30] ,
         \_18_net_[29] , \_18_net_[28] , \_18_net_[27] , \_18_net_[26] ,
         \_18_net_[25] , \_18_net_[24] , \_18_net_[23] , \_18_net_[22] ,
         \_18_net_[21] , \_18_net_[20] , \_18_net_[19] , \_18_net_[18] ,
         \_18_net_[17] , \_18_net_[16] , \_18_net_[15] , \_18_net_[14] ,
         \_18_net_[13] , \_18_net_[12] , \_18_net_[11] , \_18_net_[10] ,
         \_20_net_[31] , \_20_net_[30] , \_20_net_[29] , \_20_net_[28] ,
         \_20_net_[27] , \_20_net_[26] , \_20_net_[25] , \_20_net_[24] ,
         \_20_net_[23] , \_20_net_[22] , \_20_net_[21] , \_20_net_[20] ,
         \_20_net_[19] , \_20_net_[18] , \_20_net_[17] , \_20_net_[16] ,
         \_20_net_[15] , \_20_net_[14] , \_20_net_[13] , \_20_net_[12] ,
         \_20_net_[11] , \_22_net_[31] , \_22_net_[30] , \_22_net_[29] ,
         \_22_net_[28] , \_22_net_[27] , \_22_net_[26] , \_22_net_[25] ,
         \_22_net_[24] , \_22_net_[23] , \_22_net_[22] , \_22_net_[21] ,
         \_22_net_[20] , \_22_net_[19] , \_22_net_[18] , \_22_net_[17] ,
         \_22_net_[16] , \_22_net_[15] , \_22_net_[14] , \_22_net_[13] ,
         \_22_net_[12] , \_24_net_[31] , \_24_net_[30] , \_24_net_[29] ,
         \_24_net_[28] , \_24_net_[27] , \_24_net_[26] , \_24_net_[25] ,
         \_24_net_[24] , \_24_net_[23] , \_24_net_[22] , \_24_net_[21] ,
         \_24_net_[20] , \_24_net_[19] , \_24_net_[18] , \_24_net_[17] ,
         \_24_net_[16] , \_24_net_[15] , \_24_net_[14] , \_24_net_[13] ,
         \_26_net_[31] , \_26_net_[30] , \_26_net_[29] , \_26_net_[28] ,
         \_26_net_[27] , \_26_net_[26] , \_26_net_[25] , \_26_net_[24] ,
         \_26_net_[23] , \_26_net_[22] , \_26_net_[21] , \_26_net_[20] ,
         \_26_net_[19] , \_26_net_[18] , \_26_net_[17] , \_26_net_[16] ,
         \_26_net_[15] , \_26_net_[14] , \_28_net_[31] , \_28_net_[30] ,
         \_28_net_[29] , \_28_net_[28] , \_28_net_[27] , \_28_net_[26] ,
         \_28_net_[25] , \_28_net_[24] , \_28_net_[23] , \_28_net_[22] ,
         \_28_net_[21] , \_28_net_[20] , \_28_net_[19] , \_28_net_[18] ,
         \_28_net_[17] , \_28_net_[16] , \_28_net_[15] , \_30_net_[31] ,
         \_30_net_[30] , \_30_net_[29] , \_30_net_[28] , \_30_net_[27] ,
         \_30_net_[26] , \_30_net_[25] , \_30_net_[24] , \_30_net_[23] ,
         \_30_net_[22] , \_30_net_[21] , \_30_net_[20] , \_30_net_[19] ,
         \_30_net_[18] , \_30_net_[17] , \_30_net_[16] , \_32_net_[31] ,
         \_32_net_[30] , \_32_net_[29] , \_32_net_[28] , \_32_net_[27] ,
         \_32_net_[26] , \_32_net_[25] , \_32_net_[24] , \_32_net_[23] ,
         \_32_net_[22] , \_32_net_[21] , \_32_net_[20] , \_32_net_[19] ,
         \_32_net_[18] , \_32_net_[17] , \_34_net_[31] , \_34_net_[30] ,
         \_34_net_[29] , \_34_net_[28] , \_34_net_[27] , \_34_net_[26] ,
         \_34_net_[25] , \_34_net_[24] , \_34_net_[23] , \_34_net_[22] ,
         \_34_net_[21] , \_34_net_[20] , \_34_net_[19] , \_34_net_[18] ,
         \_36_net_[31] , \_36_net_[30] , \_36_net_[29] , \_36_net_[28] ,
         \_36_net_[27] , \_36_net_[26] , \_36_net_[25] , \_36_net_[24] ,
         \_36_net_[23] , \_36_net_[22] , \_36_net_[21] , \_36_net_[20] ,
         \_36_net_[19] , \_38_net_[31] , \_38_net_[30] , \_38_net_[29] ,
         \_38_net_[28] , \_38_net_[27] , \_38_net_[26] , \_38_net_[25] ,
         \_38_net_[24] , \_38_net_[23] , \_38_net_[22] , \_38_net_[21] ,
         \_38_net_[20] , \_40_net_[31] , \_40_net_[30] , \_40_net_[29] ,
         \_40_net_[28] , \_40_net_[27] , \_40_net_[26] , \_40_net_[25] ,
         \_40_net_[24] , \_40_net_[23] , \_40_net_[22] , \_40_net_[21] ,
         \_42_net_[31] , \_42_net_[30] , \_42_net_[29] , \_42_net_[28] ,
         \_42_net_[27] , \_42_net_[26] , \_42_net_[25] , \_42_net_[24] ,
         \_42_net_[23] , \_42_net_[22] , \_44_net_[31] , \_44_net_[30] ,
         \_44_net_[29] , \_44_net_[28] , \_44_net_[27] , \_44_net_[26] ,
         \_44_net_[25] , \_44_net_[24] , \_44_net_[23] , \_46_net_[31] ,
         \_46_net_[30] , \_46_net_[29] , \_46_net_[28] , \_46_net_[27] ,
         \_46_net_[26] , \_46_net_[25] , \_46_net_[24] , \_48_net_[31] ,
         \_48_net_[30] , \_48_net_[29] , \_48_net_[28] , \_48_net_[27] ,
         \_48_net_[26] , \_48_net_[25] , \_50_net_[31] , \_50_net_[30] ,
         \_50_net_[29] , \_50_net_[28] , \_50_net_[27] , \_50_net_[26] ,
         \_52_net_[31] , \_52_net_[30] , \_52_net_[29] , \_52_net_[28] ,
         \_52_net_[27] , \_54_net_[31] , \_54_net_[30] , \_54_net_[29] ,
         \_54_net_[28] , \_56_net_[31] , \_56_net_[30] , \_56_net_[29] ,
         \_58_net_[31] , \_58_net_[30] , \_60_net_[31] ;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30;

  ADD_N32_158 \FAINST[1].ADD_  ( .A({\_0_net_[31] , \_0_net_[30] , 
        \_0_net_[29] , \_0_net_[28] , \_0_net_[27] , \_0_net_[26] , 
        \_0_net_[25] , \_0_net_[24] , \_0_net_[23] , \_0_net_[22] , 
        \_0_net_[21] , \_0_net_[20] , \_0_net_[19] , \_0_net_[18] , 
        \_0_net_[17] , \_0_net_[16] , \_0_net_[15] , \_0_net_[14] , 
        \_0_net_[13] , \_0_net_[12] , \_0_net_[11] , \_0_net_[10] , 
        \_0_net_[9] , \_0_net_[8] , \_0_net_[7] , \_0_net_[6] , \_0_net_[5] , 
        \_0_net_[4] , \_0_net_[3] , \_0_net_[2] , \_0_net_[1] , 1'b0}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .S({
        \w[2][31] , \w[2][30] , \w[2][29] , \w[2][28] , \w[2][27] , \w[2][26] , 
        \w[2][25] , \w[2][24] , \w[2][23] , \w[2][22] , \w[2][21] , \w[2][20] , 
        \w[2][19] , \w[2][18] , \w[2][17] , \w[2][16] , \w[2][15] , \w[2][14] , 
        \w[2][13] , \w[2][12] , \w[2][11] , \w[2][10] , \w[2][9] , \w[2][8] , 
        \w[2][7] , \w[2][6] , \w[2][5] , \w[2][4] , \w[2][3] , \w[2][2] , 
        \w[2][1] , SYNOPSYS_UNCONNECTED__0}) );
  ADD_N32_157 \FAINST[2].ADD_  ( .A({\_2_net_[31] , \_2_net_[30] , 
        \_2_net_[29] , \_2_net_[28] , \_2_net_[27] , \_2_net_[26] , 
        \_2_net_[25] , \_2_net_[24] , \_2_net_[23] , \_2_net_[22] , 
        \_2_net_[21] , \_2_net_[20] , \_2_net_[19] , \_2_net_[18] , 
        \_2_net_[17] , \_2_net_[16] , \_2_net_[15] , \_2_net_[14] , 
        \_2_net_[13] , \_2_net_[12] , \_2_net_[11] , \_2_net_[10] , 
        \_2_net_[9] , \_2_net_[8] , \_2_net_[7] , \_2_net_[6] , \_2_net_[5] , 
        \_2_net_[4] , \_2_net_[3] , \_2_net_[2] , 1'b0, 1'b0}), .B({\w[2][31] , 
        \w[2][30] , \w[2][29] , \w[2][28] , \w[2][27] , \w[2][26] , \w[2][25] , 
        \w[2][24] , \w[2][23] , \w[2][22] , \w[2][21] , \w[2][20] , \w[2][19] , 
        \w[2][18] , \w[2][17] , \w[2][16] , \w[2][15] , \w[2][14] , \w[2][13] , 
        \w[2][12] , \w[2][11] , \w[2][10] , \w[2][9] , \w[2][8] , \w[2][7] , 
        \w[2][6] , \w[2][5] , \w[2][4] , \w[2][3] , \w[2][2] , \w[2][1] , 1'b0}), .CI(1'b0), .S({\w[3][31] , \w[3][30] , \w[3][29] , \w[3][28] , \w[3][27] , 
        \w[3][26] , \w[3][25] , \w[3][24] , \w[3][23] , \w[3][22] , \w[3][21] , 
        \w[3][20] , \w[3][19] , \w[3][18] , \w[3][17] , \w[3][16] , \w[3][15] , 
        \w[3][14] , \w[3][13] , \w[3][12] , \w[3][11] , \w[3][10] , \w[3][9] , 
        \w[3][8] , \w[3][7] , \w[3][6] , \w[3][5] , \w[3][4] , \w[3][3] , 
        \w[3][2] , \w[3][1] , SYNOPSYS_UNCONNECTED__1}) );
  ADD_N32_156 \FAINST[3].ADD_  ( .A({\_4_net_[31] , \_4_net_[30] , 
        \_4_net_[29] , \_4_net_[28] , \_4_net_[27] , \_4_net_[26] , 
        \_4_net_[25] , \_4_net_[24] , \_4_net_[23] , \_4_net_[22] , 
        \_4_net_[21] , \_4_net_[20] , \_4_net_[19] , \_4_net_[18] , 
        \_4_net_[17] , \_4_net_[16] , \_4_net_[15] , \_4_net_[14] , 
        \_4_net_[13] , \_4_net_[12] , \_4_net_[11] , \_4_net_[10] , 
        \_4_net_[9] , \_4_net_[8] , \_4_net_[7] , \_4_net_[6] , \_4_net_[5] , 
        \_4_net_[4] , \_4_net_[3] , 1'b0, 1'b0, 1'b0}), .B({\w[3][31] , 
        \w[3][30] , \w[3][29] , \w[3][28] , \w[3][27] , \w[3][26] , \w[3][25] , 
        \w[3][24] , \w[3][23] , \w[3][22] , \w[3][21] , \w[3][20] , \w[3][19] , 
        \w[3][18] , \w[3][17] , \w[3][16] , \w[3][15] , \w[3][14] , \w[3][13] , 
        \w[3][12] , \w[3][11] , \w[3][10] , \w[3][9] , \w[3][8] , \w[3][7] , 
        \w[3][6] , \w[3][5] , \w[3][4] , \w[3][3] , \w[3][2] , \w[3][1] , 1'b0}), .CI(1'b0), .S({\w[4][31] , \w[4][30] , \w[4][29] , \w[4][28] , \w[4][27] , 
        \w[4][26] , \w[4][25] , \w[4][24] , \w[4][23] , \w[4][22] , \w[4][21] , 
        \w[4][20] , \w[4][19] , \w[4][18] , \w[4][17] , \w[4][16] , \w[4][15] , 
        \w[4][14] , \w[4][13] , \w[4][12] , \w[4][11] , \w[4][10] , \w[4][9] , 
        \w[4][8] , \w[4][7] , \w[4][6] , \w[4][5] , \w[4][4] , \w[4][3] , 
        \w[4][2] , \w[4][1] , SYNOPSYS_UNCONNECTED__2}) );
  ADD_N32_155 \FAINST[4].ADD_  ( .A({\_6_net_[31] , \_6_net_[30] , 
        \_6_net_[29] , \_6_net_[28] , \_6_net_[27] , \_6_net_[26] , 
        \_6_net_[25] , \_6_net_[24] , \_6_net_[23] , \_6_net_[22] , 
        \_6_net_[21] , \_6_net_[20] , \_6_net_[19] , \_6_net_[18] , 
        \_6_net_[17] , \_6_net_[16] , \_6_net_[15] , \_6_net_[14] , 
        \_6_net_[13] , \_6_net_[12] , \_6_net_[11] , \_6_net_[10] , 
        \_6_net_[9] , \_6_net_[8] , \_6_net_[7] , \_6_net_[6] , \_6_net_[5] , 
        \_6_net_[4] , 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[4][31] , \w[4][30] , 
        \w[4][29] , \w[4][28] , \w[4][27] , \w[4][26] , \w[4][25] , \w[4][24] , 
        \w[4][23] , \w[4][22] , \w[4][21] , \w[4][20] , \w[4][19] , \w[4][18] , 
        \w[4][17] , \w[4][16] , \w[4][15] , \w[4][14] , \w[4][13] , \w[4][12] , 
        \w[4][11] , \w[4][10] , \w[4][9] , \w[4][8] , \w[4][7] , \w[4][6] , 
        \w[4][5] , \w[4][4] , \w[4][3] , \w[4][2] , \w[4][1] , 1'b0}), .CI(
        1'b0), .S({\w[5][31] , \w[5][30] , \w[5][29] , \w[5][28] , \w[5][27] , 
        \w[5][26] , \w[5][25] , \w[5][24] , \w[5][23] , \w[5][22] , \w[5][21] , 
        \w[5][20] , \w[5][19] , \w[5][18] , \w[5][17] , \w[5][16] , \w[5][15] , 
        \w[5][14] , \w[5][13] , \w[5][12] , \w[5][11] , \w[5][10] , \w[5][9] , 
        \w[5][8] , \w[5][7] , \w[5][6] , \w[5][5] , \w[5][4] , \w[5][3] , 
        \w[5][2] , \w[5][1] , SYNOPSYS_UNCONNECTED__3}) );
  ADD_N32_154 \FAINST[5].ADD_  ( .A({\_8_net_[31] , \_8_net_[30] , 
        \_8_net_[29] , \_8_net_[28] , \_8_net_[27] , \_8_net_[26] , 
        \_8_net_[25] , \_8_net_[24] , \_8_net_[23] , \_8_net_[22] , 
        \_8_net_[21] , \_8_net_[20] , \_8_net_[19] , \_8_net_[18] , 
        \_8_net_[17] , \_8_net_[16] , \_8_net_[15] , \_8_net_[14] , 
        \_8_net_[13] , \_8_net_[12] , \_8_net_[11] , \_8_net_[10] , 
        \_8_net_[9] , \_8_net_[8] , \_8_net_[7] , \_8_net_[6] , \_8_net_[5] , 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[5][31] , \w[5][30] , \w[5][29] , 
        \w[5][28] , \w[5][27] , \w[5][26] , \w[5][25] , \w[5][24] , \w[5][23] , 
        \w[5][22] , \w[5][21] , \w[5][20] , \w[5][19] , \w[5][18] , \w[5][17] , 
        \w[5][16] , \w[5][15] , \w[5][14] , \w[5][13] , \w[5][12] , \w[5][11] , 
        \w[5][10] , \w[5][9] , \w[5][8] , \w[5][7] , \w[5][6] , \w[5][5] , 
        \w[5][4] , \w[5][3] , \w[5][2] , \w[5][1] , 1'b0}), .CI(1'b0), .S({
        \w[6][31] , \w[6][30] , \w[6][29] , \w[6][28] , \w[6][27] , \w[6][26] , 
        \w[6][25] , \w[6][24] , \w[6][23] , \w[6][22] , \w[6][21] , \w[6][20] , 
        \w[6][19] , \w[6][18] , \w[6][17] , \w[6][16] , \w[6][15] , \w[6][14] , 
        \w[6][13] , \w[6][12] , \w[6][11] , \w[6][10] , \w[6][9] , \w[6][8] , 
        \w[6][7] , \w[6][6] , \w[6][5] , \w[6][4] , \w[6][3] , \w[6][2] , 
        \w[6][1] , SYNOPSYS_UNCONNECTED__4}) );
  ADD_N32_153 \FAINST[6].ADD_  ( .A({\_10_net_[31] , \_10_net_[30] , 
        \_10_net_[29] , \_10_net_[28] , \_10_net_[27] , \_10_net_[26] , 
        \_10_net_[25] , \_10_net_[24] , \_10_net_[23] , \_10_net_[22] , 
        \_10_net_[21] , \_10_net_[20] , \_10_net_[19] , \_10_net_[18] , 
        \_10_net_[17] , \_10_net_[16] , \_10_net_[15] , \_10_net_[14] , 
        \_10_net_[13] , \_10_net_[12] , \_10_net_[11] , \_10_net_[10] , 
        \_10_net_[9] , \_10_net_[8] , \_10_net_[7] , \_10_net_[6] , 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[6][31] , \w[6][30] , \w[6][29] , 
        \w[6][28] , \w[6][27] , \w[6][26] , \w[6][25] , \w[6][24] , \w[6][23] , 
        \w[6][22] , \w[6][21] , \w[6][20] , \w[6][19] , \w[6][18] , \w[6][17] , 
        \w[6][16] , \w[6][15] , \w[6][14] , \w[6][13] , \w[6][12] , \w[6][11] , 
        \w[6][10] , \w[6][9] , \w[6][8] , \w[6][7] , \w[6][6] , \w[6][5] , 
        \w[6][4] , \w[6][3] , \w[6][2] , \w[6][1] , 1'b0}), .CI(1'b0), .S({
        \w[7][31] , \w[7][30] , \w[7][29] , \w[7][28] , \w[7][27] , \w[7][26] , 
        \w[7][25] , \w[7][24] , \w[7][23] , \w[7][22] , \w[7][21] , \w[7][20] , 
        \w[7][19] , \w[7][18] , \w[7][17] , \w[7][16] , \w[7][15] , \w[7][14] , 
        \w[7][13] , \w[7][12] , \w[7][11] , \w[7][10] , \w[7][9] , \w[7][8] , 
        \w[7][7] , \w[7][6] , \w[7][5] , \w[7][4] , \w[7][3] , \w[7][2] , 
        \w[7][1] , SYNOPSYS_UNCONNECTED__5}) );
  ADD_N32_152 \FAINST[7].ADD_  ( .A({\_12_net_[31] , \_12_net_[30] , 
        \_12_net_[29] , \_12_net_[28] , \_12_net_[27] , \_12_net_[26] , 
        \_12_net_[25] , \_12_net_[24] , \_12_net_[23] , \_12_net_[22] , 
        \_12_net_[21] , \_12_net_[20] , \_12_net_[19] , \_12_net_[18] , 
        \_12_net_[17] , \_12_net_[16] , \_12_net_[15] , \_12_net_[14] , 
        \_12_net_[13] , \_12_net_[12] , \_12_net_[11] , \_12_net_[10] , 
        \_12_net_[9] , \_12_net_[8] , \_12_net_[7] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({\w[7][31] , \w[7][30] , \w[7][29] , \w[7][28] , 
        \w[7][27] , \w[7][26] , \w[7][25] , \w[7][24] , \w[7][23] , \w[7][22] , 
        \w[7][21] , \w[7][20] , \w[7][19] , \w[7][18] , \w[7][17] , \w[7][16] , 
        \w[7][15] , \w[7][14] , \w[7][13] , \w[7][12] , \w[7][11] , \w[7][10] , 
        \w[7][9] , \w[7][8] , \w[7][7] , \w[7][6] , \w[7][5] , \w[7][4] , 
        \w[7][3] , \w[7][2] , \w[7][1] , 1'b0}), .CI(1'b0), .S({\w[8][31] , 
        \w[8][30] , \w[8][29] , \w[8][28] , \w[8][27] , \w[8][26] , \w[8][25] , 
        \w[8][24] , \w[8][23] , \w[8][22] , \w[8][21] , \w[8][20] , \w[8][19] , 
        \w[8][18] , \w[8][17] , \w[8][16] , \w[8][15] , \w[8][14] , \w[8][13] , 
        \w[8][12] , \w[8][11] , \w[8][10] , \w[8][9] , \w[8][8] , \w[8][7] , 
        \w[8][6] , \w[8][5] , \w[8][4] , \w[8][3] , \w[8][2] , \w[8][1] , 
        SYNOPSYS_UNCONNECTED__6}) );
  ADD_N32_151 \FAINST[8].ADD_  ( .A({\_14_net_[31] , \_14_net_[30] , 
        \_14_net_[29] , \_14_net_[28] , \_14_net_[27] , \_14_net_[26] , 
        \_14_net_[25] , \_14_net_[24] , \_14_net_[23] , \_14_net_[22] , 
        \_14_net_[21] , \_14_net_[20] , \_14_net_[19] , \_14_net_[18] , 
        \_14_net_[17] , \_14_net_[16] , \_14_net_[15] , \_14_net_[14] , 
        \_14_net_[13] , \_14_net_[12] , \_14_net_[11] , \_14_net_[10] , 
        \_14_net_[9] , \_14_net_[8] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({\w[8][31] , \w[8][30] , \w[8][29] , \w[8][28] , \w[8][27] , 
        \w[8][26] , \w[8][25] , \w[8][24] , \w[8][23] , \w[8][22] , \w[8][21] , 
        \w[8][20] , \w[8][19] , \w[8][18] , \w[8][17] , \w[8][16] , \w[8][15] , 
        \w[8][14] , \w[8][13] , \w[8][12] , \w[8][11] , \w[8][10] , \w[8][9] , 
        \w[8][8] , \w[8][7] , \w[8][6] , \w[8][5] , \w[8][4] , \w[8][3] , 
        \w[8][2] , \w[8][1] , 1'b0}), .CI(1'b0), .S({\w[9][31] , \w[9][30] , 
        \w[9][29] , \w[9][28] , \w[9][27] , \w[9][26] , \w[9][25] , \w[9][24] , 
        \w[9][23] , \w[9][22] , \w[9][21] , \w[9][20] , \w[9][19] , \w[9][18] , 
        \w[9][17] , \w[9][16] , \w[9][15] , \w[9][14] , \w[9][13] , \w[9][12] , 
        \w[9][11] , \w[9][10] , \w[9][9] , \w[9][8] , \w[9][7] , \w[9][6] , 
        \w[9][5] , \w[9][4] , \w[9][3] , \w[9][2] , \w[9][1] , 
        SYNOPSYS_UNCONNECTED__7}) );
  ADD_N32_150 \FAINST[9].ADD_  ( .A({\_16_net_[31] , \_16_net_[30] , 
        \_16_net_[29] , \_16_net_[28] , \_16_net_[27] , \_16_net_[26] , 
        \_16_net_[25] , \_16_net_[24] , \_16_net_[23] , \_16_net_[22] , 
        \_16_net_[21] , \_16_net_[20] , \_16_net_[19] , \_16_net_[18] , 
        \_16_net_[17] , \_16_net_[16] , \_16_net_[15] , \_16_net_[14] , 
        \_16_net_[13] , \_16_net_[12] , \_16_net_[11] , \_16_net_[10] , 
        \_16_net_[9] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({\w[9][31] , \w[9][30] , \w[9][29] , \w[9][28] , \w[9][27] , 
        \w[9][26] , \w[9][25] , \w[9][24] , \w[9][23] , \w[9][22] , \w[9][21] , 
        \w[9][20] , \w[9][19] , \w[9][18] , \w[9][17] , \w[9][16] , \w[9][15] , 
        \w[9][14] , \w[9][13] , \w[9][12] , \w[9][11] , \w[9][10] , \w[9][9] , 
        \w[9][8] , \w[9][7] , \w[9][6] , \w[9][5] , \w[9][4] , \w[9][3] , 
        \w[9][2] , \w[9][1] , 1'b0}), .CI(1'b0), .S({\w[10][31] , \w[10][30] , 
        \w[10][29] , \w[10][28] , \w[10][27] , \w[10][26] , \w[10][25] , 
        \w[10][24] , \w[10][23] , \w[10][22] , \w[10][21] , \w[10][20] , 
        \w[10][19] , \w[10][18] , \w[10][17] , \w[10][16] , \w[10][15] , 
        \w[10][14] , \w[10][13] , \w[10][12] , \w[10][11] , \w[10][10] , 
        \w[10][9] , \w[10][8] , \w[10][7] , \w[10][6] , \w[10][5] , \w[10][4] , 
        \w[10][3] , \w[10][2] , \w[10][1] , SYNOPSYS_UNCONNECTED__8}) );
  ADD_N32_149 \FAINST[10].ADD_  ( .A({\_18_net_[31] , \_18_net_[30] , 
        \_18_net_[29] , \_18_net_[28] , \_18_net_[27] , \_18_net_[26] , 
        \_18_net_[25] , \_18_net_[24] , \_18_net_[23] , \_18_net_[22] , 
        \_18_net_[21] , \_18_net_[20] , \_18_net_[19] , \_18_net_[18] , 
        \_18_net_[17] , \_18_net_[16] , \_18_net_[15] , \_18_net_[14] , 
        \_18_net_[13] , \_18_net_[12] , \_18_net_[11] , \_18_net_[10] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[10][31] , \w[10][30] , \w[10][29] , \w[10][28] , \w[10][27] , 
        \w[10][26] , \w[10][25] , \w[10][24] , \w[10][23] , \w[10][22] , 
        \w[10][21] , \w[10][20] , \w[10][19] , \w[10][18] , \w[10][17] , 
        \w[10][16] , \w[10][15] , \w[10][14] , \w[10][13] , \w[10][12] , 
        \w[10][11] , \w[10][10] , \w[10][9] , \w[10][8] , \w[10][7] , 
        \w[10][6] , \w[10][5] , \w[10][4] , \w[10][3] , \w[10][2] , \w[10][1] , 
        1'b0}), .CI(1'b0), .S({\w[11][31] , \w[11][30] , \w[11][29] , 
        \w[11][28] , \w[11][27] , \w[11][26] , \w[11][25] , \w[11][24] , 
        \w[11][23] , \w[11][22] , \w[11][21] , \w[11][20] , \w[11][19] , 
        \w[11][18] , \w[11][17] , \w[11][16] , \w[11][15] , \w[11][14] , 
        \w[11][13] , \w[11][12] , \w[11][11] , \w[11][10] , \w[11][9] , 
        \w[11][8] , \w[11][7] , \w[11][6] , \w[11][5] , \w[11][4] , \w[11][3] , 
        \w[11][2] , \w[11][1] , SYNOPSYS_UNCONNECTED__9}) );
  ADD_N32_148 \FAINST[11].ADD_  ( .A({\_20_net_[31] , \_20_net_[30] , 
        \_20_net_[29] , \_20_net_[28] , \_20_net_[27] , \_20_net_[26] , 
        \_20_net_[25] , \_20_net_[24] , \_20_net_[23] , \_20_net_[22] , 
        \_20_net_[21] , \_20_net_[20] , \_20_net_[19] , \_20_net_[18] , 
        \_20_net_[17] , \_20_net_[16] , \_20_net_[15] , \_20_net_[14] , 
        \_20_net_[13] , \_20_net_[12] , \_20_net_[11] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[11][31] , 
        \w[11][30] , \w[11][29] , \w[11][28] , \w[11][27] , \w[11][26] , 
        \w[11][25] , \w[11][24] , \w[11][23] , \w[11][22] , \w[11][21] , 
        \w[11][20] , \w[11][19] , \w[11][18] , \w[11][17] , \w[11][16] , 
        \w[11][15] , \w[11][14] , \w[11][13] , \w[11][12] , \w[11][11] , 
        \w[11][10] , \w[11][9] , \w[11][8] , \w[11][7] , \w[11][6] , 
        \w[11][5] , \w[11][4] , \w[11][3] , \w[11][2] , \w[11][1] , 1'b0}), 
        .CI(1'b0), .S({\w[12][31] , \w[12][30] , \w[12][29] , \w[12][28] , 
        \w[12][27] , \w[12][26] , \w[12][25] , \w[12][24] , \w[12][23] , 
        \w[12][22] , \w[12][21] , \w[12][20] , \w[12][19] , \w[12][18] , 
        \w[12][17] , \w[12][16] , \w[12][15] , \w[12][14] , \w[12][13] , 
        \w[12][12] , \w[12][11] , \w[12][10] , \w[12][9] , \w[12][8] , 
        \w[12][7] , \w[12][6] , \w[12][5] , \w[12][4] , \w[12][3] , \w[12][2] , 
        \w[12][1] , SYNOPSYS_UNCONNECTED__10}) );
  ADD_N32_147 \FAINST[12].ADD_  ( .A({\_22_net_[31] , \_22_net_[30] , 
        \_22_net_[29] , \_22_net_[28] , \_22_net_[27] , \_22_net_[26] , 
        \_22_net_[25] , \_22_net_[24] , \_22_net_[23] , \_22_net_[22] , 
        \_22_net_[21] , \_22_net_[20] , \_22_net_[19] , \_22_net_[18] , 
        \_22_net_[17] , \_22_net_[16] , \_22_net_[15] , \_22_net_[14] , 
        \_22_net_[13] , \_22_net_[12] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[12][31] , \w[12][30] , 
        \w[12][29] , \w[12][28] , \w[12][27] , \w[12][26] , \w[12][25] , 
        \w[12][24] , \w[12][23] , \w[12][22] , \w[12][21] , \w[12][20] , 
        \w[12][19] , \w[12][18] , \w[12][17] , \w[12][16] , \w[12][15] , 
        \w[12][14] , \w[12][13] , \w[12][12] , \w[12][11] , \w[12][10] , 
        \w[12][9] , \w[12][8] , \w[12][7] , \w[12][6] , \w[12][5] , \w[12][4] , 
        \w[12][3] , \w[12][2] , \w[12][1] , 1'b0}), .CI(1'b0), .S({\w[13][31] , 
        \w[13][30] , \w[13][29] , \w[13][28] , \w[13][27] , \w[13][26] , 
        \w[13][25] , \w[13][24] , \w[13][23] , \w[13][22] , \w[13][21] , 
        \w[13][20] , \w[13][19] , \w[13][18] , \w[13][17] , \w[13][16] , 
        \w[13][15] , \w[13][14] , \w[13][13] , \w[13][12] , \w[13][11] , 
        \w[13][10] , \w[13][9] , \w[13][8] , \w[13][7] , \w[13][6] , 
        \w[13][5] , \w[13][4] , \w[13][3] , \w[13][2] , \w[13][1] , 
        SYNOPSYS_UNCONNECTED__11}) );
  ADD_N32_146 \FAINST[13].ADD_  ( .A({\_24_net_[31] , \_24_net_[30] , 
        \_24_net_[29] , \_24_net_[28] , \_24_net_[27] , \_24_net_[26] , 
        \_24_net_[25] , \_24_net_[24] , \_24_net_[23] , \_24_net_[22] , 
        \_24_net_[21] , \_24_net_[20] , \_24_net_[19] , \_24_net_[18] , 
        \_24_net_[17] , \_24_net_[16] , \_24_net_[15] , \_24_net_[14] , 
        \_24_net_[13] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[13][31] , \w[13][30] , \w[13][29] , 
        \w[13][28] , \w[13][27] , \w[13][26] , \w[13][25] , \w[13][24] , 
        \w[13][23] , \w[13][22] , \w[13][21] , \w[13][20] , \w[13][19] , 
        \w[13][18] , \w[13][17] , \w[13][16] , \w[13][15] , \w[13][14] , 
        \w[13][13] , \w[13][12] , \w[13][11] , \w[13][10] , \w[13][9] , 
        \w[13][8] , \w[13][7] , \w[13][6] , \w[13][5] , \w[13][4] , \w[13][3] , 
        \w[13][2] , \w[13][1] , 1'b0}), .CI(1'b0), .S({\w[14][31] , 
        \w[14][30] , \w[14][29] , \w[14][28] , \w[14][27] , \w[14][26] , 
        \w[14][25] , \w[14][24] , \w[14][23] , \w[14][22] , \w[14][21] , 
        \w[14][20] , \w[14][19] , \w[14][18] , \w[14][17] , \w[14][16] , 
        \w[14][15] , \w[14][14] , \w[14][13] , \w[14][12] , \w[14][11] , 
        \w[14][10] , \w[14][9] , \w[14][8] , \w[14][7] , \w[14][6] , 
        \w[14][5] , \w[14][4] , \w[14][3] , \w[14][2] , \w[14][1] , 
        SYNOPSYS_UNCONNECTED__12}) );
  ADD_N32_145 \FAINST[14].ADD_  ( .A({\_26_net_[31] , \_26_net_[30] , 
        \_26_net_[29] , \_26_net_[28] , \_26_net_[27] , \_26_net_[26] , 
        \_26_net_[25] , \_26_net_[24] , \_26_net_[23] , \_26_net_[22] , 
        \_26_net_[21] , \_26_net_[20] , \_26_net_[19] , \_26_net_[18] , 
        \_26_net_[17] , \_26_net_[16] , \_26_net_[15] , \_26_net_[14] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({\w[14][31] , \w[14][30] , \w[14][29] , \w[14][28] , 
        \w[14][27] , \w[14][26] , \w[14][25] , \w[14][24] , \w[14][23] , 
        \w[14][22] , \w[14][21] , \w[14][20] , \w[14][19] , \w[14][18] , 
        \w[14][17] , \w[14][16] , \w[14][15] , \w[14][14] , \w[14][13] , 
        \w[14][12] , \w[14][11] , \w[14][10] , \w[14][9] , \w[14][8] , 
        \w[14][7] , \w[14][6] , \w[14][5] , \w[14][4] , \w[14][3] , \w[14][2] , 
        \w[14][1] , 1'b0}), .CI(1'b0), .S({\w[15][31] , \w[15][30] , 
        \w[15][29] , \w[15][28] , \w[15][27] , \w[15][26] , \w[15][25] , 
        \w[15][24] , \w[15][23] , \w[15][22] , \w[15][21] , \w[15][20] , 
        \w[15][19] , \w[15][18] , \w[15][17] , \w[15][16] , \w[15][15] , 
        \w[15][14] , \w[15][13] , \w[15][12] , \w[15][11] , \w[15][10] , 
        \w[15][9] , \w[15][8] , \w[15][7] , \w[15][6] , \w[15][5] , \w[15][4] , 
        \w[15][3] , \w[15][2] , \w[15][1] , SYNOPSYS_UNCONNECTED__13}) );
  ADD_N32_144 \FAINST[15].ADD_  ( .A({\_28_net_[31] , \_28_net_[30] , 
        \_28_net_[29] , \_28_net_[28] , \_28_net_[27] , \_28_net_[26] , 
        \_28_net_[25] , \_28_net_[24] , \_28_net_[23] , \_28_net_[22] , 
        \_28_net_[21] , \_28_net_[20] , \_28_net_[19] , \_28_net_[18] , 
        \_28_net_[17] , \_28_net_[16] , \_28_net_[15] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({\w[15][31] , \w[15][30] , \w[15][29] , \w[15][28] , \w[15][27] , 
        \w[15][26] , \w[15][25] , \w[15][24] , \w[15][23] , \w[15][22] , 
        \w[15][21] , \w[15][20] , \w[15][19] , \w[15][18] , \w[15][17] , 
        \w[15][16] , \w[15][15] , \w[15][14] , \w[15][13] , \w[15][12] , 
        \w[15][11] , \w[15][10] , \w[15][9] , \w[15][8] , \w[15][7] , 
        \w[15][6] , \w[15][5] , \w[15][4] , \w[15][3] , \w[15][2] , \w[15][1] , 
        1'b0}), .CI(1'b0), .S({\w[16][31] , \w[16][30] , \w[16][29] , 
        \w[16][28] , \w[16][27] , \w[16][26] , \w[16][25] , \w[16][24] , 
        \w[16][23] , \w[16][22] , \w[16][21] , \w[16][20] , \w[16][19] , 
        \w[16][18] , \w[16][17] , \w[16][16] , \w[16][15] , \w[16][14] , 
        \w[16][13] , \w[16][12] , \w[16][11] , \w[16][10] , \w[16][9] , 
        \w[16][8] , \w[16][7] , \w[16][6] , \w[16][5] , \w[16][4] , \w[16][3] , 
        \w[16][2] , \w[16][1] , SYNOPSYS_UNCONNECTED__14}) );
  ADD_N32_143 \FAINST[16].ADD_  ( .A({\_30_net_[31] , \_30_net_[30] , 
        \_30_net_[29] , \_30_net_[28] , \_30_net_[27] , \_30_net_[26] , 
        \_30_net_[25] , \_30_net_[24] , \_30_net_[23] , \_30_net_[22] , 
        \_30_net_[21] , \_30_net_[20] , \_30_net_[19] , \_30_net_[18] , 
        \_30_net_[17] , \_30_net_[16] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[16][31] , \w[16][30] , \w[16][29] , \w[16][28] , \w[16][27] , 
        \w[16][26] , \w[16][25] , \w[16][24] , \w[16][23] , \w[16][22] , 
        \w[16][21] , \w[16][20] , \w[16][19] , \w[16][18] , \w[16][17] , 
        \w[16][16] , \w[16][15] , \w[16][14] , \w[16][13] , \w[16][12] , 
        \w[16][11] , \w[16][10] , \w[16][9] , \w[16][8] , \w[16][7] , 
        \w[16][6] , \w[16][5] , \w[16][4] , \w[16][3] , \w[16][2] , \w[16][1] , 
        1'b0}), .CI(1'b0), .S({\w[17][31] , \w[17][30] , \w[17][29] , 
        \w[17][28] , \w[17][27] , \w[17][26] , \w[17][25] , \w[17][24] , 
        \w[17][23] , \w[17][22] , \w[17][21] , \w[17][20] , \w[17][19] , 
        \w[17][18] , \w[17][17] , \w[17][16] , \w[17][15] , \w[17][14] , 
        \w[17][13] , \w[17][12] , \w[17][11] , \w[17][10] , \w[17][9] , 
        \w[17][8] , \w[17][7] , \w[17][6] , \w[17][5] , \w[17][4] , \w[17][3] , 
        \w[17][2] , \w[17][1] , SYNOPSYS_UNCONNECTED__15}) );
  ADD_N32_142 \FAINST[17].ADD_  ( .A({\_32_net_[31] , \_32_net_[30] , 
        \_32_net_[29] , \_32_net_[28] , \_32_net_[27] , \_32_net_[26] , 
        \_32_net_[25] , \_32_net_[24] , \_32_net_[23] , \_32_net_[22] , 
        \_32_net_[21] , \_32_net_[20] , \_32_net_[19] , \_32_net_[18] , 
        \_32_net_[17] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[17][31] , 
        \w[17][30] , \w[17][29] , \w[17][28] , \w[17][27] , \w[17][26] , 
        \w[17][25] , \w[17][24] , \w[17][23] , \w[17][22] , \w[17][21] , 
        \w[17][20] , \w[17][19] , \w[17][18] , \w[17][17] , \w[17][16] , 
        \w[17][15] , \w[17][14] , \w[17][13] , \w[17][12] , \w[17][11] , 
        \w[17][10] , \w[17][9] , \w[17][8] , \w[17][7] , \w[17][6] , 
        \w[17][5] , \w[17][4] , \w[17][3] , \w[17][2] , \w[17][1] , 1'b0}), 
        .CI(1'b0), .S({\w[18][31] , \w[18][30] , \w[18][29] , \w[18][28] , 
        \w[18][27] , \w[18][26] , \w[18][25] , \w[18][24] , \w[18][23] , 
        \w[18][22] , \w[18][21] , \w[18][20] , \w[18][19] , \w[18][18] , 
        \w[18][17] , \w[18][16] , \w[18][15] , \w[18][14] , \w[18][13] , 
        \w[18][12] , \w[18][11] , \w[18][10] , \w[18][9] , \w[18][8] , 
        \w[18][7] , \w[18][6] , \w[18][5] , \w[18][4] , \w[18][3] , \w[18][2] , 
        \w[18][1] , SYNOPSYS_UNCONNECTED__16}) );
  ADD_N32_141 \FAINST[18].ADD_  ( .A({\_34_net_[31] , \_34_net_[30] , 
        \_34_net_[29] , \_34_net_[28] , \_34_net_[27] , \_34_net_[26] , 
        \_34_net_[25] , \_34_net_[24] , \_34_net_[23] , \_34_net_[22] , 
        \_34_net_[21] , \_34_net_[20] , \_34_net_[19] , \_34_net_[18] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[18][31] , \w[18][30] , 
        \w[18][29] , \w[18][28] , \w[18][27] , \w[18][26] , \w[18][25] , 
        \w[18][24] , \w[18][23] , \w[18][22] , \w[18][21] , \w[18][20] , 
        \w[18][19] , \w[18][18] , \w[18][17] , \w[18][16] , \w[18][15] , 
        \w[18][14] , \w[18][13] , \w[18][12] , \w[18][11] , \w[18][10] , 
        \w[18][9] , \w[18][8] , \w[18][7] , \w[18][6] , \w[18][5] , \w[18][4] , 
        \w[18][3] , \w[18][2] , \w[18][1] , 1'b0}), .CI(1'b0), .S({\w[19][31] , 
        \w[19][30] , \w[19][29] , \w[19][28] , \w[19][27] , \w[19][26] , 
        \w[19][25] , \w[19][24] , \w[19][23] , \w[19][22] , \w[19][21] , 
        \w[19][20] , \w[19][19] , \w[19][18] , \w[19][17] , \w[19][16] , 
        \w[19][15] , \w[19][14] , \w[19][13] , \w[19][12] , \w[19][11] , 
        \w[19][10] , \w[19][9] , \w[19][8] , \w[19][7] , \w[19][6] , 
        \w[19][5] , \w[19][4] , \w[19][3] , \w[19][2] , \w[19][1] , 
        SYNOPSYS_UNCONNECTED__17}) );
  ADD_N32_140 \FAINST[19].ADD_  ( .A({\_36_net_[31] , \_36_net_[30] , 
        \_36_net_[29] , \_36_net_[28] , \_36_net_[27] , \_36_net_[26] , 
        \_36_net_[25] , \_36_net_[24] , \_36_net_[23] , \_36_net_[22] , 
        \_36_net_[21] , \_36_net_[20] , \_36_net_[19] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({\w[19][31] , \w[19][30] , \w[19][29] , 
        \w[19][28] , \w[19][27] , \w[19][26] , \w[19][25] , \w[19][24] , 
        \w[19][23] , \w[19][22] , \w[19][21] , \w[19][20] , \w[19][19] , 
        \w[19][18] , \w[19][17] , \w[19][16] , \w[19][15] , \w[19][14] , 
        \w[19][13] , \w[19][12] , \w[19][11] , \w[19][10] , \w[19][9] , 
        \w[19][8] , \w[19][7] , \w[19][6] , \w[19][5] , \w[19][4] , \w[19][3] , 
        \w[19][2] , \w[19][1] , 1'b0}), .CI(1'b0), .S({\w[20][31] , 
        \w[20][30] , \w[20][29] , \w[20][28] , \w[20][27] , \w[20][26] , 
        \w[20][25] , \w[20][24] , \w[20][23] , \w[20][22] , \w[20][21] , 
        \w[20][20] , \w[20][19] , \w[20][18] , \w[20][17] , \w[20][16] , 
        \w[20][15] , \w[20][14] , \w[20][13] , \w[20][12] , \w[20][11] , 
        \w[20][10] , \w[20][9] , \w[20][8] , \w[20][7] , \w[20][6] , 
        \w[20][5] , \w[20][4] , \w[20][3] , \w[20][2] , \w[20][1] , 
        SYNOPSYS_UNCONNECTED__18}) );
  ADD_N32_139 \FAINST[20].ADD_  ( .A({\_38_net_[31] , \_38_net_[30] , 
        \_38_net_[29] , \_38_net_[28] , \_38_net_[27] , \_38_net_[26] , 
        \_38_net_[25] , \_38_net_[24] , \_38_net_[23] , \_38_net_[22] , 
        \_38_net_[21] , \_38_net_[20] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .B({\w[20][31] , \w[20][30] , \w[20][29] , \w[20][28] , 
        \w[20][27] , \w[20][26] , \w[20][25] , \w[20][24] , \w[20][23] , 
        \w[20][22] , \w[20][21] , \w[20][20] , \w[20][19] , \w[20][18] , 
        \w[20][17] , \w[20][16] , \w[20][15] , \w[20][14] , \w[20][13] , 
        \w[20][12] , \w[20][11] , \w[20][10] , \w[20][9] , \w[20][8] , 
        \w[20][7] , \w[20][6] , \w[20][5] , \w[20][4] , \w[20][3] , \w[20][2] , 
        \w[20][1] , 1'b0}), .CI(1'b0), .S({\w[21][31] , \w[21][30] , 
        \w[21][29] , \w[21][28] , \w[21][27] , \w[21][26] , \w[21][25] , 
        \w[21][24] , \w[21][23] , \w[21][22] , \w[21][21] , \w[21][20] , 
        \w[21][19] , \w[21][18] , \w[21][17] , \w[21][16] , \w[21][15] , 
        \w[21][14] , \w[21][13] , \w[21][12] , \w[21][11] , \w[21][10] , 
        \w[21][9] , \w[21][8] , \w[21][7] , \w[21][6] , \w[21][5] , \w[21][4] , 
        \w[21][3] , \w[21][2] , \w[21][1] , SYNOPSYS_UNCONNECTED__19}) );
  ADD_N32_138 \FAINST[21].ADD_  ( .A({\_40_net_[31] , \_40_net_[30] , 
        \_40_net_[29] , \_40_net_[28] , \_40_net_[27] , \_40_net_[26] , 
        \_40_net_[25] , \_40_net_[24] , \_40_net_[23] , \_40_net_[22] , 
        \_40_net_[21] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[21][31] , \w[21][30] , \w[21][29] , \w[21][28] , \w[21][27] , 
        \w[21][26] , \w[21][25] , \w[21][24] , \w[21][23] , \w[21][22] , 
        \w[21][21] , \w[21][20] , \w[21][19] , \w[21][18] , \w[21][17] , 
        \w[21][16] , \w[21][15] , \w[21][14] , \w[21][13] , \w[21][12] , 
        \w[21][11] , \w[21][10] , \w[21][9] , \w[21][8] , \w[21][7] , 
        \w[21][6] , \w[21][5] , \w[21][4] , \w[21][3] , \w[21][2] , \w[21][1] , 
        1'b0}), .CI(1'b0), .S({\w[22][31] , \w[22][30] , \w[22][29] , 
        \w[22][28] , \w[22][27] , \w[22][26] , \w[22][25] , \w[22][24] , 
        \w[22][23] , \w[22][22] , \w[22][21] , \w[22][20] , \w[22][19] , 
        \w[22][18] , \w[22][17] , \w[22][16] , \w[22][15] , \w[22][14] , 
        \w[22][13] , \w[22][12] , \w[22][11] , \w[22][10] , \w[22][9] , 
        \w[22][8] , \w[22][7] , \w[22][6] , \w[22][5] , \w[22][4] , \w[22][3] , 
        \w[22][2] , \w[22][1] , SYNOPSYS_UNCONNECTED__20}) );
  ADD_N32_137 \FAINST[22].ADD_  ( .A({\_42_net_[31] , \_42_net_[30] , 
        \_42_net_[29] , \_42_net_[28] , \_42_net_[27] , \_42_net_[26] , 
        \_42_net_[25] , \_42_net_[24] , \_42_net_[23] , \_42_net_[22] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[22][31] , \w[22][30] , \w[22][29] , \w[22][28] , \w[22][27] , 
        \w[22][26] , \w[22][25] , \w[22][24] , \w[22][23] , \w[22][22] , 
        \w[22][21] , \w[22][20] , \w[22][19] , \w[22][18] , \w[22][17] , 
        \w[22][16] , \w[22][15] , \w[22][14] , \w[22][13] , \w[22][12] , 
        \w[22][11] , \w[22][10] , \w[22][9] , \w[22][8] , \w[22][7] , 
        \w[22][6] , \w[22][5] , \w[22][4] , \w[22][3] , \w[22][2] , \w[22][1] , 
        1'b0}), .CI(1'b0), .S({\w[23][31] , \w[23][30] , \w[23][29] , 
        \w[23][28] , \w[23][27] , \w[23][26] , \w[23][25] , \w[23][24] , 
        \w[23][23] , \w[23][22] , \w[23][21] , \w[23][20] , \w[23][19] , 
        \w[23][18] , \w[23][17] , \w[23][16] , \w[23][15] , \w[23][14] , 
        \w[23][13] , \w[23][12] , \w[23][11] , \w[23][10] , \w[23][9] , 
        \w[23][8] , \w[23][7] , \w[23][6] , \w[23][5] , \w[23][4] , \w[23][3] , 
        \w[23][2] , \w[23][1] , SYNOPSYS_UNCONNECTED__21}) );
  ADD_N32_136 \FAINST[23].ADD_  ( .A({\_44_net_[31] , \_44_net_[30] , 
        \_44_net_[29] , \_44_net_[28] , \_44_net_[27] , \_44_net_[26] , 
        \_44_net_[25] , \_44_net_[24] , \_44_net_[23] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[23][31] , 
        \w[23][30] , \w[23][29] , \w[23][28] , \w[23][27] , \w[23][26] , 
        \w[23][25] , \w[23][24] , \w[23][23] , \w[23][22] , \w[23][21] , 
        \w[23][20] , \w[23][19] , \w[23][18] , \w[23][17] , \w[23][16] , 
        \w[23][15] , \w[23][14] , \w[23][13] , \w[23][12] , \w[23][11] , 
        \w[23][10] , \w[23][9] , \w[23][8] , \w[23][7] , \w[23][6] , 
        \w[23][5] , \w[23][4] , \w[23][3] , \w[23][2] , \w[23][1] , 1'b0}), 
        .CI(1'b0), .S({\w[24][31] , \w[24][30] , \w[24][29] , \w[24][28] , 
        \w[24][27] , \w[24][26] , \w[24][25] , \w[24][24] , \w[24][23] , 
        \w[24][22] , \w[24][21] , \w[24][20] , \w[24][19] , \w[24][18] , 
        \w[24][17] , \w[24][16] , \w[24][15] , \w[24][14] , \w[24][13] , 
        \w[24][12] , \w[24][11] , \w[24][10] , \w[24][9] , \w[24][8] , 
        \w[24][7] , \w[24][6] , \w[24][5] , \w[24][4] , \w[24][3] , \w[24][2] , 
        \w[24][1] , SYNOPSYS_UNCONNECTED__22}) );
  ADD_N32_135 \FAINST[24].ADD_  ( .A({\_46_net_[31] , \_46_net_[30] , 
        \_46_net_[29] , \_46_net_[28] , \_46_net_[27] , \_46_net_[26] , 
        \_46_net_[25] , \_46_net_[24] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[24][31] , \w[24][30] , 
        \w[24][29] , \w[24][28] , \w[24][27] , \w[24][26] , \w[24][25] , 
        \w[24][24] , \w[24][23] , \w[24][22] , \w[24][21] , \w[24][20] , 
        \w[24][19] , \w[24][18] , \w[24][17] , \w[24][16] , \w[24][15] , 
        \w[24][14] , \w[24][13] , \w[24][12] , \w[24][11] , \w[24][10] , 
        \w[24][9] , \w[24][8] , \w[24][7] , \w[24][6] , \w[24][5] , \w[24][4] , 
        \w[24][3] , \w[24][2] , \w[24][1] , 1'b0}), .CI(1'b0), .S({\w[25][31] , 
        \w[25][30] , \w[25][29] , \w[25][28] , \w[25][27] , \w[25][26] , 
        \w[25][25] , \w[25][24] , \w[25][23] , \w[25][22] , \w[25][21] , 
        \w[25][20] , \w[25][19] , \w[25][18] , \w[25][17] , \w[25][16] , 
        \w[25][15] , \w[25][14] , \w[25][13] , \w[25][12] , \w[25][11] , 
        \w[25][10] , \w[25][9] , \w[25][8] , \w[25][7] , \w[25][6] , 
        \w[25][5] , \w[25][4] , \w[25][3] , \w[25][2] , \w[25][1] , 
        SYNOPSYS_UNCONNECTED__23}) );
  ADD_N32_134 \FAINST[25].ADD_  ( .A({\_48_net_[31] , \_48_net_[30] , 
        \_48_net_[29] , \_48_net_[28] , \_48_net_[27] , \_48_net_[26] , 
        \_48_net_[25] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[25][31] , \w[25][30] , \w[25][29] , 
        \w[25][28] , \w[25][27] , \w[25][26] , \w[25][25] , \w[25][24] , 
        \w[25][23] , \w[25][22] , \w[25][21] , \w[25][20] , \w[25][19] , 
        \w[25][18] , \w[25][17] , \w[25][16] , \w[25][15] , \w[25][14] , 
        \w[25][13] , \w[25][12] , \w[25][11] , \w[25][10] , \w[25][9] , 
        \w[25][8] , \w[25][7] , \w[25][6] , \w[25][5] , \w[25][4] , \w[25][3] , 
        \w[25][2] , \w[25][1] , 1'b0}), .CI(1'b0), .S({\w[26][31] , 
        \w[26][30] , \w[26][29] , \w[26][28] , \w[26][27] , \w[26][26] , 
        \w[26][25] , \w[26][24] , \w[26][23] , \w[26][22] , \w[26][21] , 
        \w[26][20] , \w[26][19] , \w[26][18] , \w[26][17] , \w[26][16] , 
        \w[26][15] , \w[26][14] , \w[26][13] , \w[26][12] , \w[26][11] , 
        \w[26][10] , \w[26][9] , \w[26][8] , \w[26][7] , \w[26][6] , 
        \w[26][5] , \w[26][4] , \w[26][3] , \w[26][2] , \w[26][1] , 
        SYNOPSYS_UNCONNECTED__24}) );
  ADD_N32_133 \FAINST[26].ADD_  ( .A({\_50_net_[31] , \_50_net_[30] , 
        \_50_net_[29] , \_50_net_[28] , \_50_net_[27] , \_50_net_[26] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({\w[26][31] , \w[26][30] , \w[26][29] , \w[26][28] , 
        \w[26][27] , \w[26][26] , \w[26][25] , \w[26][24] , \w[26][23] , 
        \w[26][22] , \w[26][21] , \w[26][20] , \w[26][19] , \w[26][18] , 
        \w[26][17] , \w[26][16] , \w[26][15] , \w[26][14] , \w[26][13] , 
        \w[26][12] , \w[26][11] , \w[26][10] , \w[26][9] , \w[26][8] , 
        \w[26][7] , \w[26][6] , \w[26][5] , \w[26][4] , \w[26][3] , \w[26][2] , 
        \w[26][1] , 1'b0}), .CI(1'b0), .S({\w[27][31] , \w[27][30] , 
        \w[27][29] , \w[27][28] , \w[27][27] , \w[27][26] , \w[27][25] , 
        \w[27][24] , \w[27][23] , \w[27][22] , \w[27][21] , \w[27][20] , 
        \w[27][19] , \w[27][18] , \w[27][17] , \w[27][16] , \w[27][15] , 
        \w[27][14] , \w[27][13] , \w[27][12] , \w[27][11] , \w[27][10] , 
        \w[27][9] , \w[27][8] , \w[27][7] , \w[27][6] , \w[27][5] , \w[27][4] , 
        \w[27][3] , \w[27][2] , \w[27][1] , SYNOPSYS_UNCONNECTED__25}) );
  ADD_N32_132 \FAINST[27].ADD_  ( .A({\_52_net_[31] , \_52_net_[30] , 
        \_52_net_[29] , \_52_net_[28] , \_52_net_[27] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({\w[27][31] , \w[27][30] , \w[27][29] , \w[27][28] , \w[27][27] , 
        \w[27][26] , \w[27][25] , \w[27][24] , \w[27][23] , \w[27][22] , 
        \w[27][21] , \w[27][20] , \w[27][19] , \w[27][18] , \w[27][17] , 
        \w[27][16] , \w[27][15] , \w[27][14] , \w[27][13] , \w[27][12] , 
        \w[27][11] , \w[27][10] , \w[27][9] , \w[27][8] , \w[27][7] , 
        \w[27][6] , \w[27][5] , \w[27][4] , \w[27][3] , \w[27][2] , \w[27][1] , 
        1'b0}), .CI(1'b0), .S({\w[28][31] , \w[28][30] , \w[28][29] , 
        \w[28][28] , \w[28][27] , \w[28][26] , \w[28][25] , \w[28][24] , 
        \w[28][23] , \w[28][22] , \w[28][21] , \w[28][20] , \w[28][19] , 
        \w[28][18] , \w[28][17] , \w[28][16] , \w[28][15] , \w[28][14] , 
        \w[28][13] , \w[28][12] , \w[28][11] , \w[28][10] , \w[28][9] , 
        \w[28][8] , \w[28][7] , \w[28][6] , \w[28][5] , \w[28][4] , \w[28][3] , 
        \w[28][2] , \w[28][1] , SYNOPSYS_UNCONNECTED__26}) );
  ADD_N32_131 \FAINST[28].ADD_  ( .A({\_54_net_[31] , \_54_net_[30] , 
        \_54_net_[29] , \_54_net_[28] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[28][31] , \w[28][30] , \w[28][29] , \w[28][28] , \w[28][27] , 
        \w[28][26] , \w[28][25] , \w[28][24] , \w[28][23] , \w[28][22] , 
        \w[28][21] , \w[28][20] , \w[28][19] , \w[28][18] , \w[28][17] , 
        \w[28][16] , \w[28][15] , \w[28][14] , \w[28][13] , \w[28][12] , 
        \w[28][11] , \w[28][10] , \w[28][9] , \w[28][8] , \w[28][7] , 
        \w[28][6] , \w[28][5] , \w[28][4] , \w[28][3] , \w[28][2] , \w[28][1] , 
        1'b0}), .CI(1'b0), .S({\w[29][31] , \w[29][30] , \w[29][29] , 
        \w[29][28] , \w[29][27] , \w[29][26] , \w[29][25] , \w[29][24] , 
        \w[29][23] , \w[29][22] , \w[29][21] , \w[29][20] , \w[29][19] , 
        \w[29][18] , \w[29][17] , \w[29][16] , \w[29][15] , \w[29][14] , 
        \w[29][13] , \w[29][12] , \w[29][11] , \w[29][10] , \w[29][9] , 
        \w[29][8] , \w[29][7] , \w[29][6] , \w[29][5] , \w[29][4] , \w[29][3] , 
        \w[29][2] , \w[29][1] , SYNOPSYS_UNCONNECTED__27}) );
  ADD_N32_130 \FAINST[29].ADD_  ( .A({\_56_net_[31] , \_56_net_[30] , 
        \_56_net_[29] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[29][31] , 
        \w[29][30] , \w[29][29] , \w[29][28] , \w[29][27] , \w[29][26] , 
        \w[29][25] , \w[29][24] , \w[29][23] , \w[29][22] , \w[29][21] , 
        \w[29][20] , \w[29][19] , \w[29][18] , \w[29][17] , \w[29][16] , 
        \w[29][15] , \w[29][14] , \w[29][13] , \w[29][12] , \w[29][11] , 
        \w[29][10] , \w[29][9] , \w[29][8] , \w[29][7] , \w[29][6] , 
        \w[29][5] , \w[29][4] , \w[29][3] , \w[29][2] , \w[29][1] , 1'b0}), 
        .CI(1'b0), .S({\w[30][31] , \w[30][30] , \w[30][29] , \w[30][28] , 
        \w[30][27] , \w[30][26] , \w[30][25] , \w[30][24] , \w[30][23] , 
        \w[30][22] , \w[30][21] , \w[30][20] , \w[30][19] , \w[30][18] , 
        \w[30][17] , \w[30][16] , \w[30][15] , \w[30][14] , \w[30][13] , 
        \w[30][12] , \w[30][11] , \w[30][10] , \w[30][9] , \w[30][8] , 
        \w[30][7] , \w[30][6] , \w[30][5] , \w[30][4] , \w[30][3] , \w[30][2] , 
        \w[30][1] , SYNOPSYS_UNCONNECTED__28}) );
  ADD_N32_129 \FAINST[30].ADD_  ( .A({\_58_net_[31] , \_58_net_[30] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[30][31] , \w[30][30] , 
        \w[30][29] , \w[30][28] , \w[30][27] , \w[30][26] , \w[30][25] , 
        \w[30][24] , \w[30][23] , \w[30][22] , \w[30][21] , \w[30][20] , 
        \w[30][19] , \w[30][18] , \w[30][17] , \w[30][16] , \w[30][15] , 
        \w[30][14] , \w[30][13] , \w[30][12] , \w[30][11] , \w[30][10] , 
        \w[30][9] , \w[30][8] , \w[30][7] , \w[30][6] , \w[30][5] , \w[30][4] , 
        \w[30][3] , \w[30][2] , \w[30][1] , 1'b0}), .CI(1'b0), .S({\w[31][31] , 
        \w[31][30] , \w[31][29] , \w[31][28] , \w[31][27] , \w[31][26] , 
        \w[31][25] , \w[31][24] , \w[31][23] , \w[31][22] , \w[31][21] , 
        \w[31][20] , \w[31][19] , \w[31][18] , \w[31][17] , \w[31][16] , 
        \w[31][15] , \w[31][14] , \w[31][13] , \w[31][12] , \w[31][11] , 
        \w[31][10] , \w[31][9] , \w[31][8] , \w[31][7] , \w[31][6] , 
        \w[31][5] , \w[31][4] , \w[31][3] , \w[31][2] , \w[31][1] , 
        SYNOPSYS_UNCONNECTED__29}) );
  ADD_N32_128 \FAINST[31].ADD_  ( .A({\_60_net_[31] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({\w[31][31] , \w[31][30] , \w[31][29] , 
        \w[31][28] , \w[31][27] , \w[31][26] , \w[31][25] , \w[31][24] , 
        \w[31][23] , \w[31][22] , \w[31][21] , \w[31][20] , \w[31][19] , 
        \w[31][18] , \w[31][17] , \w[31][16] , \w[31][15] , \w[31][14] , 
        \w[31][13] , \w[31][12] , \w[31][11] , \w[31][10] , \w[31][9] , 
        \w[31][8] , \w[31][7] , \w[31][6] , \w[31][5] , \w[31][4] , \w[31][3] , 
        \w[31][2] , \w[31][1] , 1'b0}), .CI(1'b0), .S({O[31:1], 
        SYNOPSYS_UNCONNECTED__30}) );
  AND U2 ( .A(A[5]), .B(B[4]), .Z(\_8_net_[9] ) );
  AND U3 ( .A(A[5]), .B(B[3]), .Z(\_8_net_[8] ) );
  AND U4 ( .A(A[5]), .B(B[2]), .Z(\_8_net_[7] ) );
  AND U5 ( .A(A[5]), .B(B[1]), .Z(\_8_net_[6] ) );
  AND U6 ( .A(A[5]), .B(B[0]), .Z(\_8_net_[5] ) );
  AND U7 ( .A(A[5]), .B(B[26]), .Z(\_8_net_[31] ) );
  AND U8 ( .A(A[5]), .B(B[25]), .Z(\_8_net_[30] ) );
  AND U9 ( .A(A[5]), .B(B[24]), .Z(\_8_net_[29] ) );
  AND U10 ( .A(A[5]), .B(B[23]), .Z(\_8_net_[28] ) );
  AND U11 ( .A(A[5]), .B(B[22]), .Z(\_8_net_[27] ) );
  AND U12 ( .A(A[5]), .B(B[21]), .Z(\_8_net_[26] ) );
  AND U13 ( .A(A[5]), .B(B[20]), .Z(\_8_net_[25] ) );
  AND U14 ( .A(A[5]), .B(B[19]), .Z(\_8_net_[24] ) );
  AND U15 ( .A(A[5]), .B(B[18]), .Z(\_8_net_[23] ) );
  AND U16 ( .A(A[5]), .B(B[17]), .Z(\_8_net_[22] ) );
  AND U17 ( .A(A[5]), .B(B[16]), .Z(\_8_net_[21] ) );
  AND U18 ( .A(A[5]), .B(B[15]), .Z(\_8_net_[20] ) );
  AND U19 ( .A(A[5]), .B(B[14]), .Z(\_8_net_[19] ) );
  AND U20 ( .A(A[5]), .B(B[13]), .Z(\_8_net_[18] ) );
  AND U21 ( .A(A[5]), .B(B[12]), .Z(\_8_net_[17] ) );
  AND U22 ( .A(A[5]), .B(B[11]), .Z(\_8_net_[16] ) );
  AND U23 ( .A(A[5]), .B(B[10]), .Z(\_8_net_[15] ) );
  AND U24 ( .A(A[5]), .B(B[9]), .Z(\_8_net_[14] ) );
  AND U25 ( .A(A[5]), .B(B[8]), .Z(\_8_net_[13] ) );
  AND U26 ( .A(A[5]), .B(B[7]), .Z(\_8_net_[12] ) );
  AND U27 ( .A(A[5]), .B(B[6]), .Z(\_8_net_[11] ) );
  AND U28 ( .A(A[5]), .B(B[5]), .Z(\_8_net_[10] ) );
  AND U29 ( .A(B[5]), .B(A[4]), .Z(\_6_net_[9] ) );
  AND U30 ( .A(B[4]), .B(A[4]), .Z(\_6_net_[8] ) );
  AND U31 ( .A(B[3]), .B(A[4]), .Z(\_6_net_[7] ) );
  AND U32 ( .A(B[2]), .B(A[4]), .Z(\_6_net_[6] ) );
  AND U33 ( .A(B[1]), .B(A[4]), .Z(\_6_net_[5] ) );
  AND U34 ( .A(B[0]), .B(A[4]), .Z(\_6_net_[4] ) );
  AND U35 ( .A(A[4]), .B(B[27]), .Z(\_6_net_[31] ) );
  AND U36 ( .A(B[26]), .B(A[4]), .Z(\_6_net_[30] ) );
  AND U37 ( .A(B[25]), .B(A[4]), .Z(\_6_net_[29] ) );
  AND U38 ( .A(B[24]), .B(A[4]), .Z(\_6_net_[28] ) );
  AND U39 ( .A(B[23]), .B(A[4]), .Z(\_6_net_[27] ) );
  AND U40 ( .A(B[22]), .B(A[4]), .Z(\_6_net_[26] ) );
  AND U41 ( .A(B[21]), .B(A[4]), .Z(\_6_net_[25] ) );
  AND U42 ( .A(B[20]), .B(A[4]), .Z(\_6_net_[24] ) );
  AND U43 ( .A(B[19]), .B(A[4]), .Z(\_6_net_[23] ) );
  AND U44 ( .A(B[18]), .B(A[4]), .Z(\_6_net_[22] ) );
  AND U45 ( .A(B[17]), .B(A[4]), .Z(\_6_net_[21] ) );
  AND U46 ( .A(B[16]), .B(A[4]), .Z(\_6_net_[20] ) );
  AND U47 ( .A(B[15]), .B(A[4]), .Z(\_6_net_[19] ) );
  AND U48 ( .A(B[14]), .B(A[4]), .Z(\_6_net_[18] ) );
  AND U49 ( .A(B[13]), .B(A[4]), .Z(\_6_net_[17] ) );
  AND U50 ( .A(B[12]), .B(A[4]), .Z(\_6_net_[16] ) );
  AND U51 ( .A(B[11]), .B(A[4]), .Z(\_6_net_[15] ) );
  AND U52 ( .A(B[10]), .B(A[4]), .Z(\_6_net_[14] ) );
  AND U53 ( .A(B[9]), .B(A[4]), .Z(\_6_net_[13] ) );
  AND U54 ( .A(B[8]), .B(A[4]), .Z(\_6_net_[12] ) );
  AND U55 ( .A(B[7]), .B(A[4]), .Z(\_6_net_[11] ) );
  AND U56 ( .A(B[6]), .B(A[4]), .Z(\_6_net_[10] ) );
  AND U57 ( .A(A[31]), .B(B[0]), .Z(\_60_net_[31] ) );
  AND U58 ( .A(B[1]), .B(A[30]), .Z(\_58_net_[31] ) );
  AND U59 ( .A(A[30]), .B(B[0]), .Z(\_58_net_[30] ) );
  AND U60 ( .A(B[2]), .B(A[29]), .Z(\_56_net_[31] ) );
  AND U61 ( .A(B[1]), .B(A[29]), .Z(\_56_net_[30] ) );
  AND U62 ( .A(A[29]), .B(B[0]), .Z(\_56_net_[29] ) );
  AND U63 ( .A(B[3]), .B(A[28]), .Z(\_54_net_[31] ) );
  AND U64 ( .A(B[2]), .B(A[28]), .Z(\_54_net_[30] ) );
  AND U65 ( .A(B[1]), .B(A[28]), .Z(\_54_net_[29] ) );
  AND U66 ( .A(A[28]), .B(B[0]), .Z(\_54_net_[28] ) );
  AND U67 ( .A(B[4]), .B(A[27]), .Z(\_52_net_[31] ) );
  AND U68 ( .A(B[3]), .B(A[27]), .Z(\_52_net_[30] ) );
  AND U69 ( .A(B[2]), .B(A[27]), .Z(\_52_net_[29] ) );
  AND U70 ( .A(B[1]), .B(A[27]), .Z(\_52_net_[28] ) );
  AND U71 ( .A(A[27]), .B(B[0]), .Z(\_52_net_[27] ) );
  AND U72 ( .A(B[5]), .B(A[26]), .Z(\_50_net_[31] ) );
  AND U73 ( .A(B[4]), .B(A[26]), .Z(\_50_net_[30] ) );
  AND U74 ( .A(B[3]), .B(A[26]), .Z(\_50_net_[29] ) );
  AND U75 ( .A(B[2]), .B(A[26]), .Z(\_50_net_[28] ) );
  AND U76 ( .A(B[1]), .B(A[26]), .Z(\_50_net_[27] ) );
  AND U77 ( .A(A[26]), .B(B[0]), .Z(\_50_net_[26] ) );
  AND U78 ( .A(B[6]), .B(A[3]), .Z(\_4_net_[9] ) );
  AND U79 ( .A(B[5]), .B(A[3]), .Z(\_4_net_[8] ) );
  AND U80 ( .A(B[4]), .B(A[3]), .Z(\_4_net_[7] ) );
  AND U81 ( .A(B[3]), .B(A[3]), .Z(\_4_net_[6] ) );
  AND U82 ( .A(B[2]), .B(A[3]), .Z(\_4_net_[5] ) );
  AND U83 ( .A(B[1]), .B(A[3]), .Z(\_4_net_[4] ) );
  AND U84 ( .A(B[0]), .B(A[3]), .Z(\_4_net_[3] ) );
  AND U85 ( .A(A[3]), .B(B[28]), .Z(\_4_net_[31] ) );
  AND U86 ( .A(B[27]), .B(A[3]), .Z(\_4_net_[30] ) );
  AND U87 ( .A(B[26]), .B(A[3]), .Z(\_4_net_[29] ) );
  AND U88 ( .A(B[25]), .B(A[3]), .Z(\_4_net_[28] ) );
  AND U89 ( .A(B[24]), .B(A[3]), .Z(\_4_net_[27] ) );
  AND U90 ( .A(B[23]), .B(A[3]), .Z(\_4_net_[26] ) );
  AND U91 ( .A(B[22]), .B(A[3]), .Z(\_4_net_[25] ) );
  AND U92 ( .A(B[21]), .B(A[3]), .Z(\_4_net_[24] ) );
  AND U93 ( .A(B[20]), .B(A[3]), .Z(\_4_net_[23] ) );
  AND U94 ( .A(B[19]), .B(A[3]), .Z(\_4_net_[22] ) );
  AND U95 ( .A(B[18]), .B(A[3]), .Z(\_4_net_[21] ) );
  AND U96 ( .A(B[17]), .B(A[3]), .Z(\_4_net_[20] ) );
  AND U97 ( .A(B[16]), .B(A[3]), .Z(\_4_net_[19] ) );
  AND U98 ( .A(B[15]), .B(A[3]), .Z(\_4_net_[18] ) );
  AND U99 ( .A(B[14]), .B(A[3]), .Z(\_4_net_[17] ) );
  AND U100 ( .A(B[13]), .B(A[3]), .Z(\_4_net_[16] ) );
  AND U101 ( .A(B[12]), .B(A[3]), .Z(\_4_net_[15] ) );
  AND U102 ( .A(B[11]), .B(A[3]), .Z(\_4_net_[14] ) );
  AND U103 ( .A(B[10]), .B(A[3]), .Z(\_4_net_[13] ) );
  AND U104 ( .A(B[9]), .B(A[3]), .Z(\_4_net_[12] ) );
  AND U105 ( .A(B[8]), .B(A[3]), .Z(\_4_net_[11] ) );
  AND U106 ( .A(B[7]), .B(A[3]), .Z(\_4_net_[10] ) );
  AND U107 ( .A(B[6]), .B(A[25]), .Z(\_48_net_[31] ) );
  AND U108 ( .A(B[5]), .B(A[25]), .Z(\_48_net_[30] ) );
  AND U109 ( .A(B[4]), .B(A[25]), .Z(\_48_net_[29] ) );
  AND U110 ( .A(B[3]), .B(A[25]), .Z(\_48_net_[28] ) );
  AND U111 ( .A(B[2]), .B(A[25]), .Z(\_48_net_[27] ) );
  AND U112 ( .A(B[1]), .B(A[25]), .Z(\_48_net_[26] ) );
  AND U113 ( .A(A[25]), .B(B[0]), .Z(\_48_net_[25] ) );
  AND U114 ( .A(B[7]), .B(A[24]), .Z(\_46_net_[31] ) );
  AND U115 ( .A(B[6]), .B(A[24]), .Z(\_46_net_[30] ) );
  AND U116 ( .A(B[5]), .B(A[24]), .Z(\_46_net_[29] ) );
  AND U117 ( .A(B[4]), .B(A[24]), .Z(\_46_net_[28] ) );
  AND U118 ( .A(B[3]), .B(A[24]), .Z(\_46_net_[27] ) );
  AND U119 ( .A(B[2]), .B(A[24]), .Z(\_46_net_[26] ) );
  AND U120 ( .A(B[1]), .B(A[24]), .Z(\_46_net_[25] ) );
  AND U121 ( .A(A[24]), .B(B[0]), .Z(\_46_net_[24] ) );
  AND U122 ( .A(B[8]), .B(A[23]), .Z(\_44_net_[31] ) );
  AND U123 ( .A(B[7]), .B(A[23]), .Z(\_44_net_[30] ) );
  AND U124 ( .A(B[6]), .B(A[23]), .Z(\_44_net_[29] ) );
  AND U125 ( .A(B[5]), .B(A[23]), .Z(\_44_net_[28] ) );
  AND U126 ( .A(B[4]), .B(A[23]), .Z(\_44_net_[27] ) );
  AND U127 ( .A(B[3]), .B(A[23]), .Z(\_44_net_[26] ) );
  AND U128 ( .A(B[2]), .B(A[23]), .Z(\_44_net_[25] ) );
  AND U129 ( .A(B[1]), .B(A[23]), .Z(\_44_net_[24] ) );
  AND U130 ( .A(A[23]), .B(B[0]), .Z(\_44_net_[23] ) );
  AND U131 ( .A(B[9]), .B(A[22]), .Z(\_42_net_[31] ) );
  AND U132 ( .A(B[8]), .B(A[22]), .Z(\_42_net_[30] ) );
  AND U133 ( .A(B[7]), .B(A[22]), .Z(\_42_net_[29] ) );
  AND U134 ( .A(B[6]), .B(A[22]), .Z(\_42_net_[28] ) );
  AND U135 ( .A(B[5]), .B(A[22]), .Z(\_42_net_[27] ) );
  AND U136 ( .A(B[4]), .B(A[22]), .Z(\_42_net_[26] ) );
  AND U137 ( .A(B[3]), .B(A[22]), .Z(\_42_net_[25] ) );
  AND U138 ( .A(B[2]), .B(A[22]), .Z(\_42_net_[24] ) );
  AND U139 ( .A(B[1]), .B(A[22]), .Z(\_42_net_[23] ) );
  AND U140 ( .A(A[22]), .B(B[0]), .Z(\_42_net_[22] ) );
  AND U141 ( .A(B[10]), .B(A[21]), .Z(\_40_net_[31] ) );
  AND U142 ( .A(B[9]), .B(A[21]), .Z(\_40_net_[30] ) );
  AND U143 ( .A(B[8]), .B(A[21]), .Z(\_40_net_[29] ) );
  AND U144 ( .A(B[7]), .B(A[21]), .Z(\_40_net_[28] ) );
  AND U145 ( .A(B[6]), .B(A[21]), .Z(\_40_net_[27] ) );
  AND U146 ( .A(B[5]), .B(A[21]), .Z(\_40_net_[26] ) );
  AND U147 ( .A(B[4]), .B(A[21]), .Z(\_40_net_[25] ) );
  AND U148 ( .A(B[3]), .B(A[21]), .Z(\_40_net_[24] ) );
  AND U149 ( .A(B[2]), .B(A[21]), .Z(\_40_net_[23] ) );
  AND U150 ( .A(B[1]), .B(A[21]), .Z(\_40_net_[22] ) );
  AND U151 ( .A(A[21]), .B(B[0]), .Z(\_40_net_[21] ) );
  AND U152 ( .A(B[11]), .B(A[20]), .Z(\_38_net_[31] ) );
  AND U153 ( .A(B[10]), .B(A[20]), .Z(\_38_net_[30] ) );
  AND U154 ( .A(B[9]), .B(A[20]), .Z(\_38_net_[29] ) );
  AND U155 ( .A(B[8]), .B(A[20]), .Z(\_38_net_[28] ) );
  AND U156 ( .A(B[7]), .B(A[20]), .Z(\_38_net_[27] ) );
  AND U157 ( .A(B[6]), .B(A[20]), .Z(\_38_net_[26] ) );
  AND U158 ( .A(B[5]), .B(A[20]), .Z(\_38_net_[25] ) );
  AND U159 ( .A(B[4]), .B(A[20]), .Z(\_38_net_[24] ) );
  AND U160 ( .A(B[3]), .B(A[20]), .Z(\_38_net_[23] ) );
  AND U161 ( .A(B[2]), .B(A[20]), .Z(\_38_net_[22] ) );
  AND U162 ( .A(B[1]), .B(A[20]), .Z(\_38_net_[21] ) );
  AND U163 ( .A(A[20]), .B(B[0]), .Z(\_38_net_[20] ) );
  AND U164 ( .A(B[12]), .B(A[19]), .Z(\_36_net_[31] ) );
  AND U165 ( .A(B[11]), .B(A[19]), .Z(\_36_net_[30] ) );
  AND U166 ( .A(B[10]), .B(A[19]), .Z(\_36_net_[29] ) );
  AND U167 ( .A(B[9]), .B(A[19]), .Z(\_36_net_[28] ) );
  AND U168 ( .A(B[8]), .B(A[19]), .Z(\_36_net_[27] ) );
  AND U169 ( .A(B[7]), .B(A[19]), .Z(\_36_net_[26] ) );
  AND U170 ( .A(B[6]), .B(A[19]), .Z(\_36_net_[25] ) );
  AND U171 ( .A(B[5]), .B(A[19]), .Z(\_36_net_[24] ) );
  AND U172 ( .A(B[4]), .B(A[19]), .Z(\_36_net_[23] ) );
  AND U173 ( .A(B[3]), .B(A[19]), .Z(\_36_net_[22] ) );
  AND U174 ( .A(B[2]), .B(A[19]), .Z(\_36_net_[21] ) );
  AND U175 ( .A(B[1]), .B(A[19]), .Z(\_36_net_[20] ) );
  AND U176 ( .A(A[19]), .B(B[0]), .Z(\_36_net_[19] ) );
  AND U177 ( .A(B[13]), .B(A[18]), .Z(\_34_net_[31] ) );
  AND U178 ( .A(B[12]), .B(A[18]), .Z(\_34_net_[30] ) );
  AND U179 ( .A(B[11]), .B(A[18]), .Z(\_34_net_[29] ) );
  AND U180 ( .A(B[10]), .B(A[18]), .Z(\_34_net_[28] ) );
  AND U181 ( .A(B[9]), .B(A[18]), .Z(\_34_net_[27] ) );
  AND U182 ( .A(B[8]), .B(A[18]), .Z(\_34_net_[26] ) );
  AND U183 ( .A(B[7]), .B(A[18]), .Z(\_34_net_[25] ) );
  AND U184 ( .A(B[6]), .B(A[18]), .Z(\_34_net_[24] ) );
  AND U185 ( .A(B[5]), .B(A[18]), .Z(\_34_net_[23] ) );
  AND U186 ( .A(B[4]), .B(A[18]), .Z(\_34_net_[22] ) );
  AND U187 ( .A(B[3]), .B(A[18]), .Z(\_34_net_[21] ) );
  AND U188 ( .A(B[2]), .B(A[18]), .Z(\_34_net_[20] ) );
  AND U189 ( .A(B[1]), .B(A[18]), .Z(\_34_net_[19] ) );
  AND U190 ( .A(A[18]), .B(B[0]), .Z(\_34_net_[18] ) );
  AND U191 ( .A(B[14]), .B(A[17]), .Z(\_32_net_[31] ) );
  AND U192 ( .A(B[13]), .B(A[17]), .Z(\_32_net_[30] ) );
  AND U193 ( .A(B[12]), .B(A[17]), .Z(\_32_net_[29] ) );
  AND U194 ( .A(B[11]), .B(A[17]), .Z(\_32_net_[28] ) );
  AND U195 ( .A(B[10]), .B(A[17]), .Z(\_32_net_[27] ) );
  AND U196 ( .A(B[9]), .B(A[17]), .Z(\_32_net_[26] ) );
  AND U197 ( .A(B[8]), .B(A[17]), .Z(\_32_net_[25] ) );
  AND U198 ( .A(B[7]), .B(A[17]), .Z(\_32_net_[24] ) );
  AND U199 ( .A(B[6]), .B(A[17]), .Z(\_32_net_[23] ) );
  AND U200 ( .A(B[5]), .B(A[17]), .Z(\_32_net_[22] ) );
  AND U201 ( .A(B[4]), .B(A[17]), .Z(\_32_net_[21] ) );
  AND U202 ( .A(B[3]), .B(A[17]), .Z(\_32_net_[20] ) );
  AND U203 ( .A(B[2]), .B(A[17]), .Z(\_32_net_[19] ) );
  AND U204 ( .A(B[1]), .B(A[17]), .Z(\_32_net_[18] ) );
  AND U205 ( .A(A[17]), .B(B[0]), .Z(\_32_net_[17] ) );
  AND U206 ( .A(B[15]), .B(A[16]), .Z(\_30_net_[31] ) );
  AND U207 ( .A(B[14]), .B(A[16]), .Z(\_30_net_[30] ) );
  AND U208 ( .A(B[13]), .B(A[16]), .Z(\_30_net_[29] ) );
  AND U209 ( .A(B[12]), .B(A[16]), .Z(\_30_net_[28] ) );
  AND U210 ( .A(B[11]), .B(A[16]), .Z(\_30_net_[27] ) );
  AND U211 ( .A(B[10]), .B(A[16]), .Z(\_30_net_[26] ) );
  AND U212 ( .A(B[9]), .B(A[16]), .Z(\_30_net_[25] ) );
  AND U213 ( .A(B[8]), .B(A[16]), .Z(\_30_net_[24] ) );
  AND U214 ( .A(B[7]), .B(A[16]), .Z(\_30_net_[23] ) );
  AND U215 ( .A(B[6]), .B(A[16]), .Z(\_30_net_[22] ) );
  AND U216 ( .A(B[5]), .B(A[16]), .Z(\_30_net_[21] ) );
  AND U217 ( .A(B[4]), .B(A[16]), .Z(\_30_net_[20] ) );
  AND U218 ( .A(B[3]), .B(A[16]), .Z(\_30_net_[19] ) );
  AND U219 ( .A(B[2]), .B(A[16]), .Z(\_30_net_[18] ) );
  AND U220 ( .A(B[1]), .B(A[16]), .Z(\_30_net_[17] ) );
  AND U221 ( .A(A[16]), .B(B[0]), .Z(\_30_net_[16] ) );
  AND U222 ( .A(B[7]), .B(A[2]), .Z(\_2_net_[9] ) );
  AND U223 ( .A(B[6]), .B(A[2]), .Z(\_2_net_[8] ) );
  AND U224 ( .A(B[5]), .B(A[2]), .Z(\_2_net_[7] ) );
  AND U225 ( .A(B[4]), .B(A[2]), .Z(\_2_net_[6] ) );
  AND U226 ( .A(B[3]), .B(A[2]), .Z(\_2_net_[5] ) );
  AND U227 ( .A(B[2]), .B(A[2]), .Z(\_2_net_[4] ) );
  AND U228 ( .A(B[1]), .B(A[2]), .Z(\_2_net_[3] ) );
  AND U229 ( .A(A[2]), .B(B[29]), .Z(\_2_net_[31] ) );
  AND U230 ( .A(B[28]), .B(A[2]), .Z(\_2_net_[30] ) );
  AND U231 ( .A(B[0]), .B(A[2]), .Z(\_2_net_[2] ) );
  AND U232 ( .A(B[27]), .B(A[2]), .Z(\_2_net_[29] ) );
  AND U233 ( .A(B[26]), .B(A[2]), .Z(\_2_net_[28] ) );
  AND U234 ( .A(B[25]), .B(A[2]), .Z(\_2_net_[27] ) );
  AND U235 ( .A(B[24]), .B(A[2]), .Z(\_2_net_[26] ) );
  AND U236 ( .A(B[23]), .B(A[2]), .Z(\_2_net_[25] ) );
  AND U237 ( .A(B[22]), .B(A[2]), .Z(\_2_net_[24] ) );
  AND U238 ( .A(B[21]), .B(A[2]), .Z(\_2_net_[23] ) );
  AND U239 ( .A(B[20]), .B(A[2]), .Z(\_2_net_[22] ) );
  AND U240 ( .A(B[19]), .B(A[2]), .Z(\_2_net_[21] ) );
  AND U241 ( .A(B[18]), .B(A[2]), .Z(\_2_net_[20] ) );
  AND U242 ( .A(B[17]), .B(A[2]), .Z(\_2_net_[19] ) );
  AND U243 ( .A(B[16]), .B(A[2]), .Z(\_2_net_[18] ) );
  AND U244 ( .A(B[15]), .B(A[2]), .Z(\_2_net_[17] ) );
  AND U245 ( .A(B[14]), .B(A[2]), .Z(\_2_net_[16] ) );
  AND U246 ( .A(B[13]), .B(A[2]), .Z(\_2_net_[15] ) );
  AND U247 ( .A(B[12]), .B(A[2]), .Z(\_2_net_[14] ) );
  AND U248 ( .A(B[11]), .B(A[2]), .Z(\_2_net_[13] ) );
  AND U249 ( .A(B[10]), .B(A[2]), .Z(\_2_net_[12] ) );
  AND U250 ( .A(B[9]), .B(A[2]), .Z(\_2_net_[11] ) );
  AND U251 ( .A(B[8]), .B(A[2]), .Z(\_2_net_[10] ) );
  AND U252 ( .A(B[16]), .B(A[15]), .Z(\_28_net_[31] ) );
  AND U253 ( .A(B[15]), .B(A[15]), .Z(\_28_net_[30] ) );
  AND U254 ( .A(B[14]), .B(A[15]), .Z(\_28_net_[29] ) );
  AND U255 ( .A(B[13]), .B(A[15]), .Z(\_28_net_[28] ) );
  AND U256 ( .A(B[12]), .B(A[15]), .Z(\_28_net_[27] ) );
  AND U257 ( .A(B[11]), .B(A[15]), .Z(\_28_net_[26] ) );
  AND U258 ( .A(B[10]), .B(A[15]), .Z(\_28_net_[25] ) );
  AND U259 ( .A(B[9]), .B(A[15]), .Z(\_28_net_[24] ) );
  AND U260 ( .A(B[8]), .B(A[15]), .Z(\_28_net_[23] ) );
  AND U261 ( .A(B[7]), .B(A[15]), .Z(\_28_net_[22] ) );
  AND U262 ( .A(B[6]), .B(A[15]), .Z(\_28_net_[21] ) );
  AND U263 ( .A(B[5]), .B(A[15]), .Z(\_28_net_[20] ) );
  AND U264 ( .A(B[4]), .B(A[15]), .Z(\_28_net_[19] ) );
  AND U265 ( .A(B[3]), .B(A[15]), .Z(\_28_net_[18] ) );
  AND U266 ( .A(B[2]), .B(A[15]), .Z(\_28_net_[17] ) );
  AND U267 ( .A(B[1]), .B(A[15]), .Z(\_28_net_[16] ) );
  AND U268 ( .A(A[15]), .B(B[0]), .Z(\_28_net_[15] ) );
  AND U269 ( .A(B[17]), .B(A[14]), .Z(\_26_net_[31] ) );
  AND U270 ( .A(B[16]), .B(A[14]), .Z(\_26_net_[30] ) );
  AND U271 ( .A(B[15]), .B(A[14]), .Z(\_26_net_[29] ) );
  AND U272 ( .A(B[14]), .B(A[14]), .Z(\_26_net_[28] ) );
  AND U273 ( .A(B[13]), .B(A[14]), .Z(\_26_net_[27] ) );
  AND U274 ( .A(B[12]), .B(A[14]), .Z(\_26_net_[26] ) );
  AND U275 ( .A(B[11]), .B(A[14]), .Z(\_26_net_[25] ) );
  AND U276 ( .A(B[10]), .B(A[14]), .Z(\_26_net_[24] ) );
  AND U277 ( .A(B[9]), .B(A[14]), .Z(\_26_net_[23] ) );
  AND U278 ( .A(B[8]), .B(A[14]), .Z(\_26_net_[22] ) );
  AND U279 ( .A(B[7]), .B(A[14]), .Z(\_26_net_[21] ) );
  AND U280 ( .A(B[6]), .B(A[14]), .Z(\_26_net_[20] ) );
  AND U281 ( .A(B[5]), .B(A[14]), .Z(\_26_net_[19] ) );
  AND U282 ( .A(B[4]), .B(A[14]), .Z(\_26_net_[18] ) );
  AND U283 ( .A(B[3]), .B(A[14]), .Z(\_26_net_[17] ) );
  AND U284 ( .A(B[2]), .B(A[14]), .Z(\_26_net_[16] ) );
  AND U285 ( .A(B[1]), .B(A[14]), .Z(\_26_net_[15] ) );
  AND U286 ( .A(A[14]), .B(B[0]), .Z(\_26_net_[14] ) );
  AND U287 ( .A(B[18]), .B(A[13]), .Z(\_24_net_[31] ) );
  AND U288 ( .A(B[17]), .B(A[13]), .Z(\_24_net_[30] ) );
  AND U289 ( .A(B[16]), .B(A[13]), .Z(\_24_net_[29] ) );
  AND U290 ( .A(B[15]), .B(A[13]), .Z(\_24_net_[28] ) );
  AND U291 ( .A(B[14]), .B(A[13]), .Z(\_24_net_[27] ) );
  AND U292 ( .A(B[13]), .B(A[13]), .Z(\_24_net_[26] ) );
  AND U293 ( .A(B[12]), .B(A[13]), .Z(\_24_net_[25] ) );
  AND U294 ( .A(B[11]), .B(A[13]), .Z(\_24_net_[24] ) );
  AND U295 ( .A(B[10]), .B(A[13]), .Z(\_24_net_[23] ) );
  AND U296 ( .A(B[9]), .B(A[13]), .Z(\_24_net_[22] ) );
  AND U297 ( .A(B[8]), .B(A[13]), .Z(\_24_net_[21] ) );
  AND U298 ( .A(B[7]), .B(A[13]), .Z(\_24_net_[20] ) );
  AND U299 ( .A(B[6]), .B(A[13]), .Z(\_24_net_[19] ) );
  AND U300 ( .A(B[5]), .B(A[13]), .Z(\_24_net_[18] ) );
  AND U301 ( .A(B[4]), .B(A[13]), .Z(\_24_net_[17] ) );
  AND U302 ( .A(B[3]), .B(A[13]), .Z(\_24_net_[16] ) );
  AND U303 ( .A(B[2]), .B(A[13]), .Z(\_24_net_[15] ) );
  AND U304 ( .A(B[1]), .B(A[13]), .Z(\_24_net_[14] ) );
  AND U305 ( .A(A[13]), .B(B[0]), .Z(\_24_net_[13] ) );
  AND U306 ( .A(B[19]), .B(A[12]), .Z(\_22_net_[31] ) );
  AND U307 ( .A(B[18]), .B(A[12]), .Z(\_22_net_[30] ) );
  AND U308 ( .A(B[17]), .B(A[12]), .Z(\_22_net_[29] ) );
  AND U309 ( .A(B[16]), .B(A[12]), .Z(\_22_net_[28] ) );
  AND U310 ( .A(B[15]), .B(A[12]), .Z(\_22_net_[27] ) );
  AND U311 ( .A(B[14]), .B(A[12]), .Z(\_22_net_[26] ) );
  AND U312 ( .A(B[13]), .B(A[12]), .Z(\_22_net_[25] ) );
  AND U313 ( .A(B[12]), .B(A[12]), .Z(\_22_net_[24] ) );
  AND U314 ( .A(B[11]), .B(A[12]), .Z(\_22_net_[23] ) );
  AND U315 ( .A(B[10]), .B(A[12]), .Z(\_22_net_[22] ) );
  AND U316 ( .A(B[9]), .B(A[12]), .Z(\_22_net_[21] ) );
  AND U317 ( .A(B[8]), .B(A[12]), .Z(\_22_net_[20] ) );
  AND U318 ( .A(B[7]), .B(A[12]), .Z(\_22_net_[19] ) );
  AND U319 ( .A(B[6]), .B(A[12]), .Z(\_22_net_[18] ) );
  AND U320 ( .A(B[5]), .B(A[12]), .Z(\_22_net_[17] ) );
  AND U321 ( .A(B[4]), .B(A[12]), .Z(\_22_net_[16] ) );
  AND U322 ( .A(B[3]), .B(A[12]), .Z(\_22_net_[15] ) );
  AND U323 ( .A(B[2]), .B(A[12]), .Z(\_22_net_[14] ) );
  AND U324 ( .A(B[1]), .B(A[12]), .Z(\_22_net_[13] ) );
  AND U325 ( .A(A[12]), .B(B[0]), .Z(\_22_net_[12] ) );
  AND U326 ( .A(B[20]), .B(A[11]), .Z(\_20_net_[31] ) );
  AND U327 ( .A(B[19]), .B(A[11]), .Z(\_20_net_[30] ) );
  AND U328 ( .A(B[18]), .B(A[11]), .Z(\_20_net_[29] ) );
  AND U329 ( .A(B[17]), .B(A[11]), .Z(\_20_net_[28] ) );
  AND U330 ( .A(B[16]), .B(A[11]), .Z(\_20_net_[27] ) );
  AND U331 ( .A(B[15]), .B(A[11]), .Z(\_20_net_[26] ) );
  AND U332 ( .A(B[14]), .B(A[11]), .Z(\_20_net_[25] ) );
  AND U333 ( .A(B[13]), .B(A[11]), .Z(\_20_net_[24] ) );
  AND U334 ( .A(B[12]), .B(A[11]), .Z(\_20_net_[23] ) );
  AND U335 ( .A(B[11]), .B(A[11]), .Z(\_20_net_[22] ) );
  AND U336 ( .A(B[10]), .B(A[11]), .Z(\_20_net_[21] ) );
  AND U337 ( .A(B[9]), .B(A[11]), .Z(\_20_net_[20] ) );
  AND U338 ( .A(B[8]), .B(A[11]), .Z(\_20_net_[19] ) );
  AND U339 ( .A(B[7]), .B(A[11]), .Z(\_20_net_[18] ) );
  AND U340 ( .A(B[6]), .B(A[11]), .Z(\_20_net_[17] ) );
  AND U341 ( .A(B[5]), .B(A[11]), .Z(\_20_net_[16] ) );
  AND U342 ( .A(B[4]), .B(A[11]), .Z(\_20_net_[15] ) );
  AND U343 ( .A(B[3]), .B(A[11]), .Z(\_20_net_[14] ) );
  AND U344 ( .A(B[2]), .B(A[11]), .Z(\_20_net_[13] ) );
  AND U345 ( .A(B[1]), .B(A[11]), .Z(\_20_net_[12] ) );
  AND U346 ( .A(A[11]), .B(B[0]), .Z(\_20_net_[11] ) );
  AND U347 ( .A(B[21]), .B(A[10]), .Z(\_18_net_[31] ) );
  AND U348 ( .A(B[20]), .B(A[10]), .Z(\_18_net_[30] ) );
  AND U349 ( .A(B[19]), .B(A[10]), .Z(\_18_net_[29] ) );
  AND U350 ( .A(B[18]), .B(A[10]), .Z(\_18_net_[28] ) );
  AND U351 ( .A(B[17]), .B(A[10]), .Z(\_18_net_[27] ) );
  AND U352 ( .A(B[16]), .B(A[10]), .Z(\_18_net_[26] ) );
  AND U353 ( .A(B[15]), .B(A[10]), .Z(\_18_net_[25] ) );
  AND U354 ( .A(B[14]), .B(A[10]), .Z(\_18_net_[24] ) );
  AND U355 ( .A(B[13]), .B(A[10]), .Z(\_18_net_[23] ) );
  AND U356 ( .A(B[12]), .B(A[10]), .Z(\_18_net_[22] ) );
  AND U357 ( .A(B[11]), .B(A[10]), .Z(\_18_net_[21] ) );
  AND U358 ( .A(B[10]), .B(A[10]), .Z(\_18_net_[20] ) );
  AND U359 ( .A(B[9]), .B(A[10]), .Z(\_18_net_[19] ) );
  AND U360 ( .A(B[8]), .B(A[10]), .Z(\_18_net_[18] ) );
  AND U361 ( .A(B[7]), .B(A[10]), .Z(\_18_net_[17] ) );
  AND U362 ( .A(B[6]), .B(A[10]), .Z(\_18_net_[16] ) );
  AND U363 ( .A(B[5]), .B(A[10]), .Z(\_18_net_[15] ) );
  AND U364 ( .A(B[4]), .B(A[10]), .Z(\_18_net_[14] ) );
  AND U365 ( .A(B[3]), .B(A[10]), .Z(\_18_net_[13] ) );
  AND U366 ( .A(B[2]), .B(A[10]), .Z(\_18_net_[12] ) );
  AND U367 ( .A(B[1]), .B(A[10]), .Z(\_18_net_[11] ) );
  AND U368 ( .A(A[10]), .B(B[0]), .Z(\_18_net_[10] ) );
  AND U369 ( .A(B[0]), .B(A[9]), .Z(\_16_net_[9] ) );
  AND U370 ( .A(B[22]), .B(A[9]), .Z(\_16_net_[31] ) );
  AND U371 ( .A(B[21]), .B(A[9]), .Z(\_16_net_[30] ) );
  AND U372 ( .A(B[20]), .B(A[9]), .Z(\_16_net_[29] ) );
  AND U373 ( .A(B[19]), .B(A[9]), .Z(\_16_net_[28] ) );
  AND U374 ( .A(B[18]), .B(A[9]), .Z(\_16_net_[27] ) );
  AND U375 ( .A(B[17]), .B(A[9]), .Z(\_16_net_[26] ) );
  AND U376 ( .A(B[16]), .B(A[9]), .Z(\_16_net_[25] ) );
  AND U377 ( .A(B[15]), .B(A[9]), .Z(\_16_net_[24] ) );
  AND U378 ( .A(B[14]), .B(A[9]), .Z(\_16_net_[23] ) );
  AND U379 ( .A(B[13]), .B(A[9]), .Z(\_16_net_[22] ) );
  AND U380 ( .A(B[12]), .B(A[9]), .Z(\_16_net_[21] ) );
  AND U381 ( .A(B[11]), .B(A[9]), .Z(\_16_net_[20] ) );
  AND U382 ( .A(B[10]), .B(A[9]), .Z(\_16_net_[19] ) );
  AND U383 ( .A(B[9]), .B(A[9]), .Z(\_16_net_[18] ) );
  AND U384 ( .A(B[8]), .B(A[9]), .Z(\_16_net_[17] ) );
  AND U385 ( .A(B[7]), .B(A[9]), .Z(\_16_net_[16] ) );
  AND U386 ( .A(B[6]), .B(A[9]), .Z(\_16_net_[15] ) );
  AND U387 ( .A(B[5]), .B(A[9]), .Z(\_16_net_[14] ) );
  AND U388 ( .A(B[4]), .B(A[9]), .Z(\_16_net_[13] ) );
  AND U389 ( .A(B[3]), .B(A[9]), .Z(\_16_net_[12] ) );
  AND U390 ( .A(B[2]), .B(A[9]), .Z(\_16_net_[11] ) );
  AND U391 ( .A(A[9]), .B(B[1]), .Z(\_16_net_[10] ) );
  AND U392 ( .A(B[1]), .B(A[8]), .Z(\_14_net_[9] ) );
  AND U393 ( .A(B[0]), .B(A[8]), .Z(\_14_net_[8] ) );
  AND U394 ( .A(B[23]), .B(A[8]), .Z(\_14_net_[31] ) );
  AND U395 ( .A(B[22]), .B(A[8]), .Z(\_14_net_[30] ) );
  AND U396 ( .A(B[21]), .B(A[8]), .Z(\_14_net_[29] ) );
  AND U397 ( .A(B[20]), .B(A[8]), .Z(\_14_net_[28] ) );
  AND U398 ( .A(B[19]), .B(A[8]), .Z(\_14_net_[27] ) );
  AND U399 ( .A(B[18]), .B(A[8]), .Z(\_14_net_[26] ) );
  AND U400 ( .A(B[17]), .B(A[8]), .Z(\_14_net_[25] ) );
  AND U401 ( .A(B[16]), .B(A[8]), .Z(\_14_net_[24] ) );
  AND U402 ( .A(B[15]), .B(A[8]), .Z(\_14_net_[23] ) );
  AND U403 ( .A(B[14]), .B(A[8]), .Z(\_14_net_[22] ) );
  AND U404 ( .A(B[13]), .B(A[8]), .Z(\_14_net_[21] ) );
  AND U405 ( .A(B[12]), .B(A[8]), .Z(\_14_net_[20] ) );
  AND U406 ( .A(B[11]), .B(A[8]), .Z(\_14_net_[19] ) );
  AND U407 ( .A(B[10]), .B(A[8]), .Z(\_14_net_[18] ) );
  AND U408 ( .A(B[9]), .B(A[8]), .Z(\_14_net_[17] ) );
  AND U409 ( .A(B[8]), .B(A[8]), .Z(\_14_net_[16] ) );
  AND U410 ( .A(B[7]), .B(A[8]), .Z(\_14_net_[15] ) );
  AND U411 ( .A(B[6]), .B(A[8]), .Z(\_14_net_[14] ) );
  AND U412 ( .A(B[5]), .B(A[8]), .Z(\_14_net_[13] ) );
  AND U413 ( .A(B[4]), .B(A[8]), .Z(\_14_net_[12] ) );
  AND U414 ( .A(B[3]), .B(A[8]), .Z(\_14_net_[11] ) );
  AND U415 ( .A(A[8]), .B(B[2]), .Z(\_14_net_[10] ) );
  AND U416 ( .A(B[2]), .B(A[7]), .Z(\_12_net_[9] ) );
  AND U417 ( .A(B[1]), .B(A[7]), .Z(\_12_net_[8] ) );
  AND U418 ( .A(B[0]), .B(A[7]), .Z(\_12_net_[7] ) );
  AND U419 ( .A(B[24]), .B(A[7]), .Z(\_12_net_[31] ) );
  AND U420 ( .A(B[23]), .B(A[7]), .Z(\_12_net_[30] ) );
  AND U421 ( .A(B[22]), .B(A[7]), .Z(\_12_net_[29] ) );
  AND U422 ( .A(B[21]), .B(A[7]), .Z(\_12_net_[28] ) );
  AND U423 ( .A(B[20]), .B(A[7]), .Z(\_12_net_[27] ) );
  AND U424 ( .A(B[19]), .B(A[7]), .Z(\_12_net_[26] ) );
  AND U425 ( .A(B[18]), .B(A[7]), .Z(\_12_net_[25] ) );
  AND U426 ( .A(B[17]), .B(A[7]), .Z(\_12_net_[24] ) );
  AND U427 ( .A(B[16]), .B(A[7]), .Z(\_12_net_[23] ) );
  AND U428 ( .A(B[15]), .B(A[7]), .Z(\_12_net_[22] ) );
  AND U429 ( .A(B[14]), .B(A[7]), .Z(\_12_net_[21] ) );
  AND U430 ( .A(B[13]), .B(A[7]), .Z(\_12_net_[20] ) );
  AND U431 ( .A(B[12]), .B(A[7]), .Z(\_12_net_[19] ) );
  AND U432 ( .A(B[11]), .B(A[7]), .Z(\_12_net_[18] ) );
  AND U433 ( .A(B[10]), .B(A[7]), .Z(\_12_net_[17] ) );
  AND U434 ( .A(B[9]), .B(A[7]), .Z(\_12_net_[16] ) );
  AND U435 ( .A(B[8]), .B(A[7]), .Z(\_12_net_[15] ) );
  AND U436 ( .A(B[7]), .B(A[7]), .Z(\_12_net_[14] ) );
  AND U437 ( .A(B[6]), .B(A[7]), .Z(\_12_net_[13] ) );
  AND U438 ( .A(B[5]), .B(A[7]), .Z(\_12_net_[12] ) );
  AND U439 ( .A(B[4]), .B(A[7]), .Z(\_12_net_[11] ) );
  AND U440 ( .A(A[7]), .B(B[3]), .Z(\_12_net_[10] ) );
  AND U441 ( .A(B[3]), .B(A[6]), .Z(\_10_net_[9] ) );
  AND U442 ( .A(B[2]), .B(A[6]), .Z(\_10_net_[8] ) );
  AND U443 ( .A(B[1]), .B(A[6]), .Z(\_10_net_[7] ) );
  AND U444 ( .A(B[0]), .B(A[6]), .Z(\_10_net_[6] ) );
  AND U445 ( .A(B[25]), .B(A[6]), .Z(\_10_net_[31] ) );
  AND U446 ( .A(B[24]), .B(A[6]), .Z(\_10_net_[30] ) );
  AND U447 ( .A(B[23]), .B(A[6]), .Z(\_10_net_[29] ) );
  AND U448 ( .A(B[22]), .B(A[6]), .Z(\_10_net_[28] ) );
  AND U449 ( .A(B[21]), .B(A[6]), .Z(\_10_net_[27] ) );
  AND U450 ( .A(B[20]), .B(A[6]), .Z(\_10_net_[26] ) );
  AND U451 ( .A(B[19]), .B(A[6]), .Z(\_10_net_[25] ) );
  AND U452 ( .A(B[18]), .B(A[6]), .Z(\_10_net_[24] ) );
  AND U453 ( .A(B[17]), .B(A[6]), .Z(\_10_net_[23] ) );
  AND U454 ( .A(B[16]), .B(A[6]), .Z(\_10_net_[22] ) );
  AND U455 ( .A(B[15]), .B(A[6]), .Z(\_10_net_[21] ) );
  AND U456 ( .A(B[14]), .B(A[6]), .Z(\_10_net_[20] ) );
  AND U457 ( .A(B[13]), .B(A[6]), .Z(\_10_net_[19] ) );
  AND U458 ( .A(B[12]), .B(A[6]), .Z(\_10_net_[18] ) );
  AND U459 ( .A(B[11]), .B(A[6]), .Z(\_10_net_[17] ) );
  AND U460 ( .A(B[10]), .B(A[6]), .Z(\_10_net_[16] ) );
  AND U461 ( .A(B[9]), .B(A[6]), .Z(\_10_net_[15] ) );
  AND U462 ( .A(B[8]), .B(A[6]), .Z(\_10_net_[14] ) );
  AND U463 ( .A(B[7]), .B(A[6]), .Z(\_10_net_[13] ) );
  AND U464 ( .A(B[6]), .B(A[6]), .Z(\_10_net_[12] ) );
  AND U465 ( .A(B[5]), .B(A[6]), .Z(\_10_net_[11] ) );
  AND U466 ( .A(A[6]), .B(B[4]), .Z(\_10_net_[10] ) );
  AND U467 ( .A(B[8]), .B(A[1]), .Z(\_0_net_[9] ) );
  AND U468 ( .A(B[7]), .B(A[1]), .Z(\_0_net_[8] ) );
  AND U469 ( .A(B[6]), .B(A[1]), .Z(\_0_net_[7] ) );
  AND U470 ( .A(B[5]), .B(A[1]), .Z(\_0_net_[6] ) );
  AND U471 ( .A(B[4]), .B(A[1]), .Z(\_0_net_[5] ) );
  AND U472 ( .A(B[3]), .B(A[1]), .Z(\_0_net_[4] ) );
  AND U473 ( .A(B[2]), .B(A[1]), .Z(\_0_net_[3] ) );
  AND U474 ( .A(B[30]), .B(A[1]), .Z(\_0_net_[31] ) );
  AND U475 ( .A(B[29]), .B(A[1]), .Z(\_0_net_[30] ) );
  AND U476 ( .A(B[1]), .B(A[1]), .Z(\_0_net_[2] ) );
  AND U477 ( .A(B[28]), .B(A[1]), .Z(\_0_net_[29] ) );
  AND U478 ( .A(B[27]), .B(A[1]), .Z(\_0_net_[28] ) );
  AND U479 ( .A(B[26]), .B(A[1]), .Z(\_0_net_[27] ) );
  AND U480 ( .A(B[25]), .B(A[1]), .Z(\_0_net_[26] ) );
  AND U481 ( .A(B[24]), .B(A[1]), .Z(\_0_net_[25] ) );
  AND U482 ( .A(B[23]), .B(A[1]), .Z(\_0_net_[24] ) );
  AND U483 ( .A(B[22]), .B(A[1]), .Z(\_0_net_[23] ) );
  AND U484 ( .A(B[21]), .B(A[1]), .Z(\_0_net_[22] ) );
  AND U485 ( .A(B[20]), .B(A[1]), .Z(\_0_net_[21] ) );
  AND U486 ( .A(B[19]), .B(A[1]), .Z(\_0_net_[20] ) );
  AND U487 ( .A(B[0]), .B(A[1]), .Z(\_0_net_[1] ) );
  AND U488 ( .A(B[18]), .B(A[1]), .Z(\_0_net_[19] ) );
  AND U489 ( .A(B[17]), .B(A[1]), .Z(\_0_net_[18] ) );
  AND U490 ( .A(B[16]), .B(A[1]), .Z(\_0_net_[17] ) );
  AND U491 ( .A(B[15]), .B(A[1]), .Z(\_0_net_[16] ) );
  AND U492 ( .A(B[14]), .B(A[1]), .Z(\_0_net_[15] ) );
  AND U493 ( .A(B[13]), .B(A[1]), .Z(\_0_net_[14] ) );
  AND U494 ( .A(B[12]), .B(A[1]), .Z(\_0_net_[13] ) );
  AND U495 ( .A(B[11]), .B(A[1]), .Z(\_0_net_[12] ) );
  AND U496 ( .A(B[10]), .B(A[1]), .Z(\_0_net_[11] ) );
  AND U497 ( .A(A[1]), .B(B[9]), .Z(\_0_net_[10] ) );
endmodule


module FA_4961 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_4962 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4963 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4964 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4965 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4966 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4967 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4968 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4969 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4970 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4971 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4972 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4973 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4974 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4975 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4976 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4977 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4978 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4979 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4980 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4981 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4982 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4983 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4984 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4985 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4986 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4987 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4988 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4989 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4990 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4991 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_159 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;


  FA_4991 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_4990 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_4989 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_4988 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_4987 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_4986 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_4985 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_4984 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_4983 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_4982 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_4981 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_4980 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_4979 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_4978 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_4977 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_4976 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_4975 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_4974 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_4973 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_4972 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_4971 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_4970 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_4969 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_4968 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_4967 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_4966 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_4965 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_4964 \FAINST[28].FA_  ( .A(1'b0), .B(B[28]), .CI(1'b0), .S(S[28]) );
  FA_4963 \FAINST[29].FA_  ( .A(1'b0), .B(B[29]), .CI(1'b0), .S(S[29]) );
  FA_4962 \FAINST[30].FA_  ( .A(1'b0), .B(B[30]), .CI(1'b0), .S(S[30]) );
  FA_4961 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(1'b0), .S(S[31]) );
endmodule


module FA_4993 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_4994 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_4995 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4996 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4997 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4998 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4999 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5000 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5001 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5002 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5003 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5004 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5005 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5006 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5007 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5008 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5009 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5010 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5011 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5012 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5013 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5014 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5015 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5016 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5017 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5018 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5019 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5020 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5021 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5022 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5023 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_160 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;
  wire   \C[31] ;

  FA_5023 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_5022 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_5021 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_5020 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_5019 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_5018 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_5017 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_5016 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_5015 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_5014 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_5013 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_5012 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_5011 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_5010 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_5009 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_5008 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_5007 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_5006 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_5005 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_5004 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_5003 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_5002 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_5001 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_5000 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_4999 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_4998 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_4997 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_4996 \FAINST[28].FA_  ( .A(1'b0), .B(B[28]), .CI(1'b0), .S(S[28]) );
  FA_4995 \FAINST[29].FA_  ( .A(1'b0), .B(B[29]), .CI(1'b0), .S(S[29]) );
  FA_4994 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(1'b0), .S(S[30]), .CO(
        \C[31] ) );
  FA_4993 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(\C[31] ), .S(S[31]) );
endmodule


module FA_5025 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_5026 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5027 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_5028 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5029 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5030 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5031 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5032 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5033 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5034 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5035 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5036 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5037 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5038 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5039 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5040 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5041 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5042 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5043 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5044 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5045 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5046 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5047 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5048 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5049 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5050 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5051 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5052 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5053 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5054 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5055 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_161 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_5055 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_5054 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_5053 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_5052 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_5051 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_5050 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_5049 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_5048 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_5047 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_5046 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_5045 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_5044 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_5043 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_5042 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_5041 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_5040 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_5039 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_5038 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_5037 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_5036 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_5035 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_5034 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_5033 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_5032 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_5031 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_5030 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_5029 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_5028 \FAINST[28].FA_  ( .A(1'b0), .B(B[28]), .CI(1'b0), .S(S[28]) );
  FA_5027 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(1'b0), .S(S[29]), .CO(
        C[30]) );
  FA_5026 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_5025 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_5057 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_5058 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5059 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5060 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_5061 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5062 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5063 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5064 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5065 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5066 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5067 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5068 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5069 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5070 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5071 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5072 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5073 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5074 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5075 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5076 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5077 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5078 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5079 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5080 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5081 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5082 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5083 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5084 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5085 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5086 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5087 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_162 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_5087 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_5086 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_5085 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_5084 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_5083 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_5082 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_5081 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_5080 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_5079 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_5078 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_5077 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_5076 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_5075 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_5074 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_5073 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_5072 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_5071 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_5070 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_5069 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_5068 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_5067 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_5066 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_5065 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_5064 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_5063 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_5062 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_5061 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_5060 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(1'b0), .S(S[28]), .CO(
        C[29]) );
  FA_5059 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_5058 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_5057 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_5089 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_5090 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5091 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5092 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5093 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_5094 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5095 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5096 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5097 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5098 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5099 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5104 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_163 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_5119 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_5118 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_5117 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_5116 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_5115 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_5114 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_5113 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_5112 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_5111 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_5110 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_5109 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_5108 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_5107 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_5106 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_5105 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_5104 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_5103 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_5102 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_5101 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_5100 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_5099 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_5098 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_5097 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_5096 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_5095 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_5094 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_5093 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(1'b0), .S(S[27]), .CO(
        C[28]) );
  FA_5092 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_5091 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_5090 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_5089 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_5121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_5122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_5127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5136 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_164 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_5151 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_5150 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_5149 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_5148 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_5147 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_5146 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_5145 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_5144 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_5143 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_5142 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_5141 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_5140 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_5139 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_5138 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_5137 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_5136 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_5135 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_5134 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_5133 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_5132 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_5131 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_5130 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_5129 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_5128 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_5127 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_5126 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(1'b0), .S(S[26]), .CO(
        C[27]) );
  FA_5125 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_5124 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_5123 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_5122 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_5121 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_5153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_5154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_5160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5168 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_165 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_5183 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_5182 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_5181 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_5180 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_5179 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_5178 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_5177 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_5176 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_5175 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_5174 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_5173 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_5172 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_5171 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_5170 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_5169 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_5168 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_5167 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_5166 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_5165 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_5164 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_5163 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_5162 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_5161 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_5160 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_5159 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(1'b0), .S(S[25]), .CO(
        C[26]) );
  FA_5158 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_5157 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_5156 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_5155 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_5154 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_5153 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_5185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_5186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_5193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5200 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_166 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_5215 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_5214 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_5213 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_5212 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_5211 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_5210 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_5209 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_5208 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_5207 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_5206 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_5205 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_5204 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_5203 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_5202 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_5201 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_5200 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_5199 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_5198 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_5197 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_5196 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_5195 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_5194 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_5193 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_5192 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(1'b0), .S(S[24]), .CO(
        C[25]) );
  FA_5191 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_5190 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_5189 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_5188 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_5187 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_5186 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_5185 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_5217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_5218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_5226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5232 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_167 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_5247 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_5246 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_5245 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_5244 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_5243 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_5242 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_5241 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_5240 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_5239 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_5238 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_5237 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_5236 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_5235 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_5234 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_5233 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_5232 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_5231 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_5230 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_5229 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_5228 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_5227 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_5226 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_5225 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(1'b0), .S(S[23]), .CO(
        C[24]) );
  FA_5224 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_5223 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_5222 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_5221 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_5220 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_5219 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_5218 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_5217 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_5249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_5250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_5259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5264 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_168 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_5279 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_5278 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_5277 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_5276 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_5275 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_5274 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_5273 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_5272 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_5271 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_5270 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_5269 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_5268 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_5267 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_5266 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_5265 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_5264 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_5263 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_5262 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_5261 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_5260 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_5259 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_5258 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(1'b0), .S(S[22]), .CO(
        C[23]) );
  FA_5257 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_5256 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_5255 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_5254 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_5253 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_5252 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_5251 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_5250 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_5249 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_5281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_5282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_5292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5296 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_169 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_5311 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_5310 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_5309 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_5308 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_5307 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_5306 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_5305 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_5304 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_5303 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_5302 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_5301 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_5300 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_5299 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_5298 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_5297 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_5296 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_5295 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_5294 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_5293 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_5292 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_5291 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(1'b0), .S(S[21]), .CO(
        C[22]) );
  FA_5290 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_5289 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_5288 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_5287 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_5286 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_5285 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_5284 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_5283 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_5282 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_5281 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_5313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_5314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_5325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5328 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_170 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_5343 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_5342 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_5341 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_5340 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_5339 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_5338 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_5337 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_5336 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_5335 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_5334 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_5333 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_5332 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_5331 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_5330 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_5329 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_5328 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_5327 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_5326 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_5325 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_5324 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(1'b0), .S(S[20]), .CO(
        C[21]) );
  FA_5323 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_5322 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_5321 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_5320 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_5319 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_5318 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_5317 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_5316 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_5315 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_5314 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_5313 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_5345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_5346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_5358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5360 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_171 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_5375 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_5374 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_5373 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_5372 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_5371 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_5370 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_5369 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_5368 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_5367 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_5366 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_5365 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_5364 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_5363 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_5362 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_5361 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_5360 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_5359 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_5358 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_5357 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(1'b0), .S(S[19]), .CO(
        C[20]) );
  FA_5356 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_5355 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_5354 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_5353 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_5352 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_5351 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_5350 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_5349 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_5348 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_5347 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_5346 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_5345 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_5377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_5378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_5391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5392 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_172 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_5407 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_5406 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_5405 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_5404 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_5403 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_5402 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_5401 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_5400 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_5399 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_5398 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_5397 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_5396 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_5395 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_5394 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_5393 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_5392 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_5391 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_5390 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(1'b0), .S(S[18]), .CO(
        C[19]) );
  FA_5389 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_5388 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_5387 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_5386 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_5385 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_5384 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_5383 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_5382 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_5381 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_5380 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_5379 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_5378 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_5377 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_5409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_5410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_5424 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_173 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_5439 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_5438 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_5437 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_5436 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_5435 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_5434 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_5433 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_5432 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_5431 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_5430 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_5429 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_5428 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_5427 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_5426 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_5425 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_5424 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_5423 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(1'b0), .S(S[17]), .CO(
        C[18]) );
  FA_5422 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_5421 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_5420 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_5419 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_5418 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_5417 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_5416 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_5415 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_5414 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_5413 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_5412 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_5411 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_5410 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_5409 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_5441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_5442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5456 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_5457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_174 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_5471 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_5470 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_5469 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_5468 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_5467 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_5466 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_5465 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_5464 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_5463 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_5462 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_5461 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_5460 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_5459 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_5458 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_5457 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_5456 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(1'b0), .S(S[16]), .CO(
        C[17]) );
  FA_5455 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_5454 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_5453 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_5452 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_5451 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_5450 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_5449 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_5448 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_5447 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_5446 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_5445 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_5444 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_5443 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_5442 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_5441 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_5473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_5474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5488 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_5490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_175 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_5503 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_5502 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_5501 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_5500 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_5499 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_5498 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_5497 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_5496 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_5495 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_5494 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_5493 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_5492 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_5491 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_5490 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_5489 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(1'b0), .S(S[15]), .CO(
        C[16]) );
  FA_5488 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_5487 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_5486 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_5485 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_5484 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_5483 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_5482 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_5481 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_5480 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_5479 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_5478 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_5477 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_5476 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_5475 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_5474 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_5473 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_5505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_5506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5512 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5513 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5514 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5515 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5516 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5517 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5518 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5519 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5520 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5521 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5522 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_5523 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5524 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5525 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5526 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5527 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5528 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5529 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5530 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5531 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5532 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5533 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5534 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5535 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_176 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_5535 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_5534 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_5533 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_5532 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_5531 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_5530 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_5529 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_5528 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_5527 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_5526 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_5525 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_5524 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_5523 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_5522 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(1'b0), .S(S[14]), .CO(
        C[15]) );
  FA_5521 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_5520 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_5519 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_5518 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_5517 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_5516 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_5515 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_5514 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_5513 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_5512 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_5511 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_5510 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_5509 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_5508 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_5507 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_5506 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_5505 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_5537 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_5538 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5539 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5540 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5541 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5542 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5543 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5544 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5545 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5546 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5547 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5548 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5549 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5550 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5551 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5552 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5553 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5554 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5555 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_5556 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5557 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5558 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5559 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5560 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5561 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5562 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5563 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5564 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5565 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5566 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5567 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_177 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_5567 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_5566 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_5565 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_5564 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_5563 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_5562 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_5561 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_5560 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_5559 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_5558 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_5557 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_5556 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_5555 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(1'b0), .S(S[13]), .CO(
        C[14]) );
  FA_5554 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_5553 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_5552 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_5551 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_5550 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_5549 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_5548 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_5547 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_5546 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_5545 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_5544 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_5543 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_5542 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_5541 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_5540 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_5539 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_5538 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_5537 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_5569 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_5570 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5571 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5572 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5573 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5574 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5575 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5576 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5577 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5578 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5579 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5580 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5581 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5582 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5583 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5584 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5585 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5586 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5587 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5588 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_5589 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5590 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5591 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5592 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5593 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5594 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5595 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5596 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5597 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5598 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5599 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_178 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_5599 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_5598 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_5597 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_5596 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_5595 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_5594 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_5593 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_5592 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_5591 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_5590 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_5589 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_5588 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(1'b0), .S(S[12]), .CO(
        C[13]) );
  FA_5587 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_5586 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_5585 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_5584 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_5583 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_5582 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_5581 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_5580 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_5579 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_5578 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_5577 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_5576 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_5575 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_5574 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_5573 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_5572 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_5571 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_5570 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_5569 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_5601 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_5602 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5603 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5604 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5605 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5606 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5607 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5608 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5609 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5610 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5611 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5612 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5613 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5614 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5615 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5616 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5617 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5618 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5619 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5620 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5621 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_5622 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5623 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5624 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5625 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5626 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5627 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5628 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5629 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5630 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5631 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_179 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_5631 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_5630 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_5629 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_5628 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_5627 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_5626 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_5625 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_5624 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_5623 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_5622 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_5621 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(1'b0), .S(S[11]), .CO(
        C[12]) );
  FA_5620 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_5619 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_5618 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_5617 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_5616 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_5615 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_5614 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_5613 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_5612 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_5611 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_5610 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_5609 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_5608 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_5607 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_5606 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_5605 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_5604 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_5603 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_5602 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_5601 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_5633 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_5634 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5635 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5636 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5637 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5638 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5639 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5640 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5641 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5642 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5643 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5644 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5645 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5646 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5647 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5648 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5649 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5650 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5651 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5652 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5653 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5654 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_5655 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5656 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5657 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5658 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5659 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5660 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5661 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5662 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5663 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_180 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_5663 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_5662 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_5661 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_5660 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_5659 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_5658 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_5657 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_5656 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_5655 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_5654 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(1'b0), .S(S[10]), .CO(
        C[11]) );
  FA_5653 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_5652 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_5651 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_5650 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_5649 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_5648 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_5647 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_5646 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_5645 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_5644 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_5643 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_5642 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_5641 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_5640 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_5639 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_5638 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_5637 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_5636 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_5635 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_5634 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_5633 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_5665 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_5666 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5667 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5668 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5669 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5670 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5671 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5672 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5673 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5674 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5675 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5676 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5677 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5678 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5679 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5680 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5681 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5682 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5683 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5684 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5685 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5686 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5687 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_5688 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5689 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5690 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5691 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5692 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5693 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5694 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5695 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_181 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_5695 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_5694 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_5693 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_5692 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_5691 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_5690 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_5689 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_5688 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_5687 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(1'b0), .S(S[9]), .CO(C[10]) );
  FA_5686 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_5685 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_5684 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_5683 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_5682 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_5681 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_5680 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_5679 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_5678 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_5677 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_5676 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_5675 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_5674 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_5673 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_5672 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_5671 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_5670 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_5669 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_5668 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_5667 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_5666 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_5665 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_5697 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_5698 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5699 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5700 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5701 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5702 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5703 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5704 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5705 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5706 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5707 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5708 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5709 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5710 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5711 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5712 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5713 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5714 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5715 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5716 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5717 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5718 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5719 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5720 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_5721 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5722 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5723 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5724 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5725 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5726 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5727 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_182 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_5727 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_5726 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_5725 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_5724 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_5723 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_5722 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_5721 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_5720 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(1'b0), .S(S[8]), .CO(C[9])
         );
  FA_5719 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_5718 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_5717 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_5716 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_5715 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_5714 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_5713 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_5712 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_5711 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_5710 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_5709 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_5708 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_5707 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_5706 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_5705 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_5704 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_5703 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_5702 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_5701 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_5700 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_5699 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_5698 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_5697 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_5729 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_5730 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5731 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5732 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5733 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5734 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5735 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5736 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5737 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5738 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5739 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5740 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5741 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5742 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5743 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5744 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5745 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5746 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5747 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5748 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5749 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5750 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5751 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5752 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5753 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_5754 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5755 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5756 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5757 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5758 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5759 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_183 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_5759 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_5758 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_5757 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_5756 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_5755 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_5754 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_5753 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(1'b0), .S(S[7]), .CO(C[8])
         );
  FA_5752 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_5751 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_5750 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_5749 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_5748 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_5747 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_5746 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_5745 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_5744 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_5743 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_5742 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_5741 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_5740 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_5739 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_5738 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_5737 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_5736 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_5735 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_5734 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_5733 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_5732 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_5731 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_5730 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_5729 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_5761 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_5762 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5763 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5764 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5765 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5766 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5767 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5768 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5769 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5770 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5771 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5772 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5773 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5774 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5775 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5776 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5777 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5778 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5779 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5780 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5781 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5782 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5783 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5784 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5785 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5786 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_5787 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5788 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5789 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5790 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5791 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_184 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_5791 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_5790 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_5789 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_5788 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_5787 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_5786 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(1'b0), .S(S[6]), .CO(C[7])
         );
  FA_5785 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_5784 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_5783 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_5782 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_5781 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_5780 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_5779 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_5778 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_5777 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_5776 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_5775 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_5774 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_5773 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_5772 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_5771 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_5770 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_5769 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_5768 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_5767 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_5766 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_5765 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_5764 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_5763 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_5762 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_5761 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_5793 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_5794 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5795 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5796 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5797 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5798 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5799 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5800 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5801 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5802 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5803 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5804 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5805 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5806 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5807 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5808 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5809 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5810 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5811 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5812 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5813 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5814 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5815 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5816 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5817 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5818 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5819 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_5820 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5821 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5822 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5823 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_185 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_5823 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_5822 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_5821 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_5820 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_5819 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(1'b0), .S(S[5]), .CO(C[6])
         );
  FA_5818 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_5817 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_5816 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_5815 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_5814 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_5813 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_5812 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_5811 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_5810 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_5809 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_5808 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_5807 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_5806 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_5805 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_5804 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_5803 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_5802 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_5801 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_5800 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_5799 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_5798 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_5797 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_5796 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_5795 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_5794 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_5793 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_5825 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_5826 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5827 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5828 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5829 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5830 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5831 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5832 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5833 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5834 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5835 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5836 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5837 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5838 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5839 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5840 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5841 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5842 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5843 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5844 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5845 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5846 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5847 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5848 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5849 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5850 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5851 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5852 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_5853 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5854 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5855 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_186 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_5855 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_5854 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_5853 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_5852 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(1'b0), .S(S[4]), .CO(C[5])
         );
  FA_5851 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_5850 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_5849 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_5848 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_5847 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_5846 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_5845 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_5844 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_5843 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_5842 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_5841 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_5840 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_5839 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_5838 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_5837 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_5836 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_5835 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_5834 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_5833 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_5832 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_5831 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_5830 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_5829 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_5828 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_5827 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_5826 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_5825 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_5857 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_5858 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5859 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5860 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5861 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5862 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5863 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5864 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5865 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5866 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5867 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5868 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5869 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5870 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5871 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5872 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5873 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5874 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5875 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5876 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5877 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5878 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5879 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5880 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5881 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5882 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5883 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5884 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5885 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_5886 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5887 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_187 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_5887 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_5886 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_5885 \FAINST[3].FA_  ( .A(A[3]), .B(B[3]), .CI(1'b0), .S(S[3]), .CO(C[4])
         );
  FA_5884 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_5883 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_5882 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_5881 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_5880 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_5879 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_5878 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_5877 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_5876 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_5875 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_5874 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_5873 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_5872 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_5871 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_5870 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_5869 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_5868 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_5867 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_5866 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_5865 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_5864 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_5863 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_5862 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_5861 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_5860 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_5859 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_5858 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_5857 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_5889 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_5890 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5891 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5892 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5893 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5894 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5895 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5896 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5897 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5898 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5899 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5900 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5901 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5902 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5903 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5904 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5905 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5906 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5907 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5908 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5909 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5910 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5911 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5912 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5913 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5914 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5915 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5916 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5917 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5918 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_5919 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_188 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_5919 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_5918 \FAINST[2].FA_  ( .A(A[2]), .B(B[2]), .CI(1'b0), .S(S[2]), .CO(C[3])
         );
  FA_5917 \FAINST[3].FA_  ( .A(A[3]), .B(B[3]), .CI(C[3]), .S(S[3]), .CO(C[4])
         );
  FA_5916 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_5915 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_5914 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_5913 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_5912 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_5911 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_5910 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_5909 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_5908 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_5907 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_5906 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_5905 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_5904 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_5903 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_5902 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_5901 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_5900 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_5899 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_5898 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_5897 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_5896 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_5895 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_5894 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_5893 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_5892 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_5891 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_5890 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_5889 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_5921 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_5922 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_5923 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_5924 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_5925 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_5926 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_5927 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_5928 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_5929 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_5930 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_5931 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_5932 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_5933 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_5934 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_5935 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_5936 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_5937 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_5938 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_5939 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_5940 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_5941 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_5942 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_5943 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_5944 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_5945 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_5946 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_5947 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_5948 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_5949 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_5950 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_5951 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module ADD_N32_189 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;


  FA_5951 \FAINST[1].FA_  ( .A(A[1]), .B(1'b0), .CI(1'b0), .S(S[1]) );
  FA_5950 \FAINST[2].FA_  ( .A(A[2]), .B(1'b0), .CI(1'b0), .S(S[2]) );
  FA_5949 \FAINST[3].FA_  ( .A(A[3]), .B(1'b0), .CI(1'b0), .S(S[3]) );
  FA_5948 \FAINST[4].FA_  ( .A(A[4]), .B(1'b0), .CI(1'b0), .S(S[4]) );
  FA_5947 \FAINST[5].FA_  ( .A(A[5]), .B(1'b0), .CI(1'b0), .S(S[5]) );
  FA_5946 \FAINST[6].FA_  ( .A(A[6]), .B(1'b0), .CI(1'b0), .S(S[6]) );
  FA_5945 \FAINST[7].FA_  ( .A(A[7]), .B(1'b0), .CI(1'b0), .S(S[7]) );
  FA_5944 \FAINST[8].FA_  ( .A(A[8]), .B(1'b0), .CI(1'b0), .S(S[8]) );
  FA_5943 \FAINST[9].FA_  ( .A(A[9]), .B(1'b0), .CI(1'b0), .S(S[9]) );
  FA_5942 \FAINST[10].FA_  ( .A(A[10]), .B(1'b0), .CI(1'b0), .S(S[10]) );
  FA_5941 \FAINST[11].FA_  ( .A(A[11]), .B(1'b0), .CI(1'b0), .S(S[11]) );
  FA_5940 \FAINST[12].FA_  ( .A(A[12]), .B(1'b0), .CI(1'b0), .S(S[12]) );
  FA_5939 \FAINST[13].FA_  ( .A(A[13]), .B(1'b0), .CI(1'b0), .S(S[13]) );
  FA_5938 \FAINST[14].FA_  ( .A(A[14]), .B(1'b0), .CI(1'b0), .S(S[14]) );
  FA_5937 \FAINST[15].FA_  ( .A(A[15]), .B(1'b0), .CI(1'b0), .S(S[15]) );
  FA_5936 \FAINST[16].FA_  ( .A(A[16]), .B(1'b0), .CI(1'b0), .S(S[16]) );
  FA_5935 \FAINST[17].FA_  ( .A(A[17]), .B(1'b0), .CI(1'b0), .S(S[17]) );
  FA_5934 \FAINST[18].FA_  ( .A(A[18]), .B(1'b0), .CI(1'b0), .S(S[18]) );
  FA_5933 \FAINST[19].FA_  ( .A(A[19]), .B(1'b0), .CI(1'b0), .S(S[19]) );
  FA_5932 \FAINST[20].FA_  ( .A(A[20]), .B(1'b0), .CI(1'b0), .S(S[20]) );
  FA_5931 \FAINST[21].FA_  ( .A(A[21]), .B(1'b0), .CI(1'b0), .S(S[21]) );
  FA_5930 \FAINST[22].FA_  ( .A(A[22]), .B(1'b0), .CI(1'b0), .S(S[22]) );
  FA_5929 \FAINST[23].FA_  ( .A(A[23]), .B(1'b0), .CI(1'b0), .S(S[23]) );
  FA_5928 \FAINST[24].FA_  ( .A(A[24]), .B(1'b0), .CI(1'b0), .S(S[24]) );
  FA_5927 \FAINST[25].FA_  ( .A(A[25]), .B(1'b0), .CI(1'b0), .S(S[25]) );
  FA_5926 \FAINST[26].FA_  ( .A(A[26]), .B(1'b0), .CI(1'b0), .S(S[26]) );
  FA_5925 \FAINST[27].FA_  ( .A(A[27]), .B(1'b0), .CI(1'b0), .S(S[27]) );
  FA_5924 \FAINST[28].FA_  ( .A(A[28]), .B(1'b0), .CI(1'b0), .S(S[28]) );
  FA_5923 \FAINST[29].FA_  ( .A(A[29]), .B(1'b0), .CI(1'b0), .S(S[29]) );
  FA_5922 \FAINST[30].FA_  ( .A(A[30]), .B(1'b0), .CI(1'b0), .S(S[30]) );
  FA_5921 \FAINST[31].FA_  ( .A(A[31]), .B(1'b0), .CI(1'b0), .S(S[31]) );
endmodule


module MULT_N32_6 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   \w[31][31] , \w[31][30] , \w[31][29] , \w[31][28] , \w[31][27] ,
         \w[31][26] , \w[31][25] , \w[31][24] , \w[31][23] , \w[31][22] ,
         \w[31][21] , \w[31][20] , \w[31][19] , \w[31][18] , \w[31][17] ,
         \w[31][16] , \w[31][15] , \w[31][14] , \w[31][13] , \w[31][12] ,
         \w[31][11] , \w[31][10] , \w[31][9] , \w[31][8] , \w[31][7] ,
         \w[31][6] , \w[31][5] , \w[31][4] , \w[31][3] , \w[31][2] ,
         \w[31][1] , \w[30][31] , \w[30][30] , \w[30][29] , \w[30][28] ,
         \w[30][27] , \w[30][26] , \w[30][25] , \w[30][24] , \w[30][23] ,
         \w[30][22] , \w[30][21] , \w[30][20] , \w[30][19] , \w[30][18] ,
         \w[30][17] , \w[30][16] , \w[30][15] , \w[30][14] , \w[30][13] ,
         \w[30][12] , \w[30][11] , \w[30][10] , \w[30][9] , \w[30][8] ,
         \w[30][7] , \w[30][6] , \w[30][5] , \w[30][4] , \w[30][3] ,
         \w[30][2] , \w[30][1] , \w[29][31] , \w[29][30] , \w[29][29] ,
         \w[29][28] , \w[29][27] , \w[29][26] , \w[29][25] , \w[29][24] ,
         \w[29][23] , \w[29][22] , \w[29][21] , \w[29][20] , \w[29][19] ,
         \w[29][18] , \w[29][17] , \w[29][16] , \w[29][15] , \w[29][14] ,
         \w[29][13] , \w[29][12] , \w[29][11] , \w[29][10] , \w[29][9] ,
         \w[29][8] , \w[29][7] , \w[29][6] , \w[29][5] , \w[29][4] ,
         \w[29][3] , \w[29][2] , \w[29][1] , \w[28][31] , \w[28][30] ,
         \w[28][29] , \w[28][28] , \w[28][27] , \w[28][26] , \w[28][25] ,
         \w[28][24] , \w[28][23] , \w[28][22] , \w[28][21] , \w[28][20] ,
         \w[28][19] , \w[28][18] , \w[28][17] , \w[28][16] , \w[28][15] ,
         \w[28][14] , \w[28][13] , \w[28][12] , \w[28][11] , \w[28][10] ,
         \w[28][9] , \w[28][8] , \w[28][7] , \w[28][6] , \w[28][5] ,
         \w[28][4] , \w[28][3] , \w[28][2] , \w[28][1] , \w[27][31] ,
         \w[27][30] , \w[27][29] , \w[27][28] , \w[27][27] , \w[27][26] ,
         \w[27][25] , \w[27][24] , \w[27][23] , \w[27][22] , \w[27][21] ,
         \w[27][20] , \w[27][19] , \w[27][18] , \w[27][17] , \w[27][16] ,
         \w[27][15] , \w[27][14] , \w[27][13] , \w[27][12] , \w[27][11] ,
         \w[27][10] , \w[27][9] , \w[27][8] , \w[27][7] , \w[27][6] ,
         \w[27][5] , \w[27][4] , \w[27][3] , \w[27][2] , \w[27][1] ,
         \w[26][31] , \w[26][30] , \w[26][29] , \w[26][28] , \w[26][27] ,
         \w[26][26] , \w[26][25] , \w[26][24] , \w[26][23] , \w[26][22] ,
         \w[26][21] , \w[26][20] , \w[26][19] , \w[26][18] , \w[26][17] ,
         \w[26][16] , \w[26][15] , \w[26][14] , \w[26][13] , \w[26][12] ,
         \w[26][11] , \w[26][10] , \w[26][9] , \w[26][8] , \w[26][7] ,
         \w[26][6] , \w[26][5] , \w[26][4] , \w[26][3] , \w[26][2] ,
         \w[26][1] , \w[25][31] , \w[25][30] , \w[25][29] , \w[25][28] ,
         \w[25][27] , \w[25][26] , \w[25][25] , \w[25][24] , \w[25][23] ,
         \w[25][22] , \w[25][21] , \w[25][20] , \w[25][19] , \w[25][18] ,
         \w[25][17] , \w[25][16] , \w[25][15] , \w[25][14] , \w[25][13] ,
         \w[25][12] , \w[25][11] , \w[25][10] , \w[25][9] , \w[25][8] ,
         \w[25][7] , \w[25][6] , \w[25][5] , \w[25][4] , \w[25][3] ,
         \w[25][2] , \w[25][1] , \w[24][31] , \w[24][30] , \w[24][29] ,
         \w[24][28] , \w[24][27] , \w[24][26] , \w[24][25] , \w[24][24] ,
         \w[24][23] , \w[24][22] , \w[24][21] , \w[24][20] , \w[24][19] ,
         \w[24][18] , \w[24][17] , \w[24][16] , \w[24][15] , \w[24][14] ,
         \w[24][13] , \w[24][12] , \w[24][11] , \w[24][10] , \w[24][9] ,
         \w[24][8] , \w[24][7] , \w[24][6] , \w[24][5] , \w[24][4] ,
         \w[24][3] , \w[24][2] , \w[24][1] , \w[23][31] , \w[23][30] ,
         \w[23][29] , \w[23][28] , \w[23][27] , \w[23][26] , \w[23][25] ,
         \w[23][24] , \w[23][23] , \w[23][22] , \w[23][21] , \w[23][20] ,
         \w[23][19] , \w[23][18] , \w[23][17] , \w[23][16] , \w[23][15] ,
         \w[23][14] , \w[23][13] , \w[23][12] , \w[23][11] , \w[23][10] ,
         \w[23][9] , \w[23][8] , \w[23][7] , \w[23][6] , \w[23][5] ,
         \w[23][4] , \w[23][3] , \w[23][2] , \w[23][1] , \w[22][31] ,
         \w[22][30] , \w[22][29] , \w[22][28] , \w[22][27] , \w[22][26] ,
         \w[22][25] , \w[22][24] , \w[22][23] , \w[22][22] , \w[22][21] ,
         \w[22][20] , \w[22][19] , \w[22][18] , \w[22][17] , \w[22][16] ,
         \w[22][15] , \w[22][14] , \w[22][13] , \w[22][12] , \w[22][11] ,
         \w[22][10] , \w[22][9] , \w[22][8] , \w[22][7] , \w[22][6] ,
         \w[22][5] , \w[22][4] , \w[22][3] , \w[22][2] , \w[22][1] ,
         \w[21][31] , \w[21][30] , \w[21][29] , \w[21][28] , \w[21][27] ,
         \w[21][26] , \w[21][25] , \w[21][24] , \w[21][23] , \w[21][22] ,
         \w[21][21] , \w[21][20] , \w[21][19] , \w[21][18] , \w[21][17] ,
         \w[21][16] , \w[21][15] , \w[21][14] , \w[21][13] , \w[21][12] ,
         \w[21][11] , \w[21][10] , \w[21][9] , \w[21][8] , \w[21][7] ,
         \w[21][6] , \w[21][5] , \w[21][4] , \w[21][3] , \w[21][2] ,
         \w[21][1] , \w[20][31] , \w[20][30] , \w[20][29] , \w[20][28] ,
         \w[20][27] , \w[20][26] , \w[20][25] , \w[20][24] , \w[20][23] ,
         \w[20][22] , \w[20][21] , \w[20][20] , \w[20][19] , \w[20][18] ,
         \w[20][17] , \w[20][16] , \w[20][15] , \w[20][14] , \w[20][13] ,
         \w[20][12] , \w[20][11] , \w[20][10] , \w[20][9] , \w[20][8] ,
         \w[20][7] , \w[20][6] , \w[20][5] , \w[20][4] , \w[20][3] ,
         \w[20][2] , \w[20][1] , \w[19][31] , \w[19][30] , \w[19][29] ,
         \w[19][28] , \w[19][27] , \w[19][26] , \w[19][25] , \w[19][24] ,
         \w[19][23] , \w[19][22] , \w[19][21] , \w[19][20] , \w[19][19] ,
         \w[19][18] , \w[19][17] , \w[19][16] , \w[19][15] , \w[19][14] ,
         \w[19][13] , \w[19][12] , \w[19][11] , \w[19][10] , \w[19][9] ,
         \w[19][8] , \w[19][7] , \w[19][6] , \w[19][5] , \w[19][4] ,
         \w[19][3] , \w[19][2] , \w[19][1] , \w[18][31] , \w[18][30] ,
         \w[18][29] , \w[18][28] , \w[18][27] , \w[18][26] , \w[18][25] ,
         \w[18][24] , \w[18][23] , \w[18][22] , \w[18][21] , \w[18][20] ,
         \w[18][19] , \w[18][18] , \w[18][17] , \w[18][16] , \w[18][15] ,
         \w[18][14] , \w[18][13] , \w[18][12] , \w[18][11] , \w[18][10] ,
         \w[18][9] , \w[18][8] , \w[18][7] , \w[18][6] , \w[18][5] ,
         \w[18][4] , \w[18][3] , \w[18][2] , \w[18][1] , \w[17][31] ,
         \w[17][30] , \w[17][29] , \w[17][28] , \w[17][27] , \w[17][26] ,
         \w[17][25] , \w[17][24] , \w[17][23] , \w[17][22] , \w[17][21] ,
         \w[17][20] , \w[17][19] , \w[17][18] , \w[17][17] , \w[17][16] ,
         \w[17][15] , \w[17][14] , \w[17][13] , \w[17][12] , \w[17][11] ,
         \w[17][10] , \w[17][9] , \w[17][8] , \w[17][7] , \w[17][6] ,
         \w[17][5] , \w[17][4] , \w[17][3] , \w[17][2] , \w[17][1] ,
         \w[16][31] , \w[16][30] , \w[16][29] , \w[16][28] , \w[16][27] ,
         \w[16][26] , \w[16][25] , \w[16][24] , \w[16][23] , \w[16][22] ,
         \w[16][21] , \w[16][20] , \w[16][19] , \w[16][18] , \w[16][17] ,
         \w[16][16] , \w[16][15] , \w[16][14] , \w[16][13] , \w[16][12] ,
         \w[16][11] , \w[16][10] , \w[16][9] , \w[16][8] , \w[16][7] ,
         \w[16][6] , \w[16][5] , \w[16][4] , \w[16][3] , \w[16][2] ,
         \w[16][1] , \w[15][31] , \w[15][30] , \w[15][29] , \w[15][28] ,
         \w[15][27] , \w[15][26] , \w[15][25] , \w[15][24] , \w[15][23] ,
         \w[15][22] , \w[15][21] , \w[15][20] , \w[15][19] , \w[15][18] ,
         \w[15][17] , \w[15][16] , \w[15][15] , \w[15][14] , \w[15][13] ,
         \w[15][12] , \w[15][11] , \w[15][10] , \w[15][9] , \w[15][8] ,
         \w[15][7] , \w[15][6] , \w[15][5] , \w[15][4] , \w[15][3] ,
         \w[15][2] , \w[15][1] , \w[14][31] , \w[14][30] , \w[14][29] ,
         \w[14][28] , \w[14][27] , \w[14][26] , \w[14][25] , \w[14][24] ,
         \w[14][23] , \w[14][22] , \w[14][21] , \w[14][20] , \w[14][19] ,
         \w[14][18] , \w[14][17] , \w[14][16] , \w[14][15] , \w[14][14] ,
         \w[14][13] , \w[14][12] , \w[14][11] , \w[14][10] , \w[14][9] ,
         \w[14][8] , \w[14][7] , \w[14][6] , \w[14][5] , \w[14][4] ,
         \w[14][3] , \w[14][2] , \w[14][1] , \w[13][31] , \w[13][30] ,
         \w[13][29] , \w[13][28] , \w[13][27] , \w[13][26] , \w[13][25] ,
         \w[13][24] , \w[13][23] , \w[13][22] , \w[13][21] , \w[13][20] ,
         \w[13][19] , \w[13][18] , \w[13][17] , \w[13][16] , \w[13][15] ,
         \w[13][14] , \w[13][13] , \w[13][12] , \w[13][11] , \w[13][10] ,
         \w[13][9] , \w[13][8] , \w[13][7] , \w[13][6] , \w[13][5] ,
         \w[13][4] , \w[13][3] , \w[13][2] , \w[13][1] , \w[12][31] ,
         \w[12][30] , \w[12][29] , \w[12][28] , \w[12][27] , \w[12][26] ,
         \w[12][25] , \w[12][24] , \w[12][23] , \w[12][22] , \w[12][21] ,
         \w[12][20] , \w[12][19] , \w[12][18] , \w[12][17] , \w[12][16] ,
         \w[12][15] , \w[12][14] , \w[12][13] , \w[12][12] , \w[12][11] ,
         \w[12][10] , \w[12][9] , \w[12][8] , \w[12][7] , \w[12][6] ,
         \w[12][5] , \w[12][4] , \w[12][3] , \w[12][2] , \w[12][1] ,
         \w[11][31] , \w[11][30] , \w[11][29] , \w[11][28] , \w[11][27] ,
         \w[11][26] , \w[11][25] , \w[11][24] , \w[11][23] , \w[11][22] ,
         \w[11][21] , \w[11][20] , \w[11][19] , \w[11][18] , \w[11][17] ,
         \w[11][16] , \w[11][15] , \w[11][14] , \w[11][13] , \w[11][12] ,
         \w[11][11] , \w[11][10] , \w[11][9] , \w[11][8] , \w[11][7] ,
         \w[11][6] , \w[11][5] , \w[11][4] , \w[11][3] , \w[11][2] ,
         \w[11][1] , \w[10][31] , \w[10][30] , \w[10][29] , \w[10][28] ,
         \w[10][27] , \w[10][26] , \w[10][25] , \w[10][24] , \w[10][23] ,
         \w[10][22] , \w[10][21] , \w[10][20] , \w[10][19] , \w[10][18] ,
         \w[10][17] , \w[10][16] , \w[10][15] , \w[10][14] , \w[10][13] ,
         \w[10][12] , \w[10][11] , \w[10][10] , \w[10][9] , \w[10][8] ,
         \w[10][7] , \w[10][6] , \w[10][5] , \w[10][4] , \w[10][3] ,
         \w[10][2] , \w[10][1] , \w[9][31] , \w[9][30] , \w[9][29] ,
         \w[9][28] , \w[9][27] , \w[9][26] , \w[9][25] , \w[9][24] ,
         \w[9][23] , \w[9][22] , \w[9][21] , \w[9][20] , \w[9][19] ,
         \w[9][18] , \w[9][17] , \w[9][16] , \w[9][15] , \w[9][14] ,
         \w[9][13] , \w[9][12] , \w[9][11] , \w[9][10] , \w[9][9] , \w[9][8] ,
         \w[9][7] , \w[9][6] , \w[9][5] , \w[9][4] , \w[9][3] , \w[9][2] ,
         \w[9][1] , \w[8][31] , \w[8][30] , \w[8][29] , \w[8][28] , \w[8][27] ,
         \w[8][26] , \w[8][25] , \w[8][24] , \w[8][23] , \w[8][22] ,
         \w[8][21] , \w[8][20] , \w[8][19] , \w[8][18] , \w[8][17] ,
         \w[8][16] , \w[8][15] , \w[8][14] , \w[8][13] , \w[8][12] ,
         \w[8][11] , \w[8][10] , \w[8][9] , \w[8][8] , \w[8][7] , \w[8][6] ,
         \w[8][5] , \w[8][4] , \w[8][3] , \w[8][2] , \w[8][1] , \w[7][31] ,
         \w[7][30] , \w[7][29] , \w[7][28] , \w[7][27] , \w[7][26] ,
         \w[7][25] , \w[7][24] , \w[7][23] , \w[7][22] , \w[7][21] ,
         \w[7][20] , \w[7][19] , \w[7][18] , \w[7][17] , \w[7][16] ,
         \w[7][15] , \w[7][14] , \w[7][13] , \w[7][12] , \w[7][11] ,
         \w[7][10] , \w[7][9] , \w[7][8] , \w[7][7] , \w[7][6] , \w[7][5] ,
         \w[7][4] , \w[7][3] , \w[7][2] , \w[7][1] , \w[6][31] , \w[6][30] ,
         \w[6][29] , \w[6][28] , \w[6][27] , \w[6][26] , \w[6][25] ,
         \w[6][24] , \w[6][23] , \w[6][22] , \w[6][21] , \w[6][20] ,
         \w[6][19] , \w[6][18] , \w[6][17] , \w[6][16] , \w[6][15] ,
         \w[6][14] , \w[6][13] , \w[6][12] , \w[6][11] , \w[6][10] , \w[6][9] ,
         \w[6][8] , \w[6][7] , \w[6][6] , \w[6][5] , \w[6][4] , \w[6][3] ,
         \w[6][2] , \w[6][1] , \w[5][31] , \w[5][30] , \w[5][29] , \w[5][28] ,
         \w[5][27] , \w[5][26] , \w[5][25] , \w[5][24] , \w[5][23] ,
         \w[5][22] , \w[5][21] , \w[5][20] , \w[5][19] , \w[5][18] ,
         \w[5][17] , \w[5][16] , \w[5][15] , \w[5][14] , \w[5][13] ,
         \w[5][12] , \w[5][11] , \w[5][10] , \w[5][9] , \w[5][8] , \w[5][7] ,
         \w[5][6] , \w[5][5] , \w[5][4] , \w[5][3] , \w[5][2] , \w[5][1] ,
         \w[4][31] , \w[4][30] , \w[4][29] , \w[4][28] , \w[4][27] ,
         \w[4][26] , \w[4][25] , \w[4][24] , \w[4][23] , \w[4][22] ,
         \w[4][21] , \w[4][20] , \w[4][19] , \w[4][18] , \w[4][17] ,
         \w[4][16] , \w[4][15] , \w[4][14] , \w[4][13] , \w[4][12] ,
         \w[4][11] , \w[4][10] , \w[4][9] , \w[4][8] , \w[4][7] , \w[4][6] ,
         \w[4][5] , \w[4][4] , \w[4][3] , \w[4][2] , \w[4][1] , \w[3][31] ,
         \w[3][30] , \w[3][29] , \w[3][28] , \w[3][27] , \w[3][26] ,
         \w[3][25] , \w[3][24] , \w[3][23] , \w[3][22] , \w[3][21] ,
         \w[3][20] , \w[3][19] , \w[3][18] , \w[3][17] , \w[3][16] ,
         \w[3][15] , \w[3][14] , \w[3][13] , \w[3][12] , \w[3][11] ,
         \w[3][10] , \w[3][9] , \w[3][8] , \w[3][7] , \w[3][6] , \w[3][5] ,
         \w[3][4] , \w[3][3] , \w[3][2] , \w[3][1] , \w[2][31] , \w[2][30] ,
         \w[2][29] , \w[2][28] , \w[2][27] , \w[2][26] , \w[2][25] ,
         \w[2][24] , \w[2][23] , \w[2][22] , \w[2][21] , \w[2][20] ,
         \w[2][19] , \w[2][18] , \w[2][17] , \w[2][16] , \w[2][15] ,
         \w[2][14] , \w[2][13] , \w[2][12] , \w[2][11] , \w[2][10] , \w[2][9] ,
         \w[2][8] , \w[2][7] , \w[2][6] , \w[2][5] , \w[2][4] , \w[2][3] ,
         \w[2][2] , \w[2][1] , \_0_net_[31] , \_0_net_[30] , \_0_net_[29] ,
         \_0_net_[28] , \_0_net_[27] , \_0_net_[26] , \_0_net_[25] ,
         \_0_net_[24] , \_0_net_[23] , \_0_net_[22] , \_0_net_[21] ,
         \_0_net_[20] , \_0_net_[19] , \_0_net_[18] , \_0_net_[17] ,
         \_0_net_[16] , \_0_net_[15] , \_0_net_[14] , \_0_net_[13] ,
         \_0_net_[12] , \_0_net_[11] , \_0_net_[10] , \_0_net_[9] ,
         \_0_net_[8] , \_0_net_[7] , \_0_net_[6] , \_0_net_[5] , \_0_net_[4] ,
         \_0_net_[3] , \_0_net_[2] , \_0_net_[1] , \_2_net_[31] ,
         \_2_net_[30] , \_2_net_[29] , \_2_net_[28] , \_2_net_[27] ,
         \_2_net_[26] , \_2_net_[25] , \_2_net_[24] , \_2_net_[23] ,
         \_2_net_[22] , \_2_net_[21] , \_2_net_[20] , \_2_net_[19] ,
         \_2_net_[18] , \_2_net_[17] , \_2_net_[16] , \_2_net_[15] ,
         \_2_net_[14] , \_2_net_[13] , \_2_net_[12] , \_2_net_[11] ,
         \_2_net_[10] , \_2_net_[9] , \_2_net_[8] , \_2_net_[7] , \_2_net_[6] ,
         \_2_net_[5] , \_2_net_[4] , \_2_net_[3] , \_2_net_[2] , \_4_net_[31] ,
         \_4_net_[30] , \_4_net_[29] , \_4_net_[28] , \_4_net_[27] ,
         \_4_net_[26] , \_4_net_[25] , \_4_net_[24] , \_4_net_[23] ,
         \_4_net_[22] , \_4_net_[21] , \_4_net_[20] , \_4_net_[19] ,
         \_4_net_[18] , \_4_net_[17] , \_4_net_[16] , \_4_net_[15] ,
         \_4_net_[14] , \_4_net_[13] , \_4_net_[12] , \_4_net_[11] ,
         \_4_net_[10] , \_4_net_[9] , \_4_net_[8] , \_4_net_[7] , \_4_net_[6] ,
         \_4_net_[5] , \_4_net_[4] , \_4_net_[3] , \_6_net_[31] ,
         \_6_net_[30] , \_6_net_[29] , \_6_net_[28] , \_6_net_[27] ,
         \_6_net_[26] , \_6_net_[25] , \_6_net_[24] , \_6_net_[23] ,
         \_6_net_[22] , \_6_net_[21] , \_6_net_[20] , \_6_net_[19] ,
         \_6_net_[18] , \_6_net_[17] , \_6_net_[16] , \_6_net_[15] ,
         \_6_net_[14] , \_6_net_[13] , \_6_net_[12] , \_6_net_[11] ,
         \_6_net_[10] , \_6_net_[9] , \_6_net_[8] , \_6_net_[7] , \_6_net_[6] ,
         \_6_net_[5] , \_6_net_[4] , \_8_net_[31] , \_8_net_[30] ,
         \_8_net_[29] , \_8_net_[28] , \_8_net_[27] , \_8_net_[26] ,
         \_8_net_[25] , \_8_net_[24] , \_8_net_[23] , \_8_net_[22] ,
         \_8_net_[21] , \_8_net_[20] , \_8_net_[19] , \_8_net_[18] ,
         \_8_net_[17] , \_8_net_[16] , \_8_net_[15] , \_8_net_[14] ,
         \_8_net_[13] , \_8_net_[12] , \_8_net_[11] , \_8_net_[10] ,
         \_8_net_[9] , \_8_net_[8] , \_8_net_[7] , \_8_net_[6] , \_8_net_[5] ,
         \_10_net_[31] , \_10_net_[30] , \_10_net_[29] , \_10_net_[28] ,
         \_10_net_[27] , \_10_net_[26] , \_10_net_[25] , \_10_net_[24] ,
         \_10_net_[23] , \_10_net_[22] , \_10_net_[21] , \_10_net_[20] ,
         \_10_net_[19] , \_10_net_[18] , \_10_net_[17] , \_10_net_[16] ,
         \_10_net_[15] , \_10_net_[14] , \_10_net_[13] , \_10_net_[12] ,
         \_10_net_[11] , \_10_net_[10] , \_10_net_[9] , \_10_net_[8] ,
         \_10_net_[7] , \_10_net_[6] , \_12_net_[31] , \_12_net_[30] ,
         \_12_net_[29] , \_12_net_[28] , \_12_net_[27] , \_12_net_[26] ,
         \_12_net_[25] , \_12_net_[24] , \_12_net_[23] , \_12_net_[22] ,
         \_12_net_[21] , \_12_net_[20] , \_12_net_[19] , \_12_net_[18] ,
         \_12_net_[17] , \_12_net_[16] , \_12_net_[15] , \_12_net_[14] ,
         \_12_net_[13] , \_12_net_[12] , \_12_net_[11] , \_12_net_[10] ,
         \_12_net_[9] , \_12_net_[8] , \_12_net_[7] , \_14_net_[31] ,
         \_14_net_[30] , \_14_net_[29] , \_14_net_[28] , \_14_net_[27] ,
         \_14_net_[26] , \_14_net_[25] , \_14_net_[24] , \_14_net_[23] ,
         \_14_net_[22] , \_14_net_[21] , \_14_net_[20] , \_14_net_[19] ,
         \_14_net_[18] , \_14_net_[17] , \_14_net_[16] , \_14_net_[15] ,
         \_14_net_[14] , \_14_net_[13] , \_14_net_[12] , \_14_net_[11] ,
         \_14_net_[10] , \_14_net_[9] , \_14_net_[8] , \_16_net_[31] ,
         \_16_net_[30] , \_16_net_[29] , \_16_net_[28] , \_16_net_[27] ,
         \_16_net_[26] , \_16_net_[25] , \_16_net_[24] , \_16_net_[23] ,
         \_16_net_[22] , \_16_net_[21] , \_16_net_[20] , \_16_net_[19] ,
         \_16_net_[18] , \_16_net_[17] , \_16_net_[16] , \_16_net_[15] ,
         \_16_net_[14] , \_16_net_[13] , \_16_net_[12] , \_16_net_[11] ,
         \_16_net_[10] , \_16_net_[9] , \_18_net_[31] , \_18_net_[30] ,
         \_18_net_[29] , \_18_net_[28] , \_18_net_[27] , \_18_net_[26] ,
         \_18_net_[25] , \_18_net_[24] , \_18_net_[23] , \_18_net_[22] ,
         \_18_net_[21] , \_18_net_[20] , \_18_net_[19] , \_18_net_[18] ,
         \_18_net_[17] , \_18_net_[16] , \_18_net_[15] , \_18_net_[14] ,
         \_18_net_[13] , \_18_net_[12] , \_18_net_[11] , \_18_net_[10] ,
         \_20_net_[31] , \_20_net_[30] , \_20_net_[29] , \_20_net_[28] ,
         \_20_net_[27] , \_20_net_[26] , \_20_net_[25] , \_20_net_[24] ,
         \_20_net_[23] , \_20_net_[22] , \_20_net_[21] , \_20_net_[20] ,
         \_20_net_[19] , \_20_net_[18] , \_20_net_[17] , \_20_net_[16] ,
         \_20_net_[15] , \_20_net_[14] , \_20_net_[13] , \_20_net_[12] ,
         \_20_net_[11] , \_22_net_[31] , \_22_net_[30] , \_22_net_[29] ,
         \_22_net_[28] , \_22_net_[27] , \_22_net_[26] , \_22_net_[25] ,
         \_22_net_[24] , \_22_net_[23] , \_22_net_[22] , \_22_net_[21] ,
         \_22_net_[20] , \_22_net_[19] , \_22_net_[18] , \_22_net_[17] ,
         \_22_net_[16] , \_22_net_[15] , \_22_net_[14] , \_22_net_[13] ,
         \_22_net_[12] , \_24_net_[31] , \_24_net_[30] , \_24_net_[29] ,
         \_24_net_[28] , \_24_net_[27] , \_24_net_[26] , \_24_net_[25] ,
         \_24_net_[24] , \_24_net_[23] , \_24_net_[22] , \_24_net_[21] ,
         \_24_net_[20] , \_24_net_[19] , \_24_net_[18] , \_24_net_[17] ,
         \_24_net_[16] , \_24_net_[15] , \_24_net_[14] , \_24_net_[13] ,
         \_26_net_[31] , \_26_net_[30] , \_26_net_[29] , \_26_net_[28] ,
         \_26_net_[27] , \_26_net_[26] , \_26_net_[25] , \_26_net_[24] ,
         \_26_net_[23] , \_26_net_[22] , \_26_net_[21] , \_26_net_[20] ,
         \_26_net_[19] , \_26_net_[18] , \_26_net_[17] , \_26_net_[16] ,
         \_26_net_[15] , \_26_net_[14] , \_28_net_[31] , \_28_net_[30] ,
         \_28_net_[29] , \_28_net_[28] , \_28_net_[27] , \_28_net_[26] ,
         \_28_net_[25] , \_28_net_[24] , \_28_net_[23] , \_28_net_[22] ,
         \_28_net_[21] , \_28_net_[20] , \_28_net_[19] , \_28_net_[18] ,
         \_28_net_[17] , \_28_net_[16] , \_28_net_[15] , \_30_net_[31] ,
         \_30_net_[30] , \_30_net_[29] , \_30_net_[28] , \_30_net_[27] ,
         \_30_net_[26] , \_30_net_[25] , \_30_net_[24] , \_30_net_[23] ,
         \_30_net_[22] , \_30_net_[21] , \_30_net_[20] , \_30_net_[19] ,
         \_30_net_[18] , \_30_net_[17] , \_30_net_[16] , \_32_net_[31] ,
         \_32_net_[30] , \_32_net_[29] , \_32_net_[28] , \_32_net_[27] ,
         \_32_net_[26] , \_32_net_[25] , \_32_net_[24] , \_32_net_[23] ,
         \_32_net_[22] , \_32_net_[21] , \_32_net_[20] , \_32_net_[19] ,
         \_32_net_[18] , \_32_net_[17] , \_34_net_[31] , \_34_net_[30] ,
         \_34_net_[29] , \_34_net_[28] , \_34_net_[27] , \_34_net_[26] ,
         \_34_net_[25] , \_34_net_[24] , \_34_net_[23] , \_34_net_[22] ,
         \_34_net_[21] , \_34_net_[20] , \_34_net_[19] , \_34_net_[18] ,
         \_36_net_[31] , \_36_net_[30] , \_36_net_[29] , \_36_net_[28] ,
         \_36_net_[27] , \_36_net_[26] , \_36_net_[25] , \_36_net_[24] ,
         \_36_net_[23] , \_36_net_[22] , \_36_net_[21] , \_36_net_[20] ,
         \_36_net_[19] , \_38_net_[31] , \_38_net_[30] , \_38_net_[29] ,
         \_38_net_[28] , \_38_net_[27] , \_38_net_[26] , \_38_net_[25] ,
         \_38_net_[24] , \_38_net_[23] , \_38_net_[22] , \_38_net_[21] ,
         \_38_net_[20] , \_40_net_[31] , \_40_net_[30] , \_40_net_[29] ,
         \_40_net_[28] , \_40_net_[27] , \_40_net_[26] , \_40_net_[25] ,
         \_40_net_[24] , \_40_net_[23] , \_40_net_[22] , \_40_net_[21] ,
         \_42_net_[31] , \_42_net_[30] , \_42_net_[29] , \_42_net_[28] ,
         \_42_net_[27] , \_42_net_[26] , \_42_net_[25] , \_42_net_[24] ,
         \_42_net_[23] , \_42_net_[22] , \_44_net_[31] , \_44_net_[30] ,
         \_44_net_[29] , \_44_net_[28] , \_44_net_[27] , \_44_net_[26] ,
         \_44_net_[25] , \_44_net_[24] , \_44_net_[23] , \_46_net_[31] ,
         \_46_net_[30] , \_46_net_[29] , \_46_net_[28] , \_46_net_[27] ,
         \_46_net_[26] , \_46_net_[25] , \_46_net_[24] , \_48_net_[31] ,
         \_48_net_[30] , \_48_net_[29] , \_48_net_[28] , \_48_net_[27] ,
         \_48_net_[26] , \_48_net_[25] , \_50_net_[31] , \_50_net_[30] ,
         \_50_net_[29] , \_50_net_[28] , \_50_net_[27] , \_50_net_[26] ,
         \_52_net_[31] , \_52_net_[30] , \_52_net_[29] , \_52_net_[28] ,
         \_52_net_[27] , \_54_net_[31] , \_54_net_[30] , \_54_net_[29] ,
         \_54_net_[28] , \_56_net_[31] , \_56_net_[30] , \_56_net_[29] ,
         \_58_net_[31] , \_58_net_[30] , \_60_net_[31] ;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30;

  ADD_N32_189 \FAINST[1].ADD_  ( .A({\_0_net_[31] , \_0_net_[30] , 
        \_0_net_[29] , \_0_net_[28] , \_0_net_[27] , \_0_net_[26] , 
        \_0_net_[25] , \_0_net_[24] , \_0_net_[23] , \_0_net_[22] , 
        \_0_net_[21] , \_0_net_[20] , \_0_net_[19] , \_0_net_[18] , 
        \_0_net_[17] , \_0_net_[16] , \_0_net_[15] , \_0_net_[14] , 
        \_0_net_[13] , \_0_net_[12] , \_0_net_[11] , \_0_net_[10] , 
        \_0_net_[9] , \_0_net_[8] , \_0_net_[7] , \_0_net_[6] , \_0_net_[5] , 
        \_0_net_[4] , \_0_net_[3] , \_0_net_[2] , \_0_net_[1] , 1'b0}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .S({
        \w[2][31] , \w[2][30] , \w[2][29] , \w[2][28] , \w[2][27] , \w[2][26] , 
        \w[2][25] , \w[2][24] , \w[2][23] , \w[2][22] , \w[2][21] , \w[2][20] , 
        \w[2][19] , \w[2][18] , \w[2][17] , \w[2][16] , \w[2][15] , \w[2][14] , 
        \w[2][13] , \w[2][12] , \w[2][11] , \w[2][10] , \w[2][9] , \w[2][8] , 
        \w[2][7] , \w[2][6] , \w[2][5] , \w[2][4] , \w[2][3] , \w[2][2] , 
        \w[2][1] , SYNOPSYS_UNCONNECTED__0}) );
  ADD_N32_188 \FAINST[2].ADD_  ( .A({\_2_net_[31] , \_2_net_[30] , 
        \_2_net_[29] , \_2_net_[28] , \_2_net_[27] , \_2_net_[26] , 
        \_2_net_[25] , \_2_net_[24] , \_2_net_[23] , \_2_net_[22] , 
        \_2_net_[21] , \_2_net_[20] , \_2_net_[19] , \_2_net_[18] , 
        \_2_net_[17] , \_2_net_[16] , \_2_net_[15] , \_2_net_[14] , 
        \_2_net_[13] , \_2_net_[12] , \_2_net_[11] , \_2_net_[10] , 
        \_2_net_[9] , \_2_net_[8] , \_2_net_[7] , \_2_net_[6] , \_2_net_[5] , 
        \_2_net_[4] , \_2_net_[3] , \_2_net_[2] , 1'b0, 1'b0}), .B({\w[2][31] , 
        \w[2][30] , \w[2][29] , \w[2][28] , \w[2][27] , \w[2][26] , \w[2][25] , 
        \w[2][24] , \w[2][23] , \w[2][22] , \w[2][21] , \w[2][20] , \w[2][19] , 
        \w[2][18] , \w[2][17] , \w[2][16] , \w[2][15] , \w[2][14] , \w[2][13] , 
        \w[2][12] , \w[2][11] , \w[2][10] , \w[2][9] , \w[2][8] , \w[2][7] , 
        \w[2][6] , \w[2][5] , \w[2][4] , \w[2][3] , \w[2][2] , \w[2][1] , 1'b0}), .CI(1'b0), .S({\w[3][31] , \w[3][30] , \w[3][29] , \w[3][28] , \w[3][27] , 
        \w[3][26] , \w[3][25] , \w[3][24] , \w[3][23] , \w[3][22] , \w[3][21] , 
        \w[3][20] , \w[3][19] , \w[3][18] , \w[3][17] , \w[3][16] , \w[3][15] , 
        \w[3][14] , \w[3][13] , \w[3][12] , \w[3][11] , \w[3][10] , \w[3][9] , 
        \w[3][8] , \w[3][7] , \w[3][6] , \w[3][5] , \w[3][4] , \w[3][3] , 
        \w[3][2] , \w[3][1] , SYNOPSYS_UNCONNECTED__1}) );
  ADD_N32_187 \FAINST[3].ADD_  ( .A({\_4_net_[31] , \_4_net_[30] , 
        \_4_net_[29] , \_4_net_[28] , \_4_net_[27] , \_4_net_[26] , 
        \_4_net_[25] , \_4_net_[24] , \_4_net_[23] , \_4_net_[22] , 
        \_4_net_[21] , \_4_net_[20] , \_4_net_[19] , \_4_net_[18] , 
        \_4_net_[17] , \_4_net_[16] , \_4_net_[15] , \_4_net_[14] , 
        \_4_net_[13] , \_4_net_[12] , \_4_net_[11] , \_4_net_[10] , 
        \_4_net_[9] , \_4_net_[8] , \_4_net_[7] , \_4_net_[6] , \_4_net_[5] , 
        \_4_net_[4] , \_4_net_[3] , 1'b0, 1'b0, 1'b0}), .B({\w[3][31] , 
        \w[3][30] , \w[3][29] , \w[3][28] , \w[3][27] , \w[3][26] , \w[3][25] , 
        \w[3][24] , \w[3][23] , \w[3][22] , \w[3][21] , \w[3][20] , \w[3][19] , 
        \w[3][18] , \w[3][17] , \w[3][16] , \w[3][15] , \w[3][14] , \w[3][13] , 
        \w[3][12] , \w[3][11] , \w[3][10] , \w[3][9] , \w[3][8] , \w[3][7] , 
        \w[3][6] , \w[3][5] , \w[3][4] , \w[3][3] , \w[3][2] , \w[3][1] , 1'b0}), .CI(1'b0), .S({\w[4][31] , \w[4][30] , \w[4][29] , \w[4][28] , \w[4][27] , 
        \w[4][26] , \w[4][25] , \w[4][24] , \w[4][23] , \w[4][22] , \w[4][21] , 
        \w[4][20] , \w[4][19] , \w[4][18] , \w[4][17] , \w[4][16] , \w[4][15] , 
        \w[4][14] , \w[4][13] , \w[4][12] , \w[4][11] , \w[4][10] , \w[4][9] , 
        \w[4][8] , \w[4][7] , \w[4][6] , \w[4][5] , \w[4][4] , \w[4][3] , 
        \w[4][2] , \w[4][1] , SYNOPSYS_UNCONNECTED__2}) );
  ADD_N32_186 \FAINST[4].ADD_  ( .A({\_6_net_[31] , \_6_net_[30] , 
        \_6_net_[29] , \_6_net_[28] , \_6_net_[27] , \_6_net_[26] , 
        \_6_net_[25] , \_6_net_[24] , \_6_net_[23] , \_6_net_[22] , 
        \_6_net_[21] , \_6_net_[20] , \_6_net_[19] , \_6_net_[18] , 
        \_6_net_[17] , \_6_net_[16] , \_6_net_[15] , \_6_net_[14] , 
        \_6_net_[13] , \_6_net_[12] , \_6_net_[11] , \_6_net_[10] , 
        \_6_net_[9] , \_6_net_[8] , \_6_net_[7] , \_6_net_[6] , \_6_net_[5] , 
        \_6_net_[4] , 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[4][31] , \w[4][30] , 
        \w[4][29] , \w[4][28] , \w[4][27] , \w[4][26] , \w[4][25] , \w[4][24] , 
        \w[4][23] , \w[4][22] , \w[4][21] , \w[4][20] , \w[4][19] , \w[4][18] , 
        \w[4][17] , \w[4][16] , \w[4][15] , \w[4][14] , \w[4][13] , \w[4][12] , 
        \w[4][11] , \w[4][10] , \w[4][9] , \w[4][8] , \w[4][7] , \w[4][6] , 
        \w[4][5] , \w[4][4] , \w[4][3] , \w[4][2] , \w[4][1] , 1'b0}), .CI(
        1'b0), .S({\w[5][31] , \w[5][30] , \w[5][29] , \w[5][28] , \w[5][27] , 
        \w[5][26] , \w[5][25] , \w[5][24] , \w[5][23] , \w[5][22] , \w[5][21] , 
        \w[5][20] , \w[5][19] , \w[5][18] , \w[5][17] , \w[5][16] , \w[5][15] , 
        \w[5][14] , \w[5][13] , \w[5][12] , \w[5][11] , \w[5][10] , \w[5][9] , 
        \w[5][8] , \w[5][7] , \w[5][6] , \w[5][5] , \w[5][4] , \w[5][3] , 
        \w[5][2] , \w[5][1] , SYNOPSYS_UNCONNECTED__3}) );
  ADD_N32_185 \FAINST[5].ADD_  ( .A({\_8_net_[31] , \_8_net_[30] , 
        \_8_net_[29] , \_8_net_[28] , \_8_net_[27] , \_8_net_[26] , 
        \_8_net_[25] , \_8_net_[24] , \_8_net_[23] , \_8_net_[22] , 
        \_8_net_[21] , \_8_net_[20] , \_8_net_[19] , \_8_net_[18] , 
        \_8_net_[17] , \_8_net_[16] , \_8_net_[15] , \_8_net_[14] , 
        \_8_net_[13] , \_8_net_[12] , \_8_net_[11] , \_8_net_[10] , 
        \_8_net_[9] , \_8_net_[8] , \_8_net_[7] , \_8_net_[6] , \_8_net_[5] , 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[5][31] , \w[5][30] , \w[5][29] , 
        \w[5][28] , \w[5][27] , \w[5][26] , \w[5][25] , \w[5][24] , \w[5][23] , 
        \w[5][22] , \w[5][21] , \w[5][20] , \w[5][19] , \w[5][18] , \w[5][17] , 
        \w[5][16] , \w[5][15] , \w[5][14] , \w[5][13] , \w[5][12] , \w[5][11] , 
        \w[5][10] , \w[5][9] , \w[5][8] , \w[5][7] , \w[5][6] , \w[5][5] , 
        \w[5][4] , \w[5][3] , \w[5][2] , \w[5][1] , 1'b0}), .CI(1'b0), .S({
        \w[6][31] , \w[6][30] , \w[6][29] , \w[6][28] , \w[6][27] , \w[6][26] , 
        \w[6][25] , \w[6][24] , \w[6][23] , \w[6][22] , \w[6][21] , \w[6][20] , 
        \w[6][19] , \w[6][18] , \w[6][17] , \w[6][16] , \w[6][15] , \w[6][14] , 
        \w[6][13] , \w[6][12] , \w[6][11] , \w[6][10] , \w[6][9] , \w[6][8] , 
        \w[6][7] , \w[6][6] , \w[6][5] , \w[6][4] , \w[6][3] , \w[6][2] , 
        \w[6][1] , SYNOPSYS_UNCONNECTED__4}) );
  ADD_N32_184 \FAINST[6].ADD_  ( .A({\_10_net_[31] , \_10_net_[30] , 
        \_10_net_[29] , \_10_net_[28] , \_10_net_[27] , \_10_net_[26] , 
        \_10_net_[25] , \_10_net_[24] , \_10_net_[23] , \_10_net_[22] , 
        \_10_net_[21] , \_10_net_[20] , \_10_net_[19] , \_10_net_[18] , 
        \_10_net_[17] , \_10_net_[16] , \_10_net_[15] , \_10_net_[14] , 
        \_10_net_[13] , \_10_net_[12] , \_10_net_[11] , \_10_net_[10] , 
        \_10_net_[9] , \_10_net_[8] , \_10_net_[7] , \_10_net_[6] , 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[6][31] , \w[6][30] , \w[6][29] , 
        \w[6][28] , \w[6][27] , \w[6][26] , \w[6][25] , \w[6][24] , \w[6][23] , 
        \w[6][22] , \w[6][21] , \w[6][20] , \w[6][19] , \w[6][18] , \w[6][17] , 
        \w[6][16] , \w[6][15] , \w[6][14] , \w[6][13] , \w[6][12] , \w[6][11] , 
        \w[6][10] , \w[6][9] , \w[6][8] , \w[6][7] , \w[6][6] , \w[6][5] , 
        \w[6][4] , \w[6][3] , \w[6][2] , \w[6][1] , 1'b0}), .CI(1'b0), .S({
        \w[7][31] , \w[7][30] , \w[7][29] , \w[7][28] , \w[7][27] , \w[7][26] , 
        \w[7][25] , \w[7][24] , \w[7][23] , \w[7][22] , \w[7][21] , \w[7][20] , 
        \w[7][19] , \w[7][18] , \w[7][17] , \w[7][16] , \w[7][15] , \w[7][14] , 
        \w[7][13] , \w[7][12] , \w[7][11] , \w[7][10] , \w[7][9] , \w[7][8] , 
        \w[7][7] , \w[7][6] , \w[7][5] , \w[7][4] , \w[7][3] , \w[7][2] , 
        \w[7][1] , SYNOPSYS_UNCONNECTED__5}) );
  ADD_N32_183 \FAINST[7].ADD_  ( .A({\_12_net_[31] , \_12_net_[30] , 
        \_12_net_[29] , \_12_net_[28] , \_12_net_[27] , \_12_net_[26] , 
        \_12_net_[25] , \_12_net_[24] , \_12_net_[23] , \_12_net_[22] , 
        \_12_net_[21] , \_12_net_[20] , \_12_net_[19] , \_12_net_[18] , 
        \_12_net_[17] , \_12_net_[16] , \_12_net_[15] , \_12_net_[14] , 
        \_12_net_[13] , \_12_net_[12] , \_12_net_[11] , \_12_net_[10] , 
        \_12_net_[9] , \_12_net_[8] , \_12_net_[7] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({\w[7][31] , \w[7][30] , \w[7][29] , \w[7][28] , 
        \w[7][27] , \w[7][26] , \w[7][25] , \w[7][24] , \w[7][23] , \w[7][22] , 
        \w[7][21] , \w[7][20] , \w[7][19] , \w[7][18] , \w[7][17] , \w[7][16] , 
        \w[7][15] , \w[7][14] , \w[7][13] , \w[7][12] , \w[7][11] , \w[7][10] , 
        \w[7][9] , \w[7][8] , \w[7][7] , \w[7][6] , \w[7][5] , \w[7][4] , 
        \w[7][3] , \w[7][2] , \w[7][1] , 1'b0}), .CI(1'b0), .S({\w[8][31] , 
        \w[8][30] , \w[8][29] , \w[8][28] , \w[8][27] , \w[8][26] , \w[8][25] , 
        \w[8][24] , \w[8][23] , \w[8][22] , \w[8][21] , \w[8][20] , \w[8][19] , 
        \w[8][18] , \w[8][17] , \w[8][16] , \w[8][15] , \w[8][14] , \w[8][13] , 
        \w[8][12] , \w[8][11] , \w[8][10] , \w[8][9] , \w[8][8] , \w[8][7] , 
        \w[8][6] , \w[8][5] , \w[8][4] , \w[8][3] , \w[8][2] , \w[8][1] , 
        SYNOPSYS_UNCONNECTED__6}) );
  ADD_N32_182 \FAINST[8].ADD_  ( .A({\_14_net_[31] , \_14_net_[30] , 
        \_14_net_[29] , \_14_net_[28] , \_14_net_[27] , \_14_net_[26] , 
        \_14_net_[25] , \_14_net_[24] , \_14_net_[23] , \_14_net_[22] , 
        \_14_net_[21] , \_14_net_[20] , \_14_net_[19] , \_14_net_[18] , 
        \_14_net_[17] , \_14_net_[16] , \_14_net_[15] , \_14_net_[14] , 
        \_14_net_[13] , \_14_net_[12] , \_14_net_[11] , \_14_net_[10] , 
        \_14_net_[9] , \_14_net_[8] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({\w[8][31] , \w[8][30] , \w[8][29] , \w[8][28] , \w[8][27] , 
        \w[8][26] , \w[8][25] , \w[8][24] , \w[8][23] , \w[8][22] , \w[8][21] , 
        \w[8][20] , \w[8][19] , \w[8][18] , \w[8][17] , \w[8][16] , \w[8][15] , 
        \w[8][14] , \w[8][13] , \w[8][12] , \w[8][11] , \w[8][10] , \w[8][9] , 
        \w[8][8] , \w[8][7] , \w[8][6] , \w[8][5] , \w[8][4] , \w[8][3] , 
        \w[8][2] , \w[8][1] , 1'b0}), .CI(1'b0), .S({\w[9][31] , \w[9][30] , 
        \w[9][29] , \w[9][28] , \w[9][27] , \w[9][26] , \w[9][25] , \w[9][24] , 
        \w[9][23] , \w[9][22] , \w[9][21] , \w[9][20] , \w[9][19] , \w[9][18] , 
        \w[9][17] , \w[9][16] , \w[9][15] , \w[9][14] , \w[9][13] , \w[9][12] , 
        \w[9][11] , \w[9][10] , \w[9][9] , \w[9][8] , \w[9][7] , \w[9][6] , 
        \w[9][5] , \w[9][4] , \w[9][3] , \w[9][2] , \w[9][1] , 
        SYNOPSYS_UNCONNECTED__7}) );
  ADD_N32_181 \FAINST[9].ADD_  ( .A({\_16_net_[31] , \_16_net_[30] , 
        \_16_net_[29] , \_16_net_[28] , \_16_net_[27] , \_16_net_[26] , 
        \_16_net_[25] , \_16_net_[24] , \_16_net_[23] , \_16_net_[22] , 
        \_16_net_[21] , \_16_net_[20] , \_16_net_[19] , \_16_net_[18] , 
        \_16_net_[17] , \_16_net_[16] , \_16_net_[15] , \_16_net_[14] , 
        \_16_net_[13] , \_16_net_[12] , \_16_net_[11] , \_16_net_[10] , 
        \_16_net_[9] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({\w[9][31] , \w[9][30] , \w[9][29] , \w[9][28] , \w[9][27] , 
        \w[9][26] , \w[9][25] , \w[9][24] , \w[9][23] , \w[9][22] , \w[9][21] , 
        \w[9][20] , \w[9][19] , \w[9][18] , \w[9][17] , \w[9][16] , \w[9][15] , 
        \w[9][14] , \w[9][13] , \w[9][12] , \w[9][11] , \w[9][10] , \w[9][9] , 
        \w[9][8] , \w[9][7] , \w[9][6] , \w[9][5] , \w[9][4] , \w[9][3] , 
        \w[9][2] , \w[9][1] , 1'b0}), .CI(1'b0), .S({\w[10][31] , \w[10][30] , 
        \w[10][29] , \w[10][28] , \w[10][27] , \w[10][26] , \w[10][25] , 
        \w[10][24] , \w[10][23] , \w[10][22] , \w[10][21] , \w[10][20] , 
        \w[10][19] , \w[10][18] , \w[10][17] , \w[10][16] , \w[10][15] , 
        \w[10][14] , \w[10][13] , \w[10][12] , \w[10][11] , \w[10][10] , 
        \w[10][9] , \w[10][8] , \w[10][7] , \w[10][6] , \w[10][5] , \w[10][4] , 
        \w[10][3] , \w[10][2] , \w[10][1] , SYNOPSYS_UNCONNECTED__8}) );
  ADD_N32_180 \FAINST[10].ADD_  ( .A({\_18_net_[31] , \_18_net_[30] , 
        \_18_net_[29] , \_18_net_[28] , \_18_net_[27] , \_18_net_[26] , 
        \_18_net_[25] , \_18_net_[24] , \_18_net_[23] , \_18_net_[22] , 
        \_18_net_[21] , \_18_net_[20] , \_18_net_[19] , \_18_net_[18] , 
        \_18_net_[17] , \_18_net_[16] , \_18_net_[15] , \_18_net_[14] , 
        \_18_net_[13] , \_18_net_[12] , \_18_net_[11] , \_18_net_[10] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[10][31] , \w[10][30] , \w[10][29] , \w[10][28] , \w[10][27] , 
        \w[10][26] , \w[10][25] , \w[10][24] , \w[10][23] , \w[10][22] , 
        \w[10][21] , \w[10][20] , \w[10][19] , \w[10][18] , \w[10][17] , 
        \w[10][16] , \w[10][15] , \w[10][14] , \w[10][13] , \w[10][12] , 
        \w[10][11] , \w[10][10] , \w[10][9] , \w[10][8] , \w[10][7] , 
        \w[10][6] , \w[10][5] , \w[10][4] , \w[10][3] , \w[10][2] , \w[10][1] , 
        1'b0}), .CI(1'b0), .S({\w[11][31] , \w[11][30] , \w[11][29] , 
        \w[11][28] , \w[11][27] , \w[11][26] , \w[11][25] , \w[11][24] , 
        \w[11][23] , \w[11][22] , \w[11][21] , \w[11][20] , \w[11][19] , 
        \w[11][18] , \w[11][17] , \w[11][16] , \w[11][15] , \w[11][14] , 
        \w[11][13] , \w[11][12] , \w[11][11] , \w[11][10] , \w[11][9] , 
        \w[11][8] , \w[11][7] , \w[11][6] , \w[11][5] , \w[11][4] , \w[11][3] , 
        \w[11][2] , \w[11][1] , SYNOPSYS_UNCONNECTED__9}) );
  ADD_N32_179 \FAINST[11].ADD_  ( .A({\_20_net_[31] , \_20_net_[30] , 
        \_20_net_[29] , \_20_net_[28] , \_20_net_[27] , \_20_net_[26] , 
        \_20_net_[25] , \_20_net_[24] , \_20_net_[23] , \_20_net_[22] , 
        \_20_net_[21] , \_20_net_[20] , \_20_net_[19] , \_20_net_[18] , 
        \_20_net_[17] , \_20_net_[16] , \_20_net_[15] , \_20_net_[14] , 
        \_20_net_[13] , \_20_net_[12] , \_20_net_[11] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[11][31] , 
        \w[11][30] , \w[11][29] , \w[11][28] , \w[11][27] , \w[11][26] , 
        \w[11][25] , \w[11][24] , \w[11][23] , \w[11][22] , \w[11][21] , 
        \w[11][20] , \w[11][19] , \w[11][18] , \w[11][17] , \w[11][16] , 
        \w[11][15] , \w[11][14] , \w[11][13] , \w[11][12] , \w[11][11] , 
        \w[11][10] , \w[11][9] , \w[11][8] , \w[11][7] , \w[11][6] , 
        \w[11][5] , \w[11][4] , \w[11][3] , \w[11][2] , \w[11][1] , 1'b0}), 
        .CI(1'b0), .S({\w[12][31] , \w[12][30] , \w[12][29] , \w[12][28] , 
        \w[12][27] , \w[12][26] , \w[12][25] , \w[12][24] , \w[12][23] , 
        \w[12][22] , \w[12][21] , \w[12][20] , \w[12][19] , \w[12][18] , 
        \w[12][17] , \w[12][16] , \w[12][15] , \w[12][14] , \w[12][13] , 
        \w[12][12] , \w[12][11] , \w[12][10] , \w[12][9] , \w[12][8] , 
        \w[12][7] , \w[12][6] , \w[12][5] , \w[12][4] , \w[12][3] , \w[12][2] , 
        \w[12][1] , SYNOPSYS_UNCONNECTED__10}) );
  ADD_N32_178 \FAINST[12].ADD_  ( .A({\_22_net_[31] , \_22_net_[30] , 
        \_22_net_[29] , \_22_net_[28] , \_22_net_[27] , \_22_net_[26] , 
        \_22_net_[25] , \_22_net_[24] , \_22_net_[23] , \_22_net_[22] , 
        \_22_net_[21] , \_22_net_[20] , \_22_net_[19] , \_22_net_[18] , 
        \_22_net_[17] , \_22_net_[16] , \_22_net_[15] , \_22_net_[14] , 
        \_22_net_[13] , \_22_net_[12] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[12][31] , \w[12][30] , 
        \w[12][29] , \w[12][28] , \w[12][27] , \w[12][26] , \w[12][25] , 
        \w[12][24] , \w[12][23] , \w[12][22] , \w[12][21] , \w[12][20] , 
        \w[12][19] , \w[12][18] , \w[12][17] , \w[12][16] , \w[12][15] , 
        \w[12][14] , \w[12][13] , \w[12][12] , \w[12][11] , \w[12][10] , 
        \w[12][9] , \w[12][8] , \w[12][7] , \w[12][6] , \w[12][5] , \w[12][4] , 
        \w[12][3] , \w[12][2] , \w[12][1] , 1'b0}), .CI(1'b0), .S({\w[13][31] , 
        \w[13][30] , \w[13][29] , \w[13][28] , \w[13][27] , \w[13][26] , 
        \w[13][25] , \w[13][24] , \w[13][23] , \w[13][22] , \w[13][21] , 
        \w[13][20] , \w[13][19] , \w[13][18] , \w[13][17] , \w[13][16] , 
        \w[13][15] , \w[13][14] , \w[13][13] , \w[13][12] , \w[13][11] , 
        \w[13][10] , \w[13][9] , \w[13][8] , \w[13][7] , \w[13][6] , 
        \w[13][5] , \w[13][4] , \w[13][3] , \w[13][2] , \w[13][1] , 
        SYNOPSYS_UNCONNECTED__11}) );
  ADD_N32_177 \FAINST[13].ADD_  ( .A({\_24_net_[31] , \_24_net_[30] , 
        \_24_net_[29] , \_24_net_[28] , \_24_net_[27] , \_24_net_[26] , 
        \_24_net_[25] , \_24_net_[24] , \_24_net_[23] , \_24_net_[22] , 
        \_24_net_[21] , \_24_net_[20] , \_24_net_[19] , \_24_net_[18] , 
        \_24_net_[17] , \_24_net_[16] , \_24_net_[15] , \_24_net_[14] , 
        \_24_net_[13] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[13][31] , \w[13][30] , \w[13][29] , 
        \w[13][28] , \w[13][27] , \w[13][26] , \w[13][25] , \w[13][24] , 
        \w[13][23] , \w[13][22] , \w[13][21] , \w[13][20] , \w[13][19] , 
        \w[13][18] , \w[13][17] , \w[13][16] , \w[13][15] , \w[13][14] , 
        \w[13][13] , \w[13][12] , \w[13][11] , \w[13][10] , \w[13][9] , 
        \w[13][8] , \w[13][7] , \w[13][6] , \w[13][5] , \w[13][4] , \w[13][3] , 
        \w[13][2] , \w[13][1] , 1'b0}), .CI(1'b0), .S({\w[14][31] , 
        \w[14][30] , \w[14][29] , \w[14][28] , \w[14][27] , \w[14][26] , 
        \w[14][25] , \w[14][24] , \w[14][23] , \w[14][22] , \w[14][21] , 
        \w[14][20] , \w[14][19] , \w[14][18] , \w[14][17] , \w[14][16] , 
        \w[14][15] , \w[14][14] , \w[14][13] , \w[14][12] , \w[14][11] , 
        \w[14][10] , \w[14][9] , \w[14][8] , \w[14][7] , \w[14][6] , 
        \w[14][5] , \w[14][4] , \w[14][3] , \w[14][2] , \w[14][1] , 
        SYNOPSYS_UNCONNECTED__12}) );
  ADD_N32_176 \FAINST[14].ADD_  ( .A({\_26_net_[31] , \_26_net_[30] , 
        \_26_net_[29] , \_26_net_[28] , \_26_net_[27] , \_26_net_[26] , 
        \_26_net_[25] , \_26_net_[24] , \_26_net_[23] , \_26_net_[22] , 
        \_26_net_[21] , \_26_net_[20] , \_26_net_[19] , \_26_net_[18] , 
        \_26_net_[17] , \_26_net_[16] , \_26_net_[15] , \_26_net_[14] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({\w[14][31] , \w[14][30] , \w[14][29] , \w[14][28] , 
        \w[14][27] , \w[14][26] , \w[14][25] , \w[14][24] , \w[14][23] , 
        \w[14][22] , \w[14][21] , \w[14][20] , \w[14][19] , \w[14][18] , 
        \w[14][17] , \w[14][16] , \w[14][15] , \w[14][14] , \w[14][13] , 
        \w[14][12] , \w[14][11] , \w[14][10] , \w[14][9] , \w[14][8] , 
        \w[14][7] , \w[14][6] , \w[14][5] , \w[14][4] , \w[14][3] , \w[14][2] , 
        \w[14][1] , 1'b0}), .CI(1'b0), .S({\w[15][31] , \w[15][30] , 
        \w[15][29] , \w[15][28] , \w[15][27] , \w[15][26] , \w[15][25] , 
        \w[15][24] , \w[15][23] , \w[15][22] , \w[15][21] , \w[15][20] , 
        \w[15][19] , \w[15][18] , \w[15][17] , \w[15][16] , \w[15][15] , 
        \w[15][14] , \w[15][13] , \w[15][12] , \w[15][11] , \w[15][10] , 
        \w[15][9] , \w[15][8] , \w[15][7] , \w[15][6] , \w[15][5] , \w[15][4] , 
        \w[15][3] , \w[15][2] , \w[15][1] , SYNOPSYS_UNCONNECTED__13}) );
  ADD_N32_175 \FAINST[15].ADD_  ( .A({\_28_net_[31] , \_28_net_[30] , 
        \_28_net_[29] , \_28_net_[28] , \_28_net_[27] , \_28_net_[26] , 
        \_28_net_[25] , \_28_net_[24] , \_28_net_[23] , \_28_net_[22] , 
        \_28_net_[21] , \_28_net_[20] , \_28_net_[19] , \_28_net_[18] , 
        \_28_net_[17] , \_28_net_[16] , \_28_net_[15] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({\w[15][31] , \w[15][30] , \w[15][29] , \w[15][28] , \w[15][27] , 
        \w[15][26] , \w[15][25] , \w[15][24] , \w[15][23] , \w[15][22] , 
        \w[15][21] , \w[15][20] , \w[15][19] , \w[15][18] , \w[15][17] , 
        \w[15][16] , \w[15][15] , \w[15][14] , \w[15][13] , \w[15][12] , 
        \w[15][11] , \w[15][10] , \w[15][9] , \w[15][8] , \w[15][7] , 
        \w[15][6] , \w[15][5] , \w[15][4] , \w[15][3] , \w[15][2] , \w[15][1] , 
        1'b0}), .CI(1'b0), .S({\w[16][31] , \w[16][30] , \w[16][29] , 
        \w[16][28] , \w[16][27] , \w[16][26] , \w[16][25] , \w[16][24] , 
        \w[16][23] , \w[16][22] , \w[16][21] , \w[16][20] , \w[16][19] , 
        \w[16][18] , \w[16][17] , \w[16][16] , \w[16][15] , \w[16][14] , 
        \w[16][13] , \w[16][12] , \w[16][11] , \w[16][10] , \w[16][9] , 
        \w[16][8] , \w[16][7] , \w[16][6] , \w[16][5] , \w[16][4] , \w[16][3] , 
        \w[16][2] , \w[16][1] , SYNOPSYS_UNCONNECTED__14}) );
  ADD_N32_174 \FAINST[16].ADD_  ( .A({\_30_net_[31] , \_30_net_[30] , 
        \_30_net_[29] , \_30_net_[28] , \_30_net_[27] , \_30_net_[26] , 
        \_30_net_[25] , \_30_net_[24] , \_30_net_[23] , \_30_net_[22] , 
        \_30_net_[21] , \_30_net_[20] , \_30_net_[19] , \_30_net_[18] , 
        \_30_net_[17] , \_30_net_[16] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[16][31] , \w[16][30] , \w[16][29] , \w[16][28] , \w[16][27] , 
        \w[16][26] , \w[16][25] , \w[16][24] , \w[16][23] , \w[16][22] , 
        \w[16][21] , \w[16][20] , \w[16][19] , \w[16][18] , \w[16][17] , 
        \w[16][16] , \w[16][15] , \w[16][14] , \w[16][13] , \w[16][12] , 
        \w[16][11] , \w[16][10] , \w[16][9] , \w[16][8] , \w[16][7] , 
        \w[16][6] , \w[16][5] , \w[16][4] , \w[16][3] , \w[16][2] , \w[16][1] , 
        1'b0}), .CI(1'b0), .S({\w[17][31] , \w[17][30] , \w[17][29] , 
        \w[17][28] , \w[17][27] , \w[17][26] , \w[17][25] , \w[17][24] , 
        \w[17][23] , \w[17][22] , \w[17][21] , \w[17][20] , \w[17][19] , 
        \w[17][18] , \w[17][17] , \w[17][16] , \w[17][15] , \w[17][14] , 
        \w[17][13] , \w[17][12] , \w[17][11] , \w[17][10] , \w[17][9] , 
        \w[17][8] , \w[17][7] , \w[17][6] , \w[17][5] , \w[17][4] , \w[17][3] , 
        \w[17][2] , \w[17][1] , SYNOPSYS_UNCONNECTED__15}) );
  ADD_N32_173 \FAINST[17].ADD_  ( .A({\_32_net_[31] , \_32_net_[30] , 
        \_32_net_[29] , \_32_net_[28] , \_32_net_[27] , \_32_net_[26] , 
        \_32_net_[25] , \_32_net_[24] , \_32_net_[23] , \_32_net_[22] , 
        \_32_net_[21] , \_32_net_[20] , \_32_net_[19] , \_32_net_[18] , 
        \_32_net_[17] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[17][31] , 
        \w[17][30] , \w[17][29] , \w[17][28] , \w[17][27] , \w[17][26] , 
        \w[17][25] , \w[17][24] , \w[17][23] , \w[17][22] , \w[17][21] , 
        \w[17][20] , \w[17][19] , \w[17][18] , \w[17][17] , \w[17][16] , 
        \w[17][15] , \w[17][14] , \w[17][13] , \w[17][12] , \w[17][11] , 
        \w[17][10] , \w[17][9] , \w[17][8] , \w[17][7] , \w[17][6] , 
        \w[17][5] , \w[17][4] , \w[17][3] , \w[17][2] , \w[17][1] , 1'b0}), 
        .CI(1'b0), .S({\w[18][31] , \w[18][30] , \w[18][29] , \w[18][28] , 
        \w[18][27] , \w[18][26] , \w[18][25] , \w[18][24] , \w[18][23] , 
        \w[18][22] , \w[18][21] , \w[18][20] , \w[18][19] , \w[18][18] , 
        \w[18][17] , \w[18][16] , \w[18][15] , \w[18][14] , \w[18][13] , 
        \w[18][12] , \w[18][11] , \w[18][10] , \w[18][9] , \w[18][8] , 
        \w[18][7] , \w[18][6] , \w[18][5] , \w[18][4] , \w[18][3] , \w[18][2] , 
        \w[18][1] , SYNOPSYS_UNCONNECTED__16}) );
  ADD_N32_172 \FAINST[18].ADD_  ( .A({\_34_net_[31] , \_34_net_[30] , 
        \_34_net_[29] , \_34_net_[28] , \_34_net_[27] , \_34_net_[26] , 
        \_34_net_[25] , \_34_net_[24] , \_34_net_[23] , \_34_net_[22] , 
        \_34_net_[21] , \_34_net_[20] , \_34_net_[19] , \_34_net_[18] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[18][31] , \w[18][30] , 
        \w[18][29] , \w[18][28] , \w[18][27] , \w[18][26] , \w[18][25] , 
        \w[18][24] , \w[18][23] , \w[18][22] , \w[18][21] , \w[18][20] , 
        \w[18][19] , \w[18][18] , \w[18][17] , \w[18][16] , \w[18][15] , 
        \w[18][14] , \w[18][13] , \w[18][12] , \w[18][11] , \w[18][10] , 
        \w[18][9] , \w[18][8] , \w[18][7] , \w[18][6] , \w[18][5] , \w[18][4] , 
        \w[18][3] , \w[18][2] , \w[18][1] , 1'b0}), .CI(1'b0), .S({\w[19][31] , 
        \w[19][30] , \w[19][29] , \w[19][28] , \w[19][27] , \w[19][26] , 
        \w[19][25] , \w[19][24] , \w[19][23] , \w[19][22] , \w[19][21] , 
        \w[19][20] , \w[19][19] , \w[19][18] , \w[19][17] , \w[19][16] , 
        \w[19][15] , \w[19][14] , \w[19][13] , \w[19][12] , \w[19][11] , 
        \w[19][10] , \w[19][9] , \w[19][8] , \w[19][7] , \w[19][6] , 
        \w[19][5] , \w[19][4] , \w[19][3] , \w[19][2] , \w[19][1] , 
        SYNOPSYS_UNCONNECTED__17}) );
  ADD_N32_171 \FAINST[19].ADD_  ( .A({\_36_net_[31] , \_36_net_[30] , 
        \_36_net_[29] , \_36_net_[28] , \_36_net_[27] , \_36_net_[26] , 
        \_36_net_[25] , \_36_net_[24] , \_36_net_[23] , \_36_net_[22] , 
        \_36_net_[21] , \_36_net_[20] , \_36_net_[19] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({\w[19][31] , \w[19][30] , \w[19][29] , 
        \w[19][28] , \w[19][27] , \w[19][26] , \w[19][25] , \w[19][24] , 
        \w[19][23] , \w[19][22] , \w[19][21] , \w[19][20] , \w[19][19] , 
        \w[19][18] , \w[19][17] , \w[19][16] , \w[19][15] , \w[19][14] , 
        \w[19][13] , \w[19][12] , \w[19][11] , \w[19][10] , \w[19][9] , 
        \w[19][8] , \w[19][7] , \w[19][6] , \w[19][5] , \w[19][4] , \w[19][3] , 
        \w[19][2] , \w[19][1] , 1'b0}), .CI(1'b0), .S({\w[20][31] , 
        \w[20][30] , \w[20][29] , \w[20][28] , \w[20][27] , \w[20][26] , 
        \w[20][25] , \w[20][24] , \w[20][23] , \w[20][22] , \w[20][21] , 
        \w[20][20] , \w[20][19] , \w[20][18] , \w[20][17] , \w[20][16] , 
        \w[20][15] , \w[20][14] , \w[20][13] , \w[20][12] , \w[20][11] , 
        \w[20][10] , \w[20][9] , \w[20][8] , \w[20][7] , \w[20][6] , 
        \w[20][5] , \w[20][4] , \w[20][3] , \w[20][2] , \w[20][1] , 
        SYNOPSYS_UNCONNECTED__18}) );
  ADD_N32_170 \FAINST[20].ADD_  ( .A({\_38_net_[31] , \_38_net_[30] , 
        \_38_net_[29] , \_38_net_[28] , \_38_net_[27] , \_38_net_[26] , 
        \_38_net_[25] , \_38_net_[24] , \_38_net_[23] , \_38_net_[22] , 
        \_38_net_[21] , \_38_net_[20] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .B({\w[20][31] , \w[20][30] , \w[20][29] , \w[20][28] , 
        \w[20][27] , \w[20][26] , \w[20][25] , \w[20][24] , \w[20][23] , 
        \w[20][22] , \w[20][21] , \w[20][20] , \w[20][19] , \w[20][18] , 
        \w[20][17] , \w[20][16] , \w[20][15] , \w[20][14] , \w[20][13] , 
        \w[20][12] , \w[20][11] , \w[20][10] , \w[20][9] , \w[20][8] , 
        \w[20][7] , \w[20][6] , \w[20][5] , \w[20][4] , \w[20][3] , \w[20][2] , 
        \w[20][1] , 1'b0}), .CI(1'b0), .S({\w[21][31] , \w[21][30] , 
        \w[21][29] , \w[21][28] , \w[21][27] , \w[21][26] , \w[21][25] , 
        \w[21][24] , \w[21][23] , \w[21][22] , \w[21][21] , \w[21][20] , 
        \w[21][19] , \w[21][18] , \w[21][17] , \w[21][16] , \w[21][15] , 
        \w[21][14] , \w[21][13] , \w[21][12] , \w[21][11] , \w[21][10] , 
        \w[21][9] , \w[21][8] , \w[21][7] , \w[21][6] , \w[21][5] , \w[21][4] , 
        \w[21][3] , \w[21][2] , \w[21][1] , SYNOPSYS_UNCONNECTED__19}) );
  ADD_N32_169 \FAINST[21].ADD_  ( .A({\_40_net_[31] , \_40_net_[30] , 
        \_40_net_[29] , \_40_net_[28] , \_40_net_[27] , \_40_net_[26] , 
        \_40_net_[25] , \_40_net_[24] , \_40_net_[23] , \_40_net_[22] , 
        \_40_net_[21] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[21][31] , \w[21][30] , \w[21][29] , \w[21][28] , \w[21][27] , 
        \w[21][26] , \w[21][25] , \w[21][24] , \w[21][23] , \w[21][22] , 
        \w[21][21] , \w[21][20] , \w[21][19] , \w[21][18] , \w[21][17] , 
        \w[21][16] , \w[21][15] , \w[21][14] , \w[21][13] , \w[21][12] , 
        \w[21][11] , \w[21][10] , \w[21][9] , \w[21][8] , \w[21][7] , 
        \w[21][6] , \w[21][5] , \w[21][4] , \w[21][3] , \w[21][2] , \w[21][1] , 
        1'b0}), .CI(1'b0), .S({\w[22][31] , \w[22][30] , \w[22][29] , 
        \w[22][28] , \w[22][27] , \w[22][26] , \w[22][25] , \w[22][24] , 
        \w[22][23] , \w[22][22] , \w[22][21] , \w[22][20] , \w[22][19] , 
        \w[22][18] , \w[22][17] , \w[22][16] , \w[22][15] , \w[22][14] , 
        \w[22][13] , \w[22][12] , \w[22][11] , \w[22][10] , \w[22][9] , 
        \w[22][8] , \w[22][7] , \w[22][6] , \w[22][5] , \w[22][4] , \w[22][3] , 
        \w[22][2] , \w[22][1] , SYNOPSYS_UNCONNECTED__20}) );
  ADD_N32_168 \FAINST[22].ADD_  ( .A({\_42_net_[31] , \_42_net_[30] , 
        \_42_net_[29] , \_42_net_[28] , \_42_net_[27] , \_42_net_[26] , 
        \_42_net_[25] , \_42_net_[24] , \_42_net_[23] , \_42_net_[22] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[22][31] , \w[22][30] , \w[22][29] , \w[22][28] , \w[22][27] , 
        \w[22][26] , \w[22][25] , \w[22][24] , \w[22][23] , \w[22][22] , 
        \w[22][21] , \w[22][20] , \w[22][19] , \w[22][18] , \w[22][17] , 
        \w[22][16] , \w[22][15] , \w[22][14] , \w[22][13] , \w[22][12] , 
        \w[22][11] , \w[22][10] , \w[22][9] , \w[22][8] , \w[22][7] , 
        \w[22][6] , \w[22][5] , \w[22][4] , \w[22][3] , \w[22][2] , \w[22][1] , 
        1'b0}), .CI(1'b0), .S({\w[23][31] , \w[23][30] , \w[23][29] , 
        \w[23][28] , \w[23][27] , \w[23][26] , \w[23][25] , \w[23][24] , 
        \w[23][23] , \w[23][22] , \w[23][21] , \w[23][20] , \w[23][19] , 
        \w[23][18] , \w[23][17] , \w[23][16] , \w[23][15] , \w[23][14] , 
        \w[23][13] , \w[23][12] , \w[23][11] , \w[23][10] , \w[23][9] , 
        \w[23][8] , \w[23][7] , \w[23][6] , \w[23][5] , \w[23][4] , \w[23][3] , 
        \w[23][2] , \w[23][1] , SYNOPSYS_UNCONNECTED__21}) );
  ADD_N32_167 \FAINST[23].ADD_  ( .A({\_44_net_[31] , \_44_net_[30] , 
        \_44_net_[29] , \_44_net_[28] , \_44_net_[27] , \_44_net_[26] , 
        \_44_net_[25] , \_44_net_[24] , \_44_net_[23] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[23][31] , 
        \w[23][30] , \w[23][29] , \w[23][28] , \w[23][27] , \w[23][26] , 
        \w[23][25] , \w[23][24] , \w[23][23] , \w[23][22] , \w[23][21] , 
        \w[23][20] , \w[23][19] , \w[23][18] , \w[23][17] , \w[23][16] , 
        \w[23][15] , \w[23][14] , \w[23][13] , \w[23][12] , \w[23][11] , 
        \w[23][10] , \w[23][9] , \w[23][8] , \w[23][7] , \w[23][6] , 
        \w[23][5] , \w[23][4] , \w[23][3] , \w[23][2] , \w[23][1] , 1'b0}), 
        .CI(1'b0), .S({\w[24][31] , \w[24][30] , \w[24][29] , \w[24][28] , 
        \w[24][27] , \w[24][26] , \w[24][25] , \w[24][24] , \w[24][23] , 
        \w[24][22] , \w[24][21] , \w[24][20] , \w[24][19] , \w[24][18] , 
        \w[24][17] , \w[24][16] , \w[24][15] , \w[24][14] , \w[24][13] , 
        \w[24][12] , \w[24][11] , \w[24][10] , \w[24][9] , \w[24][8] , 
        \w[24][7] , \w[24][6] , \w[24][5] , \w[24][4] , \w[24][3] , \w[24][2] , 
        \w[24][1] , SYNOPSYS_UNCONNECTED__22}) );
  ADD_N32_166 \FAINST[24].ADD_  ( .A({\_46_net_[31] , \_46_net_[30] , 
        \_46_net_[29] , \_46_net_[28] , \_46_net_[27] , \_46_net_[26] , 
        \_46_net_[25] , \_46_net_[24] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[24][31] , \w[24][30] , 
        \w[24][29] , \w[24][28] , \w[24][27] , \w[24][26] , \w[24][25] , 
        \w[24][24] , \w[24][23] , \w[24][22] , \w[24][21] , \w[24][20] , 
        \w[24][19] , \w[24][18] , \w[24][17] , \w[24][16] , \w[24][15] , 
        \w[24][14] , \w[24][13] , \w[24][12] , \w[24][11] , \w[24][10] , 
        \w[24][9] , \w[24][8] , \w[24][7] , \w[24][6] , \w[24][5] , \w[24][4] , 
        \w[24][3] , \w[24][2] , \w[24][1] , 1'b0}), .CI(1'b0), .S({\w[25][31] , 
        \w[25][30] , \w[25][29] , \w[25][28] , \w[25][27] , \w[25][26] , 
        \w[25][25] , \w[25][24] , \w[25][23] , \w[25][22] , \w[25][21] , 
        \w[25][20] , \w[25][19] , \w[25][18] , \w[25][17] , \w[25][16] , 
        \w[25][15] , \w[25][14] , \w[25][13] , \w[25][12] , \w[25][11] , 
        \w[25][10] , \w[25][9] , \w[25][8] , \w[25][7] , \w[25][6] , 
        \w[25][5] , \w[25][4] , \w[25][3] , \w[25][2] , \w[25][1] , 
        SYNOPSYS_UNCONNECTED__23}) );
  ADD_N32_165 \FAINST[25].ADD_  ( .A({\_48_net_[31] , \_48_net_[30] , 
        \_48_net_[29] , \_48_net_[28] , \_48_net_[27] , \_48_net_[26] , 
        \_48_net_[25] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[25][31] , \w[25][30] , \w[25][29] , 
        \w[25][28] , \w[25][27] , \w[25][26] , \w[25][25] , \w[25][24] , 
        \w[25][23] , \w[25][22] , \w[25][21] , \w[25][20] , \w[25][19] , 
        \w[25][18] , \w[25][17] , \w[25][16] , \w[25][15] , \w[25][14] , 
        \w[25][13] , \w[25][12] , \w[25][11] , \w[25][10] , \w[25][9] , 
        \w[25][8] , \w[25][7] , \w[25][6] , \w[25][5] , \w[25][4] , \w[25][3] , 
        \w[25][2] , \w[25][1] , 1'b0}), .CI(1'b0), .S({\w[26][31] , 
        \w[26][30] , \w[26][29] , \w[26][28] , \w[26][27] , \w[26][26] , 
        \w[26][25] , \w[26][24] , \w[26][23] , \w[26][22] , \w[26][21] , 
        \w[26][20] , \w[26][19] , \w[26][18] , \w[26][17] , \w[26][16] , 
        \w[26][15] , \w[26][14] , \w[26][13] , \w[26][12] , \w[26][11] , 
        \w[26][10] , \w[26][9] , \w[26][8] , \w[26][7] , \w[26][6] , 
        \w[26][5] , \w[26][4] , \w[26][3] , \w[26][2] , \w[26][1] , 
        SYNOPSYS_UNCONNECTED__24}) );
  ADD_N32_164 \FAINST[26].ADD_  ( .A({\_50_net_[31] , \_50_net_[30] , 
        \_50_net_[29] , \_50_net_[28] , \_50_net_[27] , \_50_net_[26] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({\w[26][31] , \w[26][30] , \w[26][29] , \w[26][28] , 
        \w[26][27] , \w[26][26] , \w[26][25] , \w[26][24] , \w[26][23] , 
        \w[26][22] , \w[26][21] , \w[26][20] , \w[26][19] , \w[26][18] , 
        \w[26][17] , \w[26][16] , \w[26][15] , \w[26][14] , \w[26][13] , 
        \w[26][12] , \w[26][11] , \w[26][10] , \w[26][9] , \w[26][8] , 
        \w[26][7] , \w[26][6] , \w[26][5] , \w[26][4] , \w[26][3] , \w[26][2] , 
        \w[26][1] , 1'b0}), .CI(1'b0), .S({\w[27][31] , \w[27][30] , 
        \w[27][29] , \w[27][28] , \w[27][27] , \w[27][26] , \w[27][25] , 
        \w[27][24] , \w[27][23] , \w[27][22] , \w[27][21] , \w[27][20] , 
        \w[27][19] , \w[27][18] , \w[27][17] , \w[27][16] , \w[27][15] , 
        \w[27][14] , \w[27][13] , \w[27][12] , \w[27][11] , \w[27][10] , 
        \w[27][9] , \w[27][8] , \w[27][7] , \w[27][6] , \w[27][5] , \w[27][4] , 
        \w[27][3] , \w[27][2] , \w[27][1] , SYNOPSYS_UNCONNECTED__25}) );
  ADD_N32_163 \FAINST[27].ADD_  ( .A({\_52_net_[31] , \_52_net_[30] , 
        \_52_net_[29] , \_52_net_[28] , \_52_net_[27] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({\w[27][31] , \w[27][30] , \w[27][29] , \w[27][28] , \w[27][27] , 
        \w[27][26] , \w[27][25] , \w[27][24] , \w[27][23] , \w[27][22] , 
        \w[27][21] , \w[27][20] , \w[27][19] , \w[27][18] , \w[27][17] , 
        \w[27][16] , \w[27][15] , \w[27][14] , \w[27][13] , \w[27][12] , 
        \w[27][11] , \w[27][10] , \w[27][9] , \w[27][8] , \w[27][7] , 
        \w[27][6] , \w[27][5] , \w[27][4] , \w[27][3] , \w[27][2] , \w[27][1] , 
        1'b0}), .CI(1'b0), .S({\w[28][31] , \w[28][30] , \w[28][29] , 
        \w[28][28] , \w[28][27] , \w[28][26] , \w[28][25] , \w[28][24] , 
        \w[28][23] , \w[28][22] , \w[28][21] , \w[28][20] , \w[28][19] , 
        \w[28][18] , \w[28][17] , \w[28][16] , \w[28][15] , \w[28][14] , 
        \w[28][13] , \w[28][12] , \w[28][11] , \w[28][10] , \w[28][9] , 
        \w[28][8] , \w[28][7] , \w[28][6] , \w[28][5] , \w[28][4] , \w[28][3] , 
        \w[28][2] , \w[28][1] , SYNOPSYS_UNCONNECTED__26}) );
  ADD_N32_162 \FAINST[28].ADD_  ( .A({\_54_net_[31] , \_54_net_[30] , 
        \_54_net_[29] , \_54_net_[28] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[28][31] , \w[28][30] , \w[28][29] , \w[28][28] , \w[28][27] , 
        \w[28][26] , \w[28][25] , \w[28][24] , \w[28][23] , \w[28][22] , 
        \w[28][21] , \w[28][20] , \w[28][19] , \w[28][18] , \w[28][17] , 
        \w[28][16] , \w[28][15] , \w[28][14] , \w[28][13] , \w[28][12] , 
        \w[28][11] , \w[28][10] , \w[28][9] , \w[28][8] , \w[28][7] , 
        \w[28][6] , \w[28][5] , \w[28][4] , \w[28][3] , \w[28][2] , \w[28][1] , 
        1'b0}), .CI(1'b0), .S({\w[29][31] , \w[29][30] , \w[29][29] , 
        \w[29][28] , \w[29][27] , \w[29][26] , \w[29][25] , \w[29][24] , 
        \w[29][23] , \w[29][22] , \w[29][21] , \w[29][20] , \w[29][19] , 
        \w[29][18] , \w[29][17] , \w[29][16] , \w[29][15] , \w[29][14] , 
        \w[29][13] , \w[29][12] , \w[29][11] , \w[29][10] , \w[29][9] , 
        \w[29][8] , \w[29][7] , \w[29][6] , \w[29][5] , \w[29][4] , \w[29][3] , 
        \w[29][2] , \w[29][1] , SYNOPSYS_UNCONNECTED__27}) );
  ADD_N32_161 \FAINST[29].ADD_  ( .A({\_56_net_[31] , \_56_net_[30] , 
        \_56_net_[29] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[29][31] , 
        \w[29][30] , \w[29][29] , \w[29][28] , \w[29][27] , \w[29][26] , 
        \w[29][25] , \w[29][24] , \w[29][23] , \w[29][22] , \w[29][21] , 
        \w[29][20] , \w[29][19] , \w[29][18] , \w[29][17] , \w[29][16] , 
        \w[29][15] , \w[29][14] , \w[29][13] , \w[29][12] , \w[29][11] , 
        \w[29][10] , \w[29][9] , \w[29][8] , \w[29][7] , \w[29][6] , 
        \w[29][5] , \w[29][4] , \w[29][3] , \w[29][2] , \w[29][1] , 1'b0}), 
        .CI(1'b0), .S({\w[30][31] , \w[30][30] , \w[30][29] , \w[30][28] , 
        \w[30][27] , \w[30][26] , \w[30][25] , \w[30][24] , \w[30][23] , 
        \w[30][22] , \w[30][21] , \w[30][20] , \w[30][19] , \w[30][18] , 
        \w[30][17] , \w[30][16] , \w[30][15] , \w[30][14] , \w[30][13] , 
        \w[30][12] , \w[30][11] , \w[30][10] , \w[30][9] , \w[30][8] , 
        \w[30][7] , \w[30][6] , \w[30][5] , \w[30][4] , \w[30][3] , \w[30][2] , 
        \w[30][1] , SYNOPSYS_UNCONNECTED__28}) );
  ADD_N32_160 \FAINST[30].ADD_  ( .A({\_58_net_[31] , \_58_net_[30] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[30][31] , \w[30][30] , 
        \w[30][29] , \w[30][28] , \w[30][27] , \w[30][26] , \w[30][25] , 
        \w[30][24] , \w[30][23] , \w[30][22] , \w[30][21] , \w[30][20] , 
        \w[30][19] , \w[30][18] , \w[30][17] , \w[30][16] , \w[30][15] , 
        \w[30][14] , \w[30][13] , \w[30][12] , \w[30][11] , \w[30][10] , 
        \w[30][9] , \w[30][8] , \w[30][7] , \w[30][6] , \w[30][5] , \w[30][4] , 
        \w[30][3] , \w[30][2] , \w[30][1] , 1'b0}), .CI(1'b0), .S({\w[31][31] , 
        \w[31][30] , \w[31][29] , \w[31][28] , \w[31][27] , \w[31][26] , 
        \w[31][25] , \w[31][24] , \w[31][23] , \w[31][22] , \w[31][21] , 
        \w[31][20] , \w[31][19] , \w[31][18] , \w[31][17] , \w[31][16] , 
        \w[31][15] , \w[31][14] , \w[31][13] , \w[31][12] , \w[31][11] , 
        \w[31][10] , \w[31][9] , \w[31][8] , \w[31][7] , \w[31][6] , 
        \w[31][5] , \w[31][4] , \w[31][3] , \w[31][2] , \w[31][1] , 
        SYNOPSYS_UNCONNECTED__29}) );
  ADD_N32_159 \FAINST[31].ADD_  ( .A({\_60_net_[31] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({\w[31][31] , \w[31][30] , \w[31][29] , 
        \w[31][28] , \w[31][27] , \w[31][26] , \w[31][25] , \w[31][24] , 
        \w[31][23] , \w[31][22] , \w[31][21] , \w[31][20] , \w[31][19] , 
        \w[31][18] , \w[31][17] , \w[31][16] , \w[31][15] , \w[31][14] , 
        \w[31][13] , \w[31][12] , \w[31][11] , \w[31][10] , \w[31][9] , 
        \w[31][8] , \w[31][7] , \w[31][6] , \w[31][5] , \w[31][4] , \w[31][3] , 
        \w[31][2] , \w[31][1] , 1'b0}), .CI(1'b0), .S({O[31:1], 
        SYNOPSYS_UNCONNECTED__30}) );
  AND U2 ( .A(A[5]), .B(B[4]), .Z(\_8_net_[9] ) );
  AND U3 ( .A(A[5]), .B(B[3]), .Z(\_8_net_[8] ) );
  AND U4 ( .A(A[5]), .B(B[2]), .Z(\_8_net_[7] ) );
  AND U5 ( .A(A[5]), .B(B[1]), .Z(\_8_net_[6] ) );
  AND U6 ( .A(A[5]), .B(B[0]), .Z(\_8_net_[5] ) );
  AND U7 ( .A(A[5]), .B(B[26]), .Z(\_8_net_[31] ) );
  AND U8 ( .A(A[5]), .B(B[25]), .Z(\_8_net_[30] ) );
  AND U9 ( .A(A[5]), .B(B[24]), .Z(\_8_net_[29] ) );
  AND U10 ( .A(A[5]), .B(B[23]), .Z(\_8_net_[28] ) );
  AND U11 ( .A(A[5]), .B(B[22]), .Z(\_8_net_[27] ) );
  AND U12 ( .A(A[5]), .B(B[21]), .Z(\_8_net_[26] ) );
  AND U13 ( .A(A[5]), .B(B[20]), .Z(\_8_net_[25] ) );
  AND U14 ( .A(A[5]), .B(B[19]), .Z(\_8_net_[24] ) );
  AND U15 ( .A(A[5]), .B(B[18]), .Z(\_8_net_[23] ) );
  AND U16 ( .A(A[5]), .B(B[17]), .Z(\_8_net_[22] ) );
  AND U17 ( .A(A[5]), .B(B[16]), .Z(\_8_net_[21] ) );
  AND U18 ( .A(A[5]), .B(B[15]), .Z(\_8_net_[20] ) );
  AND U19 ( .A(A[5]), .B(B[14]), .Z(\_8_net_[19] ) );
  AND U20 ( .A(A[5]), .B(B[13]), .Z(\_8_net_[18] ) );
  AND U21 ( .A(A[5]), .B(B[12]), .Z(\_8_net_[17] ) );
  AND U22 ( .A(A[5]), .B(B[11]), .Z(\_8_net_[16] ) );
  AND U23 ( .A(A[5]), .B(B[10]), .Z(\_8_net_[15] ) );
  AND U24 ( .A(A[5]), .B(B[9]), .Z(\_8_net_[14] ) );
  AND U25 ( .A(A[5]), .B(B[8]), .Z(\_8_net_[13] ) );
  AND U26 ( .A(A[5]), .B(B[7]), .Z(\_8_net_[12] ) );
  AND U27 ( .A(A[5]), .B(B[6]), .Z(\_8_net_[11] ) );
  AND U28 ( .A(A[5]), .B(B[5]), .Z(\_8_net_[10] ) );
  AND U29 ( .A(B[5]), .B(A[4]), .Z(\_6_net_[9] ) );
  AND U30 ( .A(B[4]), .B(A[4]), .Z(\_6_net_[8] ) );
  AND U31 ( .A(B[3]), .B(A[4]), .Z(\_6_net_[7] ) );
  AND U32 ( .A(B[2]), .B(A[4]), .Z(\_6_net_[6] ) );
  AND U33 ( .A(B[1]), .B(A[4]), .Z(\_6_net_[5] ) );
  AND U34 ( .A(B[0]), .B(A[4]), .Z(\_6_net_[4] ) );
  AND U35 ( .A(A[4]), .B(B[27]), .Z(\_6_net_[31] ) );
  AND U36 ( .A(B[26]), .B(A[4]), .Z(\_6_net_[30] ) );
  AND U37 ( .A(B[25]), .B(A[4]), .Z(\_6_net_[29] ) );
  AND U38 ( .A(B[24]), .B(A[4]), .Z(\_6_net_[28] ) );
  AND U39 ( .A(B[23]), .B(A[4]), .Z(\_6_net_[27] ) );
  AND U40 ( .A(B[22]), .B(A[4]), .Z(\_6_net_[26] ) );
  AND U41 ( .A(B[21]), .B(A[4]), .Z(\_6_net_[25] ) );
  AND U42 ( .A(B[20]), .B(A[4]), .Z(\_6_net_[24] ) );
  AND U43 ( .A(B[19]), .B(A[4]), .Z(\_6_net_[23] ) );
  AND U44 ( .A(B[18]), .B(A[4]), .Z(\_6_net_[22] ) );
  AND U45 ( .A(B[17]), .B(A[4]), .Z(\_6_net_[21] ) );
  AND U46 ( .A(B[16]), .B(A[4]), .Z(\_6_net_[20] ) );
  AND U47 ( .A(B[15]), .B(A[4]), .Z(\_6_net_[19] ) );
  AND U48 ( .A(B[14]), .B(A[4]), .Z(\_6_net_[18] ) );
  AND U49 ( .A(B[13]), .B(A[4]), .Z(\_6_net_[17] ) );
  AND U50 ( .A(B[12]), .B(A[4]), .Z(\_6_net_[16] ) );
  AND U51 ( .A(B[11]), .B(A[4]), .Z(\_6_net_[15] ) );
  AND U52 ( .A(B[10]), .B(A[4]), .Z(\_6_net_[14] ) );
  AND U53 ( .A(B[9]), .B(A[4]), .Z(\_6_net_[13] ) );
  AND U54 ( .A(B[8]), .B(A[4]), .Z(\_6_net_[12] ) );
  AND U55 ( .A(B[7]), .B(A[4]), .Z(\_6_net_[11] ) );
  AND U56 ( .A(B[6]), .B(A[4]), .Z(\_6_net_[10] ) );
  AND U57 ( .A(A[31]), .B(B[0]), .Z(\_60_net_[31] ) );
  AND U58 ( .A(B[1]), .B(A[30]), .Z(\_58_net_[31] ) );
  AND U59 ( .A(A[30]), .B(B[0]), .Z(\_58_net_[30] ) );
  AND U60 ( .A(B[2]), .B(A[29]), .Z(\_56_net_[31] ) );
  AND U61 ( .A(B[1]), .B(A[29]), .Z(\_56_net_[30] ) );
  AND U62 ( .A(A[29]), .B(B[0]), .Z(\_56_net_[29] ) );
  AND U63 ( .A(B[3]), .B(A[28]), .Z(\_54_net_[31] ) );
  AND U64 ( .A(B[2]), .B(A[28]), .Z(\_54_net_[30] ) );
  AND U65 ( .A(B[1]), .B(A[28]), .Z(\_54_net_[29] ) );
  AND U66 ( .A(A[28]), .B(B[0]), .Z(\_54_net_[28] ) );
  AND U67 ( .A(B[4]), .B(A[27]), .Z(\_52_net_[31] ) );
  AND U68 ( .A(B[3]), .B(A[27]), .Z(\_52_net_[30] ) );
  AND U69 ( .A(B[2]), .B(A[27]), .Z(\_52_net_[29] ) );
  AND U70 ( .A(B[1]), .B(A[27]), .Z(\_52_net_[28] ) );
  AND U71 ( .A(A[27]), .B(B[0]), .Z(\_52_net_[27] ) );
  AND U72 ( .A(B[5]), .B(A[26]), .Z(\_50_net_[31] ) );
  AND U73 ( .A(B[4]), .B(A[26]), .Z(\_50_net_[30] ) );
  AND U74 ( .A(B[3]), .B(A[26]), .Z(\_50_net_[29] ) );
  AND U75 ( .A(B[2]), .B(A[26]), .Z(\_50_net_[28] ) );
  AND U76 ( .A(B[1]), .B(A[26]), .Z(\_50_net_[27] ) );
  AND U77 ( .A(A[26]), .B(B[0]), .Z(\_50_net_[26] ) );
  AND U78 ( .A(B[6]), .B(A[3]), .Z(\_4_net_[9] ) );
  AND U79 ( .A(B[5]), .B(A[3]), .Z(\_4_net_[8] ) );
  AND U80 ( .A(B[4]), .B(A[3]), .Z(\_4_net_[7] ) );
  AND U81 ( .A(B[3]), .B(A[3]), .Z(\_4_net_[6] ) );
  AND U82 ( .A(B[2]), .B(A[3]), .Z(\_4_net_[5] ) );
  AND U83 ( .A(B[1]), .B(A[3]), .Z(\_4_net_[4] ) );
  AND U84 ( .A(B[0]), .B(A[3]), .Z(\_4_net_[3] ) );
  AND U85 ( .A(A[3]), .B(B[28]), .Z(\_4_net_[31] ) );
  AND U86 ( .A(B[27]), .B(A[3]), .Z(\_4_net_[30] ) );
  AND U87 ( .A(B[26]), .B(A[3]), .Z(\_4_net_[29] ) );
  AND U88 ( .A(B[25]), .B(A[3]), .Z(\_4_net_[28] ) );
  AND U89 ( .A(B[24]), .B(A[3]), .Z(\_4_net_[27] ) );
  AND U90 ( .A(B[23]), .B(A[3]), .Z(\_4_net_[26] ) );
  AND U91 ( .A(B[22]), .B(A[3]), .Z(\_4_net_[25] ) );
  AND U92 ( .A(B[21]), .B(A[3]), .Z(\_4_net_[24] ) );
  AND U93 ( .A(B[20]), .B(A[3]), .Z(\_4_net_[23] ) );
  AND U94 ( .A(B[19]), .B(A[3]), .Z(\_4_net_[22] ) );
  AND U95 ( .A(B[18]), .B(A[3]), .Z(\_4_net_[21] ) );
  AND U96 ( .A(B[17]), .B(A[3]), .Z(\_4_net_[20] ) );
  AND U97 ( .A(B[16]), .B(A[3]), .Z(\_4_net_[19] ) );
  AND U98 ( .A(B[15]), .B(A[3]), .Z(\_4_net_[18] ) );
  AND U99 ( .A(B[14]), .B(A[3]), .Z(\_4_net_[17] ) );
  AND U100 ( .A(B[13]), .B(A[3]), .Z(\_4_net_[16] ) );
  AND U101 ( .A(B[12]), .B(A[3]), .Z(\_4_net_[15] ) );
  AND U102 ( .A(B[11]), .B(A[3]), .Z(\_4_net_[14] ) );
  AND U103 ( .A(B[10]), .B(A[3]), .Z(\_4_net_[13] ) );
  AND U104 ( .A(B[9]), .B(A[3]), .Z(\_4_net_[12] ) );
  AND U105 ( .A(B[8]), .B(A[3]), .Z(\_4_net_[11] ) );
  AND U106 ( .A(B[7]), .B(A[3]), .Z(\_4_net_[10] ) );
  AND U107 ( .A(B[6]), .B(A[25]), .Z(\_48_net_[31] ) );
  AND U108 ( .A(B[5]), .B(A[25]), .Z(\_48_net_[30] ) );
  AND U109 ( .A(B[4]), .B(A[25]), .Z(\_48_net_[29] ) );
  AND U110 ( .A(B[3]), .B(A[25]), .Z(\_48_net_[28] ) );
  AND U111 ( .A(B[2]), .B(A[25]), .Z(\_48_net_[27] ) );
  AND U112 ( .A(B[1]), .B(A[25]), .Z(\_48_net_[26] ) );
  AND U113 ( .A(A[25]), .B(B[0]), .Z(\_48_net_[25] ) );
  AND U114 ( .A(B[7]), .B(A[24]), .Z(\_46_net_[31] ) );
  AND U115 ( .A(B[6]), .B(A[24]), .Z(\_46_net_[30] ) );
  AND U116 ( .A(B[5]), .B(A[24]), .Z(\_46_net_[29] ) );
  AND U117 ( .A(B[4]), .B(A[24]), .Z(\_46_net_[28] ) );
  AND U118 ( .A(B[3]), .B(A[24]), .Z(\_46_net_[27] ) );
  AND U119 ( .A(B[2]), .B(A[24]), .Z(\_46_net_[26] ) );
  AND U120 ( .A(B[1]), .B(A[24]), .Z(\_46_net_[25] ) );
  AND U121 ( .A(A[24]), .B(B[0]), .Z(\_46_net_[24] ) );
  AND U122 ( .A(B[8]), .B(A[23]), .Z(\_44_net_[31] ) );
  AND U123 ( .A(B[7]), .B(A[23]), .Z(\_44_net_[30] ) );
  AND U124 ( .A(B[6]), .B(A[23]), .Z(\_44_net_[29] ) );
  AND U125 ( .A(B[5]), .B(A[23]), .Z(\_44_net_[28] ) );
  AND U126 ( .A(B[4]), .B(A[23]), .Z(\_44_net_[27] ) );
  AND U127 ( .A(B[3]), .B(A[23]), .Z(\_44_net_[26] ) );
  AND U128 ( .A(B[2]), .B(A[23]), .Z(\_44_net_[25] ) );
  AND U129 ( .A(B[1]), .B(A[23]), .Z(\_44_net_[24] ) );
  AND U130 ( .A(A[23]), .B(B[0]), .Z(\_44_net_[23] ) );
  AND U131 ( .A(B[9]), .B(A[22]), .Z(\_42_net_[31] ) );
  AND U132 ( .A(B[8]), .B(A[22]), .Z(\_42_net_[30] ) );
  AND U133 ( .A(B[7]), .B(A[22]), .Z(\_42_net_[29] ) );
  AND U134 ( .A(B[6]), .B(A[22]), .Z(\_42_net_[28] ) );
  AND U135 ( .A(B[5]), .B(A[22]), .Z(\_42_net_[27] ) );
  AND U136 ( .A(B[4]), .B(A[22]), .Z(\_42_net_[26] ) );
  AND U137 ( .A(B[3]), .B(A[22]), .Z(\_42_net_[25] ) );
  AND U138 ( .A(B[2]), .B(A[22]), .Z(\_42_net_[24] ) );
  AND U139 ( .A(B[1]), .B(A[22]), .Z(\_42_net_[23] ) );
  AND U140 ( .A(A[22]), .B(B[0]), .Z(\_42_net_[22] ) );
  AND U141 ( .A(B[10]), .B(A[21]), .Z(\_40_net_[31] ) );
  AND U142 ( .A(B[9]), .B(A[21]), .Z(\_40_net_[30] ) );
  AND U143 ( .A(B[8]), .B(A[21]), .Z(\_40_net_[29] ) );
  AND U144 ( .A(B[7]), .B(A[21]), .Z(\_40_net_[28] ) );
  AND U145 ( .A(B[6]), .B(A[21]), .Z(\_40_net_[27] ) );
  AND U146 ( .A(B[5]), .B(A[21]), .Z(\_40_net_[26] ) );
  AND U147 ( .A(B[4]), .B(A[21]), .Z(\_40_net_[25] ) );
  AND U148 ( .A(B[3]), .B(A[21]), .Z(\_40_net_[24] ) );
  AND U149 ( .A(B[2]), .B(A[21]), .Z(\_40_net_[23] ) );
  AND U150 ( .A(B[1]), .B(A[21]), .Z(\_40_net_[22] ) );
  AND U151 ( .A(A[21]), .B(B[0]), .Z(\_40_net_[21] ) );
  AND U152 ( .A(B[11]), .B(A[20]), .Z(\_38_net_[31] ) );
  AND U153 ( .A(B[10]), .B(A[20]), .Z(\_38_net_[30] ) );
  AND U154 ( .A(B[9]), .B(A[20]), .Z(\_38_net_[29] ) );
  AND U155 ( .A(B[8]), .B(A[20]), .Z(\_38_net_[28] ) );
  AND U156 ( .A(B[7]), .B(A[20]), .Z(\_38_net_[27] ) );
  AND U157 ( .A(B[6]), .B(A[20]), .Z(\_38_net_[26] ) );
  AND U158 ( .A(B[5]), .B(A[20]), .Z(\_38_net_[25] ) );
  AND U159 ( .A(B[4]), .B(A[20]), .Z(\_38_net_[24] ) );
  AND U160 ( .A(B[3]), .B(A[20]), .Z(\_38_net_[23] ) );
  AND U161 ( .A(B[2]), .B(A[20]), .Z(\_38_net_[22] ) );
  AND U162 ( .A(B[1]), .B(A[20]), .Z(\_38_net_[21] ) );
  AND U163 ( .A(A[20]), .B(B[0]), .Z(\_38_net_[20] ) );
  AND U164 ( .A(B[12]), .B(A[19]), .Z(\_36_net_[31] ) );
  AND U165 ( .A(B[11]), .B(A[19]), .Z(\_36_net_[30] ) );
  AND U166 ( .A(B[10]), .B(A[19]), .Z(\_36_net_[29] ) );
  AND U167 ( .A(B[9]), .B(A[19]), .Z(\_36_net_[28] ) );
  AND U168 ( .A(B[8]), .B(A[19]), .Z(\_36_net_[27] ) );
  AND U169 ( .A(B[7]), .B(A[19]), .Z(\_36_net_[26] ) );
  AND U170 ( .A(B[6]), .B(A[19]), .Z(\_36_net_[25] ) );
  AND U171 ( .A(B[5]), .B(A[19]), .Z(\_36_net_[24] ) );
  AND U172 ( .A(B[4]), .B(A[19]), .Z(\_36_net_[23] ) );
  AND U173 ( .A(B[3]), .B(A[19]), .Z(\_36_net_[22] ) );
  AND U174 ( .A(B[2]), .B(A[19]), .Z(\_36_net_[21] ) );
  AND U175 ( .A(B[1]), .B(A[19]), .Z(\_36_net_[20] ) );
  AND U176 ( .A(A[19]), .B(B[0]), .Z(\_36_net_[19] ) );
  AND U177 ( .A(B[13]), .B(A[18]), .Z(\_34_net_[31] ) );
  AND U178 ( .A(B[12]), .B(A[18]), .Z(\_34_net_[30] ) );
  AND U179 ( .A(B[11]), .B(A[18]), .Z(\_34_net_[29] ) );
  AND U180 ( .A(B[10]), .B(A[18]), .Z(\_34_net_[28] ) );
  AND U181 ( .A(B[9]), .B(A[18]), .Z(\_34_net_[27] ) );
  AND U182 ( .A(B[8]), .B(A[18]), .Z(\_34_net_[26] ) );
  AND U183 ( .A(B[7]), .B(A[18]), .Z(\_34_net_[25] ) );
  AND U184 ( .A(B[6]), .B(A[18]), .Z(\_34_net_[24] ) );
  AND U185 ( .A(B[5]), .B(A[18]), .Z(\_34_net_[23] ) );
  AND U186 ( .A(B[4]), .B(A[18]), .Z(\_34_net_[22] ) );
  AND U187 ( .A(B[3]), .B(A[18]), .Z(\_34_net_[21] ) );
  AND U188 ( .A(B[2]), .B(A[18]), .Z(\_34_net_[20] ) );
  AND U189 ( .A(B[1]), .B(A[18]), .Z(\_34_net_[19] ) );
  AND U190 ( .A(A[18]), .B(B[0]), .Z(\_34_net_[18] ) );
  AND U191 ( .A(B[14]), .B(A[17]), .Z(\_32_net_[31] ) );
  AND U192 ( .A(B[13]), .B(A[17]), .Z(\_32_net_[30] ) );
  AND U193 ( .A(B[12]), .B(A[17]), .Z(\_32_net_[29] ) );
  AND U194 ( .A(B[11]), .B(A[17]), .Z(\_32_net_[28] ) );
  AND U195 ( .A(B[10]), .B(A[17]), .Z(\_32_net_[27] ) );
  AND U196 ( .A(B[9]), .B(A[17]), .Z(\_32_net_[26] ) );
  AND U197 ( .A(B[8]), .B(A[17]), .Z(\_32_net_[25] ) );
  AND U198 ( .A(B[7]), .B(A[17]), .Z(\_32_net_[24] ) );
  AND U199 ( .A(B[6]), .B(A[17]), .Z(\_32_net_[23] ) );
  AND U200 ( .A(B[5]), .B(A[17]), .Z(\_32_net_[22] ) );
  AND U201 ( .A(B[4]), .B(A[17]), .Z(\_32_net_[21] ) );
  AND U202 ( .A(B[3]), .B(A[17]), .Z(\_32_net_[20] ) );
  AND U203 ( .A(B[2]), .B(A[17]), .Z(\_32_net_[19] ) );
  AND U204 ( .A(B[1]), .B(A[17]), .Z(\_32_net_[18] ) );
  AND U205 ( .A(A[17]), .B(B[0]), .Z(\_32_net_[17] ) );
  AND U206 ( .A(B[15]), .B(A[16]), .Z(\_30_net_[31] ) );
  AND U207 ( .A(B[14]), .B(A[16]), .Z(\_30_net_[30] ) );
  AND U208 ( .A(B[13]), .B(A[16]), .Z(\_30_net_[29] ) );
  AND U209 ( .A(B[12]), .B(A[16]), .Z(\_30_net_[28] ) );
  AND U210 ( .A(B[11]), .B(A[16]), .Z(\_30_net_[27] ) );
  AND U211 ( .A(B[10]), .B(A[16]), .Z(\_30_net_[26] ) );
  AND U212 ( .A(B[9]), .B(A[16]), .Z(\_30_net_[25] ) );
  AND U213 ( .A(B[8]), .B(A[16]), .Z(\_30_net_[24] ) );
  AND U214 ( .A(B[7]), .B(A[16]), .Z(\_30_net_[23] ) );
  AND U215 ( .A(B[6]), .B(A[16]), .Z(\_30_net_[22] ) );
  AND U216 ( .A(B[5]), .B(A[16]), .Z(\_30_net_[21] ) );
  AND U217 ( .A(B[4]), .B(A[16]), .Z(\_30_net_[20] ) );
  AND U218 ( .A(B[3]), .B(A[16]), .Z(\_30_net_[19] ) );
  AND U219 ( .A(B[2]), .B(A[16]), .Z(\_30_net_[18] ) );
  AND U220 ( .A(B[1]), .B(A[16]), .Z(\_30_net_[17] ) );
  AND U221 ( .A(A[16]), .B(B[0]), .Z(\_30_net_[16] ) );
  AND U222 ( .A(B[7]), .B(A[2]), .Z(\_2_net_[9] ) );
  AND U223 ( .A(B[6]), .B(A[2]), .Z(\_2_net_[8] ) );
  AND U224 ( .A(B[5]), .B(A[2]), .Z(\_2_net_[7] ) );
  AND U225 ( .A(B[4]), .B(A[2]), .Z(\_2_net_[6] ) );
  AND U226 ( .A(B[3]), .B(A[2]), .Z(\_2_net_[5] ) );
  AND U227 ( .A(B[2]), .B(A[2]), .Z(\_2_net_[4] ) );
  AND U228 ( .A(B[1]), .B(A[2]), .Z(\_2_net_[3] ) );
  AND U229 ( .A(A[2]), .B(B[29]), .Z(\_2_net_[31] ) );
  AND U230 ( .A(B[28]), .B(A[2]), .Z(\_2_net_[30] ) );
  AND U231 ( .A(B[0]), .B(A[2]), .Z(\_2_net_[2] ) );
  AND U232 ( .A(B[27]), .B(A[2]), .Z(\_2_net_[29] ) );
  AND U233 ( .A(B[26]), .B(A[2]), .Z(\_2_net_[28] ) );
  AND U234 ( .A(B[25]), .B(A[2]), .Z(\_2_net_[27] ) );
  AND U235 ( .A(B[24]), .B(A[2]), .Z(\_2_net_[26] ) );
  AND U236 ( .A(B[23]), .B(A[2]), .Z(\_2_net_[25] ) );
  AND U237 ( .A(B[22]), .B(A[2]), .Z(\_2_net_[24] ) );
  AND U238 ( .A(B[21]), .B(A[2]), .Z(\_2_net_[23] ) );
  AND U239 ( .A(B[20]), .B(A[2]), .Z(\_2_net_[22] ) );
  AND U240 ( .A(B[19]), .B(A[2]), .Z(\_2_net_[21] ) );
  AND U241 ( .A(B[18]), .B(A[2]), .Z(\_2_net_[20] ) );
  AND U242 ( .A(B[17]), .B(A[2]), .Z(\_2_net_[19] ) );
  AND U243 ( .A(B[16]), .B(A[2]), .Z(\_2_net_[18] ) );
  AND U244 ( .A(B[15]), .B(A[2]), .Z(\_2_net_[17] ) );
  AND U245 ( .A(B[14]), .B(A[2]), .Z(\_2_net_[16] ) );
  AND U246 ( .A(B[13]), .B(A[2]), .Z(\_2_net_[15] ) );
  AND U247 ( .A(B[12]), .B(A[2]), .Z(\_2_net_[14] ) );
  AND U248 ( .A(B[11]), .B(A[2]), .Z(\_2_net_[13] ) );
  AND U249 ( .A(B[10]), .B(A[2]), .Z(\_2_net_[12] ) );
  AND U250 ( .A(B[9]), .B(A[2]), .Z(\_2_net_[11] ) );
  AND U251 ( .A(B[8]), .B(A[2]), .Z(\_2_net_[10] ) );
  AND U252 ( .A(B[16]), .B(A[15]), .Z(\_28_net_[31] ) );
  AND U253 ( .A(B[15]), .B(A[15]), .Z(\_28_net_[30] ) );
  AND U254 ( .A(B[14]), .B(A[15]), .Z(\_28_net_[29] ) );
  AND U255 ( .A(B[13]), .B(A[15]), .Z(\_28_net_[28] ) );
  AND U256 ( .A(B[12]), .B(A[15]), .Z(\_28_net_[27] ) );
  AND U257 ( .A(B[11]), .B(A[15]), .Z(\_28_net_[26] ) );
  AND U258 ( .A(B[10]), .B(A[15]), .Z(\_28_net_[25] ) );
  AND U259 ( .A(B[9]), .B(A[15]), .Z(\_28_net_[24] ) );
  AND U260 ( .A(B[8]), .B(A[15]), .Z(\_28_net_[23] ) );
  AND U261 ( .A(B[7]), .B(A[15]), .Z(\_28_net_[22] ) );
  AND U262 ( .A(B[6]), .B(A[15]), .Z(\_28_net_[21] ) );
  AND U263 ( .A(B[5]), .B(A[15]), .Z(\_28_net_[20] ) );
  AND U264 ( .A(B[4]), .B(A[15]), .Z(\_28_net_[19] ) );
  AND U265 ( .A(B[3]), .B(A[15]), .Z(\_28_net_[18] ) );
  AND U266 ( .A(B[2]), .B(A[15]), .Z(\_28_net_[17] ) );
  AND U267 ( .A(B[1]), .B(A[15]), .Z(\_28_net_[16] ) );
  AND U268 ( .A(A[15]), .B(B[0]), .Z(\_28_net_[15] ) );
  AND U269 ( .A(B[17]), .B(A[14]), .Z(\_26_net_[31] ) );
  AND U270 ( .A(B[16]), .B(A[14]), .Z(\_26_net_[30] ) );
  AND U271 ( .A(B[15]), .B(A[14]), .Z(\_26_net_[29] ) );
  AND U272 ( .A(B[14]), .B(A[14]), .Z(\_26_net_[28] ) );
  AND U273 ( .A(B[13]), .B(A[14]), .Z(\_26_net_[27] ) );
  AND U274 ( .A(B[12]), .B(A[14]), .Z(\_26_net_[26] ) );
  AND U275 ( .A(B[11]), .B(A[14]), .Z(\_26_net_[25] ) );
  AND U276 ( .A(B[10]), .B(A[14]), .Z(\_26_net_[24] ) );
  AND U277 ( .A(B[9]), .B(A[14]), .Z(\_26_net_[23] ) );
  AND U278 ( .A(B[8]), .B(A[14]), .Z(\_26_net_[22] ) );
  AND U279 ( .A(B[7]), .B(A[14]), .Z(\_26_net_[21] ) );
  AND U280 ( .A(B[6]), .B(A[14]), .Z(\_26_net_[20] ) );
  AND U281 ( .A(B[5]), .B(A[14]), .Z(\_26_net_[19] ) );
  AND U282 ( .A(B[4]), .B(A[14]), .Z(\_26_net_[18] ) );
  AND U283 ( .A(B[3]), .B(A[14]), .Z(\_26_net_[17] ) );
  AND U284 ( .A(B[2]), .B(A[14]), .Z(\_26_net_[16] ) );
  AND U285 ( .A(B[1]), .B(A[14]), .Z(\_26_net_[15] ) );
  AND U286 ( .A(A[14]), .B(B[0]), .Z(\_26_net_[14] ) );
  AND U287 ( .A(B[18]), .B(A[13]), .Z(\_24_net_[31] ) );
  AND U288 ( .A(B[17]), .B(A[13]), .Z(\_24_net_[30] ) );
  AND U289 ( .A(B[16]), .B(A[13]), .Z(\_24_net_[29] ) );
  AND U290 ( .A(B[15]), .B(A[13]), .Z(\_24_net_[28] ) );
  AND U291 ( .A(B[14]), .B(A[13]), .Z(\_24_net_[27] ) );
  AND U292 ( .A(B[13]), .B(A[13]), .Z(\_24_net_[26] ) );
  AND U293 ( .A(B[12]), .B(A[13]), .Z(\_24_net_[25] ) );
  AND U294 ( .A(B[11]), .B(A[13]), .Z(\_24_net_[24] ) );
  AND U295 ( .A(B[10]), .B(A[13]), .Z(\_24_net_[23] ) );
  AND U296 ( .A(B[9]), .B(A[13]), .Z(\_24_net_[22] ) );
  AND U297 ( .A(B[8]), .B(A[13]), .Z(\_24_net_[21] ) );
  AND U298 ( .A(B[7]), .B(A[13]), .Z(\_24_net_[20] ) );
  AND U299 ( .A(B[6]), .B(A[13]), .Z(\_24_net_[19] ) );
  AND U300 ( .A(B[5]), .B(A[13]), .Z(\_24_net_[18] ) );
  AND U301 ( .A(B[4]), .B(A[13]), .Z(\_24_net_[17] ) );
  AND U302 ( .A(B[3]), .B(A[13]), .Z(\_24_net_[16] ) );
  AND U303 ( .A(B[2]), .B(A[13]), .Z(\_24_net_[15] ) );
  AND U304 ( .A(B[1]), .B(A[13]), .Z(\_24_net_[14] ) );
  AND U305 ( .A(A[13]), .B(B[0]), .Z(\_24_net_[13] ) );
  AND U306 ( .A(B[19]), .B(A[12]), .Z(\_22_net_[31] ) );
  AND U307 ( .A(B[18]), .B(A[12]), .Z(\_22_net_[30] ) );
  AND U308 ( .A(B[17]), .B(A[12]), .Z(\_22_net_[29] ) );
  AND U309 ( .A(B[16]), .B(A[12]), .Z(\_22_net_[28] ) );
  AND U310 ( .A(B[15]), .B(A[12]), .Z(\_22_net_[27] ) );
  AND U311 ( .A(B[14]), .B(A[12]), .Z(\_22_net_[26] ) );
  AND U312 ( .A(B[13]), .B(A[12]), .Z(\_22_net_[25] ) );
  AND U313 ( .A(B[12]), .B(A[12]), .Z(\_22_net_[24] ) );
  AND U314 ( .A(B[11]), .B(A[12]), .Z(\_22_net_[23] ) );
  AND U315 ( .A(B[10]), .B(A[12]), .Z(\_22_net_[22] ) );
  AND U316 ( .A(B[9]), .B(A[12]), .Z(\_22_net_[21] ) );
  AND U317 ( .A(B[8]), .B(A[12]), .Z(\_22_net_[20] ) );
  AND U318 ( .A(B[7]), .B(A[12]), .Z(\_22_net_[19] ) );
  AND U319 ( .A(B[6]), .B(A[12]), .Z(\_22_net_[18] ) );
  AND U320 ( .A(B[5]), .B(A[12]), .Z(\_22_net_[17] ) );
  AND U321 ( .A(B[4]), .B(A[12]), .Z(\_22_net_[16] ) );
  AND U322 ( .A(B[3]), .B(A[12]), .Z(\_22_net_[15] ) );
  AND U323 ( .A(B[2]), .B(A[12]), .Z(\_22_net_[14] ) );
  AND U324 ( .A(B[1]), .B(A[12]), .Z(\_22_net_[13] ) );
  AND U325 ( .A(A[12]), .B(B[0]), .Z(\_22_net_[12] ) );
  AND U326 ( .A(B[20]), .B(A[11]), .Z(\_20_net_[31] ) );
  AND U327 ( .A(B[19]), .B(A[11]), .Z(\_20_net_[30] ) );
  AND U328 ( .A(B[18]), .B(A[11]), .Z(\_20_net_[29] ) );
  AND U329 ( .A(B[17]), .B(A[11]), .Z(\_20_net_[28] ) );
  AND U330 ( .A(B[16]), .B(A[11]), .Z(\_20_net_[27] ) );
  AND U331 ( .A(B[15]), .B(A[11]), .Z(\_20_net_[26] ) );
  AND U332 ( .A(B[14]), .B(A[11]), .Z(\_20_net_[25] ) );
  AND U333 ( .A(B[13]), .B(A[11]), .Z(\_20_net_[24] ) );
  AND U334 ( .A(B[12]), .B(A[11]), .Z(\_20_net_[23] ) );
  AND U335 ( .A(B[11]), .B(A[11]), .Z(\_20_net_[22] ) );
  AND U336 ( .A(B[10]), .B(A[11]), .Z(\_20_net_[21] ) );
  AND U337 ( .A(B[9]), .B(A[11]), .Z(\_20_net_[20] ) );
  AND U338 ( .A(B[8]), .B(A[11]), .Z(\_20_net_[19] ) );
  AND U339 ( .A(B[7]), .B(A[11]), .Z(\_20_net_[18] ) );
  AND U340 ( .A(B[6]), .B(A[11]), .Z(\_20_net_[17] ) );
  AND U341 ( .A(B[5]), .B(A[11]), .Z(\_20_net_[16] ) );
  AND U342 ( .A(B[4]), .B(A[11]), .Z(\_20_net_[15] ) );
  AND U343 ( .A(B[3]), .B(A[11]), .Z(\_20_net_[14] ) );
  AND U344 ( .A(B[2]), .B(A[11]), .Z(\_20_net_[13] ) );
  AND U345 ( .A(B[1]), .B(A[11]), .Z(\_20_net_[12] ) );
  AND U346 ( .A(A[11]), .B(B[0]), .Z(\_20_net_[11] ) );
  AND U347 ( .A(B[21]), .B(A[10]), .Z(\_18_net_[31] ) );
  AND U348 ( .A(B[20]), .B(A[10]), .Z(\_18_net_[30] ) );
  AND U349 ( .A(B[19]), .B(A[10]), .Z(\_18_net_[29] ) );
  AND U350 ( .A(B[18]), .B(A[10]), .Z(\_18_net_[28] ) );
  AND U351 ( .A(B[17]), .B(A[10]), .Z(\_18_net_[27] ) );
  AND U352 ( .A(B[16]), .B(A[10]), .Z(\_18_net_[26] ) );
  AND U353 ( .A(B[15]), .B(A[10]), .Z(\_18_net_[25] ) );
  AND U354 ( .A(B[14]), .B(A[10]), .Z(\_18_net_[24] ) );
  AND U355 ( .A(B[13]), .B(A[10]), .Z(\_18_net_[23] ) );
  AND U356 ( .A(B[12]), .B(A[10]), .Z(\_18_net_[22] ) );
  AND U357 ( .A(B[11]), .B(A[10]), .Z(\_18_net_[21] ) );
  AND U358 ( .A(B[10]), .B(A[10]), .Z(\_18_net_[20] ) );
  AND U359 ( .A(B[9]), .B(A[10]), .Z(\_18_net_[19] ) );
  AND U360 ( .A(B[8]), .B(A[10]), .Z(\_18_net_[18] ) );
  AND U361 ( .A(B[7]), .B(A[10]), .Z(\_18_net_[17] ) );
  AND U362 ( .A(B[6]), .B(A[10]), .Z(\_18_net_[16] ) );
  AND U363 ( .A(B[5]), .B(A[10]), .Z(\_18_net_[15] ) );
  AND U364 ( .A(B[4]), .B(A[10]), .Z(\_18_net_[14] ) );
  AND U365 ( .A(B[3]), .B(A[10]), .Z(\_18_net_[13] ) );
  AND U366 ( .A(B[2]), .B(A[10]), .Z(\_18_net_[12] ) );
  AND U367 ( .A(B[1]), .B(A[10]), .Z(\_18_net_[11] ) );
  AND U368 ( .A(A[10]), .B(B[0]), .Z(\_18_net_[10] ) );
  AND U369 ( .A(B[0]), .B(A[9]), .Z(\_16_net_[9] ) );
  AND U370 ( .A(B[22]), .B(A[9]), .Z(\_16_net_[31] ) );
  AND U371 ( .A(B[21]), .B(A[9]), .Z(\_16_net_[30] ) );
  AND U372 ( .A(B[20]), .B(A[9]), .Z(\_16_net_[29] ) );
  AND U373 ( .A(B[19]), .B(A[9]), .Z(\_16_net_[28] ) );
  AND U374 ( .A(B[18]), .B(A[9]), .Z(\_16_net_[27] ) );
  AND U375 ( .A(B[17]), .B(A[9]), .Z(\_16_net_[26] ) );
  AND U376 ( .A(B[16]), .B(A[9]), .Z(\_16_net_[25] ) );
  AND U377 ( .A(B[15]), .B(A[9]), .Z(\_16_net_[24] ) );
  AND U378 ( .A(B[14]), .B(A[9]), .Z(\_16_net_[23] ) );
  AND U379 ( .A(B[13]), .B(A[9]), .Z(\_16_net_[22] ) );
  AND U380 ( .A(B[12]), .B(A[9]), .Z(\_16_net_[21] ) );
  AND U381 ( .A(B[11]), .B(A[9]), .Z(\_16_net_[20] ) );
  AND U382 ( .A(B[10]), .B(A[9]), .Z(\_16_net_[19] ) );
  AND U383 ( .A(B[9]), .B(A[9]), .Z(\_16_net_[18] ) );
  AND U384 ( .A(B[8]), .B(A[9]), .Z(\_16_net_[17] ) );
  AND U385 ( .A(B[7]), .B(A[9]), .Z(\_16_net_[16] ) );
  AND U386 ( .A(B[6]), .B(A[9]), .Z(\_16_net_[15] ) );
  AND U387 ( .A(B[5]), .B(A[9]), .Z(\_16_net_[14] ) );
  AND U388 ( .A(B[4]), .B(A[9]), .Z(\_16_net_[13] ) );
  AND U389 ( .A(B[3]), .B(A[9]), .Z(\_16_net_[12] ) );
  AND U390 ( .A(B[2]), .B(A[9]), .Z(\_16_net_[11] ) );
  AND U391 ( .A(A[9]), .B(B[1]), .Z(\_16_net_[10] ) );
  AND U392 ( .A(B[1]), .B(A[8]), .Z(\_14_net_[9] ) );
  AND U393 ( .A(B[0]), .B(A[8]), .Z(\_14_net_[8] ) );
  AND U394 ( .A(B[23]), .B(A[8]), .Z(\_14_net_[31] ) );
  AND U395 ( .A(B[22]), .B(A[8]), .Z(\_14_net_[30] ) );
  AND U396 ( .A(B[21]), .B(A[8]), .Z(\_14_net_[29] ) );
  AND U397 ( .A(B[20]), .B(A[8]), .Z(\_14_net_[28] ) );
  AND U398 ( .A(B[19]), .B(A[8]), .Z(\_14_net_[27] ) );
  AND U399 ( .A(B[18]), .B(A[8]), .Z(\_14_net_[26] ) );
  AND U400 ( .A(B[17]), .B(A[8]), .Z(\_14_net_[25] ) );
  AND U401 ( .A(B[16]), .B(A[8]), .Z(\_14_net_[24] ) );
  AND U402 ( .A(B[15]), .B(A[8]), .Z(\_14_net_[23] ) );
  AND U403 ( .A(B[14]), .B(A[8]), .Z(\_14_net_[22] ) );
  AND U404 ( .A(B[13]), .B(A[8]), .Z(\_14_net_[21] ) );
  AND U405 ( .A(B[12]), .B(A[8]), .Z(\_14_net_[20] ) );
  AND U406 ( .A(B[11]), .B(A[8]), .Z(\_14_net_[19] ) );
  AND U407 ( .A(B[10]), .B(A[8]), .Z(\_14_net_[18] ) );
  AND U408 ( .A(B[9]), .B(A[8]), .Z(\_14_net_[17] ) );
  AND U409 ( .A(B[8]), .B(A[8]), .Z(\_14_net_[16] ) );
  AND U410 ( .A(B[7]), .B(A[8]), .Z(\_14_net_[15] ) );
  AND U411 ( .A(B[6]), .B(A[8]), .Z(\_14_net_[14] ) );
  AND U412 ( .A(B[5]), .B(A[8]), .Z(\_14_net_[13] ) );
  AND U413 ( .A(B[4]), .B(A[8]), .Z(\_14_net_[12] ) );
  AND U414 ( .A(B[3]), .B(A[8]), .Z(\_14_net_[11] ) );
  AND U415 ( .A(A[8]), .B(B[2]), .Z(\_14_net_[10] ) );
  AND U416 ( .A(B[2]), .B(A[7]), .Z(\_12_net_[9] ) );
  AND U417 ( .A(B[1]), .B(A[7]), .Z(\_12_net_[8] ) );
  AND U418 ( .A(B[0]), .B(A[7]), .Z(\_12_net_[7] ) );
  AND U419 ( .A(B[24]), .B(A[7]), .Z(\_12_net_[31] ) );
  AND U420 ( .A(B[23]), .B(A[7]), .Z(\_12_net_[30] ) );
  AND U421 ( .A(B[22]), .B(A[7]), .Z(\_12_net_[29] ) );
  AND U422 ( .A(B[21]), .B(A[7]), .Z(\_12_net_[28] ) );
  AND U423 ( .A(B[20]), .B(A[7]), .Z(\_12_net_[27] ) );
  AND U424 ( .A(B[19]), .B(A[7]), .Z(\_12_net_[26] ) );
  AND U425 ( .A(B[18]), .B(A[7]), .Z(\_12_net_[25] ) );
  AND U426 ( .A(B[17]), .B(A[7]), .Z(\_12_net_[24] ) );
  AND U427 ( .A(B[16]), .B(A[7]), .Z(\_12_net_[23] ) );
  AND U428 ( .A(B[15]), .B(A[7]), .Z(\_12_net_[22] ) );
  AND U429 ( .A(B[14]), .B(A[7]), .Z(\_12_net_[21] ) );
  AND U430 ( .A(B[13]), .B(A[7]), .Z(\_12_net_[20] ) );
  AND U431 ( .A(B[12]), .B(A[7]), .Z(\_12_net_[19] ) );
  AND U432 ( .A(B[11]), .B(A[7]), .Z(\_12_net_[18] ) );
  AND U433 ( .A(B[10]), .B(A[7]), .Z(\_12_net_[17] ) );
  AND U434 ( .A(B[9]), .B(A[7]), .Z(\_12_net_[16] ) );
  AND U435 ( .A(B[8]), .B(A[7]), .Z(\_12_net_[15] ) );
  AND U436 ( .A(B[7]), .B(A[7]), .Z(\_12_net_[14] ) );
  AND U437 ( .A(B[6]), .B(A[7]), .Z(\_12_net_[13] ) );
  AND U438 ( .A(B[5]), .B(A[7]), .Z(\_12_net_[12] ) );
  AND U439 ( .A(B[4]), .B(A[7]), .Z(\_12_net_[11] ) );
  AND U440 ( .A(A[7]), .B(B[3]), .Z(\_12_net_[10] ) );
  AND U441 ( .A(B[3]), .B(A[6]), .Z(\_10_net_[9] ) );
  AND U442 ( .A(B[2]), .B(A[6]), .Z(\_10_net_[8] ) );
  AND U443 ( .A(B[1]), .B(A[6]), .Z(\_10_net_[7] ) );
  AND U444 ( .A(B[0]), .B(A[6]), .Z(\_10_net_[6] ) );
  AND U445 ( .A(B[25]), .B(A[6]), .Z(\_10_net_[31] ) );
  AND U446 ( .A(B[24]), .B(A[6]), .Z(\_10_net_[30] ) );
  AND U447 ( .A(B[23]), .B(A[6]), .Z(\_10_net_[29] ) );
  AND U448 ( .A(B[22]), .B(A[6]), .Z(\_10_net_[28] ) );
  AND U449 ( .A(B[21]), .B(A[6]), .Z(\_10_net_[27] ) );
  AND U450 ( .A(B[20]), .B(A[6]), .Z(\_10_net_[26] ) );
  AND U451 ( .A(B[19]), .B(A[6]), .Z(\_10_net_[25] ) );
  AND U452 ( .A(B[18]), .B(A[6]), .Z(\_10_net_[24] ) );
  AND U453 ( .A(B[17]), .B(A[6]), .Z(\_10_net_[23] ) );
  AND U454 ( .A(B[16]), .B(A[6]), .Z(\_10_net_[22] ) );
  AND U455 ( .A(B[15]), .B(A[6]), .Z(\_10_net_[21] ) );
  AND U456 ( .A(B[14]), .B(A[6]), .Z(\_10_net_[20] ) );
  AND U457 ( .A(B[13]), .B(A[6]), .Z(\_10_net_[19] ) );
  AND U458 ( .A(B[12]), .B(A[6]), .Z(\_10_net_[18] ) );
  AND U459 ( .A(B[11]), .B(A[6]), .Z(\_10_net_[17] ) );
  AND U460 ( .A(B[10]), .B(A[6]), .Z(\_10_net_[16] ) );
  AND U461 ( .A(B[9]), .B(A[6]), .Z(\_10_net_[15] ) );
  AND U462 ( .A(B[8]), .B(A[6]), .Z(\_10_net_[14] ) );
  AND U463 ( .A(B[7]), .B(A[6]), .Z(\_10_net_[13] ) );
  AND U464 ( .A(B[6]), .B(A[6]), .Z(\_10_net_[12] ) );
  AND U465 ( .A(B[5]), .B(A[6]), .Z(\_10_net_[11] ) );
  AND U466 ( .A(A[6]), .B(B[4]), .Z(\_10_net_[10] ) );
  AND U467 ( .A(B[8]), .B(A[1]), .Z(\_0_net_[9] ) );
  AND U468 ( .A(B[7]), .B(A[1]), .Z(\_0_net_[8] ) );
  AND U469 ( .A(B[6]), .B(A[1]), .Z(\_0_net_[7] ) );
  AND U470 ( .A(B[5]), .B(A[1]), .Z(\_0_net_[6] ) );
  AND U471 ( .A(B[4]), .B(A[1]), .Z(\_0_net_[5] ) );
  AND U472 ( .A(B[3]), .B(A[1]), .Z(\_0_net_[4] ) );
  AND U473 ( .A(B[2]), .B(A[1]), .Z(\_0_net_[3] ) );
  AND U474 ( .A(B[30]), .B(A[1]), .Z(\_0_net_[31] ) );
  AND U475 ( .A(B[29]), .B(A[1]), .Z(\_0_net_[30] ) );
  AND U476 ( .A(B[1]), .B(A[1]), .Z(\_0_net_[2] ) );
  AND U477 ( .A(B[28]), .B(A[1]), .Z(\_0_net_[29] ) );
  AND U478 ( .A(B[27]), .B(A[1]), .Z(\_0_net_[28] ) );
  AND U479 ( .A(B[26]), .B(A[1]), .Z(\_0_net_[27] ) );
  AND U480 ( .A(B[25]), .B(A[1]), .Z(\_0_net_[26] ) );
  AND U481 ( .A(B[24]), .B(A[1]), .Z(\_0_net_[25] ) );
  AND U482 ( .A(B[23]), .B(A[1]), .Z(\_0_net_[24] ) );
  AND U483 ( .A(B[22]), .B(A[1]), .Z(\_0_net_[23] ) );
  AND U484 ( .A(B[21]), .B(A[1]), .Z(\_0_net_[22] ) );
  AND U485 ( .A(B[20]), .B(A[1]), .Z(\_0_net_[21] ) );
  AND U486 ( .A(B[19]), .B(A[1]), .Z(\_0_net_[20] ) );
  AND U487 ( .A(B[0]), .B(A[1]), .Z(\_0_net_[1] ) );
  AND U488 ( .A(B[18]), .B(A[1]), .Z(\_0_net_[19] ) );
  AND U489 ( .A(B[17]), .B(A[1]), .Z(\_0_net_[18] ) );
  AND U490 ( .A(B[16]), .B(A[1]), .Z(\_0_net_[17] ) );
  AND U491 ( .A(B[15]), .B(A[1]), .Z(\_0_net_[16] ) );
  AND U492 ( .A(B[14]), .B(A[1]), .Z(\_0_net_[15] ) );
  AND U493 ( .A(B[13]), .B(A[1]), .Z(\_0_net_[14] ) );
  AND U494 ( .A(B[12]), .B(A[1]), .Z(\_0_net_[13] ) );
  AND U495 ( .A(B[11]), .B(A[1]), .Z(\_0_net_[12] ) );
  AND U496 ( .A(B[10]), .B(A[1]), .Z(\_0_net_[11] ) );
  AND U497 ( .A(A[1]), .B(B[9]), .Z(\_0_net_[10] ) );
endmodule


module FA_5953 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_5954 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5955 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5956 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5957 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5958 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5959 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5960 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5961 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5962 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5963 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5964 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5965 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5966 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5967 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5968 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5969 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5970 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5971 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5972 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5973 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5974 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5975 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5976 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5977 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5978 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5979 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5980 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5981 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5982 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5983 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_190 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;


  FA_5983 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_5982 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_5981 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_5980 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_5979 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_5978 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_5977 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_5976 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_5975 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_5974 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_5973 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_5972 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_5971 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_5970 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_5969 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_5968 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_5967 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_5966 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_5965 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_5964 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_5963 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_5962 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_5961 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_5960 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_5959 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_5958 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_5957 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_5956 \FAINST[28].FA_  ( .A(1'b0), .B(B[28]), .CI(1'b0), .S(S[28]) );
  FA_5955 \FAINST[29].FA_  ( .A(1'b0), .B(B[29]), .CI(1'b0), .S(S[29]) );
  FA_5954 \FAINST[30].FA_  ( .A(1'b0), .B(B[30]), .CI(1'b0), .S(S[30]) );
  FA_5953 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(1'b0), .S(S[31]) );
endmodule


module FA_5985 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_5986 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_5987 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5988 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5989 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5990 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5991 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5992 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5993 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5994 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5995 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5996 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5997 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5998 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5999 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6000 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6001 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6002 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6003 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6004 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6005 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6006 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6007 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6008 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6009 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6010 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6011 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6012 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6013 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6014 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6015 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_191 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;
  wire   \C[31] ;

  FA_6015 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_6014 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_6013 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_6012 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_6011 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_6010 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_6009 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_6008 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_6007 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_6006 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_6005 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_6004 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_6003 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_6002 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_6001 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_6000 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_5999 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_5998 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_5997 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_5996 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_5995 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_5994 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_5993 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_5992 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_5991 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_5990 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_5989 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_5988 \FAINST[28].FA_  ( .A(1'b0), .B(B[28]), .CI(1'b0), .S(S[28]) );
  FA_5987 \FAINST[29].FA_  ( .A(1'b0), .B(B[29]), .CI(1'b0), .S(S[29]) );
  FA_5986 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(1'b0), .S(S[30]), .CO(
        \C[31] ) );
  FA_5985 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(\C[31] ), .S(S[31]) );
endmodule


module FA_6017 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_6018 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6019 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_6020 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6021 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6022 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6023 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6024 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6025 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6026 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6027 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6028 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6029 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6030 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6031 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6032 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6033 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6034 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6035 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6036 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6037 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6038 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6039 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6040 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6041 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6042 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6043 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6044 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6045 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6046 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6047 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_192 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_6047 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_6046 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_6045 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_6044 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_6043 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_6042 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_6041 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_6040 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_6039 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_6038 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_6037 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_6036 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_6035 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_6034 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_6033 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_6032 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_6031 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_6030 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_6029 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_6028 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_6027 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_6026 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_6025 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_6024 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_6023 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_6022 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_6021 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_6020 \FAINST[28].FA_  ( .A(1'b0), .B(B[28]), .CI(1'b0), .S(S[28]) );
  FA_6019 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(1'b0), .S(S[29]), .CO(
        C[30]) );
  FA_6018 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_6017 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_6049 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_6050 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6051 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6052 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_6053 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6054 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6055 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6056 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6057 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6058 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6059 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6060 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6061 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6062 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6063 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6064 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6065 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6066 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6067 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6068 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6069 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6070 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6071 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6072 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6073 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6074 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6075 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6076 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6077 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6078 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6079 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_193 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_6079 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_6078 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_6077 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_6076 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_6075 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_6074 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_6073 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_6072 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_6071 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_6070 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_6069 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_6068 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_6067 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_6066 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_6065 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_6064 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_6063 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_6062 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_6061 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_6060 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_6059 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_6058 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_6057 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_6056 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_6055 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_6054 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_6053 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_6052 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(1'b0), .S(S[28]), .CO(
        C[29]) );
  FA_6051 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_6050 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_6049 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_6081 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_6082 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6083 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6084 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6085 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_6086 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6087 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6088 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6089 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6090 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6091 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6092 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6093 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6094 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6095 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6096 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6097 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6098 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6099 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6104 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_194 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_6111 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_6110 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_6109 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_6108 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_6107 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_6106 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_6105 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_6104 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_6103 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_6102 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_6101 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_6100 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_6099 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_6098 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_6097 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_6096 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_6095 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_6094 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_6093 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_6092 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_6091 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_6090 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_6089 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_6088 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_6087 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_6086 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_6085 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(1'b0), .S(S[27]), .CO(
        C[28]) );
  FA_6084 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_6083 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_6082 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_6081 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_6113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_6114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_6119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6120 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6136 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_195 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_6143 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_6142 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_6141 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_6140 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_6139 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_6138 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_6137 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_6136 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_6135 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_6134 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_6133 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_6132 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_6131 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_6130 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_6129 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_6128 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_6127 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_6126 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_6125 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_6124 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_6123 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_6122 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_6121 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_6120 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_6119 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_6118 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(1'b0), .S(S[26]), .CO(
        C[27]) );
  FA_6117 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_6116 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_6115 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_6114 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_6113 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_6145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_6146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_6152 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6168 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_196 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_6175 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_6174 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_6173 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_6172 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_6171 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_6170 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_6169 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_6168 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_6167 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_6166 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_6165 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_6164 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_6163 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_6162 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_6161 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_6160 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_6159 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_6158 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_6157 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_6156 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_6155 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_6154 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_6153 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_6152 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_6151 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(1'b0), .S(S[25]), .CO(
        C[26]) );
  FA_6150 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_6149 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_6148 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_6147 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_6146 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_6145 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_6177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_6178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6184 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_6185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6200 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_197 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_6207 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_6206 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_6205 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_6204 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_6203 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_6202 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_6201 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_6200 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_6199 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_6198 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_6197 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_6196 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_6195 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_6194 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_6193 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_6192 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_6191 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_6190 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_6189 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_6188 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_6187 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_6186 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_6185 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_6184 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(1'b0), .S(S[24]), .CO(
        C[25]) );
  FA_6183 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_6182 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_6181 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_6180 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_6179 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_6178 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_6177 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_6209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_6210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6216 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_6218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6232 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_198 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_6239 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_6238 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_6237 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_6236 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_6235 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_6234 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_6233 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_6232 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_6231 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_6230 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_6229 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_6228 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_6227 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_6226 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_6225 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_6224 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_6223 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_6222 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_6221 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_6220 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_6219 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_6218 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_6217 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(1'b0), .S(S[23]), .CO(
        C[24]) );
  FA_6216 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_6215 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_6214 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_6213 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_6212 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_6211 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_6210 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_6209 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_6241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_6242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6248 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_6251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6264 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_199 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_6271 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_6270 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_6269 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_6268 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_6267 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_6266 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_6265 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_6264 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_6263 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_6262 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_6261 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_6260 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_6259 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_6258 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_6257 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_6256 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_6255 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_6254 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_6253 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_6252 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_6251 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_6250 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(1'b0), .S(S[22]), .CO(
        C[23]) );
  FA_6249 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_6248 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_6247 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_6246 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_6245 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_6244 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_6243 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_6242 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_6241 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_6273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_6274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6280 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_6284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6296 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_200 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_6303 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_6302 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_6301 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_6300 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_6299 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_6298 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_6297 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_6296 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_6295 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_6294 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_6293 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_6292 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_6291 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_6290 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_6289 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_6288 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_6287 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_6286 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_6285 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_6284 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_6283 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(1'b0), .S(S[21]), .CO(
        C[22]) );
  FA_6282 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_6281 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_6280 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_6279 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_6278 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_6277 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_6276 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_6275 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_6274 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_6273 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_6305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_6306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6312 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_6317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6328 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_201 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_6335 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_6334 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_6333 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_6332 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_6331 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_6330 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_6329 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_6328 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_6327 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_6326 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_6325 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_6324 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_6323 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_6322 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_6321 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_6320 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_6319 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_6318 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_6317 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_6316 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(1'b0), .S(S[20]), .CO(
        C[21]) );
  FA_6315 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_6314 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_6313 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_6312 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_6311 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_6310 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_6309 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_6308 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_6307 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_6306 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_6305 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_6337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_6338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6344 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_6350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6360 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_202 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_6367 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_6366 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_6365 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_6364 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_6363 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_6362 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_6361 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_6360 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_6359 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_6358 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_6357 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_6356 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_6355 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_6354 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_6353 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_6352 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_6351 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_6350 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_6349 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(1'b0), .S(S[19]), .CO(
        C[20]) );
  FA_6348 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_6347 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_6346 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_6345 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_6344 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_6343 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_6342 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_6341 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_6340 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_6339 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_6338 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_6337 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_6369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_6370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6376 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_6383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6392 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_203 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_6399 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_6398 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_6397 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_6396 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_6395 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_6394 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_6393 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_6392 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_6391 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_6390 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_6389 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_6388 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_6387 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_6386 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_6385 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_6384 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_6383 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_6382 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(1'b0), .S(S[18]), .CO(
        C[19]) );
  FA_6381 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_6380 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_6379 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_6378 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_6377 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_6376 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_6375 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_6374 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_6373 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_6372 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_6371 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_6370 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_6369 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_6401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_6402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6408 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_6416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6424 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_204 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_6431 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_6430 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_6429 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_6428 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_6427 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_6426 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_6425 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_6424 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_6423 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_6422 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_6421 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_6420 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_6419 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_6418 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_6417 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_6416 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_6415 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(1'b0), .S(S[17]), .CO(
        C[18]) );
  FA_6414 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_6413 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_6412 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_6411 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_6410 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_6409 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_6408 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_6407 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_6406 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_6405 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_6404 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_6403 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_6402 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_6401 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_6433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_6434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6440 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_6449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6456 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_205 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_6463 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_6462 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_6461 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_6460 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_6459 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_6458 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_6457 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_6456 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_6455 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_6454 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_6453 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_6452 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_6451 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_6450 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_6449 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_6448 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(1'b0), .S(S[16]), .CO(
        C[17]) );
  FA_6447 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_6446 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_6445 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_6444 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_6443 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_6442 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_6441 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_6440 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_6439 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_6438 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_6437 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_6436 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_6435 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_6434 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_6433 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_6465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_6466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6472 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_6482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6488 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_206 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_6495 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_6494 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_6493 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_6492 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_6491 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_6490 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_6489 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_6488 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_6487 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_6486 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_6485 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_6484 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_6483 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_6482 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_6481 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(1'b0), .S(S[15]), .CO(
        C[16]) );
  FA_6480 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_6479 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_6478 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_6477 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_6476 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_6475 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_6474 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_6473 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_6472 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_6471 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_6470 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_6469 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_6468 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_6467 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_6466 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_6465 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_6497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_6498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6504 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6512 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6513 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6514 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_6515 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6516 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6517 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6518 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6519 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6520 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6521 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6522 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6523 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6524 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6525 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6526 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6527 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_207 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_6527 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_6526 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_6525 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_6524 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_6523 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_6522 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_6521 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_6520 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_6519 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_6518 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_6517 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_6516 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_6515 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_6514 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(1'b0), .S(S[14]), .CO(
        C[15]) );
  FA_6513 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_6512 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_6511 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_6510 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_6509 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_6508 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_6507 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_6506 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_6505 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_6504 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_6503 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_6502 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_6501 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_6500 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_6499 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_6498 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_6497 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_6529 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_6530 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6531 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6532 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6533 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6534 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6535 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6536 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6537 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6538 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6539 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6540 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6541 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6542 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6543 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6544 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6545 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6546 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6547 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_6548 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6549 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6550 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6551 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6552 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6553 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6554 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6555 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6556 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6557 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6558 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6559 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_208 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_6559 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_6558 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_6557 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_6556 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_6555 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_6554 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_6553 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_6552 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_6551 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_6550 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_6549 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_6548 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_6547 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(1'b0), .S(S[13]), .CO(
        C[14]) );
  FA_6546 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_6545 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_6544 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_6543 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_6542 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_6541 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_6540 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_6539 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_6538 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_6537 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_6536 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_6535 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_6534 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_6533 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_6532 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_6531 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_6530 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_6529 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_6561 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_6562 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6563 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6564 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6565 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6566 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6567 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6568 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6569 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6570 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6571 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6572 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6573 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6574 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6575 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6576 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6577 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6578 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6579 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6580 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_6581 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6582 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6583 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6584 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6585 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6586 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6587 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6588 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6589 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6590 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6591 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_209 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_6591 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_6590 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_6589 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_6588 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_6587 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_6586 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_6585 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_6584 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_6583 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_6582 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_6581 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_6580 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(1'b0), .S(S[12]), .CO(
        C[13]) );
  FA_6579 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_6578 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_6577 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_6576 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_6575 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_6574 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_6573 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_6572 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_6571 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_6570 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_6569 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_6568 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_6567 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_6566 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_6565 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_6564 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_6563 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_6562 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_6561 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_6593 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_6594 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6595 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6596 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6597 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6598 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6599 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6600 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6601 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6602 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6603 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6604 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6605 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6606 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6607 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6608 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6609 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6610 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6611 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6612 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6613 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_6614 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6615 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6616 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6617 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6618 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6619 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6620 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6621 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6622 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6623 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_210 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_6623 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_6622 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_6621 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_6620 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_6619 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_6618 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_6617 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_6616 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_6615 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_6614 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_6613 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(1'b0), .S(S[11]), .CO(
        C[12]) );
  FA_6612 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_6611 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_6610 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_6609 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_6608 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_6607 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_6606 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_6605 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_6604 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_6603 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_6602 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_6601 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_6600 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_6599 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_6598 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_6597 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_6596 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_6595 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_6594 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_6593 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_6625 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_6626 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6627 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6628 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6629 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6630 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6631 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6632 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6633 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6634 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6635 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6636 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6637 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6638 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6639 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6640 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6641 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6642 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6643 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6644 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6645 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6646 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_6647 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6648 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6649 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6650 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6651 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6652 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6653 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6654 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6655 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_211 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_6655 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_6654 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_6653 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_6652 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_6651 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_6650 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_6649 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_6648 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_6647 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_6646 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(1'b0), .S(S[10]), .CO(
        C[11]) );
  FA_6645 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_6644 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_6643 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_6642 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_6641 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_6640 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_6639 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_6638 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_6637 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_6636 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_6635 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_6634 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_6633 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_6632 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_6631 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_6630 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_6629 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_6628 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_6627 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_6626 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_6625 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_6657 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_6658 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6659 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6660 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6661 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6662 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6663 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6664 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6665 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6666 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6667 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6668 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6669 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6670 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6671 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6672 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6673 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6674 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6675 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6676 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6677 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6678 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6679 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_6680 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6681 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6682 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6683 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6684 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6685 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6686 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6687 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_212 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_6687 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_6686 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_6685 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_6684 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_6683 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_6682 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_6681 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_6680 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_6679 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(1'b0), .S(S[9]), .CO(C[10]) );
  FA_6678 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_6677 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_6676 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_6675 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_6674 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_6673 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_6672 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_6671 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_6670 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_6669 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_6668 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_6667 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_6666 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_6665 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_6664 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_6663 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_6662 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_6661 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_6660 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_6659 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_6658 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_6657 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_6689 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_6690 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6691 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6692 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6693 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6694 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6695 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6696 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6697 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6698 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6699 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6700 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6701 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6702 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6703 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6704 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6705 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6706 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6707 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6708 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6709 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6710 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6711 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6712 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_6713 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6714 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6715 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6716 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6717 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6718 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6719 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_213 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_6719 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_6718 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_6717 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_6716 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_6715 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_6714 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_6713 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_6712 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(1'b0), .S(S[8]), .CO(C[9])
         );
  FA_6711 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_6710 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_6709 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_6708 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_6707 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_6706 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_6705 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_6704 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_6703 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_6702 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_6701 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_6700 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_6699 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_6698 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_6697 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_6696 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_6695 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_6694 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_6693 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_6692 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_6691 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_6690 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_6689 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_6721 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_6722 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6723 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6724 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6725 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6726 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6727 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6728 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6729 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6730 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6731 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6732 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6733 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6734 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6735 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6736 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6737 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6738 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6739 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6740 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6741 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6742 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6743 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6744 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6745 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_6746 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6747 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6748 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6749 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6750 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6751 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_214 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_6751 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_6750 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_6749 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_6748 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_6747 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_6746 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_6745 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(1'b0), .S(S[7]), .CO(C[8])
         );
  FA_6744 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_6743 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_6742 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_6741 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_6740 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_6739 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_6738 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_6737 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_6736 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_6735 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_6734 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_6733 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_6732 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_6731 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_6730 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_6729 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_6728 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_6727 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_6726 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_6725 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_6724 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_6723 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_6722 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_6721 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_6753 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_6754 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6755 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6756 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6757 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6758 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6759 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6760 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6761 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6762 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6763 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6764 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6765 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6766 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6767 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6768 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6769 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6770 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6771 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6772 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6773 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6774 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6775 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6776 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6777 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6778 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_6779 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6780 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6781 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6782 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6783 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_215 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_6783 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_6782 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_6781 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_6780 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_6779 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_6778 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(1'b0), .S(S[6]), .CO(C[7])
         );
  FA_6777 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_6776 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_6775 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_6774 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_6773 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_6772 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_6771 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_6770 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_6769 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_6768 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_6767 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_6766 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_6765 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_6764 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_6763 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_6762 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_6761 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_6760 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_6759 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_6758 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_6757 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_6756 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_6755 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_6754 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_6753 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_6785 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_6786 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6787 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6788 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6789 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6790 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6791 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6792 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6793 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6794 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6795 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6796 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6797 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6798 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6799 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6800 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6801 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6802 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6803 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6804 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6805 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6806 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6807 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6808 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6809 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6810 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6811 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_6812 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6813 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6814 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6815 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_216 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_6815 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_6814 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_6813 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_6812 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_6811 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(1'b0), .S(S[5]), .CO(C[6])
         );
  FA_6810 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_6809 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_6808 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_6807 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_6806 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_6805 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_6804 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_6803 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_6802 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_6801 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_6800 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_6799 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_6798 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_6797 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_6796 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_6795 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_6794 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_6793 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_6792 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_6791 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_6790 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_6789 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_6788 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_6787 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_6786 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_6785 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_6817 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_6818 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6819 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6820 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6821 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6822 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6823 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6824 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6825 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6826 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6827 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6828 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6829 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6830 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6831 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6832 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6833 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6834 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6835 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6836 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6837 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6838 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6839 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6840 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6841 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6842 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6843 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6844 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_6845 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6846 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6847 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_217 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_6847 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_6846 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_6845 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_6844 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(1'b0), .S(S[4]), .CO(C[5])
         );
  FA_6843 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_6842 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_6841 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_6840 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_6839 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_6838 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_6837 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_6836 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_6835 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_6834 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_6833 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_6832 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_6831 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_6830 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_6829 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_6828 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_6827 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_6826 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_6825 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_6824 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_6823 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_6822 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_6821 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_6820 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_6819 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_6818 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_6817 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_6849 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_6850 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6851 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6852 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6853 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6854 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6855 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6856 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6857 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6858 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6859 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6860 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6861 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6862 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6863 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6864 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6865 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6866 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6867 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6868 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6869 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6870 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6871 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6872 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6873 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6874 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6875 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6876 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6877 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_6878 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6879 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_218 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_6879 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_6878 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_6877 \FAINST[3].FA_  ( .A(A[3]), .B(B[3]), .CI(1'b0), .S(S[3]), .CO(C[4])
         );
  FA_6876 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_6875 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_6874 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_6873 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_6872 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_6871 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_6870 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_6869 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_6868 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_6867 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_6866 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_6865 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_6864 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_6863 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_6862 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_6861 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_6860 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_6859 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_6858 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_6857 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_6856 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_6855 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_6854 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_6853 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_6852 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_6851 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_6850 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_6849 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_6881 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_6882 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6883 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6884 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6885 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6886 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6887 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6888 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6889 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6890 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6891 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6892 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6893 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6894 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6895 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6896 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6897 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6898 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6899 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6900 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6901 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6902 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6903 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6904 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6905 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6906 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6907 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6908 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6909 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6910 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_6911 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_219 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_6911 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_6910 \FAINST[2].FA_  ( .A(A[2]), .B(B[2]), .CI(1'b0), .S(S[2]), .CO(C[3])
         );
  FA_6909 \FAINST[3].FA_  ( .A(A[3]), .B(B[3]), .CI(C[3]), .S(S[3]), .CO(C[4])
         );
  FA_6908 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_6907 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_6906 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_6905 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_6904 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_6903 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_6902 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_6901 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_6900 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_6899 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_6898 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_6897 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_6896 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_6895 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_6894 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_6893 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_6892 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_6891 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_6890 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_6889 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_6888 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_6887 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_6886 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_6885 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_6884 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_6883 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_6882 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_6881 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_6913 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_6914 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_6915 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_6916 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_6917 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_6918 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_6919 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_6920 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_6921 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_6922 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_6923 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_6924 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_6925 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_6926 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_6927 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_6928 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_6929 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_6930 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_6931 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_6932 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_6933 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_6934 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_6935 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_6936 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_6937 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_6938 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_6939 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_6940 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_6941 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_6942 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_6943 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module ADD_N32_220 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;


  FA_6943 \FAINST[1].FA_  ( .A(A[1]), .B(1'b0), .CI(1'b0), .S(S[1]) );
  FA_6942 \FAINST[2].FA_  ( .A(A[2]), .B(1'b0), .CI(1'b0), .S(S[2]) );
  FA_6941 \FAINST[3].FA_  ( .A(A[3]), .B(1'b0), .CI(1'b0), .S(S[3]) );
  FA_6940 \FAINST[4].FA_  ( .A(A[4]), .B(1'b0), .CI(1'b0), .S(S[4]) );
  FA_6939 \FAINST[5].FA_  ( .A(A[5]), .B(1'b0), .CI(1'b0), .S(S[5]) );
  FA_6938 \FAINST[6].FA_  ( .A(A[6]), .B(1'b0), .CI(1'b0), .S(S[6]) );
  FA_6937 \FAINST[7].FA_  ( .A(A[7]), .B(1'b0), .CI(1'b0), .S(S[7]) );
  FA_6936 \FAINST[8].FA_  ( .A(A[8]), .B(1'b0), .CI(1'b0), .S(S[8]) );
  FA_6935 \FAINST[9].FA_  ( .A(A[9]), .B(1'b0), .CI(1'b0), .S(S[9]) );
  FA_6934 \FAINST[10].FA_  ( .A(A[10]), .B(1'b0), .CI(1'b0), .S(S[10]) );
  FA_6933 \FAINST[11].FA_  ( .A(A[11]), .B(1'b0), .CI(1'b0), .S(S[11]) );
  FA_6932 \FAINST[12].FA_  ( .A(A[12]), .B(1'b0), .CI(1'b0), .S(S[12]) );
  FA_6931 \FAINST[13].FA_  ( .A(A[13]), .B(1'b0), .CI(1'b0), .S(S[13]) );
  FA_6930 \FAINST[14].FA_  ( .A(A[14]), .B(1'b0), .CI(1'b0), .S(S[14]) );
  FA_6929 \FAINST[15].FA_  ( .A(A[15]), .B(1'b0), .CI(1'b0), .S(S[15]) );
  FA_6928 \FAINST[16].FA_  ( .A(A[16]), .B(1'b0), .CI(1'b0), .S(S[16]) );
  FA_6927 \FAINST[17].FA_  ( .A(A[17]), .B(1'b0), .CI(1'b0), .S(S[17]) );
  FA_6926 \FAINST[18].FA_  ( .A(A[18]), .B(1'b0), .CI(1'b0), .S(S[18]) );
  FA_6925 \FAINST[19].FA_  ( .A(A[19]), .B(1'b0), .CI(1'b0), .S(S[19]) );
  FA_6924 \FAINST[20].FA_  ( .A(A[20]), .B(1'b0), .CI(1'b0), .S(S[20]) );
  FA_6923 \FAINST[21].FA_  ( .A(A[21]), .B(1'b0), .CI(1'b0), .S(S[21]) );
  FA_6922 \FAINST[22].FA_  ( .A(A[22]), .B(1'b0), .CI(1'b0), .S(S[22]) );
  FA_6921 \FAINST[23].FA_  ( .A(A[23]), .B(1'b0), .CI(1'b0), .S(S[23]) );
  FA_6920 \FAINST[24].FA_  ( .A(A[24]), .B(1'b0), .CI(1'b0), .S(S[24]) );
  FA_6919 \FAINST[25].FA_  ( .A(A[25]), .B(1'b0), .CI(1'b0), .S(S[25]) );
  FA_6918 \FAINST[26].FA_  ( .A(A[26]), .B(1'b0), .CI(1'b0), .S(S[26]) );
  FA_6917 \FAINST[27].FA_  ( .A(A[27]), .B(1'b0), .CI(1'b0), .S(S[27]) );
  FA_6916 \FAINST[28].FA_  ( .A(A[28]), .B(1'b0), .CI(1'b0), .S(S[28]) );
  FA_6915 \FAINST[29].FA_  ( .A(A[29]), .B(1'b0), .CI(1'b0), .S(S[29]) );
  FA_6914 \FAINST[30].FA_  ( .A(A[30]), .B(1'b0), .CI(1'b0), .S(S[30]) );
  FA_6913 \FAINST[31].FA_  ( .A(A[31]), .B(1'b0), .CI(1'b0), .S(S[31]) );
endmodule


module MULT_N32_7 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   \w[31][31] , \w[31][30] , \w[31][29] , \w[31][28] , \w[31][27] ,
         \w[31][26] , \w[31][25] , \w[31][24] , \w[31][23] , \w[31][22] ,
         \w[31][21] , \w[31][20] , \w[31][19] , \w[31][18] , \w[31][17] ,
         \w[31][16] , \w[31][15] , \w[31][14] , \w[31][13] , \w[31][12] ,
         \w[31][11] , \w[31][10] , \w[31][9] , \w[31][8] , \w[31][7] ,
         \w[31][6] , \w[31][5] , \w[31][4] , \w[31][3] , \w[31][2] ,
         \w[31][1] , \w[30][31] , \w[30][30] , \w[30][29] , \w[30][28] ,
         \w[30][27] , \w[30][26] , \w[30][25] , \w[30][24] , \w[30][23] ,
         \w[30][22] , \w[30][21] , \w[30][20] , \w[30][19] , \w[30][18] ,
         \w[30][17] , \w[30][16] , \w[30][15] , \w[30][14] , \w[30][13] ,
         \w[30][12] , \w[30][11] , \w[30][10] , \w[30][9] , \w[30][8] ,
         \w[30][7] , \w[30][6] , \w[30][5] , \w[30][4] , \w[30][3] ,
         \w[30][2] , \w[30][1] , \w[29][31] , \w[29][30] , \w[29][29] ,
         \w[29][28] , \w[29][27] , \w[29][26] , \w[29][25] , \w[29][24] ,
         \w[29][23] , \w[29][22] , \w[29][21] , \w[29][20] , \w[29][19] ,
         \w[29][18] , \w[29][17] , \w[29][16] , \w[29][15] , \w[29][14] ,
         \w[29][13] , \w[29][12] , \w[29][11] , \w[29][10] , \w[29][9] ,
         \w[29][8] , \w[29][7] , \w[29][6] , \w[29][5] , \w[29][4] ,
         \w[29][3] , \w[29][2] , \w[29][1] , \w[28][31] , \w[28][30] ,
         \w[28][29] , \w[28][28] , \w[28][27] , \w[28][26] , \w[28][25] ,
         \w[28][24] , \w[28][23] , \w[28][22] , \w[28][21] , \w[28][20] ,
         \w[28][19] , \w[28][18] , \w[28][17] , \w[28][16] , \w[28][15] ,
         \w[28][14] , \w[28][13] , \w[28][12] , \w[28][11] , \w[28][10] ,
         \w[28][9] , \w[28][8] , \w[28][7] , \w[28][6] , \w[28][5] ,
         \w[28][4] , \w[28][3] , \w[28][2] , \w[28][1] , \w[27][31] ,
         \w[27][30] , \w[27][29] , \w[27][28] , \w[27][27] , \w[27][26] ,
         \w[27][25] , \w[27][24] , \w[27][23] , \w[27][22] , \w[27][21] ,
         \w[27][20] , \w[27][19] , \w[27][18] , \w[27][17] , \w[27][16] ,
         \w[27][15] , \w[27][14] , \w[27][13] , \w[27][12] , \w[27][11] ,
         \w[27][10] , \w[27][9] , \w[27][8] , \w[27][7] , \w[27][6] ,
         \w[27][5] , \w[27][4] , \w[27][3] , \w[27][2] , \w[27][1] ,
         \w[26][31] , \w[26][30] , \w[26][29] , \w[26][28] , \w[26][27] ,
         \w[26][26] , \w[26][25] , \w[26][24] , \w[26][23] , \w[26][22] ,
         \w[26][21] , \w[26][20] , \w[26][19] , \w[26][18] , \w[26][17] ,
         \w[26][16] , \w[26][15] , \w[26][14] , \w[26][13] , \w[26][12] ,
         \w[26][11] , \w[26][10] , \w[26][9] , \w[26][8] , \w[26][7] ,
         \w[26][6] , \w[26][5] , \w[26][4] , \w[26][3] , \w[26][2] ,
         \w[26][1] , \w[25][31] , \w[25][30] , \w[25][29] , \w[25][28] ,
         \w[25][27] , \w[25][26] , \w[25][25] , \w[25][24] , \w[25][23] ,
         \w[25][22] , \w[25][21] , \w[25][20] , \w[25][19] , \w[25][18] ,
         \w[25][17] , \w[25][16] , \w[25][15] , \w[25][14] , \w[25][13] ,
         \w[25][12] , \w[25][11] , \w[25][10] , \w[25][9] , \w[25][8] ,
         \w[25][7] , \w[25][6] , \w[25][5] , \w[25][4] , \w[25][3] ,
         \w[25][2] , \w[25][1] , \w[24][31] , \w[24][30] , \w[24][29] ,
         \w[24][28] , \w[24][27] , \w[24][26] , \w[24][25] , \w[24][24] ,
         \w[24][23] , \w[24][22] , \w[24][21] , \w[24][20] , \w[24][19] ,
         \w[24][18] , \w[24][17] , \w[24][16] , \w[24][15] , \w[24][14] ,
         \w[24][13] , \w[24][12] , \w[24][11] , \w[24][10] , \w[24][9] ,
         \w[24][8] , \w[24][7] , \w[24][6] , \w[24][5] , \w[24][4] ,
         \w[24][3] , \w[24][2] , \w[24][1] , \w[23][31] , \w[23][30] ,
         \w[23][29] , \w[23][28] , \w[23][27] , \w[23][26] , \w[23][25] ,
         \w[23][24] , \w[23][23] , \w[23][22] , \w[23][21] , \w[23][20] ,
         \w[23][19] , \w[23][18] , \w[23][17] , \w[23][16] , \w[23][15] ,
         \w[23][14] , \w[23][13] , \w[23][12] , \w[23][11] , \w[23][10] ,
         \w[23][9] , \w[23][8] , \w[23][7] , \w[23][6] , \w[23][5] ,
         \w[23][4] , \w[23][3] , \w[23][2] , \w[23][1] , \w[22][31] ,
         \w[22][30] , \w[22][29] , \w[22][28] , \w[22][27] , \w[22][26] ,
         \w[22][25] , \w[22][24] , \w[22][23] , \w[22][22] , \w[22][21] ,
         \w[22][20] , \w[22][19] , \w[22][18] , \w[22][17] , \w[22][16] ,
         \w[22][15] , \w[22][14] , \w[22][13] , \w[22][12] , \w[22][11] ,
         \w[22][10] , \w[22][9] , \w[22][8] , \w[22][7] , \w[22][6] ,
         \w[22][5] , \w[22][4] , \w[22][3] , \w[22][2] , \w[22][1] ,
         \w[21][31] , \w[21][30] , \w[21][29] , \w[21][28] , \w[21][27] ,
         \w[21][26] , \w[21][25] , \w[21][24] , \w[21][23] , \w[21][22] ,
         \w[21][21] , \w[21][20] , \w[21][19] , \w[21][18] , \w[21][17] ,
         \w[21][16] , \w[21][15] , \w[21][14] , \w[21][13] , \w[21][12] ,
         \w[21][11] , \w[21][10] , \w[21][9] , \w[21][8] , \w[21][7] ,
         \w[21][6] , \w[21][5] , \w[21][4] , \w[21][3] , \w[21][2] ,
         \w[21][1] , \w[20][31] , \w[20][30] , \w[20][29] , \w[20][28] ,
         \w[20][27] , \w[20][26] , \w[20][25] , \w[20][24] , \w[20][23] ,
         \w[20][22] , \w[20][21] , \w[20][20] , \w[20][19] , \w[20][18] ,
         \w[20][17] , \w[20][16] , \w[20][15] , \w[20][14] , \w[20][13] ,
         \w[20][12] , \w[20][11] , \w[20][10] , \w[20][9] , \w[20][8] ,
         \w[20][7] , \w[20][6] , \w[20][5] , \w[20][4] , \w[20][3] ,
         \w[20][2] , \w[20][1] , \w[19][31] , \w[19][30] , \w[19][29] ,
         \w[19][28] , \w[19][27] , \w[19][26] , \w[19][25] , \w[19][24] ,
         \w[19][23] , \w[19][22] , \w[19][21] , \w[19][20] , \w[19][19] ,
         \w[19][18] , \w[19][17] , \w[19][16] , \w[19][15] , \w[19][14] ,
         \w[19][13] , \w[19][12] , \w[19][11] , \w[19][10] , \w[19][9] ,
         \w[19][8] , \w[19][7] , \w[19][6] , \w[19][5] , \w[19][4] ,
         \w[19][3] , \w[19][2] , \w[19][1] , \w[18][31] , \w[18][30] ,
         \w[18][29] , \w[18][28] , \w[18][27] , \w[18][26] , \w[18][25] ,
         \w[18][24] , \w[18][23] , \w[18][22] , \w[18][21] , \w[18][20] ,
         \w[18][19] , \w[18][18] , \w[18][17] , \w[18][16] , \w[18][15] ,
         \w[18][14] , \w[18][13] , \w[18][12] , \w[18][11] , \w[18][10] ,
         \w[18][9] , \w[18][8] , \w[18][7] , \w[18][6] , \w[18][5] ,
         \w[18][4] , \w[18][3] , \w[18][2] , \w[18][1] , \w[17][31] ,
         \w[17][30] , \w[17][29] , \w[17][28] , \w[17][27] , \w[17][26] ,
         \w[17][25] , \w[17][24] , \w[17][23] , \w[17][22] , \w[17][21] ,
         \w[17][20] , \w[17][19] , \w[17][18] , \w[17][17] , \w[17][16] ,
         \w[17][15] , \w[17][14] , \w[17][13] , \w[17][12] , \w[17][11] ,
         \w[17][10] , \w[17][9] , \w[17][8] , \w[17][7] , \w[17][6] ,
         \w[17][5] , \w[17][4] , \w[17][3] , \w[17][2] , \w[17][1] ,
         \w[16][31] , \w[16][30] , \w[16][29] , \w[16][28] , \w[16][27] ,
         \w[16][26] , \w[16][25] , \w[16][24] , \w[16][23] , \w[16][22] ,
         \w[16][21] , \w[16][20] , \w[16][19] , \w[16][18] , \w[16][17] ,
         \w[16][16] , \w[16][15] , \w[16][14] , \w[16][13] , \w[16][12] ,
         \w[16][11] , \w[16][10] , \w[16][9] , \w[16][8] , \w[16][7] ,
         \w[16][6] , \w[16][5] , \w[16][4] , \w[16][3] , \w[16][2] ,
         \w[16][1] , \w[15][31] , \w[15][30] , \w[15][29] , \w[15][28] ,
         \w[15][27] , \w[15][26] , \w[15][25] , \w[15][24] , \w[15][23] ,
         \w[15][22] , \w[15][21] , \w[15][20] , \w[15][19] , \w[15][18] ,
         \w[15][17] , \w[15][16] , \w[15][15] , \w[15][14] , \w[15][13] ,
         \w[15][12] , \w[15][11] , \w[15][10] , \w[15][9] , \w[15][8] ,
         \w[15][7] , \w[15][6] , \w[15][5] , \w[15][4] , \w[15][3] ,
         \w[15][2] , \w[15][1] , \w[14][31] , \w[14][30] , \w[14][29] ,
         \w[14][28] , \w[14][27] , \w[14][26] , \w[14][25] , \w[14][24] ,
         \w[14][23] , \w[14][22] , \w[14][21] , \w[14][20] , \w[14][19] ,
         \w[14][18] , \w[14][17] , \w[14][16] , \w[14][15] , \w[14][14] ,
         \w[14][13] , \w[14][12] , \w[14][11] , \w[14][10] , \w[14][9] ,
         \w[14][8] , \w[14][7] , \w[14][6] , \w[14][5] , \w[14][4] ,
         \w[14][3] , \w[14][2] , \w[14][1] , \w[13][31] , \w[13][30] ,
         \w[13][29] , \w[13][28] , \w[13][27] , \w[13][26] , \w[13][25] ,
         \w[13][24] , \w[13][23] , \w[13][22] , \w[13][21] , \w[13][20] ,
         \w[13][19] , \w[13][18] , \w[13][17] , \w[13][16] , \w[13][15] ,
         \w[13][14] , \w[13][13] , \w[13][12] , \w[13][11] , \w[13][10] ,
         \w[13][9] , \w[13][8] , \w[13][7] , \w[13][6] , \w[13][5] ,
         \w[13][4] , \w[13][3] , \w[13][2] , \w[13][1] , \w[12][31] ,
         \w[12][30] , \w[12][29] , \w[12][28] , \w[12][27] , \w[12][26] ,
         \w[12][25] , \w[12][24] , \w[12][23] , \w[12][22] , \w[12][21] ,
         \w[12][20] , \w[12][19] , \w[12][18] , \w[12][17] , \w[12][16] ,
         \w[12][15] , \w[12][14] , \w[12][13] , \w[12][12] , \w[12][11] ,
         \w[12][10] , \w[12][9] , \w[12][8] , \w[12][7] , \w[12][6] ,
         \w[12][5] , \w[12][4] , \w[12][3] , \w[12][2] , \w[12][1] ,
         \w[11][31] , \w[11][30] , \w[11][29] , \w[11][28] , \w[11][27] ,
         \w[11][26] , \w[11][25] , \w[11][24] , \w[11][23] , \w[11][22] ,
         \w[11][21] , \w[11][20] , \w[11][19] , \w[11][18] , \w[11][17] ,
         \w[11][16] , \w[11][15] , \w[11][14] , \w[11][13] , \w[11][12] ,
         \w[11][11] , \w[11][10] , \w[11][9] , \w[11][8] , \w[11][7] ,
         \w[11][6] , \w[11][5] , \w[11][4] , \w[11][3] , \w[11][2] ,
         \w[11][1] , \w[10][31] , \w[10][30] , \w[10][29] , \w[10][28] ,
         \w[10][27] , \w[10][26] , \w[10][25] , \w[10][24] , \w[10][23] ,
         \w[10][22] , \w[10][21] , \w[10][20] , \w[10][19] , \w[10][18] ,
         \w[10][17] , \w[10][16] , \w[10][15] , \w[10][14] , \w[10][13] ,
         \w[10][12] , \w[10][11] , \w[10][10] , \w[10][9] , \w[10][8] ,
         \w[10][7] , \w[10][6] , \w[10][5] , \w[10][4] , \w[10][3] ,
         \w[10][2] , \w[10][1] , \w[9][31] , \w[9][30] , \w[9][29] ,
         \w[9][28] , \w[9][27] , \w[9][26] , \w[9][25] , \w[9][24] ,
         \w[9][23] , \w[9][22] , \w[9][21] , \w[9][20] , \w[9][19] ,
         \w[9][18] , \w[9][17] , \w[9][16] , \w[9][15] , \w[9][14] ,
         \w[9][13] , \w[9][12] , \w[9][11] , \w[9][10] , \w[9][9] , \w[9][8] ,
         \w[9][7] , \w[9][6] , \w[9][5] , \w[9][4] , \w[9][3] , \w[9][2] ,
         \w[9][1] , \w[8][31] , \w[8][30] , \w[8][29] , \w[8][28] , \w[8][27] ,
         \w[8][26] , \w[8][25] , \w[8][24] , \w[8][23] , \w[8][22] ,
         \w[8][21] , \w[8][20] , \w[8][19] , \w[8][18] , \w[8][17] ,
         \w[8][16] , \w[8][15] , \w[8][14] , \w[8][13] , \w[8][12] ,
         \w[8][11] , \w[8][10] , \w[8][9] , \w[8][8] , \w[8][7] , \w[8][6] ,
         \w[8][5] , \w[8][4] , \w[8][3] , \w[8][2] , \w[8][1] , \w[7][31] ,
         \w[7][30] , \w[7][29] , \w[7][28] , \w[7][27] , \w[7][26] ,
         \w[7][25] , \w[7][24] , \w[7][23] , \w[7][22] , \w[7][21] ,
         \w[7][20] , \w[7][19] , \w[7][18] , \w[7][17] , \w[7][16] ,
         \w[7][15] , \w[7][14] , \w[7][13] , \w[7][12] , \w[7][11] ,
         \w[7][10] , \w[7][9] , \w[7][8] , \w[7][7] , \w[7][6] , \w[7][5] ,
         \w[7][4] , \w[7][3] , \w[7][2] , \w[7][1] , \w[6][31] , \w[6][30] ,
         \w[6][29] , \w[6][28] , \w[6][27] , \w[6][26] , \w[6][25] ,
         \w[6][24] , \w[6][23] , \w[6][22] , \w[6][21] , \w[6][20] ,
         \w[6][19] , \w[6][18] , \w[6][17] , \w[6][16] , \w[6][15] ,
         \w[6][14] , \w[6][13] , \w[6][12] , \w[6][11] , \w[6][10] , \w[6][9] ,
         \w[6][8] , \w[6][7] , \w[6][6] , \w[6][5] , \w[6][4] , \w[6][3] ,
         \w[6][2] , \w[6][1] , \w[5][31] , \w[5][30] , \w[5][29] , \w[5][28] ,
         \w[5][27] , \w[5][26] , \w[5][25] , \w[5][24] , \w[5][23] ,
         \w[5][22] , \w[5][21] , \w[5][20] , \w[5][19] , \w[5][18] ,
         \w[5][17] , \w[5][16] , \w[5][15] , \w[5][14] , \w[5][13] ,
         \w[5][12] , \w[5][11] , \w[5][10] , \w[5][9] , \w[5][8] , \w[5][7] ,
         \w[5][6] , \w[5][5] , \w[5][4] , \w[5][3] , \w[5][2] , \w[5][1] ,
         \w[4][31] , \w[4][30] , \w[4][29] , \w[4][28] , \w[4][27] ,
         \w[4][26] , \w[4][25] , \w[4][24] , \w[4][23] , \w[4][22] ,
         \w[4][21] , \w[4][20] , \w[4][19] , \w[4][18] , \w[4][17] ,
         \w[4][16] , \w[4][15] , \w[4][14] , \w[4][13] , \w[4][12] ,
         \w[4][11] , \w[4][10] , \w[4][9] , \w[4][8] , \w[4][7] , \w[4][6] ,
         \w[4][5] , \w[4][4] , \w[4][3] , \w[4][2] , \w[4][1] , \w[3][31] ,
         \w[3][30] , \w[3][29] , \w[3][28] , \w[3][27] , \w[3][26] ,
         \w[3][25] , \w[3][24] , \w[3][23] , \w[3][22] , \w[3][21] ,
         \w[3][20] , \w[3][19] , \w[3][18] , \w[3][17] , \w[3][16] ,
         \w[3][15] , \w[3][14] , \w[3][13] , \w[3][12] , \w[3][11] ,
         \w[3][10] , \w[3][9] , \w[3][8] , \w[3][7] , \w[3][6] , \w[3][5] ,
         \w[3][4] , \w[3][3] , \w[3][2] , \w[3][1] , \w[2][31] , \w[2][30] ,
         \w[2][29] , \w[2][28] , \w[2][27] , \w[2][26] , \w[2][25] ,
         \w[2][24] , \w[2][23] , \w[2][22] , \w[2][21] , \w[2][20] ,
         \w[2][19] , \w[2][18] , \w[2][17] , \w[2][16] , \w[2][15] ,
         \w[2][14] , \w[2][13] , \w[2][12] , \w[2][11] , \w[2][10] , \w[2][9] ,
         \w[2][8] , \w[2][7] , \w[2][6] , \w[2][5] , \w[2][4] , \w[2][3] ,
         \w[2][2] , \w[2][1] , \_0_net_[31] , \_0_net_[30] , \_0_net_[29] ,
         \_0_net_[28] , \_0_net_[27] , \_0_net_[26] , \_0_net_[25] ,
         \_0_net_[24] , \_0_net_[23] , \_0_net_[22] , \_0_net_[21] ,
         \_0_net_[20] , \_0_net_[19] , \_0_net_[18] , \_0_net_[17] ,
         \_0_net_[16] , \_0_net_[15] , \_0_net_[14] , \_0_net_[13] ,
         \_0_net_[12] , \_0_net_[11] , \_0_net_[10] , \_0_net_[9] ,
         \_0_net_[8] , \_0_net_[7] , \_0_net_[6] , \_0_net_[5] , \_0_net_[4] ,
         \_0_net_[3] , \_0_net_[2] , \_0_net_[1] , \_2_net_[31] ,
         \_2_net_[30] , \_2_net_[29] , \_2_net_[28] , \_2_net_[27] ,
         \_2_net_[26] , \_2_net_[25] , \_2_net_[24] , \_2_net_[23] ,
         \_2_net_[22] , \_2_net_[21] , \_2_net_[20] , \_2_net_[19] ,
         \_2_net_[18] , \_2_net_[17] , \_2_net_[16] , \_2_net_[15] ,
         \_2_net_[14] , \_2_net_[13] , \_2_net_[12] , \_2_net_[11] ,
         \_2_net_[10] , \_2_net_[9] , \_2_net_[8] , \_2_net_[7] , \_2_net_[6] ,
         \_2_net_[5] , \_2_net_[4] , \_2_net_[3] , \_2_net_[2] , \_4_net_[31] ,
         \_4_net_[30] , \_4_net_[29] , \_4_net_[28] , \_4_net_[27] ,
         \_4_net_[26] , \_4_net_[25] , \_4_net_[24] , \_4_net_[23] ,
         \_4_net_[22] , \_4_net_[21] , \_4_net_[20] , \_4_net_[19] ,
         \_4_net_[18] , \_4_net_[17] , \_4_net_[16] , \_4_net_[15] ,
         \_4_net_[14] , \_4_net_[13] , \_4_net_[12] , \_4_net_[11] ,
         \_4_net_[10] , \_4_net_[9] , \_4_net_[8] , \_4_net_[7] , \_4_net_[6] ,
         \_4_net_[5] , \_4_net_[4] , \_4_net_[3] , \_6_net_[31] ,
         \_6_net_[30] , \_6_net_[29] , \_6_net_[28] , \_6_net_[27] ,
         \_6_net_[26] , \_6_net_[25] , \_6_net_[24] , \_6_net_[23] ,
         \_6_net_[22] , \_6_net_[21] , \_6_net_[20] , \_6_net_[19] ,
         \_6_net_[18] , \_6_net_[17] , \_6_net_[16] , \_6_net_[15] ,
         \_6_net_[14] , \_6_net_[13] , \_6_net_[12] , \_6_net_[11] ,
         \_6_net_[10] , \_6_net_[9] , \_6_net_[8] , \_6_net_[7] , \_6_net_[6] ,
         \_6_net_[5] , \_6_net_[4] , \_8_net_[31] , \_8_net_[30] ,
         \_8_net_[29] , \_8_net_[28] , \_8_net_[27] , \_8_net_[26] ,
         \_8_net_[25] , \_8_net_[24] , \_8_net_[23] , \_8_net_[22] ,
         \_8_net_[21] , \_8_net_[20] , \_8_net_[19] , \_8_net_[18] ,
         \_8_net_[17] , \_8_net_[16] , \_8_net_[15] , \_8_net_[14] ,
         \_8_net_[13] , \_8_net_[12] , \_8_net_[11] , \_8_net_[10] ,
         \_8_net_[9] , \_8_net_[8] , \_8_net_[7] , \_8_net_[6] , \_8_net_[5] ,
         \_10_net_[31] , \_10_net_[30] , \_10_net_[29] , \_10_net_[28] ,
         \_10_net_[27] , \_10_net_[26] , \_10_net_[25] , \_10_net_[24] ,
         \_10_net_[23] , \_10_net_[22] , \_10_net_[21] , \_10_net_[20] ,
         \_10_net_[19] , \_10_net_[18] , \_10_net_[17] , \_10_net_[16] ,
         \_10_net_[15] , \_10_net_[14] , \_10_net_[13] , \_10_net_[12] ,
         \_10_net_[11] , \_10_net_[10] , \_10_net_[9] , \_10_net_[8] ,
         \_10_net_[7] , \_10_net_[6] , \_12_net_[31] , \_12_net_[30] ,
         \_12_net_[29] , \_12_net_[28] , \_12_net_[27] , \_12_net_[26] ,
         \_12_net_[25] , \_12_net_[24] , \_12_net_[23] , \_12_net_[22] ,
         \_12_net_[21] , \_12_net_[20] , \_12_net_[19] , \_12_net_[18] ,
         \_12_net_[17] , \_12_net_[16] , \_12_net_[15] , \_12_net_[14] ,
         \_12_net_[13] , \_12_net_[12] , \_12_net_[11] , \_12_net_[10] ,
         \_12_net_[9] , \_12_net_[8] , \_12_net_[7] , \_14_net_[31] ,
         \_14_net_[30] , \_14_net_[29] , \_14_net_[28] , \_14_net_[27] ,
         \_14_net_[26] , \_14_net_[25] , \_14_net_[24] , \_14_net_[23] ,
         \_14_net_[22] , \_14_net_[21] , \_14_net_[20] , \_14_net_[19] ,
         \_14_net_[18] , \_14_net_[17] , \_14_net_[16] , \_14_net_[15] ,
         \_14_net_[14] , \_14_net_[13] , \_14_net_[12] , \_14_net_[11] ,
         \_14_net_[10] , \_14_net_[9] , \_14_net_[8] , \_16_net_[31] ,
         \_16_net_[30] , \_16_net_[29] , \_16_net_[28] , \_16_net_[27] ,
         \_16_net_[26] , \_16_net_[25] , \_16_net_[24] , \_16_net_[23] ,
         \_16_net_[22] , \_16_net_[21] , \_16_net_[20] , \_16_net_[19] ,
         \_16_net_[18] , \_16_net_[17] , \_16_net_[16] , \_16_net_[15] ,
         \_16_net_[14] , \_16_net_[13] , \_16_net_[12] , \_16_net_[11] ,
         \_16_net_[10] , \_16_net_[9] , \_18_net_[31] , \_18_net_[30] ,
         \_18_net_[29] , \_18_net_[28] , \_18_net_[27] , \_18_net_[26] ,
         \_18_net_[25] , \_18_net_[24] , \_18_net_[23] , \_18_net_[22] ,
         \_18_net_[21] , \_18_net_[20] , \_18_net_[19] , \_18_net_[18] ,
         \_18_net_[17] , \_18_net_[16] , \_18_net_[15] , \_18_net_[14] ,
         \_18_net_[13] , \_18_net_[12] , \_18_net_[11] , \_18_net_[10] ,
         \_20_net_[31] , \_20_net_[30] , \_20_net_[29] , \_20_net_[28] ,
         \_20_net_[27] , \_20_net_[26] , \_20_net_[25] , \_20_net_[24] ,
         \_20_net_[23] , \_20_net_[22] , \_20_net_[21] , \_20_net_[20] ,
         \_20_net_[19] , \_20_net_[18] , \_20_net_[17] , \_20_net_[16] ,
         \_20_net_[15] , \_20_net_[14] , \_20_net_[13] , \_20_net_[12] ,
         \_20_net_[11] , \_22_net_[31] , \_22_net_[30] , \_22_net_[29] ,
         \_22_net_[28] , \_22_net_[27] , \_22_net_[26] , \_22_net_[25] ,
         \_22_net_[24] , \_22_net_[23] , \_22_net_[22] , \_22_net_[21] ,
         \_22_net_[20] , \_22_net_[19] , \_22_net_[18] , \_22_net_[17] ,
         \_22_net_[16] , \_22_net_[15] , \_22_net_[14] , \_22_net_[13] ,
         \_22_net_[12] , \_24_net_[31] , \_24_net_[30] , \_24_net_[29] ,
         \_24_net_[28] , \_24_net_[27] , \_24_net_[26] , \_24_net_[25] ,
         \_24_net_[24] , \_24_net_[23] , \_24_net_[22] , \_24_net_[21] ,
         \_24_net_[20] , \_24_net_[19] , \_24_net_[18] , \_24_net_[17] ,
         \_24_net_[16] , \_24_net_[15] , \_24_net_[14] , \_24_net_[13] ,
         \_26_net_[31] , \_26_net_[30] , \_26_net_[29] , \_26_net_[28] ,
         \_26_net_[27] , \_26_net_[26] , \_26_net_[25] , \_26_net_[24] ,
         \_26_net_[23] , \_26_net_[22] , \_26_net_[21] , \_26_net_[20] ,
         \_26_net_[19] , \_26_net_[18] , \_26_net_[17] , \_26_net_[16] ,
         \_26_net_[15] , \_26_net_[14] , \_28_net_[31] , \_28_net_[30] ,
         \_28_net_[29] , \_28_net_[28] , \_28_net_[27] , \_28_net_[26] ,
         \_28_net_[25] , \_28_net_[24] , \_28_net_[23] , \_28_net_[22] ,
         \_28_net_[21] , \_28_net_[20] , \_28_net_[19] , \_28_net_[18] ,
         \_28_net_[17] , \_28_net_[16] , \_28_net_[15] , \_30_net_[31] ,
         \_30_net_[30] , \_30_net_[29] , \_30_net_[28] , \_30_net_[27] ,
         \_30_net_[26] , \_30_net_[25] , \_30_net_[24] , \_30_net_[23] ,
         \_30_net_[22] , \_30_net_[21] , \_30_net_[20] , \_30_net_[19] ,
         \_30_net_[18] , \_30_net_[17] , \_30_net_[16] , \_32_net_[31] ,
         \_32_net_[30] , \_32_net_[29] , \_32_net_[28] , \_32_net_[27] ,
         \_32_net_[26] , \_32_net_[25] , \_32_net_[24] , \_32_net_[23] ,
         \_32_net_[22] , \_32_net_[21] , \_32_net_[20] , \_32_net_[19] ,
         \_32_net_[18] , \_32_net_[17] , \_34_net_[31] , \_34_net_[30] ,
         \_34_net_[29] , \_34_net_[28] , \_34_net_[27] , \_34_net_[26] ,
         \_34_net_[25] , \_34_net_[24] , \_34_net_[23] , \_34_net_[22] ,
         \_34_net_[21] , \_34_net_[20] , \_34_net_[19] , \_34_net_[18] ,
         \_36_net_[31] , \_36_net_[30] , \_36_net_[29] , \_36_net_[28] ,
         \_36_net_[27] , \_36_net_[26] , \_36_net_[25] , \_36_net_[24] ,
         \_36_net_[23] , \_36_net_[22] , \_36_net_[21] , \_36_net_[20] ,
         \_36_net_[19] , \_38_net_[31] , \_38_net_[30] , \_38_net_[29] ,
         \_38_net_[28] , \_38_net_[27] , \_38_net_[26] , \_38_net_[25] ,
         \_38_net_[24] , \_38_net_[23] , \_38_net_[22] , \_38_net_[21] ,
         \_38_net_[20] , \_40_net_[31] , \_40_net_[30] , \_40_net_[29] ,
         \_40_net_[28] , \_40_net_[27] , \_40_net_[26] , \_40_net_[25] ,
         \_40_net_[24] , \_40_net_[23] , \_40_net_[22] , \_40_net_[21] ,
         \_42_net_[31] , \_42_net_[30] , \_42_net_[29] , \_42_net_[28] ,
         \_42_net_[27] , \_42_net_[26] , \_42_net_[25] , \_42_net_[24] ,
         \_42_net_[23] , \_42_net_[22] , \_44_net_[31] , \_44_net_[30] ,
         \_44_net_[29] , \_44_net_[28] , \_44_net_[27] , \_44_net_[26] ,
         \_44_net_[25] , \_44_net_[24] , \_44_net_[23] , \_46_net_[31] ,
         \_46_net_[30] , \_46_net_[29] , \_46_net_[28] , \_46_net_[27] ,
         \_46_net_[26] , \_46_net_[25] , \_46_net_[24] , \_48_net_[31] ,
         \_48_net_[30] , \_48_net_[29] , \_48_net_[28] , \_48_net_[27] ,
         \_48_net_[26] , \_48_net_[25] , \_50_net_[31] , \_50_net_[30] ,
         \_50_net_[29] , \_50_net_[28] , \_50_net_[27] , \_50_net_[26] ,
         \_52_net_[31] , \_52_net_[30] , \_52_net_[29] , \_52_net_[28] ,
         \_52_net_[27] , \_54_net_[31] , \_54_net_[30] , \_54_net_[29] ,
         \_54_net_[28] , \_56_net_[31] , \_56_net_[30] , \_56_net_[29] ,
         \_58_net_[31] , \_58_net_[30] , \_60_net_[31] ;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30;

  ADD_N32_220 \FAINST[1].ADD_  ( .A({\_0_net_[31] , \_0_net_[30] , 
        \_0_net_[29] , \_0_net_[28] , \_0_net_[27] , \_0_net_[26] , 
        \_0_net_[25] , \_0_net_[24] , \_0_net_[23] , \_0_net_[22] , 
        \_0_net_[21] , \_0_net_[20] , \_0_net_[19] , \_0_net_[18] , 
        \_0_net_[17] , \_0_net_[16] , \_0_net_[15] , \_0_net_[14] , 
        \_0_net_[13] , \_0_net_[12] , \_0_net_[11] , \_0_net_[10] , 
        \_0_net_[9] , \_0_net_[8] , \_0_net_[7] , \_0_net_[6] , \_0_net_[5] , 
        \_0_net_[4] , \_0_net_[3] , \_0_net_[2] , \_0_net_[1] , 1'b0}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .S({
        \w[2][31] , \w[2][30] , \w[2][29] , \w[2][28] , \w[2][27] , \w[2][26] , 
        \w[2][25] , \w[2][24] , \w[2][23] , \w[2][22] , \w[2][21] , \w[2][20] , 
        \w[2][19] , \w[2][18] , \w[2][17] , \w[2][16] , \w[2][15] , \w[2][14] , 
        \w[2][13] , \w[2][12] , \w[2][11] , \w[2][10] , \w[2][9] , \w[2][8] , 
        \w[2][7] , \w[2][6] , \w[2][5] , \w[2][4] , \w[2][3] , \w[2][2] , 
        \w[2][1] , SYNOPSYS_UNCONNECTED__0}) );
  ADD_N32_219 \FAINST[2].ADD_  ( .A({\_2_net_[31] , \_2_net_[30] , 
        \_2_net_[29] , \_2_net_[28] , \_2_net_[27] , \_2_net_[26] , 
        \_2_net_[25] , \_2_net_[24] , \_2_net_[23] , \_2_net_[22] , 
        \_2_net_[21] , \_2_net_[20] , \_2_net_[19] , \_2_net_[18] , 
        \_2_net_[17] , \_2_net_[16] , \_2_net_[15] , \_2_net_[14] , 
        \_2_net_[13] , \_2_net_[12] , \_2_net_[11] , \_2_net_[10] , 
        \_2_net_[9] , \_2_net_[8] , \_2_net_[7] , \_2_net_[6] , \_2_net_[5] , 
        \_2_net_[4] , \_2_net_[3] , \_2_net_[2] , 1'b0, 1'b0}), .B({\w[2][31] , 
        \w[2][30] , \w[2][29] , \w[2][28] , \w[2][27] , \w[2][26] , \w[2][25] , 
        \w[2][24] , \w[2][23] , \w[2][22] , \w[2][21] , \w[2][20] , \w[2][19] , 
        \w[2][18] , \w[2][17] , \w[2][16] , \w[2][15] , \w[2][14] , \w[2][13] , 
        \w[2][12] , \w[2][11] , \w[2][10] , \w[2][9] , \w[2][8] , \w[2][7] , 
        \w[2][6] , \w[2][5] , \w[2][4] , \w[2][3] , \w[2][2] , \w[2][1] , 1'b0}), .CI(1'b0), .S({\w[3][31] , \w[3][30] , \w[3][29] , \w[3][28] , \w[3][27] , 
        \w[3][26] , \w[3][25] , \w[3][24] , \w[3][23] , \w[3][22] , \w[3][21] , 
        \w[3][20] , \w[3][19] , \w[3][18] , \w[3][17] , \w[3][16] , \w[3][15] , 
        \w[3][14] , \w[3][13] , \w[3][12] , \w[3][11] , \w[3][10] , \w[3][9] , 
        \w[3][8] , \w[3][7] , \w[3][6] , \w[3][5] , \w[3][4] , \w[3][3] , 
        \w[3][2] , \w[3][1] , SYNOPSYS_UNCONNECTED__1}) );
  ADD_N32_218 \FAINST[3].ADD_  ( .A({\_4_net_[31] , \_4_net_[30] , 
        \_4_net_[29] , \_4_net_[28] , \_4_net_[27] , \_4_net_[26] , 
        \_4_net_[25] , \_4_net_[24] , \_4_net_[23] , \_4_net_[22] , 
        \_4_net_[21] , \_4_net_[20] , \_4_net_[19] , \_4_net_[18] , 
        \_4_net_[17] , \_4_net_[16] , \_4_net_[15] , \_4_net_[14] , 
        \_4_net_[13] , \_4_net_[12] , \_4_net_[11] , \_4_net_[10] , 
        \_4_net_[9] , \_4_net_[8] , \_4_net_[7] , \_4_net_[6] , \_4_net_[5] , 
        \_4_net_[4] , \_4_net_[3] , 1'b0, 1'b0, 1'b0}), .B({\w[3][31] , 
        \w[3][30] , \w[3][29] , \w[3][28] , \w[3][27] , \w[3][26] , \w[3][25] , 
        \w[3][24] , \w[3][23] , \w[3][22] , \w[3][21] , \w[3][20] , \w[3][19] , 
        \w[3][18] , \w[3][17] , \w[3][16] , \w[3][15] , \w[3][14] , \w[3][13] , 
        \w[3][12] , \w[3][11] , \w[3][10] , \w[3][9] , \w[3][8] , \w[3][7] , 
        \w[3][6] , \w[3][5] , \w[3][4] , \w[3][3] , \w[3][2] , \w[3][1] , 1'b0}), .CI(1'b0), .S({\w[4][31] , \w[4][30] , \w[4][29] , \w[4][28] , \w[4][27] , 
        \w[4][26] , \w[4][25] , \w[4][24] , \w[4][23] , \w[4][22] , \w[4][21] , 
        \w[4][20] , \w[4][19] , \w[4][18] , \w[4][17] , \w[4][16] , \w[4][15] , 
        \w[4][14] , \w[4][13] , \w[4][12] , \w[4][11] , \w[4][10] , \w[4][9] , 
        \w[4][8] , \w[4][7] , \w[4][6] , \w[4][5] , \w[4][4] , \w[4][3] , 
        \w[4][2] , \w[4][1] , SYNOPSYS_UNCONNECTED__2}) );
  ADD_N32_217 \FAINST[4].ADD_  ( .A({\_6_net_[31] , \_6_net_[30] , 
        \_6_net_[29] , \_6_net_[28] , \_6_net_[27] , \_6_net_[26] , 
        \_6_net_[25] , \_6_net_[24] , \_6_net_[23] , \_6_net_[22] , 
        \_6_net_[21] , \_6_net_[20] , \_6_net_[19] , \_6_net_[18] , 
        \_6_net_[17] , \_6_net_[16] , \_6_net_[15] , \_6_net_[14] , 
        \_6_net_[13] , \_6_net_[12] , \_6_net_[11] , \_6_net_[10] , 
        \_6_net_[9] , \_6_net_[8] , \_6_net_[7] , \_6_net_[6] , \_6_net_[5] , 
        \_6_net_[4] , 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[4][31] , \w[4][30] , 
        \w[4][29] , \w[4][28] , \w[4][27] , \w[4][26] , \w[4][25] , \w[4][24] , 
        \w[4][23] , \w[4][22] , \w[4][21] , \w[4][20] , \w[4][19] , \w[4][18] , 
        \w[4][17] , \w[4][16] , \w[4][15] , \w[4][14] , \w[4][13] , \w[4][12] , 
        \w[4][11] , \w[4][10] , \w[4][9] , \w[4][8] , \w[4][7] , \w[4][6] , 
        \w[4][5] , \w[4][4] , \w[4][3] , \w[4][2] , \w[4][1] , 1'b0}), .CI(
        1'b0), .S({\w[5][31] , \w[5][30] , \w[5][29] , \w[5][28] , \w[5][27] , 
        \w[5][26] , \w[5][25] , \w[5][24] , \w[5][23] , \w[5][22] , \w[5][21] , 
        \w[5][20] , \w[5][19] , \w[5][18] , \w[5][17] , \w[5][16] , \w[5][15] , 
        \w[5][14] , \w[5][13] , \w[5][12] , \w[5][11] , \w[5][10] , \w[5][9] , 
        \w[5][8] , \w[5][7] , \w[5][6] , \w[5][5] , \w[5][4] , \w[5][3] , 
        \w[5][2] , \w[5][1] , SYNOPSYS_UNCONNECTED__3}) );
  ADD_N32_216 \FAINST[5].ADD_  ( .A({\_8_net_[31] , \_8_net_[30] , 
        \_8_net_[29] , \_8_net_[28] , \_8_net_[27] , \_8_net_[26] , 
        \_8_net_[25] , \_8_net_[24] , \_8_net_[23] , \_8_net_[22] , 
        \_8_net_[21] , \_8_net_[20] , \_8_net_[19] , \_8_net_[18] , 
        \_8_net_[17] , \_8_net_[16] , \_8_net_[15] , \_8_net_[14] , 
        \_8_net_[13] , \_8_net_[12] , \_8_net_[11] , \_8_net_[10] , 
        \_8_net_[9] , \_8_net_[8] , \_8_net_[7] , \_8_net_[6] , \_8_net_[5] , 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[5][31] , \w[5][30] , \w[5][29] , 
        \w[5][28] , \w[5][27] , \w[5][26] , \w[5][25] , \w[5][24] , \w[5][23] , 
        \w[5][22] , \w[5][21] , \w[5][20] , \w[5][19] , \w[5][18] , \w[5][17] , 
        \w[5][16] , \w[5][15] , \w[5][14] , \w[5][13] , \w[5][12] , \w[5][11] , 
        \w[5][10] , \w[5][9] , \w[5][8] , \w[5][7] , \w[5][6] , \w[5][5] , 
        \w[5][4] , \w[5][3] , \w[5][2] , \w[5][1] , 1'b0}), .CI(1'b0), .S({
        \w[6][31] , \w[6][30] , \w[6][29] , \w[6][28] , \w[6][27] , \w[6][26] , 
        \w[6][25] , \w[6][24] , \w[6][23] , \w[6][22] , \w[6][21] , \w[6][20] , 
        \w[6][19] , \w[6][18] , \w[6][17] , \w[6][16] , \w[6][15] , \w[6][14] , 
        \w[6][13] , \w[6][12] , \w[6][11] , \w[6][10] , \w[6][9] , \w[6][8] , 
        \w[6][7] , \w[6][6] , \w[6][5] , \w[6][4] , \w[6][3] , \w[6][2] , 
        \w[6][1] , SYNOPSYS_UNCONNECTED__4}) );
  ADD_N32_215 \FAINST[6].ADD_  ( .A({\_10_net_[31] , \_10_net_[30] , 
        \_10_net_[29] , \_10_net_[28] , \_10_net_[27] , \_10_net_[26] , 
        \_10_net_[25] , \_10_net_[24] , \_10_net_[23] , \_10_net_[22] , 
        \_10_net_[21] , \_10_net_[20] , \_10_net_[19] , \_10_net_[18] , 
        \_10_net_[17] , \_10_net_[16] , \_10_net_[15] , \_10_net_[14] , 
        \_10_net_[13] , \_10_net_[12] , \_10_net_[11] , \_10_net_[10] , 
        \_10_net_[9] , \_10_net_[8] , \_10_net_[7] , \_10_net_[6] , 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[6][31] , \w[6][30] , \w[6][29] , 
        \w[6][28] , \w[6][27] , \w[6][26] , \w[6][25] , \w[6][24] , \w[6][23] , 
        \w[6][22] , \w[6][21] , \w[6][20] , \w[6][19] , \w[6][18] , \w[6][17] , 
        \w[6][16] , \w[6][15] , \w[6][14] , \w[6][13] , \w[6][12] , \w[6][11] , 
        \w[6][10] , \w[6][9] , \w[6][8] , \w[6][7] , \w[6][6] , \w[6][5] , 
        \w[6][4] , \w[6][3] , \w[6][2] , \w[6][1] , 1'b0}), .CI(1'b0), .S({
        \w[7][31] , \w[7][30] , \w[7][29] , \w[7][28] , \w[7][27] , \w[7][26] , 
        \w[7][25] , \w[7][24] , \w[7][23] , \w[7][22] , \w[7][21] , \w[7][20] , 
        \w[7][19] , \w[7][18] , \w[7][17] , \w[7][16] , \w[7][15] , \w[7][14] , 
        \w[7][13] , \w[7][12] , \w[7][11] , \w[7][10] , \w[7][9] , \w[7][8] , 
        \w[7][7] , \w[7][6] , \w[7][5] , \w[7][4] , \w[7][3] , \w[7][2] , 
        \w[7][1] , SYNOPSYS_UNCONNECTED__5}) );
  ADD_N32_214 \FAINST[7].ADD_  ( .A({\_12_net_[31] , \_12_net_[30] , 
        \_12_net_[29] , \_12_net_[28] , \_12_net_[27] , \_12_net_[26] , 
        \_12_net_[25] , \_12_net_[24] , \_12_net_[23] , \_12_net_[22] , 
        \_12_net_[21] , \_12_net_[20] , \_12_net_[19] , \_12_net_[18] , 
        \_12_net_[17] , \_12_net_[16] , \_12_net_[15] , \_12_net_[14] , 
        \_12_net_[13] , \_12_net_[12] , \_12_net_[11] , \_12_net_[10] , 
        \_12_net_[9] , \_12_net_[8] , \_12_net_[7] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({\w[7][31] , \w[7][30] , \w[7][29] , \w[7][28] , 
        \w[7][27] , \w[7][26] , \w[7][25] , \w[7][24] , \w[7][23] , \w[7][22] , 
        \w[7][21] , \w[7][20] , \w[7][19] , \w[7][18] , \w[7][17] , \w[7][16] , 
        \w[7][15] , \w[7][14] , \w[7][13] , \w[7][12] , \w[7][11] , \w[7][10] , 
        \w[7][9] , \w[7][8] , \w[7][7] , \w[7][6] , \w[7][5] , \w[7][4] , 
        \w[7][3] , \w[7][2] , \w[7][1] , 1'b0}), .CI(1'b0), .S({\w[8][31] , 
        \w[8][30] , \w[8][29] , \w[8][28] , \w[8][27] , \w[8][26] , \w[8][25] , 
        \w[8][24] , \w[8][23] , \w[8][22] , \w[8][21] , \w[8][20] , \w[8][19] , 
        \w[8][18] , \w[8][17] , \w[8][16] , \w[8][15] , \w[8][14] , \w[8][13] , 
        \w[8][12] , \w[8][11] , \w[8][10] , \w[8][9] , \w[8][8] , \w[8][7] , 
        \w[8][6] , \w[8][5] , \w[8][4] , \w[8][3] , \w[8][2] , \w[8][1] , 
        SYNOPSYS_UNCONNECTED__6}) );
  ADD_N32_213 \FAINST[8].ADD_  ( .A({\_14_net_[31] , \_14_net_[30] , 
        \_14_net_[29] , \_14_net_[28] , \_14_net_[27] , \_14_net_[26] , 
        \_14_net_[25] , \_14_net_[24] , \_14_net_[23] , \_14_net_[22] , 
        \_14_net_[21] , \_14_net_[20] , \_14_net_[19] , \_14_net_[18] , 
        \_14_net_[17] , \_14_net_[16] , \_14_net_[15] , \_14_net_[14] , 
        \_14_net_[13] , \_14_net_[12] , \_14_net_[11] , \_14_net_[10] , 
        \_14_net_[9] , \_14_net_[8] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({\w[8][31] , \w[8][30] , \w[8][29] , \w[8][28] , \w[8][27] , 
        \w[8][26] , \w[8][25] , \w[8][24] , \w[8][23] , \w[8][22] , \w[8][21] , 
        \w[8][20] , \w[8][19] , \w[8][18] , \w[8][17] , \w[8][16] , \w[8][15] , 
        \w[8][14] , \w[8][13] , \w[8][12] , \w[8][11] , \w[8][10] , \w[8][9] , 
        \w[8][8] , \w[8][7] , \w[8][6] , \w[8][5] , \w[8][4] , \w[8][3] , 
        \w[8][2] , \w[8][1] , 1'b0}), .CI(1'b0), .S({\w[9][31] , \w[9][30] , 
        \w[9][29] , \w[9][28] , \w[9][27] , \w[9][26] , \w[9][25] , \w[9][24] , 
        \w[9][23] , \w[9][22] , \w[9][21] , \w[9][20] , \w[9][19] , \w[9][18] , 
        \w[9][17] , \w[9][16] , \w[9][15] , \w[9][14] , \w[9][13] , \w[9][12] , 
        \w[9][11] , \w[9][10] , \w[9][9] , \w[9][8] , \w[9][7] , \w[9][6] , 
        \w[9][5] , \w[9][4] , \w[9][3] , \w[9][2] , \w[9][1] , 
        SYNOPSYS_UNCONNECTED__7}) );
  ADD_N32_212 \FAINST[9].ADD_  ( .A({\_16_net_[31] , \_16_net_[30] , 
        \_16_net_[29] , \_16_net_[28] , \_16_net_[27] , \_16_net_[26] , 
        \_16_net_[25] , \_16_net_[24] , \_16_net_[23] , \_16_net_[22] , 
        \_16_net_[21] , \_16_net_[20] , \_16_net_[19] , \_16_net_[18] , 
        \_16_net_[17] , \_16_net_[16] , \_16_net_[15] , \_16_net_[14] , 
        \_16_net_[13] , \_16_net_[12] , \_16_net_[11] , \_16_net_[10] , 
        \_16_net_[9] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({\w[9][31] , \w[9][30] , \w[9][29] , \w[9][28] , \w[9][27] , 
        \w[9][26] , \w[9][25] , \w[9][24] , \w[9][23] , \w[9][22] , \w[9][21] , 
        \w[9][20] , \w[9][19] , \w[9][18] , \w[9][17] , \w[9][16] , \w[9][15] , 
        \w[9][14] , \w[9][13] , \w[9][12] , \w[9][11] , \w[9][10] , \w[9][9] , 
        \w[9][8] , \w[9][7] , \w[9][6] , \w[9][5] , \w[9][4] , \w[9][3] , 
        \w[9][2] , \w[9][1] , 1'b0}), .CI(1'b0), .S({\w[10][31] , \w[10][30] , 
        \w[10][29] , \w[10][28] , \w[10][27] , \w[10][26] , \w[10][25] , 
        \w[10][24] , \w[10][23] , \w[10][22] , \w[10][21] , \w[10][20] , 
        \w[10][19] , \w[10][18] , \w[10][17] , \w[10][16] , \w[10][15] , 
        \w[10][14] , \w[10][13] , \w[10][12] , \w[10][11] , \w[10][10] , 
        \w[10][9] , \w[10][8] , \w[10][7] , \w[10][6] , \w[10][5] , \w[10][4] , 
        \w[10][3] , \w[10][2] , \w[10][1] , SYNOPSYS_UNCONNECTED__8}) );
  ADD_N32_211 \FAINST[10].ADD_  ( .A({\_18_net_[31] , \_18_net_[30] , 
        \_18_net_[29] , \_18_net_[28] , \_18_net_[27] , \_18_net_[26] , 
        \_18_net_[25] , \_18_net_[24] , \_18_net_[23] , \_18_net_[22] , 
        \_18_net_[21] , \_18_net_[20] , \_18_net_[19] , \_18_net_[18] , 
        \_18_net_[17] , \_18_net_[16] , \_18_net_[15] , \_18_net_[14] , 
        \_18_net_[13] , \_18_net_[12] , \_18_net_[11] , \_18_net_[10] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[10][31] , \w[10][30] , \w[10][29] , \w[10][28] , \w[10][27] , 
        \w[10][26] , \w[10][25] , \w[10][24] , \w[10][23] , \w[10][22] , 
        \w[10][21] , \w[10][20] , \w[10][19] , \w[10][18] , \w[10][17] , 
        \w[10][16] , \w[10][15] , \w[10][14] , \w[10][13] , \w[10][12] , 
        \w[10][11] , \w[10][10] , \w[10][9] , \w[10][8] , \w[10][7] , 
        \w[10][6] , \w[10][5] , \w[10][4] , \w[10][3] , \w[10][2] , \w[10][1] , 
        1'b0}), .CI(1'b0), .S({\w[11][31] , \w[11][30] , \w[11][29] , 
        \w[11][28] , \w[11][27] , \w[11][26] , \w[11][25] , \w[11][24] , 
        \w[11][23] , \w[11][22] , \w[11][21] , \w[11][20] , \w[11][19] , 
        \w[11][18] , \w[11][17] , \w[11][16] , \w[11][15] , \w[11][14] , 
        \w[11][13] , \w[11][12] , \w[11][11] , \w[11][10] , \w[11][9] , 
        \w[11][8] , \w[11][7] , \w[11][6] , \w[11][5] , \w[11][4] , \w[11][3] , 
        \w[11][2] , \w[11][1] , SYNOPSYS_UNCONNECTED__9}) );
  ADD_N32_210 \FAINST[11].ADD_  ( .A({\_20_net_[31] , \_20_net_[30] , 
        \_20_net_[29] , \_20_net_[28] , \_20_net_[27] , \_20_net_[26] , 
        \_20_net_[25] , \_20_net_[24] , \_20_net_[23] , \_20_net_[22] , 
        \_20_net_[21] , \_20_net_[20] , \_20_net_[19] , \_20_net_[18] , 
        \_20_net_[17] , \_20_net_[16] , \_20_net_[15] , \_20_net_[14] , 
        \_20_net_[13] , \_20_net_[12] , \_20_net_[11] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[11][31] , 
        \w[11][30] , \w[11][29] , \w[11][28] , \w[11][27] , \w[11][26] , 
        \w[11][25] , \w[11][24] , \w[11][23] , \w[11][22] , \w[11][21] , 
        \w[11][20] , \w[11][19] , \w[11][18] , \w[11][17] , \w[11][16] , 
        \w[11][15] , \w[11][14] , \w[11][13] , \w[11][12] , \w[11][11] , 
        \w[11][10] , \w[11][9] , \w[11][8] , \w[11][7] , \w[11][6] , 
        \w[11][5] , \w[11][4] , \w[11][3] , \w[11][2] , \w[11][1] , 1'b0}), 
        .CI(1'b0), .S({\w[12][31] , \w[12][30] , \w[12][29] , \w[12][28] , 
        \w[12][27] , \w[12][26] , \w[12][25] , \w[12][24] , \w[12][23] , 
        \w[12][22] , \w[12][21] , \w[12][20] , \w[12][19] , \w[12][18] , 
        \w[12][17] , \w[12][16] , \w[12][15] , \w[12][14] , \w[12][13] , 
        \w[12][12] , \w[12][11] , \w[12][10] , \w[12][9] , \w[12][8] , 
        \w[12][7] , \w[12][6] , \w[12][5] , \w[12][4] , \w[12][3] , \w[12][2] , 
        \w[12][1] , SYNOPSYS_UNCONNECTED__10}) );
  ADD_N32_209 \FAINST[12].ADD_  ( .A({\_22_net_[31] , \_22_net_[30] , 
        \_22_net_[29] , \_22_net_[28] , \_22_net_[27] , \_22_net_[26] , 
        \_22_net_[25] , \_22_net_[24] , \_22_net_[23] , \_22_net_[22] , 
        \_22_net_[21] , \_22_net_[20] , \_22_net_[19] , \_22_net_[18] , 
        \_22_net_[17] , \_22_net_[16] , \_22_net_[15] , \_22_net_[14] , 
        \_22_net_[13] , \_22_net_[12] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[12][31] , \w[12][30] , 
        \w[12][29] , \w[12][28] , \w[12][27] , \w[12][26] , \w[12][25] , 
        \w[12][24] , \w[12][23] , \w[12][22] , \w[12][21] , \w[12][20] , 
        \w[12][19] , \w[12][18] , \w[12][17] , \w[12][16] , \w[12][15] , 
        \w[12][14] , \w[12][13] , \w[12][12] , \w[12][11] , \w[12][10] , 
        \w[12][9] , \w[12][8] , \w[12][7] , \w[12][6] , \w[12][5] , \w[12][4] , 
        \w[12][3] , \w[12][2] , \w[12][1] , 1'b0}), .CI(1'b0), .S({\w[13][31] , 
        \w[13][30] , \w[13][29] , \w[13][28] , \w[13][27] , \w[13][26] , 
        \w[13][25] , \w[13][24] , \w[13][23] , \w[13][22] , \w[13][21] , 
        \w[13][20] , \w[13][19] , \w[13][18] , \w[13][17] , \w[13][16] , 
        \w[13][15] , \w[13][14] , \w[13][13] , \w[13][12] , \w[13][11] , 
        \w[13][10] , \w[13][9] , \w[13][8] , \w[13][7] , \w[13][6] , 
        \w[13][5] , \w[13][4] , \w[13][3] , \w[13][2] , \w[13][1] , 
        SYNOPSYS_UNCONNECTED__11}) );
  ADD_N32_208 \FAINST[13].ADD_  ( .A({\_24_net_[31] , \_24_net_[30] , 
        \_24_net_[29] , \_24_net_[28] , \_24_net_[27] , \_24_net_[26] , 
        \_24_net_[25] , \_24_net_[24] , \_24_net_[23] , \_24_net_[22] , 
        \_24_net_[21] , \_24_net_[20] , \_24_net_[19] , \_24_net_[18] , 
        \_24_net_[17] , \_24_net_[16] , \_24_net_[15] , \_24_net_[14] , 
        \_24_net_[13] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[13][31] , \w[13][30] , \w[13][29] , 
        \w[13][28] , \w[13][27] , \w[13][26] , \w[13][25] , \w[13][24] , 
        \w[13][23] , \w[13][22] , \w[13][21] , \w[13][20] , \w[13][19] , 
        \w[13][18] , \w[13][17] , \w[13][16] , \w[13][15] , \w[13][14] , 
        \w[13][13] , \w[13][12] , \w[13][11] , \w[13][10] , \w[13][9] , 
        \w[13][8] , \w[13][7] , \w[13][6] , \w[13][5] , \w[13][4] , \w[13][3] , 
        \w[13][2] , \w[13][1] , 1'b0}), .CI(1'b0), .S({\w[14][31] , 
        \w[14][30] , \w[14][29] , \w[14][28] , \w[14][27] , \w[14][26] , 
        \w[14][25] , \w[14][24] , \w[14][23] , \w[14][22] , \w[14][21] , 
        \w[14][20] , \w[14][19] , \w[14][18] , \w[14][17] , \w[14][16] , 
        \w[14][15] , \w[14][14] , \w[14][13] , \w[14][12] , \w[14][11] , 
        \w[14][10] , \w[14][9] , \w[14][8] , \w[14][7] , \w[14][6] , 
        \w[14][5] , \w[14][4] , \w[14][3] , \w[14][2] , \w[14][1] , 
        SYNOPSYS_UNCONNECTED__12}) );
  ADD_N32_207 \FAINST[14].ADD_  ( .A({\_26_net_[31] , \_26_net_[30] , 
        \_26_net_[29] , \_26_net_[28] , \_26_net_[27] , \_26_net_[26] , 
        \_26_net_[25] , \_26_net_[24] , \_26_net_[23] , \_26_net_[22] , 
        \_26_net_[21] , \_26_net_[20] , \_26_net_[19] , \_26_net_[18] , 
        \_26_net_[17] , \_26_net_[16] , \_26_net_[15] , \_26_net_[14] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({\w[14][31] , \w[14][30] , \w[14][29] , \w[14][28] , 
        \w[14][27] , \w[14][26] , \w[14][25] , \w[14][24] , \w[14][23] , 
        \w[14][22] , \w[14][21] , \w[14][20] , \w[14][19] , \w[14][18] , 
        \w[14][17] , \w[14][16] , \w[14][15] , \w[14][14] , \w[14][13] , 
        \w[14][12] , \w[14][11] , \w[14][10] , \w[14][9] , \w[14][8] , 
        \w[14][7] , \w[14][6] , \w[14][5] , \w[14][4] , \w[14][3] , \w[14][2] , 
        \w[14][1] , 1'b0}), .CI(1'b0), .S({\w[15][31] , \w[15][30] , 
        \w[15][29] , \w[15][28] , \w[15][27] , \w[15][26] , \w[15][25] , 
        \w[15][24] , \w[15][23] , \w[15][22] , \w[15][21] , \w[15][20] , 
        \w[15][19] , \w[15][18] , \w[15][17] , \w[15][16] , \w[15][15] , 
        \w[15][14] , \w[15][13] , \w[15][12] , \w[15][11] , \w[15][10] , 
        \w[15][9] , \w[15][8] , \w[15][7] , \w[15][6] , \w[15][5] , \w[15][4] , 
        \w[15][3] , \w[15][2] , \w[15][1] , SYNOPSYS_UNCONNECTED__13}) );
  ADD_N32_206 \FAINST[15].ADD_  ( .A({\_28_net_[31] , \_28_net_[30] , 
        \_28_net_[29] , \_28_net_[28] , \_28_net_[27] , \_28_net_[26] , 
        \_28_net_[25] , \_28_net_[24] , \_28_net_[23] , \_28_net_[22] , 
        \_28_net_[21] , \_28_net_[20] , \_28_net_[19] , \_28_net_[18] , 
        \_28_net_[17] , \_28_net_[16] , \_28_net_[15] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({\w[15][31] , \w[15][30] , \w[15][29] , \w[15][28] , \w[15][27] , 
        \w[15][26] , \w[15][25] , \w[15][24] , \w[15][23] , \w[15][22] , 
        \w[15][21] , \w[15][20] , \w[15][19] , \w[15][18] , \w[15][17] , 
        \w[15][16] , \w[15][15] , \w[15][14] , \w[15][13] , \w[15][12] , 
        \w[15][11] , \w[15][10] , \w[15][9] , \w[15][8] , \w[15][7] , 
        \w[15][6] , \w[15][5] , \w[15][4] , \w[15][3] , \w[15][2] , \w[15][1] , 
        1'b0}), .CI(1'b0), .S({\w[16][31] , \w[16][30] , \w[16][29] , 
        \w[16][28] , \w[16][27] , \w[16][26] , \w[16][25] , \w[16][24] , 
        \w[16][23] , \w[16][22] , \w[16][21] , \w[16][20] , \w[16][19] , 
        \w[16][18] , \w[16][17] , \w[16][16] , \w[16][15] , \w[16][14] , 
        \w[16][13] , \w[16][12] , \w[16][11] , \w[16][10] , \w[16][9] , 
        \w[16][8] , \w[16][7] , \w[16][6] , \w[16][5] , \w[16][4] , \w[16][3] , 
        \w[16][2] , \w[16][1] , SYNOPSYS_UNCONNECTED__14}) );
  ADD_N32_205 \FAINST[16].ADD_  ( .A({\_30_net_[31] , \_30_net_[30] , 
        \_30_net_[29] , \_30_net_[28] , \_30_net_[27] , \_30_net_[26] , 
        \_30_net_[25] , \_30_net_[24] , \_30_net_[23] , \_30_net_[22] , 
        \_30_net_[21] , \_30_net_[20] , \_30_net_[19] , \_30_net_[18] , 
        \_30_net_[17] , \_30_net_[16] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[16][31] , \w[16][30] , \w[16][29] , \w[16][28] , \w[16][27] , 
        \w[16][26] , \w[16][25] , \w[16][24] , \w[16][23] , \w[16][22] , 
        \w[16][21] , \w[16][20] , \w[16][19] , \w[16][18] , \w[16][17] , 
        \w[16][16] , \w[16][15] , \w[16][14] , \w[16][13] , \w[16][12] , 
        \w[16][11] , \w[16][10] , \w[16][9] , \w[16][8] , \w[16][7] , 
        \w[16][6] , \w[16][5] , \w[16][4] , \w[16][3] , \w[16][2] , \w[16][1] , 
        1'b0}), .CI(1'b0), .S({\w[17][31] , \w[17][30] , \w[17][29] , 
        \w[17][28] , \w[17][27] , \w[17][26] , \w[17][25] , \w[17][24] , 
        \w[17][23] , \w[17][22] , \w[17][21] , \w[17][20] , \w[17][19] , 
        \w[17][18] , \w[17][17] , \w[17][16] , \w[17][15] , \w[17][14] , 
        \w[17][13] , \w[17][12] , \w[17][11] , \w[17][10] , \w[17][9] , 
        \w[17][8] , \w[17][7] , \w[17][6] , \w[17][5] , \w[17][4] , \w[17][3] , 
        \w[17][2] , \w[17][1] , SYNOPSYS_UNCONNECTED__15}) );
  ADD_N32_204 \FAINST[17].ADD_  ( .A({\_32_net_[31] , \_32_net_[30] , 
        \_32_net_[29] , \_32_net_[28] , \_32_net_[27] , \_32_net_[26] , 
        \_32_net_[25] , \_32_net_[24] , \_32_net_[23] , \_32_net_[22] , 
        \_32_net_[21] , \_32_net_[20] , \_32_net_[19] , \_32_net_[18] , 
        \_32_net_[17] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[17][31] , 
        \w[17][30] , \w[17][29] , \w[17][28] , \w[17][27] , \w[17][26] , 
        \w[17][25] , \w[17][24] , \w[17][23] , \w[17][22] , \w[17][21] , 
        \w[17][20] , \w[17][19] , \w[17][18] , \w[17][17] , \w[17][16] , 
        \w[17][15] , \w[17][14] , \w[17][13] , \w[17][12] , \w[17][11] , 
        \w[17][10] , \w[17][9] , \w[17][8] , \w[17][7] , \w[17][6] , 
        \w[17][5] , \w[17][4] , \w[17][3] , \w[17][2] , \w[17][1] , 1'b0}), 
        .CI(1'b0), .S({\w[18][31] , \w[18][30] , \w[18][29] , \w[18][28] , 
        \w[18][27] , \w[18][26] , \w[18][25] , \w[18][24] , \w[18][23] , 
        \w[18][22] , \w[18][21] , \w[18][20] , \w[18][19] , \w[18][18] , 
        \w[18][17] , \w[18][16] , \w[18][15] , \w[18][14] , \w[18][13] , 
        \w[18][12] , \w[18][11] , \w[18][10] , \w[18][9] , \w[18][8] , 
        \w[18][7] , \w[18][6] , \w[18][5] , \w[18][4] , \w[18][3] , \w[18][2] , 
        \w[18][1] , SYNOPSYS_UNCONNECTED__16}) );
  ADD_N32_203 \FAINST[18].ADD_  ( .A({\_34_net_[31] , \_34_net_[30] , 
        \_34_net_[29] , \_34_net_[28] , \_34_net_[27] , \_34_net_[26] , 
        \_34_net_[25] , \_34_net_[24] , \_34_net_[23] , \_34_net_[22] , 
        \_34_net_[21] , \_34_net_[20] , \_34_net_[19] , \_34_net_[18] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[18][31] , \w[18][30] , 
        \w[18][29] , \w[18][28] , \w[18][27] , \w[18][26] , \w[18][25] , 
        \w[18][24] , \w[18][23] , \w[18][22] , \w[18][21] , \w[18][20] , 
        \w[18][19] , \w[18][18] , \w[18][17] , \w[18][16] , \w[18][15] , 
        \w[18][14] , \w[18][13] , \w[18][12] , \w[18][11] , \w[18][10] , 
        \w[18][9] , \w[18][8] , \w[18][7] , \w[18][6] , \w[18][5] , \w[18][4] , 
        \w[18][3] , \w[18][2] , \w[18][1] , 1'b0}), .CI(1'b0), .S({\w[19][31] , 
        \w[19][30] , \w[19][29] , \w[19][28] , \w[19][27] , \w[19][26] , 
        \w[19][25] , \w[19][24] , \w[19][23] , \w[19][22] , \w[19][21] , 
        \w[19][20] , \w[19][19] , \w[19][18] , \w[19][17] , \w[19][16] , 
        \w[19][15] , \w[19][14] , \w[19][13] , \w[19][12] , \w[19][11] , 
        \w[19][10] , \w[19][9] , \w[19][8] , \w[19][7] , \w[19][6] , 
        \w[19][5] , \w[19][4] , \w[19][3] , \w[19][2] , \w[19][1] , 
        SYNOPSYS_UNCONNECTED__17}) );
  ADD_N32_202 \FAINST[19].ADD_  ( .A({\_36_net_[31] , \_36_net_[30] , 
        \_36_net_[29] , \_36_net_[28] , \_36_net_[27] , \_36_net_[26] , 
        \_36_net_[25] , \_36_net_[24] , \_36_net_[23] , \_36_net_[22] , 
        \_36_net_[21] , \_36_net_[20] , \_36_net_[19] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({\w[19][31] , \w[19][30] , \w[19][29] , 
        \w[19][28] , \w[19][27] , \w[19][26] , \w[19][25] , \w[19][24] , 
        \w[19][23] , \w[19][22] , \w[19][21] , \w[19][20] , \w[19][19] , 
        \w[19][18] , \w[19][17] , \w[19][16] , \w[19][15] , \w[19][14] , 
        \w[19][13] , \w[19][12] , \w[19][11] , \w[19][10] , \w[19][9] , 
        \w[19][8] , \w[19][7] , \w[19][6] , \w[19][5] , \w[19][4] , \w[19][3] , 
        \w[19][2] , \w[19][1] , 1'b0}), .CI(1'b0), .S({\w[20][31] , 
        \w[20][30] , \w[20][29] , \w[20][28] , \w[20][27] , \w[20][26] , 
        \w[20][25] , \w[20][24] , \w[20][23] , \w[20][22] , \w[20][21] , 
        \w[20][20] , \w[20][19] , \w[20][18] , \w[20][17] , \w[20][16] , 
        \w[20][15] , \w[20][14] , \w[20][13] , \w[20][12] , \w[20][11] , 
        \w[20][10] , \w[20][9] , \w[20][8] , \w[20][7] , \w[20][6] , 
        \w[20][5] , \w[20][4] , \w[20][3] , \w[20][2] , \w[20][1] , 
        SYNOPSYS_UNCONNECTED__18}) );
  ADD_N32_201 \FAINST[20].ADD_  ( .A({\_38_net_[31] , \_38_net_[30] , 
        \_38_net_[29] , \_38_net_[28] , \_38_net_[27] , \_38_net_[26] , 
        \_38_net_[25] , \_38_net_[24] , \_38_net_[23] , \_38_net_[22] , 
        \_38_net_[21] , \_38_net_[20] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .B({\w[20][31] , \w[20][30] , \w[20][29] , \w[20][28] , 
        \w[20][27] , \w[20][26] , \w[20][25] , \w[20][24] , \w[20][23] , 
        \w[20][22] , \w[20][21] , \w[20][20] , \w[20][19] , \w[20][18] , 
        \w[20][17] , \w[20][16] , \w[20][15] , \w[20][14] , \w[20][13] , 
        \w[20][12] , \w[20][11] , \w[20][10] , \w[20][9] , \w[20][8] , 
        \w[20][7] , \w[20][6] , \w[20][5] , \w[20][4] , \w[20][3] , \w[20][2] , 
        \w[20][1] , 1'b0}), .CI(1'b0), .S({\w[21][31] , \w[21][30] , 
        \w[21][29] , \w[21][28] , \w[21][27] , \w[21][26] , \w[21][25] , 
        \w[21][24] , \w[21][23] , \w[21][22] , \w[21][21] , \w[21][20] , 
        \w[21][19] , \w[21][18] , \w[21][17] , \w[21][16] , \w[21][15] , 
        \w[21][14] , \w[21][13] , \w[21][12] , \w[21][11] , \w[21][10] , 
        \w[21][9] , \w[21][8] , \w[21][7] , \w[21][6] , \w[21][5] , \w[21][4] , 
        \w[21][3] , \w[21][2] , \w[21][1] , SYNOPSYS_UNCONNECTED__19}) );
  ADD_N32_200 \FAINST[21].ADD_  ( .A({\_40_net_[31] , \_40_net_[30] , 
        \_40_net_[29] , \_40_net_[28] , \_40_net_[27] , \_40_net_[26] , 
        \_40_net_[25] , \_40_net_[24] , \_40_net_[23] , \_40_net_[22] , 
        \_40_net_[21] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[21][31] , \w[21][30] , \w[21][29] , \w[21][28] , \w[21][27] , 
        \w[21][26] , \w[21][25] , \w[21][24] , \w[21][23] , \w[21][22] , 
        \w[21][21] , \w[21][20] , \w[21][19] , \w[21][18] , \w[21][17] , 
        \w[21][16] , \w[21][15] , \w[21][14] , \w[21][13] , \w[21][12] , 
        \w[21][11] , \w[21][10] , \w[21][9] , \w[21][8] , \w[21][7] , 
        \w[21][6] , \w[21][5] , \w[21][4] , \w[21][3] , \w[21][2] , \w[21][1] , 
        1'b0}), .CI(1'b0), .S({\w[22][31] , \w[22][30] , \w[22][29] , 
        \w[22][28] , \w[22][27] , \w[22][26] , \w[22][25] , \w[22][24] , 
        \w[22][23] , \w[22][22] , \w[22][21] , \w[22][20] , \w[22][19] , 
        \w[22][18] , \w[22][17] , \w[22][16] , \w[22][15] , \w[22][14] , 
        \w[22][13] , \w[22][12] , \w[22][11] , \w[22][10] , \w[22][9] , 
        \w[22][8] , \w[22][7] , \w[22][6] , \w[22][5] , \w[22][4] , \w[22][3] , 
        \w[22][2] , \w[22][1] , SYNOPSYS_UNCONNECTED__20}) );
  ADD_N32_199 \FAINST[22].ADD_  ( .A({\_42_net_[31] , \_42_net_[30] , 
        \_42_net_[29] , \_42_net_[28] , \_42_net_[27] , \_42_net_[26] , 
        \_42_net_[25] , \_42_net_[24] , \_42_net_[23] , \_42_net_[22] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[22][31] , \w[22][30] , \w[22][29] , \w[22][28] , \w[22][27] , 
        \w[22][26] , \w[22][25] , \w[22][24] , \w[22][23] , \w[22][22] , 
        \w[22][21] , \w[22][20] , \w[22][19] , \w[22][18] , \w[22][17] , 
        \w[22][16] , \w[22][15] , \w[22][14] , \w[22][13] , \w[22][12] , 
        \w[22][11] , \w[22][10] , \w[22][9] , \w[22][8] , \w[22][7] , 
        \w[22][6] , \w[22][5] , \w[22][4] , \w[22][3] , \w[22][2] , \w[22][1] , 
        1'b0}), .CI(1'b0), .S({\w[23][31] , \w[23][30] , \w[23][29] , 
        \w[23][28] , \w[23][27] , \w[23][26] , \w[23][25] , \w[23][24] , 
        \w[23][23] , \w[23][22] , \w[23][21] , \w[23][20] , \w[23][19] , 
        \w[23][18] , \w[23][17] , \w[23][16] , \w[23][15] , \w[23][14] , 
        \w[23][13] , \w[23][12] , \w[23][11] , \w[23][10] , \w[23][9] , 
        \w[23][8] , \w[23][7] , \w[23][6] , \w[23][5] , \w[23][4] , \w[23][3] , 
        \w[23][2] , \w[23][1] , SYNOPSYS_UNCONNECTED__21}) );
  ADD_N32_198 \FAINST[23].ADD_  ( .A({\_44_net_[31] , \_44_net_[30] , 
        \_44_net_[29] , \_44_net_[28] , \_44_net_[27] , \_44_net_[26] , 
        \_44_net_[25] , \_44_net_[24] , \_44_net_[23] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[23][31] , 
        \w[23][30] , \w[23][29] , \w[23][28] , \w[23][27] , \w[23][26] , 
        \w[23][25] , \w[23][24] , \w[23][23] , \w[23][22] , \w[23][21] , 
        \w[23][20] , \w[23][19] , \w[23][18] , \w[23][17] , \w[23][16] , 
        \w[23][15] , \w[23][14] , \w[23][13] , \w[23][12] , \w[23][11] , 
        \w[23][10] , \w[23][9] , \w[23][8] , \w[23][7] , \w[23][6] , 
        \w[23][5] , \w[23][4] , \w[23][3] , \w[23][2] , \w[23][1] , 1'b0}), 
        .CI(1'b0), .S({\w[24][31] , \w[24][30] , \w[24][29] , \w[24][28] , 
        \w[24][27] , \w[24][26] , \w[24][25] , \w[24][24] , \w[24][23] , 
        \w[24][22] , \w[24][21] , \w[24][20] , \w[24][19] , \w[24][18] , 
        \w[24][17] , \w[24][16] , \w[24][15] , \w[24][14] , \w[24][13] , 
        \w[24][12] , \w[24][11] , \w[24][10] , \w[24][9] , \w[24][8] , 
        \w[24][7] , \w[24][6] , \w[24][5] , \w[24][4] , \w[24][3] , \w[24][2] , 
        \w[24][1] , SYNOPSYS_UNCONNECTED__22}) );
  ADD_N32_197 \FAINST[24].ADD_  ( .A({\_46_net_[31] , \_46_net_[30] , 
        \_46_net_[29] , \_46_net_[28] , \_46_net_[27] , \_46_net_[26] , 
        \_46_net_[25] , \_46_net_[24] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[24][31] , \w[24][30] , 
        \w[24][29] , \w[24][28] , \w[24][27] , \w[24][26] , \w[24][25] , 
        \w[24][24] , \w[24][23] , \w[24][22] , \w[24][21] , \w[24][20] , 
        \w[24][19] , \w[24][18] , \w[24][17] , \w[24][16] , \w[24][15] , 
        \w[24][14] , \w[24][13] , \w[24][12] , \w[24][11] , \w[24][10] , 
        \w[24][9] , \w[24][8] , \w[24][7] , \w[24][6] , \w[24][5] , \w[24][4] , 
        \w[24][3] , \w[24][2] , \w[24][1] , 1'b0}), .CI(1'b0), .S({\w[25][31] , 
        \w[25][30] , \w[25][29] , \w[25][28] , \w[25][27] , \w[25][26] , 
        \w[25][25] , \w[25][24] , \w[25][23] , \w[25][22] , \w[25][21] , 
        \w[25][20] , \w[25][19] , \w[25][18] , \w[25][17] , \w[25][16] , 
        \w[25][15] , \w[25][14] , \w[25][13] , \w[25][12] , \w[25][11] , 
        \w[25][10] , \w[25][9] , \w[25][8] , \w[25][7] , \w[25][6] , 
        \w[25][5] , \w[25][4] , \w[25][3] , \w[25][2] , \w[25][1] , 
        SYNOPSYS_UNCONNECTED__23}) );
  ADD_N32_196 \FAINST[25].ADD_  ( .A({\_48_net_[31] , \_48_net_[30] , 
        \_48_net_[29] , \_48_net_[28] , \_48_net_[27] , \_48_net_[26] , 
        \_48_net_[25] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[25][31] , \w[25][30] , \w[25][29] , 
        \w[25][28] , \w[25][27] , \w[25][26] , \w[25][25] , \w[25][24] , 
        \w[25][23] , \w[25][22] , \w[25][21] , \w[25][20] , \w[25][19] , 
        \w[25][18] , \w[25][17] , \w[25][16] , \w[25][15] , \w[25][14] , 
        \w[25][13] , \w[25][12] , \w[25][11] , \w[25][10] , \w[25][9] , 
        \w[25][8] , \w[25][7] , \w[25][6] , \w[25][5] , \w[25][4] , \w[25][3] , 
        \w[25][2] , \w[25][1] , 1'b0}), .CI(1'b0), .S({\w[26][31] , 
        \w[26][30] , \w[26][29] , \w[26][28] , \w[26][27] , \w[26][26] , 
        \w[26][25] , \w[26][24] , \w[26][23] , \w[26][22] , \w[26][21] , 
        \w[26][20] , \w[26][19] , \w[26][18] , \w[26][17] , \w[26][16] , 
        \w[26][15] , \w[26][14] , \w[26][13] , \w[26][12] , \w[26][11] , 
        \w[26][10] , \w[26][9] , \w[26][8] , \w[26][7] , \w[26][6] , 
        \w[26][5] , \w[26][4] , \w[26][3] , \w[26][2] , \w[26][1] , 
        SYNOPSYS_UNCONNECTED__24}) );
  ADD_N32_195 \FAINST[26].ADD_  ( .A({\_50_net_[31] , \_50_net_[30] , 
        \_50_net_[29] , \_50_net_[28] , \_50_net_[27] , \_50_net_[26] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({\w[26][31] , \w[26][30] , \w[26][29] , \w[26][28] , 
        \w[26][27] , \w[26][26] , \w[26][25] , \w[26][24] , \w[26][23] , 
        \w[26][22] , \w[26][21] , \w[26][20] , \w[26][19] , \w[26][18] , 
        \w[26][17] , \w[26][16] , \w[26][15] , \w[26][14] , \w[26][13] , 
        \w[26][12] , \w[26][11] , \w[26][10] , \w[26][9] , \w[26][8] , 
        \w[26][7] , \w[26][6] , \w[26][5] , \w[26][4] , \w[26][3] , \w[26][2] , 
        \w[26][1] , 1'b0}), .CI(1'b0), .S({\w[27][31] , \w[27][30] , 
        \w[27][29] , \w[27][28] , \w[27][27] , \w[27][26] , \w[27][25] , 
        \w[27][24] , \w[27][23] , \w[27][22] , \w[27][21] , \w[27][20] , 
        \w[27][19] , \w[27][18] , \w[27][17] , \w[27][16] , \w[27][15] , 
        \w[27][14] , \w[27][13] , \w[27][12] , \w[27][11] , \w[27][10] , 
        \w[27][9] , \w[27][8] , \w[27][7] , \w[27][6] , \w[27][5] , \w[27][4] , 
        \w[27][3] , \w[27][2] , \w[27][1] , SYNOPSYS_UNCONNECTED__25}) );
  ADD_N32_194 \FAINST[27].ADD_  ( .A({\_52_net_[31] , \_52_net_[30] , 
        \_52_net_[29] , \_52_net_[28] , \_52_net_[27] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({\w[27][31] , \w[27][30] , \w[27][29] , \w[27][28] , \w[27][27] , 
        \w[27][26] , \w[27][25] , \w[27][24] , \w[27][23] , \w[27][22] , 
        \w[27][21] , \w[27][20] , \w[27][19] , \w[27][18] , \w[27][17] , 
        \w[27][16] , \w[27][15] , \w[27][14] , \w[27][13] , \w[27][12] , 
        \w[27][11] , \w[27][10] , \w[27][9] , \w[27][8] , \w[27][7] , 
        \w[27][6] , \w[27][5] , \w[27][4] , \w[27][3] , \w[27][2] , \w[27][1] , 
        1'b0}), .CI(1'b0), .S({\w[28][31] , \w[28][30] , \w[28][29] , 
        \w[28][28] , \w[28][27] , \w[28][26] , \w[28][25] , \w[28][24] , 
        \w[28][23] , \w[28][22] , \w[28][21] , \w[28][20] , \w[28][19] , 
        \w[28][18] , \w[28][17] , \w[28][16] , \w[28][15] , \w[28][14] , 
        \w[28][13] , \w[28][12] , \w[28][11] , \w[28][10] , \w[28][9] , 
        \w[28][8] , \w[28][7] , \w[28][6] , \w[28][5] , \w[28][4] , \w[28][3] , 
        \w[28][2] , \w[28][1] , SYNOPSYS_UNCONNECTED__26}) );
  ADD_N32_193 \FAINST[28].ADD_  ( .A({\_54_net_[31] , \_54_net_[30] , 
        \_54_net_[29] , \_54_net_[28] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[28][31] , \w[28][30] , \w[28][29] , \w[28][28] , \w[28][27] , 
        \w[28][26] , \w[28][25] , \w[28][24] , \w[28][23] , \w[28][22] , 
        \w[28][21] , \w[28][20] , \w[28][19] , \w[28][18] , \w[28][17] , 
        \w[28][16] , \w[28][15] , \w[28][14] , \w[28][13] , \w[28][12] , 
        \w[28][11] , \w[28][10] , \w[28][9] , \w[28][8] , \w[28][7] , 
        \w[28][6] , \w[28][5] , \w[28][4] , \w[28][3] , \w[28][2] , \w[28][1] , 
        1'b0}), .CI(1'b0), .S({\w[29][31] , \w[29][30] , \w[29][29] , 
        \w[29][28] , \w[29][27] , \w[29][26] , \w[29][25] , \w[29][24] , 
        \w[29][23] , \w[29][22] , \w[29][21] , \w[29][20] , \w[29][19] , 
        \w[29][18] , \w[29][17] , \w[29][16] , \w[29][15] , \w[29][14] , 
        \w[29][13] , \w[29][12] , \w[29][11] , \w[29][10] , \w[29][9] , 
        \w[29][8] , \w[29][7] , \w[29][6] , \w[29][5] , \w[29][4] , \w[29][3] , 
        \w[29][2] , \w[29][1] , SYNOPSYS_UNCONNECTED__27}) );
  ADD_N32_192 \FAINST[29].ADD_  ( .A({\_56_net_[31] , \_56_net_[30] , 
        \_56_net_[29] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[29][31] , 
        \w[29][30] , \w[29][29] , \w[29][28] , \w[29][27] , \w[29][26] , 
        \w[29][25] , \w[29][24] , \w[29][23] , \w[29][22] , \w[29][21] , 
        \w[29][20] , \w[29][19] , \w[29][18] , \w[29][17] , \w[29][16] , 
        \w[29][15] , \w[29][14] , \w[29][13] , \w[29][12] , \w[29][11] , 
        \w[29][10] , \w[29][9] , \w[29][8] , \w[29][7] , \w[29][6] , 
        \w[29][5] , \w[29][4] , \w[29][3] , \w[29][2] , \w[29][1] , 1'b0}), 
        .CI(1'b0), .S({\w[30][31] , \w[30][30] , \w[30][29] , \w[30][28] , 
        \w[30][27] , \w[30][26] , \w[30][25] , \w[30][24] , \w[30][23] , 
        \w[30][22] , \w[30][21] , \w[30][20] , \w[30][19] , \w[30][18] , 
        \w[30][17] , \w[30][16] , \w[30][15] , \w[30][14] , \w[30][13] , 
        \w[30][12] , \w[30][11] , \w[30][10] , \w[30][9] , \w[30][8] , 
        \w[30][7] , \w[30][6] , \w[30][5] , \w[30][4] , \w[30][3] , \w[30][2] , 
        \w[30][1] , SYNOPSYS_UNCONNECTED__28}) );
  ADD_N32_191 \FAINST[30].ADD_  ( .A({\_58_net_[31] , \_58_net_[30] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[30][31] , \w[30][30] , 
        \w[30][29] , \w[30][28] , \w[30][27] , \w[30][26] , \w[30][25] , 
        \w[30][24] , \w[30][23] , \w[30][22] , \w[30][21] , \w[30][20] , 
        \w[30][19] , \w[30][18] , \w[30][17] , \w[30][16] , \w[30][15] , 
        \w[30][14] , \w[30][13] , \w[30][12] , \w[30][11] , \w[30][10] , 
        \w[30][9] , \w[30][8] , \w[30][7] , \w[30][6] , \w[30][5] , \w[30][4] , 
        \w[30][3] , \w[30][2] , \w[30][1] , 1'b0}), .CI(1'b0), .S({\w[31][31] , 
        \w[31][30] , \w[31][29] , \w[31][28] , \w[31][27] , \w[31][26] , 
        \w[31][25] , \w[31][24] , \w[31][23] , \w[31][22] , \w[31][21] , 
        \w[31][20] , \w[31][19] , \w[31][18] , \w[31][17] , \w[31][16] , 
        \w[31][15] , \w[31][14] , \w[31][13] , \w[31][12] , \w[31][11] , 
        \w[31][10] , \w[31][9] , \w[31][8] , \w[31][7] , \w[31][6] , 
        \w[31][5] , \w[31][4] , \w[31][3] , \w[31][2] , \w[31][1] , 
        SYNOPSYS_UNCONNECTED__29}) );
  ADD_N32_190 \FAINST[31].ADD_  ( .A({\_60_net_[31] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({\w[31][31] , \w[31][30] , \w[31][29] , 
        \w[31][28] , \w[31][27] , \w[31][26] , \w[31][25] , \w[31][24] , 
        \w[31][23] , \w[31][22] , \w[31][21] , \w[31][20] , \w[31][19] , 
        \w[31][18] , \w[31][17] , \w[31][16] , \w[31][15] , \w[31][14] , 
        \w[31][13] , \w[31][12] , \w[31][11] , \w[31][10] , \w[31][9] , 
        \w[31][8] , \w[31][7] , \w[31][6] , \w[31][5] , \w[31][4] , \w[31][3] , 
        \w[31][2] , \w[31][1] , 1'b0}), .CI(1'b0), .S({O[31:1], 
        SYNOPSYS_UNCONNECTED__30}) );
  AND U2 ( .A(A[5]), .B(B[4]), .Z(\_8_net_[9] ) );
  AND U3 ( .A(A[5]), .B(B[3]), .Z(\_8_net_[8] ) );
  AND U4 ( .A(A[5]), .B(B[2]), .Z(\_8_net_[7] ) );
  AND U5 ( .A(A[5]), .B(B[1]), .Z(\_8_net_[6] ) );
  AND U6 ( .A(A[5]), .B(B[0]), .Z(\_8_net_[5] ) );
  AND U7 ( .A(A[5]), .B(B[26]), .Z(\_8_net_[31] ) );
  AND U8 ( .A(A[5]), .B(B[25]), .Z(\_8_net_[30] ) );
  AND U9 ( .A(A[5]), .B(B[24]), .Z(\_8_net_[29] ) );
  AND U10 ( .A(A[5]), .B(B[23]), .Z(\_8_net_[28] ) );
  AND U11 ( .A(A[5]), .B(B[22]), .Z(\_8_net_[27] ) );
  AND U12 ( .A(A[5]), .B(B[21]), .Z(\_8_net_[26] ) );
  AND U13 ( .A(A[5]), .B(B[20]), .Z(\_8_net_[25] ) );
  AND U14 ( .A(A[5]), .B(B[19]), .Z(\_8_net_[24] ) );
  AND U15 ( .A(A[5]), .B(B[18]), .Z(\_8_net_[23] ) );
  AND U16 ( .A(A[5]), .B(B[17]), .Z(\_8_net_[22] ) );
  AND U17 ( .A(A[5]), .B(B[16]), .Z(\_8_net_[21] ) );
  AND U18 ( .A(A[5]), .B(B[15]), .Z(\_8_net_[20] ) );
  AND U19 ( .A(A[5]), .B(B[14]), .Z(\_8_net_[19] ) );
  AND U20 ( .A(A[5]), .B(B[13]), .Z(\_8_net_[18] ) );
  AND U21 ( .A(A[5]), .B(B[12]), .Z(\_8_net_[17] ) );
  AND U22 ( .A(A[5]), .B(B[11]), .Z(\_8_net_[16] ) );
  AND U23 ( .A(A[5]), .B(B[10]), .Z(\_8_net_[15] ) );
  AND U24 ( .A(A[5]), .B(B[9]), .Z(\_8_net_[14] ) );
  AND U25 ( .A(A[5]), .B(B[8]), .Z(\_8_net_[13] ) );
  AND U26 ( .A(A[5]), .B(B[7]), .Z(\_8_net_[12] ) );
  AND U27 ( .A(A[5]), .B(B[6]), .Z(\_8_net_[11] ) );
  AND U28 ( .A(A[5]), .B(B[5]), .Z(\_8_net_[10] ) );
  AND U29 ( .A(B[5]), .B(A[4]), .Z(\_6_net_[9] ) );
  AND U30 ( .A(B[4]), .B(A[4]), .Z(\_6_net_[8] ) );
  AND U31 ( .A(B[3]), .B(A[4]), .Z(\_6_net_[7] ) );
  AND U32 ( .A(B[2]), .B(A[4]), .Z(\_6_net_[6] ) );
  AND U33 ( .A(B[1]), .B(A[4]), .Z(\_6_net_[5] ) );
  AND U34 ( .A(B[0]), .B(A[4]), .Z(\_6_net_[4] ) );
  AND U35 ( .A(A[4]), .B(B[27]), .Z(\_6_net_[31] ) );
  AND U36 ( .A(B[26]), .B(A[4]), .Z(\_6_net_[30] ) );
  AND U37 ( .A(B[25]), .B(A[4]), .Z(\_6_net_[29] ) );
  AND U38 ( .A(B[24]), .B(A[4]), .Z(\_6_net_[28] ) );
  AND U39 ( .A(B[23]), .B(A[4]), .Z(\_6_net_[27] ) );
  AND U40 ( .A(B[22]), .B(A[4]), .Z(\_6_net_[26] ) );
  AND U41 ( .A(B[21]), .B(A[4]), .Z(\_6_net_[25] ) );
  AND U42 ( .A(B[20]), .B(A[4]), .Z(\_6_net_[24] ) );
  AND U43 ( .A(B[19]), .B(A[4]), .Z(\_6_net_[23] ) );
  AND U44 ( .A(B[18]), .B(A[4]), .Z(\_6_net_[22] ) );
  AND U45 ( .A(B[17]), .B(A[4]), .Z(\_6_net_[21] ) );
  AND U46 ( .A(B[16]), .B(A[4]), .Z(\_6_net_[20] ) );
  AND U47 ( .A(B[15]), .B(A[4]), .Z(\_6_net_[19] ) );
  AND U48 ( .A(B[14]), .B(A[4]), .Z(\_6_net_[18] ) );
  AND U49 ( .A(B[13]), .B(A[4]), .Z(\_6_net_[17] ) );
  AND U50 ( .A(B[12]), .B(A[4]), .Z(\_6_net_[16] ) );
  AND U51 ( .A(B[11]), .B(A[4]), .Z(\_6_net_[15] ) );
  AND U52 ( .A(B[10]), .B(A[4]), .Z(\_6_net_[14] ) );
  AND U53 ( .A(B[9]), .B(A[4]), .Z(\_6_net_[13] ) );
  AND U54 ( .A(B[8]), .B(A[4]), .Z(\_6_net_[12] ) );
  AND U55 ( .A(B[7]), .B(A[4]), .Z(\_6_net_[11] ) );
  AND U56 ( .A(B[6]), .B(A[4]), .Z(\_6_net_[10] ) );
  AND U57 ( .A(A[31]), .B(B[0]), .Z(\_60_net_[31] ) );
  AND U58 ( .A(B[1]), .B(A[30]), .Z(\_58_net_[31] ) );
  AND U59 ( .A(A[30]), .B(B[0]), .Z(\_58_net_[30] ) );
  AND U60 ( .A(B[2]), .B(A[29]), .Z(\_56_net_[31] ) );
  AND U61 ( .A(B[1]), .B(A[29]), .Z(\_56_net_[30] ) );
  AND U62 ( .A(A[29]), .B(B[0]), .Z(\_56_net_[29] ) );
  AND U63 ( .A(B[3]), .B(A[28]), .Z(\_54_net_[31] ) );
  AND U64 ( .A(B[2]), .B(A[28]), .Z(\_54_net_[30] ) );
  AND U65 ( .A(B[1]), .B(A[28]), .Z(\_54_net_[29] ) );
  AND U66 ( .A(A[28]), .B(B[0]), .Z(\_54_net_[28] ) );
  AND U67 ( .A(B[4]), .B(A[27]), .Z(\_52_net_[31] ) );
  AND U68 ( .A(B[3]), .B(A[27]), .Z(\_52_net_[30] ) );
  AND U69 ( .A(B[2]), .B(A[27]), .Z(\_52_net_[29] ) );
  AND U70 ( .A(B[1]), .B(A[27]), .Z(\_52_net_[28] ) );
  AND U71 ( .A(A[27]), .B(B[0]), .Z(\_52_net_[27] ) );
  AND U72 ( .A(B[5]), .B(A[26]), .Z(\_50_net_[31] ) );
  AND U73 ( .A(B[4]), .B(A[26]), .Z(\_50_net_[30] ) );
  AND U74 ( .A(B[3]), .B(A[26]), .Z(\_50_net_[29] ) );
  AND U75 ( .A(B[2]), .B(A[26]), .Z(\_50_net_[28] ) );
  AND U76 ( .A(B[1]), .B(A[26]), .Z(\_50_net_[27] ) );
  AND U77 ( .A(A[26]), .B(B[0]), .Z(\_50_net_[26] ) );
  AND U78 ( .A(B[6]), .B(A[3]), .Z(\_4_net_[9] ) );
  AND U79 ( .A(B[5]), .B(A[3]), .Z(\_4_net_[8] ) );
  AND U80 ( .A(B[4]), .B(A[3]), .Z(\_4_net_[7] ) );
  AND U81 ( .A(B[3]), .B(A[3]), .Z(\_4_net_[6] ) );
  AND U82 ( .A(B[2]), .B(A[3]), .Z(\_4_net_[5] ) );
  AND U83 ( .A(B[1]), .B(A[3]), .Z(\_4_net_[4] ) );
  AND U84 ( .A(B[0]), .B(A[3]), .Z(\_4_net_[3] ) );
  AND U85 ( .A(A[3]), .B(B[28]), .Z(\_4_net_[31] ) );
  AND U86 ( .A(B[27]), .B(A[3]), .Z(\_4_net_[30] ) );
  AND U87 ( .A(B[26]), .B(A[3]), .Z(\_4_net_[29] ) );
  AND U88 ( .A(B[25]), .B(A[3]), .Z(\_4_net_[28] ) );
  AND U89 ( .A(B[24]), .B(A[3]), .Z(\_4_net_[27] ) );
  AND U90 ( .A(B[23]), .B(A[3]), .Z(\_4_net_[26] ) );
  AND U91 ( .A(B[22]), .B(A[3]), .Z(\_4_net_[25] ) );
  AND U92 ( .A(B[21]), .B(A[3]), .Z(\_4_net_[24] ) );
  AND U93 ( .A(B[20]), .B(A[3]), .Z(\_4_net_[23] ) );
  AND U94 ( .A(B[19]), .B(A[3]), .Z(\_4_net_[22] ) );
  AND U95 ( .A(B[18]), .B(A[3]), .Z(\_4_net_[21] ) );
  AND U96 ( .A(B[17]), .B(A[3]), .Z(\_4_net_[20] ) );
  AND U97 ( .A(B[16]), .B(A[3]), .Z(\_4_net_[19] ) );
  AND U98 ( .A(B[15]), .B(A[3]), .Z(\_4_net_[18] ) );
  AND U99 ( .A(B[14]), .B(A[3]), .Z(\_4_net_[17] ) );
  AND U100 ( .A(B[13]), .B(A[3]), .Z(\_4_net_[16] ) );
  AND U101 ( .A(B[12]), .B(A[3]), .Z(\_4_net_[15] ) );
  AND U102 ( .A(B[11]), .B(A[3]), .Z(\_4_net_[14] ) );
  AND U103 ( .A(B[10]), .B(A[3]), .Z(\_4_net_[13] ) );
  AND U104 ( .A(B[9]), .B(A[3]), .Z(\_4_net_[12] ) );
  AND U105 ( .A(B[8]), .B(A[3]), .Z(\_4_net_[11] ) );
  AND U106 ( .A(B[7]), .B(A[3]), .Z(\_4_net_[10] ) );
  AND U107 ( .A(B[6]), .B(A[25]), .Z(\_48_net_[31] ) );
  AND U108 ( .A(B[5]), .B(A[25]), .Z(\_48_net_[30] ) );
  AND U109 ( .A(B[4]), .B(A[25]), .Z(\_48_net_[29] ) );
  AND U110 ( .A(B[3]), .B(A[25]), .Z(\_48_net_[28] ) );
  AND U111 ( .A(B[2]), .B(A[25]), .Z(\_48_net_[27] ) );
  AND U112 ( .A(B[1]), .B(A[25]), .Z(\_48_net_[26] ) );
  AND U113 ( .A(A[25]), .B(B[0]), .Z(\_48_net_[25] ) );
  AND U114 ( .A(B[7]), .B(A[24]), .Z(\_46_net_[31] ) );
  AND U115 ( .A(B[6]), .B(A[24]), .Z(\_46_net_[30] ) );
  AND U116 ( .A(B[5]), .B(A[24]), .Z(\_46_net_[29] ) );
  AND U117 ( .A(B[4]), .B(A[24]), .Z(\_46_net_[28] ) );
  AND U118 ( .A(B[3]), .B(A[24]), .Z(\_46_net_[27] ) );
  AND U119 ( .A(B[2]), .B(A[24]), .Z(\_46_net_[26] ) );
  AND U120 ( .A(B[1]), .B(A[24]), .Z(\_46_net_[25] ) );
  AND U121 ( .A(A[24]), .B(B[0]), .Z(\_46_net_[24] ) );
  AND U122 ( .A(B[8]), .B(A[23]), .Z(\_44_net_[31] ) );
  AND U123 ( .A(B[7]), .B(A[23]), .Z(\_44_net_[30] ) );
  AND U124 ( .A(B[6]), .B(A[23]), .Z(\_44_net_[29] ) );
  AND U125 ( .A(B[5]), .B(A[23]), .Z(\_44_net_[28] ) );
  AND U126 ( .A(B[4]), .B(A[23]), .Z(\_44_net_[27] ) );
  AND U127 ( .A(B[3]), .B(A[23]), .Z(\_44_net_[26] ) );
  AND U128 ( .A(B[2]), .B(A[23]), .Z(\_44_net_[25] ) );
  AND U129 ( .A(B[1]), .B(A[23]), .Z(\_44_net_[24] ) );
  AND U130 ( .A(A[23]), .B(B[0]), .Z(\_44_net_[23] ) );
  AND U131 ( .A(B[9]), .B(A[22]), .Z(\_42_net_[31] ) );
  AND U132 ( .A(B[8]), .B(A[22]), .Z(\_42_net_[30] ) );
  AND U133 ( .A(B[7]), .B(A[22]), .Z(\_42_net_[29] ) );
  AND U134 ( .A(B[6]), .B(A[22]), .Z(\_42_net_[28] ) );
  AND U135 ( .A(B[5]), .B(A[22]), .Z(\_42_net_[27] ) );
  AND U136 ( .A(B[4]), .B(A[22]), .Z(\_42_net_[26] ) );
  AND U137 ( .A(B[3]), .B(A[22]), .Z(\_42_net_[25] ) );
  AND U138 ( .A(B[2]), .B(A[22]), .Z(\_42_net_[24] ) );
  AND U139 ( .A(B[1]), .B(A[22]), .Z(\_42_net_[23] ) );
  AND U140 ( .A(A[22]), .B(B[0]), .Z(\_42_net_[22] ) );
  AND U141 ( .A(B[10]), .B(A[21]), .Z(\_40_net_[31] ) );
  AND U142 ( .A(B[9]), .B(A[21]), .Z(\_40_net_[30] ) );
  AND U143 ( .A(B[8]), .B(A[21]), .Z(\_40_net_[29] ) );
  AND U144 ( .A(B[7]), .B(A[21]), .Z(\_40_net_[28] ) );
  AND U145 ( .A(B[6]), .B(A[21]), .Z(\_40_net_[27] ) );
  AND U146 ( .A(B[5]), .B(A[21]), .Z(\_40_net_[26] ) );
  AND U147 ( .A(B[4]), .B(A[21]), .Z(\_40_net_[25] ) );
  AND U148 ( .A(B[3]), .B(A[21]), .Z(\_40_net_[24] ) );
  AND U149 ( .A(B[2]), .B(A[21]), .Z(\_40_net_[23] ) );
  AND U150 ( .A(B[1]), .B(A[21]), .Z(\_40_net_[22] ) );
  AND U151 ( .A(A[21]), .B(B[0]), .Z(\_40_net_[21] ) );
  AND U152 ( .A(B[11]), .B(A[20]), .Z(\_38_net_[31] ) );
  AND U153 ( .A(B[10]), .B(A[20]), .Z(\_38_net_[30] ) );
  AND U154 ( .A(B[9]), .B(A[20]), .Z(\_38_net_[29] ) );
  AND U155 ( .A(B[8]), .B(A[20]), .Z(\_38_net_[28] ) );
  AND U156 ( .A(B[7]), .B(A[20]), .Z(\_38_net_[27] ) );
  AND U157 ( .A(B[6]), .B(A[20]), .Z(\_38_net_[26] ) );
  AND U158 ( .A(B[5]), .B(A[20]), .Z(\_38_net_[25] ) );
  AND U159 ( .A(B[4]), .B(A[20]), .Z(\_38_net_[24] ) );
  AND U160 ( .A(B[3]), .B(A[20]), .Z(\_38_net_[23] ) );
  AND U161 ( .A(B[2]), .B(A[20]), .Z(\_38_net_[22] ) );
  AND U162 ( .A(B[1]), .B(A[20]), .Z(\_38_net_[21] ) );
  AND U163 ( .A(A[20]), .B(B[0]), .Z(\_38_net_[20] ) );
  AND U164 ( .A(B[12]), .B(A[19]), .Z(\_36_net_[31] ) );
  AND U165 ( .A(B[11]), .B(A[19]), .Z(\_36_net_[30] ) );
  AND U166 ( .A(B[10]), .B(A[19]), .Z(\_36_net_[29] ) );
  AND U167 ( .A(B[9]), .B(A[19]), .Z(\_36_net_[28] ) );
  AND U168 ( .A(B[8]), .B(A[19]), .Z(\_36_net_[27] ) );
  AND U169 ( .A(B[7]), .B(A[19]), .Z(\_36_net_[26] ) );
  AND U170 ( .A(B[6]), .B(A[19]), .Z(\_36_net_[25] ) );
  AND U171 ( .A(B[5]), .B(A[19]), .Z(\_36_net_[24] ) );
  AND U172 ( .A(B[4]), .B(A[19]), .Z(\_36_net_[23] ) );
  AND U173 ( .A(B[3]), .B(A[19]), .Z(\_36_net_[22] ) );
  AND U174 ( .A(B[2]), .B(A[19]), .Z(\_36_net_[21] ) );
  AND U175 ( .A(B[1]), .B(A[19]), .Z(\_36_net_[20] ) );
  AND U176 ( .A(A[19]), .B(B[0]), .Z(\_36_net_[19] ) );
  AND U177 ( .A(B[13]), .B(A[18]), .Z(\_34_net_[31] ) );
  AND U178 ( .A(B[12]), .B(A[18]), .Z(\_34_net_[30] ) );
  AND U179 ( .A(B[11]), .B(A[18]), .Z(\_34_net_[29] ) );
  AND U180 ( .A(B[10]), .B(A[18]), .Z(\_34_net_[28] ) );
  AND U181 ( .A(B[9]), .B(A[18]), .Z(\_34_net_[27] ) );
  AND U182 ( .A(B[8]), .B(A[18]), .Z(\_34_net_[26] ) );
  AND U183 ( .A(B[7]), .B(A[18]), .Z(\_34_net_[25] ) );
  AND U184 ( .A(B[6]), .B(A[18]), .Z(\_34_net_[24] ) );
  AND U185 ( .A(B[5]), .B(A[18]), .Z(\_34_net_[23] ) );
  AND U186 ( .A(B[4]), .B(A[18]), .Z(\_34_net_[22] ) );
  AND U187 ( .A(B[3]), .B(A[18]), .Z(\_34_net_[21] ) );
  AND U188 ( .A(B[2]), .B(A[18]), .Z(\_34_net_[20] ) );
  AND U189 ( .A(B[1]), .B(A[18]), .Z(\_34_net_[19] ) );
  AND U190 ( .A(A[18]), .B(B[0]), .Z(\_34_net_[18] ) );
  AND U191 ( .A(B[14]), .B(A[17]), .Z(\_32_net_[31] ) );
  AND U192 ( .A(B[13]), .B(A[17]), .Z(\_32_net_[30] ) );
  AND U193 ( .A(B[12]), .B(A[17]), .Z(\_32_net_[29] ) );
  AND U194 ( .A(B[11]), .B(A[17]), .Z(\_32_net_[28] ) );
  AND U195 ( .A(B[10]), .B(A[17]), .Z(\_32_net_[27] ) );
  AND U196 ( .A(B[9]), .B(A[17]), .Z(\_32_net_[26] ) );
  AND U197 ( .A(B[8]), .B(A[17]), .Z(\_32_net_[25] ) );
  AND U198 ( .A(B[7]), .B(A[17]), .Z(\_32_net_[24] ) );
  AND U199 ( .A(B[6]), .B(A[17]), .Z(\_32_net_[23] ) );
  AND U200 ( .A(B[5]), .B(A[17]), .Z(\_32_net_[22] ) );
  AND U201 ( .A(B[4]), .B(A[17]), .Z(\_32_net_[21] ) );
  AND U202 ( .A(B[3]), .B(A[17]), .Z(\_32_net_[20] ) );
  AND U203 ( .A(B[2]), .B(A[17]), .Z(\_32_net_[19] ) );
  AND U204 ( .A(B[1]), .B(A[17]), .Z(\_32_net_[18] ) );
  AND U205 ( .A(A[17]), .B(B[0]), .Z(\_32_net_[17] ) );
  AND U206 ( .A(B[15]), .B(A[16]), .Z(\_30_net_[31] ) );
  AND U207 ( .A(B[14]), .B(A[16]), .Z(\_30_net_[30] ) );
  AND U208 ( .A(B[13]), .B(A[16]), .Z(\_30_net_[29] ) );
  AND U209 ( .A(B[12]), .B(A[16]), .Z(\_30_net_[28] ) );
  AND U210 ( .A(B[11]), .B(A[16]), .Z(\_30_net_[27] ) );
  AND U211 ( .A(B[10]), .B(A[16]), .Z(\_30_net_[26] ) );
  AND U212 ( .A(B[9]), .B(A[16]), .Z(\_30_net_[25] ) );
  AND U213 ( .A(B[8]), .B(A[16]), .Z(\_30_net_[24] ) );
  AND U214 ( .A(B[7]), .B(A[16]), .Z(\_30_net_[23] ) );
  AND U215 ( .A(B[6]), .B(A[16]), .Z(\_30_net_[22] ) );
  AND U216 ( .A(B[5]), .B(A[16]), .Z(\_30_net_[21] ) );
  AND U217 ( .A(B[4]), .B(A[16]), .Z(\_30_net_[20] ) );
  AND U218 ( .A(B[3]), .B(A[16]), .Z(\_30_net_[19] ) );
  AND U219 ( .A(B[2]), .B(A[16]), .Z(\_30_net_[18] ) );
  AND U220 ( .A(B[1]), .B(A[16]), .Z(\_30_net_[17] ) );
  AND U221 ( .A(A[16]), .B(B[0]), .Z(\_30_net_[16] ) );
  AND U222 ( .A(B[7]), .B(A[2]), .Z(\_2_net_[9] ) );
  AND U223 ( .A(B[6]), .B(A[2]), .Z(\_2_net_[8] ) );
  AND U224 ( .A(B[5]), .B(A[2]), .Z(\_2_net_[7] ) );
  AND U225 ( .A(B[4]), .B(A[2]), .Z(\_2_net_[6] ) );
  AND U226 ( .A(B[3]), .B(A[2]), .Z(\_2_net_[5] ) );
  AND U227 ( .A(B[2]), .B(A[2]), .Z(\_2_net_[4] ) );
  AND U228 ( .A(B[1]), .B(A[2]), .Z(\_2_net_[3] ) );
  AND U229 ( .A(A[2]), .B(B[29]), .Z(\_2_net_[31] ) );
  AND U230 ( .A(B[28]), .B(A[2]), .Z(\_2_net_[30] ) );
  AND U231 ( .A(B[0]), .B(A[2]), .Z(\_2_net_[2] ) );
  AND U232 ( .A(B[27]), .B(A[2]), .Z(\_2_net_[29] ) );
  AND U233 ( .A(B[26]), .B(A[2]), .Z(\_2_net_[28] ) );
  AND U234 ( .A(B[25]), .B(A[2]), .Z(\_2_net_[27] ) );
  AND U235 ( .A(B[24]), .B(A[2]), .Z(\_2_net_[26] ) );
  AND U236 ( .A(B[23]), .B(A[2]), .Z(\_2_net_[25] ) );
  AND U237 ( .A(B[22]), .B(A[2]), .Z(\_2_net_[24] ) );
  AND U238 ( .A(B[21]), .B(A[2]), .Z(\_2_net_[23] ) );
  AND U239 ( .A(B[20]), .B(A[2]), .Z(\_2_net_[22] ) );
  AND U240 ( .A(B[19]), .B(A[2]), .Z(\_2_net_[21] ) );
  AND U241 ( .A(B[18]), .B(A[2]), .Z(\_2_net_[20] ) );
  AND U242 ( .A(B[17]), .B(A[2]), .Z(\_2_net_[19] ) );
  AND U243 ( .A(B[16]), .B(A[2]), .Z(\_2_net_[18] ) );
  AND U244 ( .A(B[15]), .B(A[2]), .Z(\_2_net_[17] ) );
  AND U245 ( .A(B[14]), .B(A[2]), .Z(\_2_net_[16] ) );
  AND U246 ( .A(B[13]), .B(A[2]), .Z(\_2_net_[15] ) );
  AND U247 ( .A(B[12]), .B(A[2]), .Z(\_2_net_[14] ) );
  AND U248 ( .A(B[11]), .B(A[2]), .Z(\_2_net_[13] ) );
  AND U249 ( .A(B[10]), .B(A[2]), .Z(\_2_net_[12] ) );
  AND U250 ( .A(B[9]), .B(A[2]), .Z(\_2_net_[11] ) );
  AND U251 ( .A(B[8]), .B(A[2]), .Z(\_2_net_[10] ) );
  AND U252 ( .A(B[16]), .B(A[15]), .Z(\_28_net_[31] ) );
  AND U253 ( .A(B[15]), .B(A[15]), .Z(\_28_net_[30] ) );
  AND U254 ( .A(B[14]), .B(A[15]), .Z(\_28_net_[29] ) );
  AND U255 ( .A(B[13]), .B(A[15]), .Z(\_28_net_[28] ) );
  AND U256 ( .A(B[12]), .B(A[15]), .Z(\_28_net_[27] ) );
  AND U257 ( .A(B[11]), .B(A[15]), .Z(\_28_net_[26] ) );
  AND U258 ( .A(B[10]), .B(A[15]), .Z(\_28_net_[25] ) );
  AND U259 ( .A(B[9]), .B(A[15]), .Z(\_28_net_[24] ) );
  AND U260 ( .A(B[8]), .B(A[15]), .Z(\_28_net_[23] ) );
  AND U261 ( .A(B[7]), .B(A[15]), .Z(\_28_net_[22] ) );
  AND U262 ( .A(B[6]), .B(A[15]), .Z(\_28_net_[21] ) );
  AND U263 ( .A(B[5]), .B(A[15]), .Z(\_28_net_[20] ) );
  AND U264 ( .A(B[4]), .B(A[15]), .Z(\_28_net_[19] ) );
  AND U265 ( .A(B[3]), .B(A[15]), .Z(\_28_net_[18] ) );
  AND U266 ( .A(B[2]), .B(A[15]), .Z(\_28_net_[17] ) );
  AND U267 ( .A(B[1]), .B(A[15]), .Z(\_28_net_[16] ) );
  AND U268 ( .A(A[15]), .B(B[0]), .Z(\_28_net_[15] ) );
  AND U269 ( .A(B[17]), .B(A[14]), .Z(\_26_net_[31] ) );
  AND U270 ( .A(B[16]), .B(A[14]), .Z(\_26_net_[30] ) );
  AND U271 ( .A(B[15]), .B(A[14]), .Z(\_26_net_[29] ) );
  AND U272 ( .A(B[14]), .B(A[14]), .Z(\_26_net_[28] ) );
  AND U273 ( .A(B[13]), .B(A[14]), .Z(\_26_net_[27] ) );
  AND U274 ( .A(B[12]), .B(A[14]), .Z(\_26_net_[26] ) );
  AND U275 ( .A(B[11]), .B(A[14]), .Z(\_26_net_[25] ) );
  AND U276 ( .A(B[10]), .B(A[14]), .Z(\_26_net_[24] ) );
  AND U277 ( .A(B[9]), .B(A[14]), .Z(\_26_net_[23] ) );
  AND U278 ( .A(B[8]), .B(A[14]), .Z(\_26_net_[22] ) );
  AND U279 ( .A(B[7]), .B(A[14]), .Z(\_26_net_[21] ) );
  AND U280 ( .A(B[6]), .B(A[14]), .Z(\_26_net_[20] ) );
  AND U281 ( .A(B[5]), .B(A[14]), .Z(\_26_net_[19] ) );
  AND U282 ( .A(B[4]), .B(A[14]), .Z(\_26_net_[18] ) );
  AND U283 ( .A(B[3]), .B(A[14]), .Z(\_26_net_[17] ) );
  AND U284 ( .A(B[2]), .B(A[14]), .Z(\_26_net_[16] ) );
  AND U285 ( .A(B[1]), .B(A[14]), .Z(\_26_net_[15] ) );
  AND U286 ( .A(A[14]), .B(B[0]), .Z(\_26_net_[14] ) );
  AND U287 ( .A(B[18]), .B(A[13]), .Z(\_24_net_[31] ) );
  AND U288 ( .A(B[17]), .B(A[13]), .Z(\_24_net_[30] ) );
  AND U289 ( .A(B[16]), .B(A[13]), .Z(\_24_net_[29] ) );
  AND U290 ( .A(B[15]), .B(A[13]), .Z(\_24_net_[28] ) );
  AND U291 ( .A(B[14]), .B(A[13]), .Z(\_24_net_[27] ) );
  AND U292 ( .A(B[13]), .B(A[13]), .Z(\_24_net_[26] ) );
  AND U293 ( .A(B[12]), .B(A[13]), .Z(\_24_net_[25] ) );
  AND U294 ( .A(B[11]), .B(A[13]), .Z(\_24_net_[24] ) );
  AND U295 ( .A(B[10]), .B(A[13]), .Z(\_24_net_[23] ) );
  AND U296 ( .A(B[9]), .B(A[13]), .Z(\_24_net_[22] ) );
  AND U297 ( .A(B[8]), .B(A[13]), .Z(\_24_net_[21] ) );
  AND U298 ( .A(B[7]), .B(A[13]), .Z(\_24_net_[20] ) );
  AND U299 ( .A(B[6]), .B(A[13]), .Z(\_24_net_[19] ) );
  AND U300 ( .A(B[5]), .B(A[13]), .Z(\_24_net_[18] ) );
  AND U301 ( .A(B[4]), .B(A[13]), .Z(\_24_net_[17] ) );
  AND U302 ( .A(B[3]), .B(A[13]), .Z(\_24_net_[16] ) );
  AND U303 ( .A(B[2]), .B(A[13]), .Z(\_24_net_[15] ) );
  AND U304 ( .A(B[1]), .B(A[13]), .Z(\_24_net_[14] ) );
  AND U305 ( .A(A[13]), .B(B[0]), .Z(\_24_net_[13] ) );
  AND U306 ( .A(B[19]), .B(A[12]), .Z(\_22_net_[31] ) );
  AND U307 ( .A(B[18]), .B(A[12]), .Z(\_22_net_[30] ) );
  AND U308 ( .A(B[17]), .B(A[12]), .Z(\_22_net_[29] ) );
  AND U309 ( .A(B[16]), .B(A[12]), .Z(\_22_net_[28] ) );
  AND U310 ( .A(B[15]), .B(A[12]), .Z(\_22_net_[27] ) );
  AND U311 ( .A(B[14]), .B(A[12]), .Z(\_22_net_[26] ) );
  AND U312 ( .A(B[13]), .B(A[12]), .Z(\_22_net_[25] ) );
  AND U313 ( .A(B[12]), .B(A[12]), .Z(\_22_net_[24] ) );
  AND U314 ( .A(B[11]), .B(A[12]), .Z(\_22_net_[23] ) );
  AND U315 ( .A(B[10]), .B(A[12]), .Z(\_22_net_[22] ) );
  AND U316 ( .A(B[9]), .B(A[12]), .Z(\_22_net_[21] ) );
  AND U317 ( .A(B[8]), .B(A[12]), .Z(\_22_net_[20] ) );
  AND U318 ( .A(B[7]), .B(A[12]), .Z(\_22_net_[19] ) );
  AND U319 ( .A(B[6]), .B(A[12]), .Z(\_22_net_[18] ) );
  AND U320 ( .A(B[5]), .B(A[12]), .Z(\_22_net_[17] ) );
  AND U321 ( .A(B[4]), .B(A[12]), .Z(\_22_net_[16] ) );
  AND U322 ( .A(B[3]), .B(A[12]), .Z(\_22_net_[15] ) );
  AND U323 ( .A(B[2]), .B(A[12]), .Z(\_22_net_[14] ) );
  AND U324 ( .A(B[1]), .B(A[12]), .Z(\_22_net_[13] ) );
  AND U325 ( .A(A[12]), .B(B[0]), .Z(\_22_net_[12] ) );
  AND U326 ( .A(B[20]), .B(A[11]), .Z(\_20_net_[31] ) );
  AND U327 ( .A(B[19]), .B(A[11]), .Z(\_20_net_[30] ) );
  AND U328 ( .A(B[18]), .B(A[11]), .Z(\_20_net_[29] ) );
  AND U329 ( .A(B[17]), .B(A[11]), .Z(\_20_net_[28] ) );
  AND U330 ( .A(B[16]), .B(A[11]), .Z(\_20_net_[27] ) );
  AND U331 ( .A(B[15]), .B(A[11]), .Z(\_20_net_[26] ) );
  AND U332 ( .A(B[14]), .B(A[11]), .Z(\_20_net_[25] ) );
  AND U333 ( .A(B[13]), .B(A[11]), .Z(\_20_net_[24] ) );
  AND U334 ( .A(B[12]), .B(A[11]), .Z(\_20_net_[23] ) );
  AND U335 ( .A(B[11]), .B(A[11]), .Z(\_20_net_[22] ) );
  AND U336 ( .A(B[10]), .B(A[11]), .Z(\_20_net_[21] ) );
  AND U337 ( .A(B[9]), .B(A[11]), .Z(\_20_net_[20] ) );
  AND U338 ( .A(B[8]), .B(A[11]), .Z(\_20_net_[19] ) );
  AND U339 ( .A(B[7]), .B(A[11]), .Z(\_20_net_[18] ) );
  AND U340 ( .A(B[6]), .B(A[11]), .Z(\_20_net_[17] ) );
  AND U341 ( .A(B[5]), .B(A[11]), .Z(\_20_net_[16] ) );
  AND U342 ( .A(B[4]), .B(A[11]), .Z(\_20_net_[15] ) );
  AND U343 ( .A(B[3]), .B(A[11]), .Z(\_20_net_[14] ) );
  AND U344 ( .A(B[2]), .B(A[11]), .Z(\_20_net_[13] ) );
  AND U345 ( .A(B[1]), .B(A[11]), .Z(\_20_net_[12] ) );
  AND U346 ( .A(A[11]), .B(B[0]), .Z(\_20_net_[11] ) );
  AND U347 ( .A(B[21]), .B(A[10]), .Z(\_18_net_[31] ) );
  AND U348 ( .A(B[20]), .B(A[10]), .Z(\_18_net_[30] ) );
  AND U349 ( .A(B[19]), .B(A[10]), .Z(\_18_net_[29] ) );
  AND U350 ( .A(B[18]), .B(A[10]), .Z(\_18_net_[28] ) );
  AND U351 ( .A(B[17]), .B(A[10]), .Z(\_18_net_[27] ) );
  AND U352 ( .A(B[16]), .B(A[10]), .Z(\_18_net_[26] ) );
  AND U353 ( .A(B[15]), .B(A[10]), .Z(\_18_net_[25] ) );
  AND U354 ( .A(B[14]), .B(A[10]), .Z(\_18_net_[24] ) );
  AND U355 ( .A(B[13]), .B(A[10]), .Z(\_18_net_[23] ) );
  AND U356 ( .A(B[12]), .B(A[10]), .Z(\_18_net_[22] ) );
  AND U357 ( .A(B[11]), .B(A[10]), .Z(\_18_net_[21] ) );
  AND U358 ( .A(B[10]), .B(A[10]), .Z(\_18_net_[20] ) );
  AND U359 ( .A(B[9]), .B(A[10]), .Z(\_18_net_[19] ) );
  AND U360 ( .A(B[8]), .B(A[10]), .Z(\_18_net_[18] ) );
  AND U361 ( .A(B[7]), .B(A[10]), .Z(\_18_net_[17] ) );
  AND U362 ( .A(B[6]), .B(A[10]), .Z(\_18_net_[16] ) );
  AND U363 ( .A(B[5]), .B(A[10]), .Z(\_18_net_[15] ) );
  AND U364 ( .A(B[4]), .B(A[10]), .Z(\_18_net_[14] ) );
  AND U365 ( .A(B[3]), .B(A[10]), .Z(\_18_net_[13] ) );
  AND U366 ( .A(B[2]), .B(A[10]), .Z(\_18_net_[12] ) );
  AND U367 ( .A(B[1]), .B(A[10]), .Z(\_18_net_[11] ) );
  AND U368 ( .A(A[10]), .B(B[0]), .Z(\_18_net_[10] ) );
  AND U369 ( .A(B[0]), .B(A[9]), .Z(\_16_net_[9] ) );
  AND U370 ( .A(B[22]), .B(A[9]), .Z(\_16_net_[31] ) );
  AND U371 ( .A(B[21]), .B(A[9]), .Z(\_16_net_[30] ) );
  AND U372 ( .A(B[20]), .B(A[9]), .Z(\_16_net_[29] ) );
  AND U373 ( .A(B[19]), .B(A[9]), .Z(\_16_net_[28] ) );
  AND U374 ( .A(B[18]), .B(A[9]), .Z(\_16_net_[27] ) );
  AND U375 ( .A(B[17]), .B(A[9]), .Z(\_16_net_[26] ) );
  AND U376 ( .A(B[16]), .B(A[9]), .Z(\_16_net_[25] ) );
  AND U377 ( .A(B[15]), .B(A[9]), .Z(\_16_net_[24] ) );
  AND U378 ( .A(B[14]), .B(A[9]), .Z(\_16_net_[23] ) );
  AND U379 ( .A(B[13]), .B(A[9]), .Z(\_16_net_[22] ) );
  AND U380 ( .A(B[12]), .B(A[9]), .Z(\_16_net_[21] ) );
  AND U381 ( .A(B[11]), .B(A[9]), .Z(\_16_net_[20] ) );
  AND U382 ( .A(B[10]), .B(A[9]), .Z(\_16_net_[19] ) );
  AND U383 ( .A(B[9]), .B(A[9]), .Z(\_16_net_[18] ) );
  AND U384 ( .A(B[8]), .B(A[9]), .Z(\_16_net_[17] ) );
  AND U385 ( .A(B[7]), .B(A[9]), .Z(\_16_net_[16] ) );
  AND U386 ( .A(B[6]), .B(A[9]), .Z(\_16_net_[15] ) );
  AND U387 ( .A(B[5]), .B(A[9]), .Z(\_16_net_[14] ) );
  AND U388 ( .A(B[4]), .B(A[9]), .Z(\_16_net_[13] ) );
  AND U389 ( .A(B[3]), .B(A[9]), .Z(\_16_net_[12] ) );
  AND U390 ( .A(B[2]), .B(A[9]), .Z(\_16_net_[11] ) );
  AND U391 ( .A(A[9]), .B(B[1]), .Z(\_16_net_[10] ) );
  AND U392 ( .A(B[1]), .B(A[8]), .Z(\_14_net_[9] ) );
  AND U393 ( .A(B[0]), .B(A[8]), .Z(\_14_net_[8] ) );
  AND U394 ( .A(B[23]), .B(A[8]), .Z(\_14_net_[31] ) );
  AND U395 ( .A(B[22]), .B(A[8]), .Z(\_14_net_[30] ) );
  AND U396 ( .A(B[21]), .B(A[8]), .Z(\_14_net_[29] ) );
  AND U397 ( .A(B[20]), .B(A[8]), .Z(\_14_net_[28] ) );
  AND U398 ( .A(B[19]), .B(A[8]), .Z(\_14_net_[27] ) );
  AND U399 ( .A(B[18]), .B(A[8]), .Z(\_14_net_[26] ) );
  AND U400 ( .A(B[17]), .B(A[8]), .Z(\_14_net_[25] ) );
  AND U401 ( .A(B[16]), .B(A[8]), .Z(\_14_net_[24] ) );
  AND U402 ( .A(B[15]), .B(A[8]), .Z(\_14_net_[23] ) );
  AND U403 ( .A(B[14]), .B(A[8]), .Z(\_14_net_[22] ) );
  AND U404 ( .A(B[13]), .B(A[8]), .Z(\_14_net_[21] ) );
  AND U405 ( .A(B[12]), .B(A[8]), .Z(\_14_net_[20] ) );
  AND U406 ( .A(B[11]), .B(A[8]), .Z(\_14_net_[19] ) );
  AND U407 ( .A(B[10]), .B(A[8]), .Z(\_14_net_[18] ) );
  AND U408 ( .A(B[9]), .B(A[8]), .Z(\_14_net_[17] ) );
  AND U409 ( .A(B[8]), .B(A[8]), .Z(\_14_net_[16] ) );
  AND U410 ( .A(B[7]), .B(A[8]), .Z(\_14_net_[15] ) );
  AND U411 ( .A(B[6]), .B(A[8]), .Z(\_14_net_[14] ) );
  AND U412 ( .A(B[5]), .B(A[8]), .Z(\_14_net_[13] ) );
  AND U413 ( .A(B[4]), .B(A[8]), .Z(\_14_net_[12] ) );
  AND U414 ( .A(B[3]), .B(A[8]), .Z(\_14_net_[11] ) );
  AND U415 ( .A(A[8]), .B(B[2]), .Z(\_14_net_[10] ) );
  AND U416 ( .A(B[2]), .B(A[7]), .Z(\_12_net_[9] ) );
  AND U417 ( .A(B[1]), .B(A[7]), .Z(\_12_net_[8] ) );
  AND U418 ( .A(B[0]), .B(A[7]), .Z(\_12_net_[7] ) );
  AND U419 ( .A(B[24]), .B(A[7]), .Z(\_12_net_[31] ) );
  AND U420 ( .A(B[23]), .B(A[7]), .Z(\_12_net_[30] ) );
  AND U421 ( .A(B[22]), .B(A[7]), .Z(\_12_net_[29] ) );
  AND U422 ( .A(B[21]), .B(A[7]), .Z(\_12_net_[28] ) );
  AND U423 ( .A(B[20]), .B(A[7]), .Z(\_12_net_[27] ) );
  AND U424 ( .A(B[19]), .B(A[7]), .Z(\_12_net_[26] ) );
  AND U425 ( .A(B[18]), .B(A[7]), .Z(\_12_net_[25] ) );
  AND U426 ( .A(B[17]), .B(A[7]), .Z(\_12_net_[24] ) );
  AND U427 ( .A(B[16]), .B(A[7]), .Z(\_12_net_[23] ) );
  AND U428 ( .A(B[15]), .B(A[7]), .Z(\_12_net_[22] ) );
  AND U429 ( .A(B[14]), .B(A[7]), .Z(\_12_net_[21] ) );
  AND U430 ( .A(B[13]), .B(A[7]), .Z(\_12_net_[20] ) );
  AND U431 ( .A(B[12]), .B(A[7]), .Z(\_12_net_[19] ) );
  AND U432 ( .A(B[11]), .B(A[7]), .Z(\_12_net_[18] ) );
  AND U433 ( .A(B[10]), .B(A[7]), .Z(\_12_net_[17] ) );
  AND U434 ( .A(B[9]), .B(A[7]), .Z(\_12_net_[16] ) );
  AND U435 ( .A(B[8]), .B(A[7]), .Z(\_12_net_[15] ) );
  AND U436 ( .A(B[7]), .B(A[7]), .Z(\_12_net_[14] ) );
  AND U437 ( .A(B[6]), .B(A[7]), .Z(\_12_net_[13] ) );
  AND U438 ( .A(B[5]), .B(A[7]), .Z(\_12_net_[12] ) );
  AND U439 ( .A(B[4]), .B(A[7]), .Z(\_12_net_[11] ) );
  AND U440 ( .A(A[7]), .B(B[3]), .Z(\_12_net_[10] ) );
  AND U441 ( .A(B[3]), .B(A[6]), .Z(\_10_net_[9] ) );
  AND U442 ( .A(B[2]), .B(A[6]), .Z(\_10_net_[8] ) );
  AND U443 ( .A(B[1]), .B(A[6]), .Z(\_10_net_[7] ) );
  AND U444 ( .A(B[0]), .B(A[6]), .Z(\_10_net_[6] ) );
  AND U445 ( .A(B[25]), .B(A[6]), .Z(\_10_net_[31] ) );
  AND U446 ( .A(B[24]), .B(A[6]), .Z(\_10_net_[30] ) );
  AND U447 ( .A(B[23]), .B(A[6]), .Z(\_10_net_[29] ) );
  AND U448 ( .A(B[22]), .B(A[6]), .Z(\_10_net_[28] ) );
  AND U449 ( .A(B[21]), .B(A[6]), .Z(\_10_net_[27] ) );
  AND U450 ( .A(B[20]), .B(A[6]), .Z(\_10_net_[26] ) );
  AND U451 ( .A(B[19]), .B(A[6]), .Z(\_10_net_[25] ) );
  AND U452 ( .A(B[18]), .B(A[6]), .Z(\_10_net_[24] ) );
  AND U453 ( .A(B[17]), .B(A[6]), .Z(\_10_net_[23] ) );
  AND U454 ( .A(B[16]), .B(A[6]), .Z(\_10_net_[22] ) );
  AND U455 ( .A(B[15]), .B(A[6]), .Z(\_10_net_[21] ) );
  AND U456 ( .A(B[14]), .B(A[6]), .Z(\_10_net_[20] ) );
  AND U457 ( .A(B[13]), .B(A[6]), .Z(\_10_net_[19] ) );
  AND U458 ( .A(B[12]), .B(A[6]), .Z(\_10_net_[18] ) );
  AND U459 ( .A(B[11]), .B(A[6]), .Z(\_10_net_[17] ) );
  AND U460 ( .A(B[10]), .B(A[6]), .Z(\_10_net_[16] ) );
  AND U461 ( .A(B[9]), .B(A[6]), .Z(\_10_net_[15] ) );
  AND U462 ( .A(B[8]), .B(A[6]), .Z(\_10_net_[14] ) );
  AND U463 ( .A(B[7]), .B(A[6]), .Z(\_10_net_[13] ) );
  AND U464 ( .A(B[6]), .B(A[6]), .Z(\_10_net_[12] ) );
  AND U465 ( .A(B[5]), .B(A[6]), .Z(\_10_net_[11] ) );
  AND U466 ( .A(A[6]), .B(B[4]), .Z(\_10_net_[10] ) );
  AND U467 ( .A(B[8]), .B(A[1]), .Z(\_0_net_[9] ) );
  AND U468 ( .A(B[7]), .B(A[1]), .Z(\_0_net_[8] ) );
  AND U469 ( .A(B[6]), .B(A[1]), .Z(\_0_net_[7] ) );
  AND U470 ( .A(B[5]), .B(A[1]), .Z(\_0_net_[6] ) );
  AND U471 ( .A(B[4]), .B(A[1]), .Z(\_0_net_[5] ) );
  AND U472 ( .A(B[3]), .B(A[1]), .Z(\_0_net_[4] ) );
  AND U473 ( .A(B[2]), .B(A[1]), .Z(\_0_net_[3] ) );
  AND U474 ( .A(B[30]), .B(A[1]), .Z(\_0_net_[31] ) );
  AND U475 ( .A(B[29]), .B(A[1]), .Z(\_0_net_[30] ) );
  AND U476 ( .A(B[1]), .B(A[1]), .Z(\_0_net_[2] ) );
  AND U477 ( .A(B[28]), .B(A[1]), .Z(\_0_net_[29] ) );
  AND U478 ( .A(B[27]), .B(A[1]), .Z(\_0_net_[28] ) );
  AND U479 ( .A(B[26]), .B(A[1]), .Z(\_0_net_[27] ) );
  AND U480 ( .A(B[25]), .B(A[1]), .Z(\_0_net_[26] ) );
  AND U481 ( .A(B[24]), .B(A[1]), .Z(\_0_net_[25] ) );
  AND U482 ( .A(B[23]), .B(A[1]), .Z(\_0_net_[24] ) );
  AND U483 ( .A(B[22]), .B(A[1]), .Z(\_0_net_[23] ) );
  AND U484 ( .A(B[21]), .B(A[1]), .Z(\_0_net_[22] ) );
  AND U485 ( .A(B[20]), .B(A[1]), .Z(\_0_net_[21] ) );
  AND U486 ( .A(B[19]), .B(A[1]), .Z(\_0_net_[20] ) );
  AND U487 ( .A(B[0]), .B(A[1]), .Z(\_0_net_[1] ) );
  AND U488 ( .A(B[18]), .B(A[1]), .Z(\_0_net_[19] ) );
  AND U489 ( .A(B[17]), .B(A[1]), .Z(\_0_net_[18] ) );
  AND U490 ( .A(B[16]), .B(A[1]), .Z(\_0_net_[17] ) );
  AND U491 ( .A(B[15]), .B(A[1]), .Z(\_0_net_[16] ) );
  AND U492 ( .A(B[14]), .B(A[1]), .Z(\_0_net_[15] ) );
  AND U493 ( .A(B[13]), .B(A[1]), .Z(\_0_net_[14] ) );
  AND U494 ( .A(B[12]), .B(A[1]), .Z(\_0_net_[13] ) );
  AND U495 ( .A(B[11]), .B(A[1]), .Z(\_0_net_[12] ) );
  AND U496 ( .A(B[10]), .B(A[1]), .Z(\_0_net_[11] ) );
  AND U497 ( .A(A[1]), .B(B[9]), .Z(\_0_net_[10] ) );
endmodule


module FA_7937 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_7938 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7939 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7940 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7941 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7942 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7943 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7944 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7945 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7946 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7947 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7948 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7949 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7950 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7951 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7952 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7953 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7954 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7955 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7956 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7957 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7958 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7959 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7960 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7961 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7962 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7963 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7964 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7965 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7966 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7967 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module ADD_N32_252 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_7967 \FAINST[1].FA_  ( .A(A[1]), .B(B[1]), .CI(1'b0), .S(S[1]), .CO(C[2])
         );
  FA_7966 \FAINST[2].FA_  ( .A(A[2]), .B(B[2]), .CI(C[2]), .S(S[2]), .CO(C[3])
         );
  FA_7965 \FAINST[3].FA_  ( .A(A[3]), .B(B[3]), .CI(C[3]), .S(S[3]), .CO(C[4])
         );
  FA_7964 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_7963 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_7962 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_7961 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_7960 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_7959 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_7958 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_7957 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_7956 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_7955 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_7954 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_7953 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_7952 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_7951 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_7950 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_7949 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_7948 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_7947 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_7946 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_7945 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_7944 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_7943 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_7942 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_7941 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_7940 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_7939 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_7938 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_7937 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_7969 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_7970 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7971 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7972 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7973 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7974 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7975 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7976 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7977 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7978 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7979 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7980 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7981 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7982 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7983 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7984 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7985 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7986 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7987 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7988 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7989 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7990 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7991 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7992 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7993 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7994 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7995 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7996 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7997 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7998 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7999 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module ADD_N32_253 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_7999 \FAINST[1].FA_  ( .A(A[1]), .B(B[1]), .CI(1'b0), .S(S[1]), .CO(C[2])
         );
  FA_7998 \FAINST[2].FA_  ( .A(A[2]), .B(B[2]), .CI(C[2]), .S(S[2]), .CO(C[3])
         );
  FA_7997 \FAINST[3].FA_  ( .A(A[3]), .B(B[3]), .CI(C[3]), .S(S[3]), .CO(C[4])
         );
  FA_7996 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_7995 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_7994 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_7993 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_7992 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_7991 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_7990 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_7989 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_7988 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_7987 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_7986 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_7985 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_7984 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_7983 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_7982 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_7981 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_7980 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_7979 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_7978 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_7977 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_7976 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_7975 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_7974 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_7973 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_7972 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_7971 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_7970 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_7969 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_8001 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_8002 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8003 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8004 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8005 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8006 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8007 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8008 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8009 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8010 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8011 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8012 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8013 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8014 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8015 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8016 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8017 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8018 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8019 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8020 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8021 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8022 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8023 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8024 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8025 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8026 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8027 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8028 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8029 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8030 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8031 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module ADD_N32_254 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_8031 \FAINST[1].FA_  ( .A(A[1]), .B(B[1]), .CI(1'b0), .S(S[1]), .CO(C[2])
         );
  FA_8030 \FAINST[2].FA_  ( .A(A[2]), .B(B[2]), .CI(C[2]), .S(S[2]), .CO(C[3])
         );
  FA_8029 \FAINST[3].FA_  ( .A(A[3]), .B(B[3]), .CI(C[3]), .S(S[3]), .CO(C[4])
         );
  FA_8028 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_8027 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_8026 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_8025 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_8024 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_8023 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_8022 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_8021 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_8020 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_8019 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_8018 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_8017 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_8016 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_8015 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_8014 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_8013 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_8012 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_8011 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_8010 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_8009 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_8008 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_8007 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_8006 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_8005 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_8004 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_8003 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_8002 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_8001 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_8033 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_8034 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8035 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8036 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8037 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8038 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8039 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8040 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8041 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8042 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8043 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8044 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8045 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8046 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8047 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8048 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8049 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8050 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8051 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8052 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8053 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8054 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8055 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8056 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8057 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8058 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8059 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8060 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8061 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8062 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8063 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module ADD_N32_255 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_8063 \FAINST[1].FA_  ( .A(A[1]), .B(B[1]), .CI(1'b0), .S(S[1]), .CO(C[2])
         );
  FA_8062 \FAINST[2].FA_  ( .A(A[2]), .B(B[2]), .CI(C[2]), .S(S[2]), .CO(C[3])
         );
  FA_8061 \FAINST[3].FA_  ( .A(A[3]), .B(B[3]), .CI(C[3]), .S(S[3]), .CO(C[4])
         );
  FA_8060 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_8059 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_8058 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_8057 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_8056 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_8055 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_8054 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_8053 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_8052 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_8051 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_8050 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_8049 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_8048 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_8047 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_8046 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_8045 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_8044 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_8043 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_8042 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_8041 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_8040 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_8039 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_8038 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_8037 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_8036 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_8035 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_8034 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_8033 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module matrixMult_N_M_2_N5_M32 ( clk, rst, x, y, o );
  input [159:0] x;
  input [159:0] y;
  output [31:0] o;
  input clk, rst;
  wire   \xyi[4][31] , \xyi[4][30] , \xyi[4][29] , \xyi[4][28] , \xyi[4][27] ,
         \xyi[4][26] , \xyi[4][25] , \xyi[4][24] , \xyi[4][23] , \xyi[4][22] ,
         \xyi[4][21] , \xyi[4][20] , \xyi[4][19] , \xyi[4][18] , \xyi[4][17] ,
         \xyi[4][16] , \xyi[4][15] , \xyi[4][14] , \xyi[4][13] , \xyi[4][12] ,
         \xyi[4][11] , \xyi[4][10] , \xyi[4][9] , \xyi[4][8] , \xyi[4][7] ,
         \xyi[4][6] , \xyi[4][5] , \xyi[4][4] , \xyi[4][3] , \xyi[4][2] ,
         \xyi[4][1] , \xyi[3][31] , \xyi[3][30] , \xyi[3][29] , \xyi[3][28] ,
         \xyi[3][27] , \xyi[3][26] , \xyi[3][25] , \xyi[3][24] , \xyi[3][23] ,
         \xyi[3][22] , \xyi[3][21] , \xyi[3][20] , \xyi[3][19] , \xyi[3][18] ,
         \xyi[3][17] , \xyi[3][16] , \xyi[3][15] , \xyi[3][14] , \xyi[3][13] ,
         \xyi[3][12] , \xyi[3][11] , \xyi[3][10] , \xyi[3][9] , \xyi[3][8] ,
         \xyi[3][7] , \xyi[3][6] , \xyi[3][5] , \xyi[3][4] , \xyi[3][3] ,
         \xyi[3][2] , \xyi[3][1] , \xyi[2][31] , \xyi[2][30] , \xyi[2][29] ,
         \xyi[2][28] , \xyi[2][27] , \xyi[2][26] , \xyi[2][25] , \xyi[2][24] ,
         \xyi[2][23] , \xyi[2][22] , \xyi[2][21] , \xyi[2][20] , \xyi[2][19] ,
         \xyi[2][18] , \xyi[2][17] , \xyi[2][16] , \xyi[2][15] , \xyi[2][14] ,
         \xyi[2][13] , \xyi[2][12] , \xyi[2][11] , \xyi[2][10] , \xyi[2][9] ,
         \xyi[2][8] , \xyi[2][7] , \xyi[2][6] , \xyi[2][5] , \xyi[2][4] ,
         \xyi[2][3] , \xyi[2][2] , \xyi[2][1] , \xyi[1][31] , \xyi[1][30] ,
         \xyi[1][29] , \xyi[1][28] , \xyi[1][27] , \xyi[1][26] , \xyi[1][25] ,
         \xyi[1][24] , \xyi[1][23] , \xyi[1][22] , \xyi[1][21] , \xyi[1][20] ,
         \xyi[1][19] , \xyi[1][18] , \xyi[1][17] , \xyi[1][16] , \xyi[1][15] ,
         \xyi[1][14] , \xyi[1][13] , \xyi[1][12] , \xyi[1][11] , \xyi[1][10] ,
         \xyi[1][9] , \xyi[1][8] , \xyi[1][7] , \xyi[1][6] , \xyi[1][5] ,
         \xyi[1][4] , \xyi[1][3] , \xyi[1][2] , \xyi[1][1] , \xyi[0][31] ,
         \xyi[0][30] , \xyi[0][29] , \xyi[0][28] , \xyi[0][27] , \xyi[0][26] ,
         \xyi[0][25] , \xyi[0][24] , \xyi[0][23] , \xyi[0][22] , \xyi[0][21] ,
         \xyi[0][20] , \xyi[0][19] , \xyi[0][18] , \xyi[0][17] , \xyi[0][16] ,
         \xyi[0][15] , \xyi[0][14] , \xyi[0][13] , \xyi[0][12] , \xyi[0][11] ,
         \xyi[0][10] , \xyi[0][9] , \xyi[0][8] , \xyi[0][7] , \xyi[0][6] ,
         \xyi[0][5] , \xyi[0][4] , \xyi[0][3] , \xyi[0][2] , \xyi[0][1] ,
         \oi[5][31] , \oi[5][30] , \oi[5][29] , \oi[5][28] , \oi[5][27] ,
         \oi[5][26] , \oi[5][25] , \oi[5][24] , \oi[5][23] , \oi[5][22] ,
         \oi[5][21] , \oi[5][20] , \oi[5][19] , \oi[5][18] , \oi[5][17] ,
         \oi[5][16] , \oi[5][15] , \oi[5][14] , \oi[5][13] , \oi[5][12] ,
         \oi[5][11] , \oi[5][10] , \oi[5][9] , \oi[5][8] , \oi[5][7] ,
         \oi[5][6] , \oi[5][5] , \oi[5][4] , \oi[5][3] , \oi[5][2] ,
         \oi[5][1] , \oi[4][31] , \oi[4][30] , \oi[4][29] , \oi[4][28] ,
         \oi[4][27] , \oi[4][26] , \oi[4][25] , \oi[4][24] , \oi[4][23] ,
         \oi[4][22] , \oi[4][21] , \oi[4][20] , \oi[4][19] , \oi[4][18] ,
         \oi[4][17] , \oi[4][16] , \oi[4][15] , \oi[4][14] , \oi[4][13] ,
         \oi[4][12] , \oi[4][11] , \oi[4][10] , \oi[4][9] , \oi[4][8] ,
         \oi[4][7] , \oi[4][6] , \oi[4][5] , \oi[4][4] , \oi[4][3] ,
         \oi[4][2] , \oi[4][1] , \oi[3][31] , \oi[3][30] , \oi[3][29] ,
         \oi[3][28] , \oi[3][27] , \oi[3][26] , \oi[3][25] , \oi[3][24] ,
         \oi[3][23] , \oi[3][22] , \oi[3][21] , \oi[3][20] , \oi[3][19] ,
         \oi[3][18] , \oi[3][17] , \oi[3][16] , \oi[3][15] , \oi[3][14] ,
         \oi[3][13] , \oi[3][12] , \oi[3][11] , \oi[3][10] , \oi[3][9] ,
         \oi[3][8] , \oi[3][7] , \oi[3][6] , \oi[3][5] , \oi[3][4] ,
         \oi[3][3] , \oi[3][2] , \oi[3][1] , \oi[2][31] , \oi[2][30] ,
         \oi[2][29] , \oi[2][28] , \oi[2][27] , \oi[2][26] , \oi[2][25] ,
         \oi[2][24] , \oi[2][23] , \oi[2][22] , \oi[2][21] , \oi[2][20] ,
         \oi[2][19] , \oi[2][18] , \oi[2][17] , \oi[2][16] , \oi[2][15] ,
         \oi[2][14] , \oi[2][13] , \oi[2][12] , \oi[2][11] , \oi[2][10] ,
         \oi[2][9] , \oi[2][8] , \oi[2][7] , \oi[2][6] , \oi[2][5] ,
         \oi[2][4] , \oi[2][3] , \oi[2][2] , \oi[2][1] , \oi[1][31] ,
         \oi[1][30] , \oi[1][29] , \oi[1][28] , \oi[1][27] , \oi[1][26] ,
         \oi[1][25] , \oi[1][24] , \oi[1][23] , \oi[1][22] , \oi[1][21] ,
         \oi[1][20] , \oi[1][19] , \oi[1][18] , \oi[1][17] , \oi[1][16] ,
         \oi[1][15] , \oi[1][14] , \oi[1][13] , \oi[1][12] , \oi[1][11] ,
         \oi[1][10] , \oi[1][9] , \oi[1][8] , \oi[1][7] , \oi[1][6] ,
         \oi[1][5] , \oi[1][4] , \oi[1][3] , \oi[1][2] , \oi[1][1] ;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9;
  assign o[0] = 1'b0;

  MULT_N32_3 \MMULT_ROW[0].MULT_  ( .A({x[31:1], 1'b0}), .B({1'b0, y[30:0]}), 
        .O({\xyi[0][31] , \xyi[0][30] , \xyi[0][29] , \xyi[0][28] , 
        \xyi[0][27] , \xyi[0][26] , \xyi[0][25] , \xyi[0][24] , \xyi[0][23] , 
        \xyi[0][22] , \xyi[0][21] , \xyi[0][20] , \xyi[0][19] , \xyi[0][18] , 
        \xyi[0][17] , \xyi[0][16] , \xyi[0][15] , \xyi[0][14] , \xyi[0][13] , 
        \xyi[0][12] , \xyi[0][11] , \xyi[0][10] , \xyi[0][9] , \xyi[0][8] , 
        \xyi[0][7] , \xyi[0][6] , \xyi[0][5] , \xyi[0][4] , \xyi[0][3] , 
        \xyi[0][2] , \xyi[0][1] , SYNOPSYS_UNCONNECTED__0}) );
  MULT_N32_7 \MMULT_ROW[1].MULT_  ( .A({x[63:33], 1'b0}), .B({1'b0, y[62:32]}), 
        .O({\xyi[1][31] , \xyi[1][30] , \xyi[1][29] , \xyi[1][28] , 
        \xyi[1][27] , \xyi[1][26] , \xyi[1][25] , \xyi[1][24] , \xyi[1][23] , 
        \xyi[1][22] , \xyi[1][21] , \xyi[1][20] , \xyi[1][19] , \xyi[1][18] , 
        \xyi[1][17] , \xyi[1][16] , \xyi[1][15] , \xyi[1][14] , \xyi[1][13] , 
        \xyi[1][12] , \xyi[1][11] , \xyi[1][10] , \xyi[1][9] , \xyi[1][8] , 
        \xyi[1][7] , \xyi[1][6] , \xyi[1][5] , \xyi[1][4] , \xyi[1][3] , 
        \xyi[1][2] , \xyi[1][1] , SYNOPSYS_UNCONNECTED__1}) );
  MULT_N32_6 \MMULT_ROW[2].MULT_  ( .A({x[95:65], 1'b0}), .B({1'b0, y[94:64]}), 
        .O({\xyi[2][31] , \xyi[2][30] , \xyi[2][29] , \xyi[2][28] , 
        \xyi[2][27] , \xyi[2][26] , \xyi[2][25] , \xyi[2][24] , \xyi[2][23] , 
        \xyi[2][22] , \xyi[2][21] , \xyi[2][20] , \xyi[2][19] , \xyi[2][18] , 
        \xyi[2][17] , \xyi[2][16] , \xyi[2][15] , \xyi[2][14] , \xyi[2][13] , 
        \xyi[2][12] , \xyi[2][11] , \xyi[2][10] , \xyi[2][9] , \xyi[2][8] , 
        \xyi[2][7] , \xyi[2][6] , \xyi[2][5] , \xyi[2][4] , \xyi[2][3] , 
        \xyi[2][2] , \xyi[2][1] , SYNOPSYS_UNCONNECTED__2}) );
  MULT_N32_5 \MMULT_ROW[3].MULT_  ( .A({x[127:97], 1'b0}), .B({1'b0, y[126:96]}), .O({\xyi[3][31] , \xyi[3][30] , \xyi[3][29] , \xyi[3][28] , \xyi[3][27] , 
        \xyi[3][26] , \xyi[3][25] , \xyi[3][24] , \xyi[3][23] , \xyi[3][22] , 
        \xyi[3][21] , \xyi[3][20] , \xyi[3][19] , \xyi[3][18] , \xyi[3][17] , 
        \xyi[3][16] , \xyi[3][15] , \xyi[3][14] , \xyi[3][13] , \xyi[3][12] , 
        \xyi[3][11] , \xyi[3][10] , \xyi[3][9] , \xyi[3][8] , \xyi[3][7] , 
        \xyi[3][6] , \xyi[3][5] , \xyi[3][4] , \xyi[3][3] , \xyi[3][2] , 
        \xyi[3][1] , SYNOPSYS_UNCONNECTED__3}) );
  MULT_N32_4 \MMULT_ROW[4].MULT_  ( .A({x[159:129], 1'b0}), .B({1'b0, 
        y[158:128]}), .O({\xyi[4][31] , \xyi[4][30] , \xyi[4][29] , 
        \xyi[4][28] , \xyi[4][27] , \xyi[4][26] , \xyi[4][25] , \xyi[4][24] , 
        \xyi[4][23] , \xyi[4][22] , \xyi[4][21] , \xyi[4][20] , \xyi[4][19] , 
        \xyi[4][18] , \xyi[4][17] , \xyi[4][16] , \xyi[4][15] , \xyi[4][14] , 
        \xyi[4][13] , \xyi[4][12] , \xyi[4][11] , \xyi[4][10] , \xyi[4][9] , 
        \xyi[4][8] , \xyi[4][7] , \xyi[4][6] , \xyi[4][5] , \xyi[4][4] , 
        \xyi[4][3] , \xyi[4][2] , \xyi[4][1] , SYNOPSYS_UNCONNECTED__4}) );
  ADD_N32_96 \ADD_ROW[0].ADD_  ( .A({\xyi[0][31] , \xyi[0][30] , \xyi[0][29] , 
        \xyi[0][28] , \xyi[0][27] , \xyi[0][26] , \xyi[0][25] , \xyi[0][24] , 
        \xyi[0][23] , \xyi[0][22] , \xyi[0][21] , \xyi[0][20] , \xyi[0][19] , 
        \xyi[0][18] , \xyi[0][17] , \xyi[0][16] , \xyi[0][15] , \xyi[0][14] , 
        \xyi[0][13] , \xyi[0][12] , \xyi[0][11] , \xyi[0][10] , \xyi[0][9] , 
        \xyi[0][8] , \xyi[0][7] , \xyi[0][6] , \xyi[0][5] , \xyi[0][4] , 
        \xyi[0][3] , \xyi[0][2] , \xyi[0][1] , 1'b0}), .B({o[31:1], 1'b0}), 
        .CI(1'b0), .S({\oi[1][31] , \oi[1][30] , \oi[1][29] , \oi[1][28] , 
        \oi[1][27] , \oi[1][26] , \oi[1][25] , \oi[1][24] , \oi[1][23] , 
        \oi[1][22] , \oi[1][21] , \oi[1][20] , \oi[1][19] , \oi[1][18] , 
        \oi[1][17] , \oi[1][16] , \oi[1][15] , \oi[1][14] , \oi[1][13] , 
        \oi[1][12] , \oi[1][11] , \oi[1][10] , \oi[1][9] , \oi[1][8] , 
        \oi[1][7] , \oi[1][6] , \oi[1][5] , \oi[1][4] , \oi[1][3] , \oi[1][2] , 
        \oi[1][1] , SYNOPSYS_UNCONNECTED__5}) );
  ADD_N32_255 \ADD_ROW[1].ADD_  ( .A({\xyi[1][31] , \xyi[1][30] , \xyi[1][29] , 
        \xyi[1][28] , \xyi[1][27] , \xyi[1][26] , \xyi[1][25] , \xyi[1][24] , 
        \xyi[1][23] , \xyi[1][22] , \xyi[1][21] , \xyi[1][20] , \xyi[1][19] , 
        \xyi[1][18] , \xyi[1][17] , \xyi[1][16] , \xyi[1][15] , \xyi[1][14] , 
        \xyi[1][13] , \xyi[1][12] , \xyi[1][11] , \xyi[1][10] , \xyi[1][9] , 
        \xyi[1][8] , \xyi[1][7] , \xyi[1][6] , \xyi[1][5] , \xyi[1][4] , 
        \xyi[1][3] , \xyi[1][2] , \xyi[1][1] , 1'b0}), .B({\oi[1][31] , 
        \oi[1][30] , \oi[1][29] , \oi[1][28] , \oi[1][27] , \oi[1][26] , 
        \oi[1][25] , \oi[1][24] , \oi[1][23] , \oi[1][22] , \oi[1][21] , 
        \oi[1][20] , \oi[1][19] , \oi[1][18] , \oi[1][17] , \oi[1][16] , 
        \oi[1][15] , \oi[1][14] , \oi[1][13] , \oi[1][12] , \oi[1][11] , 
        \oi[1][10] , \oi[1][9] , \oi[1][8] , \oi[1][7] , \oi[1][6] , 
        \oi[1][5] , \oi[1][4] , \oi[1][3] , \oi[1][2] , \oi[1][1] , 1'b0}), 
        .CI(1'b0), .S({\oi[2][31] , \oi[2][30] , \oi[2][29] , \oi[2][28] , 
        \oi[2][27] , \oi[2][26] , \oi[2][25] , \oi[2][24] , \oi[2][23] , 
        \oi[2][22] , \oi[2][21] , \oi[2][20] , \oi[2][19] , \oi[2][18] , 
        \oi[2][17] , \oi[2][16] , \oi[2][15] , \oi[2][14] , \oi[2][13] , 
        \oi[2][12] , \oi[2][11] , \oi[2][10] , \oi[2][9] , \oi[2][8] , 
        \oi[2][7] , \oi[2][6] , \oi[2][5] , \oi[2][4] , \oi[2][3] , \oi[2][2] , 
        \oi[2][1] , SYNOPSYS_UNCONNECTED__6}) );
  ADD_N32_254 \ADD_ROW[2].ADD_  ( .A({\xyi[2][31] , \xyi[2][30] , \xyi[2][29] , 
        \xyi[2][28] , \xyi[2][27] , \xyi[2][26] , \xyi[2][25] , \xyi[2][24] , 
        \xyi[2][23] , \xyi[2][22] , \xyi[2][21] , \xyi[2][20] , \xyi[2][19] , 
        \xyi[2][18] , \xyi[2][17] , \xyi[2][16] , \xyi[2][15] , \xyi[2][14] , 
        \xyi[2][13] , \xyi[2][12] , \xyi[2][11] , \xyi[2][10] , \xyi[2][9] , 
        \xyi[2][8] , \xyi[2][7] , \xyi[2][6] , \xyi[2][5] , \xyi[2][4] , 
        \xyi[2][3] , \xyi[2][2] , \xyi[2][1] , 1'b0}), .B({\oi[2][31] , 
        \oi[2][30] , \oi[2][29] , \oi[2][28] , \oi[2][27] , \oi[2][26] , 
        \oi[2][25] , \oi[2][24] , \oi[2][23] , \oi[2][22] , \oi[2][21] , 
        \oi[2][20] , \oi[2][19] , \oi[2][18] , \oi[2][17] , \oi[2][16] , 
        \oi[2][15] , \oi[2][14] , \oi[2][13] , \oi[2][12] , \oi[2][11] , 
        \oi[2][10] , \oi[2][9] , \oi[2][8] , \oi[2][7] , \oi[2][6] , 
        \oi[2][5] , \oi[2][4] , \oi[2][3] , \oi[2][2] , \oi[2][1] , 1'b0}), 
        .CI(1'b0), .S({\oi[3][31] , \oi[3][30] , \oi[3][29] , \oi[3][28] , 
        \oi[3][27] , \oi[3][26] , \oi[3][25] , \oi[3][24] , \oi[3][23] , 
        \oi[3][22] , \oi[3][21] , \oi[3][20] , \oi[3][19] , \oi[3][18] , 
        \oi[3][17] , \oi[3][16] , \oi[3][15] , \oi[3][14] , \oi[3][13] , 
        \oi[3][12] , \oi[3][11] , \oi[3][10] , \oi[3][9] , \oi[3][8] , 
        \oi[3][7] , \oi[3][6] , \oi[3][5] , \oi[3][4] , \oi[3][3] , \oi[3][2] , 
        \oi[3][1] , SYNOPSYS_UNCONNECTED__7}) );
  ADD_N32_253 \ADD_ROW[3].ADD_  ( .A({\xyi[3][31] , \xyi[3][30] , \xyi[3][29] , 
        \xyi[3][28] , \xyi[3][27] , \xyi[3][26] , \xyi[3][25] , \xyi[3][24] , 
        \xyi[3][23] , \xyi[3][22] , \xyi[3][21] , \xyi[3][20] , \xyi[3][19] , 
        \xyi[3][18] , \xyi[3][17] , \xyi[3][16] , \xyi[3][15] , \xyi[3][14] , 
        \xyi[3][13] , \xyi[3][12] , \xyi[3][11] , \xyi[3][10] , \xyi[3][9] , 
        \xyi[3][8] , \xyi[3][7] , \xyi[3][6] , \xyi[3][5] , \xyi[3][4] , 
        \xyi[3][3] , \xyi[3][2] , \xyi[3][1] , 1'b0}), .B({\oi[3][31] , 
        \oi[3][30] , \oi[3][29] , \oi[3][28] , \oi[3][27] , \oi[3][26] , 
        \oi[3][25] , \oi[3][24] , \oi[3][23] , \oi[3][22] , \oi[3][21] , 
        \oi[3][20] , \oi[3][19] , \oi[3][18] , \oi[3][17] , \oi[3][16] , 
        \oi[3][15] , \oi[3][14] , \oi[3][13] , \oi[3][12] , \oi[3][11] , 
        \oi[3][10] , \oi[3][9] , \oi[3][8] , \oi[3][7] , \oi[3][6] , 
        \oi[3][5] , \oi[3][4] , \oi[3][3] , \oi[3][2] , \oi[3][1] , 1'b0}), 
        .CI(1'b0), .S({\oi[4][31] , \oi[4][30] , \oi[4][29] , \oi[4][28] , 
        \oi[4][27] , \oi[4][26] , \oi[4][25] , \oi[4][24] , \oi[4][23] , 
        \oi[4][22] , \oi[4][21] , \oi[4][20] , \oi[4][19] , \oi[4][18] , 
        \oi[4][17] , \oi[4][16] , \oi[4][15] , \oi[4][14] , \oi[4][13] , 
        \oi[4][12] , \oi[4][11] , \oi[4][10] , \oi[4][9] , \oi[4][8] , 
        \oi[4][7] , \oi[4][6] , \oi[4][5] , \oi[4][4] , \oi[4][3] , \oi[4][2] , 
        \oi[4][1] , SYNOPSYS_UNCONNECTED__8}) );
  ADD_N32_252 \ADD_ROW[4].ADD_  ( .A({\xyi[4][31] , \xyi[4][30] , \xyi[4][29] , 
        \xyi[4][28] , \xyi[4][27] , \xyi[4][26] , \xyi[4][25] , \xyi[4][24] , 
        \xyi[4][23] , \xyi[4][22] , \xyi[4][21] , \xyi[4][20] , \xyi[4][19] , 
        \xyi[4][18] , \xyi[4][17] , \xyi[4][16] , \xyi[4][15] , \xyi[4][14] , 
        \xyi[4][13] , \xyi[4][12] , \xyi[4][11] , \xyi[4][10] , \xyi[4][9] , 
        \xyi[4][8] , \xyi[4][7] , \xyi[4][6] , \xyi[4][5] , \xyi[4][4] , 
        \xyi[4][3] , \xyi[4][2] , \xyi[4][1] , 1'b0}), .B({\oi[4][31] , 
        \oi[4][30] , \oi[4][29] , \oi[4][28] , \oi[4][27] , \oi[4][26] , 
        \oi[4][25] , \oi[4][24] , \oi[4][23] , \oi[4][22] , \oi[4][21] , 
        \oi[4][20] , \oi[4][19] , \oi[4][18] , \oi[4][17] , \oi[4][16] , 
        \oi[4][15] , \oi[4][14] , \oi[4][13] , \oi[4][12] , \oi[4][11] , 
        \oi[4][10] , \oi[4][9] , \oi[4][8] , \oi[4][7] , \oi[4][6] , 
        \oi[4][5] , \oi[4][4] , \oi[4][3] , \oi[4][2] , \oi[4][1] , 1'b0}), 
        .CI(1'b0), .S({\oi[5][31] , \oi[5][30] , \oi[5][29] , \oi[5][28] , 
        \oi[5][27] , \oi[5][26] , \oi[5][25] , \oi[5][24] , \oi[5][23] , 
        \oi[5][22] , \oi[5][21] , \oi[5][20] , \oi[5][19] , \oi[5][18] , 
        \oi[5][17] , \oi[5][16] , \oi[5][15] , \oi[5][14] , \oi[5][13] , 
        \oi[5][12] , \oi[5][11] , \oi[5][10] , \oi[5][9] , \oi[5][8] , 
        \oi[5][7] , \oi[5][6] , \oi[5][5] , \oi[5][4] , \oi[5][3] , \oi[5][2] , 
        \oi[5][1] , SYNOPSYS_UNCONNECTED__9}) );
  DFF \o_reg[1]  ( .D(\oi[5][1] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[1]) );
  DFF \o_reg[2]  ( .D(\oi[5][2] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[2]) );
  DFF \o_reg[3]  ( .D(\oi[5][3] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[3]) );
  DFF \o_reg[4]  ( .D(\oi[5][4] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[4]) );
  DFF \o_reg[5]  ( .D(\oi[5][5] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[5]) );
  DFF \o_reg[6]  ( .D(\oi[5][6] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[6]) );
  DFF \o_reg[7]  ( .D(\oi[5][7] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[7]) );
  DFF \o_reg[8]  ( .D(\oi[5][8] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[8]) );
  DFF \o_reg[9]  ( .D(\oi[5][9] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[9]) );
  DFF \o_reg[10]  ( .D(\oi[5][10] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[10])
         );
  DFF \o_reg[11]  ( .D(\oi[5][11] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[11])
         );
  DFF \o_reg[12]  ( .D(\oi[5][12] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[12])
         );
  DFF \o_reg[13]  ( .D(\oi[5][13] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[13])
         );
  DFF \o_reg[14]  ( .D(\oi[5][14] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[14])
         );
  DFF \o_reg[15]  ( .D(\oi[5][15] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[15])
         );
  DFF \o_reg[16]  ( .D(\oi[5][16] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[16])
         );
  DFF \o_reg[17]  ( .D(\oi[5][17] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[17])
         );
  DFF \o_reg[18]  ( .D(\oi[5][18] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[18])
         );
  DFF \o_reg[19]  ( .D(\oi[5][19] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[19])
         );
  DFF \o_reg[20]  ( .D(\oi[5][20] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[20])
         );
  DFF \o_reg[21]  ( .D(\oi[5][21] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[21])
         );
  DFF \o_reg[22]  ( .D(\oi[5][22] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[22])
         );
  DFF \o_reg[23]  ( .D(\oi[5][23] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[23])
         );
  DFF \o_reg[24]  ( .D(\oi[5][24] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[24])
         );
  DFF \o_reg[25]  ( .D(\oi[5][25] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[25])
         );
  DFF \o_reg[26]  ( .D(\oi[5][26] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[26])
         );
  DFF \o_reg[27]  ( .D(\oi[5][27] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[27])
         );
  DFF \o_reg[28]  ( .D(\oi[5][28] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[28])
         );
  DFF \o_reg[29]  ( .D(\oi[5][29] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[29])
         );
  DFF \o_reg[30]  ( .D(\oi[5][30] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[30])
         );
  DFF \o_reg[31]  ( .D(\oi[5][31] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[31])
         );
endmodule

