
module FA_1024 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  AND U1 ( .A(A), .B(B), .Z(CO) );
  XOR U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_2047 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2046 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2045 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2044 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2043 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2042 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2041 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2040 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2039 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2038 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2037 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2036 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2035 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2034 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2033 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2032 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2031 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2030 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2029 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2028 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2027 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2026 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2025 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2024 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2023 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2022 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2021 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2020 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2019 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2018 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2017 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2016 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2015 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2014 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2013 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2012 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2011 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2010 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2009 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2008 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2007 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2006 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2005 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2004 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2003 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2002 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2001 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2000 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1999 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1998 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1997 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1996 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1995 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1994 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1993 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1992 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1991 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1990 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1989 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1988 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1987 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1986 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1985 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1984 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1983 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1982 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1981 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1980 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1979 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1978 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1977 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1976 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1975 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1974 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1973 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1972 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1971 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1970 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1969 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1968 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1967 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1966 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1965 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1964 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1963 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1962 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1961 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1960 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1959 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1958 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1957 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1956 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1955 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1954 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1953 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1952 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1951 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1950 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1949 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1948 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1947 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1946 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1945 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1944 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1943 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1942 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1941 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1940 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1939 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1938 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1937 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1936 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1935 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1934 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1933 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1932 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1931 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1930 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1929 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1928 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1927 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1926 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1925 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1924 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1923 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1922 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1921 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1920 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1919 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1918 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1917 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1916 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1915 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1914 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1913 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1912 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1911 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1910 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1909 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1908 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1907 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1906 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1905 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1904 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1903 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1902 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1901 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1900 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1899 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1898 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1897 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1896 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1895 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1894 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1893 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1892 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1891 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1890 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1889 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1888 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1887 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1886 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1885 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1884 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1883 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1882 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1881 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1880 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1879 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1878 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1877 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1876 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1875 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1874 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1873 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1872 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1871 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1870 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1869 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1868 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1867 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1866 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1865 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1864 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1863 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1862 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1861 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1860 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1859 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1858 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1857 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1856 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1855 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1854 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1853 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1852 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1851 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1850 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1849 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1848 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1847 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1846 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1845 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1844 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1843 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1842 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1841 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1840 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1839 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1838 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1837 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1836 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1835 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1834 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1833 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1832 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1831 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1830 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1829 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1828 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1827 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1826 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1825 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1824 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1823 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1822 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1821 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1820 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1819 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1818 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1817 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1816 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1815 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1814 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1813 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1812 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1811 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1810 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1809 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1808 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1807 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1806 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1805 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1804 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1803 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1802 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1801 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1800 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1799 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1798 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1797 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1796 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1795 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1794 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1793 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1792 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1791 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1790 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1789 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1788 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1787 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1786 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1785 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1784 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1783 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1782 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1781 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1780 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1779 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1778 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1777 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1776 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1775 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1774 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1773 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1772 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1771 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1770 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1769 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1768 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1767 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1766 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1765 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1764 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1763 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1762 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1761 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1760 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1759 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1758 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1757 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1756 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1755 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1754 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1753 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1752 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1751 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1750 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1749 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1748 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1747 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1746 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1745 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1744 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1743 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1742 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1741 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1740 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1739 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1738 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1737 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1736 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1735 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1734 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1733 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1732 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1731 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1730 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1729 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1728 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1727 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1726 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1725 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1724 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1723 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1722 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1721 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1720 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1719 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1718 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1717 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1716 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1715 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1714 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1713 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1712 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1711 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1710 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1709 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1708 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1707 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1706 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1705 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1704 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1703 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1702 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1701 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1700 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1699 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1698 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1697 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1696 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1695 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1694 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1693 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1692 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1691 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1690 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1689 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1688 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1687 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1686 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1685 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1684 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1683 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1682 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1681 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1680 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1679 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1678 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1677 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1676 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1675 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1674 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1673 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1672 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1671 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1670 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1669 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1668 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1667 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1666 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1665 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1664 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1663 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1662 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1661 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1660 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1659 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1658 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1657 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1656 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1655 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1654 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1653 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1652 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1651 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1650 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1649 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1648 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1647 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1646 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1645 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1644 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1643 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1642 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1641 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1640 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1639 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1638 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1637 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1636 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1635 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1634 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1633 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1632 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1631 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1630 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1629 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1628 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1627 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1626 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1625 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1624 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1623 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1622 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1621 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1620 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1619 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1618 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1617 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1616 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1615 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1614 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1613 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1612 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1611 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1610 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1609 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1608 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1607 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1606 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1605 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1604 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1603 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1602 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1601 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1600 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1599 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1598 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1597 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1596 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1595 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1594 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1593 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1592 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1591 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1590 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1589 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1588 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1587 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1586 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1585 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1584 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1583 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1582 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1581 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1580 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1579 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1578 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1577 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1576 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1575 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1574 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1573 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1572 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1571 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1570 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1569 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1568 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1567 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1566 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1565 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1564 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1563 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1562 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1561 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1560 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1559 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1558 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1557 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1556 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1555 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1554 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1553 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1552 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1551 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1550 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1549 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1548 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1547 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1546 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1545 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1544 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1543 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1542 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1541 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1540 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1539 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1538 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1537 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1536 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1535 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1534 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1533 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1532 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1531 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1530 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1529 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1528 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1527 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1526 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1525 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1524 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1523 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1522 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1521 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1520 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1519 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1518 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1517 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1516 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1515 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1514 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1513 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1512 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1504 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1488 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1472 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1456 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1440 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1424 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1408 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1392 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1376 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1360 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1344 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1328 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1312 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1296 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1280 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1264 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1248 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1232 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1216 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1200 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1184 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1168 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1152 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1136 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1120 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1104 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1099 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1098 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1097 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1096 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1095 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1094 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1093 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1092 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1091 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1090 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1089 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1088 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1087 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1086 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1085 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1084 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1083 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1082 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1081 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1080 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1079 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1078 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1077 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1076 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1075 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1074 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1073 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1072 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1071 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1070 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1069 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1068 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1067 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1066 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1065 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1064 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1063 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1062 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1061 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1060 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1059 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1058 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1057 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1056 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1055 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1054 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1053 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1052 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1051 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1050 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1049 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1048 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1047 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1046 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1045 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1044 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1043 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1042 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1041 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1040 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1039 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1038 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1037 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1036 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1035 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1034 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1033 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1032 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1031 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1030 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1029 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1028 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1027 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1026 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  XOR U2 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_1025 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N1024_1 ( A, B, CI, S, CO );
  input [1023:0] A;
  input [1023:0] B;
  output [1023:0] S;
  input CI;
  output CO;

  wire   [1023:1] C;

  FA_1024 \FA_INST_0[0].FA_INST_1[0].FA_  ( .A(A[0]), .B(B[0]), .CI(1'b0), .S(
        S[0]), .CO(C[1]) );
  FA_2047 \FA_INST_0[0].FA_INST_1[1].FA_  ( .A(A[1]), .B(B[1]), .CI(C[1]), .S(
        S[1]), .CO(C[2]) );
  FA_2046 \FA_INST_0[0].FA_INST_1[2].FA_  ( .A(A[2]), .B(B[2]), .CI(C[2]), .S(
        S[2]), .CO(C[3]) );
  FA_2045 \FA_INST_0[0].FA_INST_1[3].FA_  ( .A(A[3]), .B(B[3]), .CI(C[3]), .S(
        S[3]), .CO(C[4]) );
  FA_2044 \FA_INST_0[0].FA_INST_1[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(
        S[4]), .CO(C[5]) );
  FA_2043 \FA_INST_0[0].FA_INST_1[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(
        S[5]), .CO(C[6]) );
  FA_2042 \FA_INST_0[0].FA_INST_1[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(
        S[6]), .CO(C[7]) );
  FA_2041 \FA_INST_0[0].FA_INST_1[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(
        S[7]), .CO(C[8]) );
  FA_2040 \FA_INST_0[0].FA_INST_1[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(
        S[8]), .CO(C[9]) );
  FA_2039 \FA_INST_0[0].FA_INST_1[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(
        S[9]), .CO(C[10]) );
  FA_2038 \FA_INST_0[0].FA_INST_1[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), 
        .S(S[10]), .CO(C[11]) );
  FA_2037 \FA_INST_0[0].FA_INST_1[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), 
        .S(S[11]), .CO(C[12]) );
  FA_2036 \FA_INST_0[0].FA_INST_1[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), 
        .S(S[12]), .CO(C[13]) );
  FA_2035 \FA_INST_0[0].FA_INST_1[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), 
        .S(S[13]), .CO(C[14]) );
  FA_2034 \FA_INST_0[0].FA_INST_1[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), 
        .S(S[14]), .CO(C[15]) );
  FA_2033 \FA_INST_0[0].FA_INST_1[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), 
        .S(S[15]), .CO(C[16]) );
  FA_2032 \FA_INST_0[0].FA_INST_1[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), 
        .S(S[16]), .CO(C[17]) );
  FA_2031 \FA_INST_0[0].FA_INST_1[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), 
        .S(S[17]), .CO(C[18]) );
  FA_2030 \FA_INST_0[0].FA_INST_1[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), 
        .S(S[18]), .CO(C[19]) );
  FA_2029 \FA_INST_0[0].FA_INST_1[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), 
        .S(S[19]), .CO(C[20]) );
  FA_2028 \FA_INST_0[0].FA_INST_1[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), 
        .S(S[20]), .CO(C[21]) );
  FA_2027 \FA_INST_0[0].FA_INST_1[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), 
        .S(S[21]), .CO(C[22]) );
  FA_2026 \FA_INST_0[0].FA_INST_1[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), 
        .S(S[22]), .CO(C[23]) );
  FA_2025 \FA_INST_0[0].FA_INST_1[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), 
        .S(S[23]), .CO(C[24]) );
  FA_2024 \FA_INST_0[0].FA_INST_1[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), 
        .S(S[24]), .CO(C[25]) );
  FA_2023 \FA_INST_0[0].FA_INST_1[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), 
        .S(S[25]), .CO(C[26]) );
  FA_2022 \FA_INST_0[0].FA_INST_1[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), 
        .S(S[26]), .CO(C[27]) );
  FA_2021 \FA_INST_0[0].FA_INST_1[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), 
        .S(S[27]), .CO(C[28]) );
  FA_2020 \FA_INST_0[0].FA_INST_1[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), 
        .S(S[28]), .CO(C[29]) );
  FA_2019 \FA_INST_0[0].FA_INST_1[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), 
        .S(S[29]), .CO(C[30]) );
  FA_2018 \FA_INST_0[0].FA_INST_1[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), 
        .S(S[30]), .CO(C[31]) );
  FA_2017 \FA_INST_0[0].FA_INST_1[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), 
        .S(S[31]), .CO(C[32]) );
  FA_2016 \FA_INST_0[0].FA_INST_1[32].FA_  ( .A(A[32]), .B(B[32]), .CI(C[32]), 
        .S(S[32]), .CO(C[33]) );
  FA_2015 \FA_INST_0[0].FA_INST_1[33].FA_  ( .A(A[33]), .B(B[33]), .CI(C[33]), 
        .S(S[33]), .CO(C[34]) );
  FA_2014 \FA_INST_0[0].FA_INST_1[34].FA_  ( .A(A[34]), .B(B[34]), .CI(C[34]), 
        .S(S[34]), .CO(C[35]) );
  FA_2013 \FA_INST_0[0].FA_INST_1[35].FA_  ( .A(A[35]), .B(B[35]), .CI(C[35]), 
        .S(S[35]), .CO(C[36]) );
  FA_2012 \FA_INST_0[0].FA_INST_1[36].FA_  ( .A(A[36]), .B(B[36]), .CI(C[36]), 
        .S(S[36]), .CO(C[37]) );
  FA_2011 \FA_INST_0[0].FA_INST_1[37].FA_  ( .A(A[37]), .B(B[37]), .CI(C[37]), 
        .S(S[37]), .CO(C[38]) );
  FA_2010 \FA_INST_0[0].FA_INST_1[38].FA_  ( .A(A[38]), .B(B[38]), .CI(C[38]), 
        .S(S[38]), .CO(C[39]) );
  FA_2009 \FA_INST_0[0].FA_INST_1[39].FA_  ( .A(A[39]), .B(B[39]), .CI(C[39]), 
        .S(S[39]), .CO(C[40]) );
  FA_2008 \FA_INST_0[0].FA_INST_1[40].FA_  ( .A(A[40]), .B(B[40]), .CI(C[40]), 
        .S(S[40]), .CO(C[41]) );
  FA_2007 \FA_INST_0[0].FA_INST_1[41].FA_  ( .A(A[41]), .B(B[41]), .CI(C[41]), 
        .S(S[41]), .CO(C[42]) );
  FA_2006 \FA_INST_0[0].FA_INST_1[42].FA_  ( .A(A[42]), .B(B[42]), .CI(C[42]), 
        .S(S[42]), .CO(C[43]) );
  FA_2005 \FA_INST_0[0].FA_INST_1[43].FA_  ( .A(A[43]), .B(B[43]), .CI(C[43]), 
        .S(S[43]), .CO(C[44]) );
  FA_2004 \FA_INST_0[0].FA_INST_1[44].FA_  ( .A(A[44]), .B(B[44]), .CI(C[44]), 
        .S(S[44]), .CO(C[45]) );
  FA_2003 \FA_INST_0[0].FA_INST_1[45].FA_  ( .A(A[45]), .B(B[45]), .CI(C[45]), 
        .S(S[45]), .CO(C[46]) );
  FA_2002 \FA_INST_0[0].FA_INST_1[46].FA_  ( .A(A[46]), .B(B[46]), .CI(C[46]), 
        .S(S[46]), .CO(C[47]) );
  FA_2001 \FA_INST_0[0].FA_INST_1[47].FA_  ( .A(A[47]), .B(B[47]), .CI(C[47]), 
        .S(S[47]), .CO(C[48]) );
  FA_2000 \FA_INST_0[0].FA_INST_1[48].FA_  ( .A(A[48]), .B(B[48]), .CI(C[48]), 
        .S(S[48]), .CO(C[49]) );
  FA_1999 \FA_INST_0[0].FA_INST_1[49].FA_  ( .A(A[49]), .B(B[49]), .CI(C[49]), 
        .S(S[49]), .CO(C[50]) );
  FA_1998 \FA_INST_0[0].FA_INST_1[50].FA_  ( .A(A[50]), .B(B[50]), .CI(C[50]), 
        .S(S[50]), .CO(C[51]) );
  FA_1997 \FA_INST_0[0].FA_INST_1[51].FA_  ( .A(A[51]), .B(B[51]), .CI(C[51]), 
        .S(S[51]), .CO(C[52]) );
  FA_1996 \FA_INST_0[0].FA_INST_1[52].FA_  ( .A(A[52]), .B(B[52]), .CI(C[52]), 
        .S(S[52]), .CO(C[53]) );
  FA_1995 \FA_INST_0[0].FA_INST_1[53].FA_  ( .A(A[53]), .B(B[53]), .CI(C[53]), 
        .S(S[53]), .CO(C[54]) );
  FA_1994 \FA_INST_0[0].FA_INST_1[54].FA_  ( .A(A[54]), .B(B[54]), .CI(C[54]), 
        .S(S[54]), .CO(C[55]) );
  FA_1993 \FA_INST_0[0].FA_INST_1[55].FA_  ( .A(A[55]), .B(B[55]), .CI(C[55]), 
        .S(S[55]), .CO(C[56]) );
  FA_1992 \FA_INST_0[0].FA_INST_1[56].FA_  ( .A(A[56]), .B(B[56]), .CI(C[56]), 
        .S(S[56]), .CO(C[57]) );
  FA_1991 \FA_INST_0[0].FA_INST_1[57].FA_  ( .A(A[57]), .B(B[57]), .CI(C[57]), 
        .S(S[57]), .CO(C[58]) );
  FA_1990 \FA_INST_0[0].FA_INST_1[58].FA_  ( .A(A[58]), .B(B[58]), .CI(C[58]), 
        .S(S[58]), .CO(C[59]) );
  FA_1989 \FA_INST_0[0].FA_INST_1[59].FA_  ( .A(A[59]), .B(B[59]), .CI(C[59]), 
        .S(S[59]), .CO(C[60]) );
  FA_1988 \FA_INST_0[0].FA_INST_1[60].FA_  ( .A(A[60]), .B(B[60]), .CI(C[60]), 
        .S(S[60]), .CO(C[61]) );
  FA_1987 \FA_INST_0[0].FA_INST_1[61].FA_  ( .A(A[61]), .B(B[61]), .CI(C[61]), 
        .S(S[61]), .CO(C[62]) );
  FA_1986 \FA_INST_0[0].FA_INST_1[62].FA_  ( .A(A[62]), .B(B[62]), .CI(C[62]), 
        .S(S[62]), .CO(C[63]) );
  FA_1985 \FA_INST_0[0].FA_INST_1[63].FA_  ( .A(A[63]), .B(B[63]), .CI(C[63]), 
        .S(S[63]), .CO(C[64]) );
  FA_1984 \FA_INST_0[0].FA_INST_1[64].FA_  ( .A(A[64]), .B(B[64]), .CI(C[64]), 
        .S(S[64]), .CO(C[65]) );
  FA_1983 \FA_INST_0[0].FA_INST_1[65].FA_  ( .A(A[65]), .B(B[65]), .CI(C[65]), 
        .S(S[65]), .CO(C[66]) );
  FA_1982 \FA_INST_0[0].FA_INST_1[66].FA_  ( .A(A[66]), .B(B[66]), .CI(C[66]), 
        .S(S[66]), .CO(C[67]) );
  FA_1981 \FA_INST_0[0].FA_INST_1[67].FA_  ( .A(A[67]), .B(B[67]), .CI(C[67]), 
        .S(S[67]), .CO(C[68]) );
  FA_1980 \FA_INST_0[0].FA_INST_1[68].FA_  ( .A(A[68]), .B(B[68]), .CI(C[68]), 
        .S(S[68]), .CO(C[69]) );
  FA_1979 \FA_INST_0[0].FA_INST_1[69].FA_  ( .A(A[69]), .B(B[69]), .CI(C[69]), 
        .S(S[69]), .CO(C[70]) );
  FA_1978 \FA_INST_0[0].FA_INST_1[70].FA_  ( .A(A[70]), .B(B[70]), .CI(C[70]), 
        .S(S[70]), .CO(C[71]) );
  FA_1977 \FA_INST_0[0].FA_INST_1[71].FA_  ( .A(A[71]), .B(B[71]), .CI(C[71]), 
        .S(S[71]), .CO(C[72]) );
  FA_1976 \FA_INST_0[0].FA_INST_1[72].FA_  ( .A(A[72]), .B(B[72]), .CI(C[72]), 
        .S(S[72]), .CO(C[73]) );
  FA_1975 \FA_INST_0[0].FA_INST_1[73].FA_  ( .A(A[73]), .B(B[73]), .CI(C[73]), 
        .S(S[73]), .CO(C[74]) );
  FA_1974 \FA_INST_0[0].FA_INST_1[74].FA_  ( .A(A[74]), .B(B[74]), .CI(C[74]), 
        .S(S[74]), .CO(C[75]) );
  FA_1973 \FA_INST_0[0].FA_INST_1[75].FA_  ( .A(A[75]), .B(B[75]), .CI(C[75]), 
        .S(S[75]), .CO(C[76]) );
  FA_1972 \FA_INST_0[0].FA_INST_1[76].FA_  ( .A(A[76]), .B(B[76]), .CI(C[76]), 
        .S(S[76]), .CO(C[77]) );
  FA_1971 \FA_INST_0[0].FA_INST_1[77].FA_  ( .A(A[77]), .B(B[77]), .CI(C[77]), 
        .S(S[77]), .CO(C[78]) );
  FA_1970 \FA_INST_0[0].FA_INST_1[78].FA_  ( .A(A[78]), .B(B[78]), .CI(C[78]), 
        .S(S[78]), .CO(C[79]) );
  FA_1969 \FA_INST_0[0].FA_INST_1[79].FA_  ( .A(A[79]), .B(B[79]), .CI(C[79]), 
        .S(S[79]), .CO(C[80]) );
  FA_1968 \FA_INST_0[0].FA_INST_1[80].FA_  ( .A(A[80]), .B(B[80]), .CI(C[80]), 
        .S(S[80]), .CO(C[81]) );
  FA_1967 \FA_INST_0[0].FA_INST_1[81].FA_  ( .A(A[81]), .B(B[81]), .CI(C[81]), 
        .S(S[81]), .CO(C[82]) );
  FA_1966 \FA_INST_0[0].FA_INST_1[82].FA_  ( .A(A[82]), .B(B[82]), .CI(C[82]), 
        .S(S[82]), .CO(C[83]) );
  FA_1965 \FA_INST_0[0].FA_INST_1[83].FA_  ( .A(A[83]), .B(B[83]), .CI(C[83]), 
        .S(S[83]), .CO(C[84]) );
  FA_1964 \FA_INST_0[0].FA_INST_1[84].FA_  ( .A(A[84]), .B(B[84]), .CI(C[84]), 
        .S(S[84]), .CO(C[85]) );
  FA_1963 \FA_INST_0[0].FA_INST_1[85].FA_  ( .A(A[85]), .B(B[85]), .CI(C[85]), 
        .S(S[85]), .CO(C[86]) );
  FA_1962 \FA_INST_0[0].FA_INST_1[86].FA_  ( .A(A[86]), .B(B[86]), .CI(C[86]), 
        .S(S[86]), .CO(C[87]) );
  FA_1961 \FA_INST_0[0].FA_INST_1[87].FA_  ( .A(A[87]), .B(B[87]), .CI(C[87]), 
        .S(S[87]), .CO(C[88]) );
  FA_1960 \FA_INST_0[0].FA_INST_1[88].FA_  ( .A(A[88]), .B(B[88]), .CI(C[88]), 
        .S(S[88]), .CO(C[89]) );
  FA_1959 \FA_INST_0[0].FA_INST_1[89].FA_  ( .A(A[89]), .B(B[89]), .CI(C[89]), 
        .S(S[89]), .CO(C[90]) );
  FA_1958 \FA_INST_0[0].FA_INST_1[90].FA_  ( .A(A[90]), .B(B[90]), .CI(C[90]), 
        .S(S[90]), .CO(C[91]) );
  FA_1957 \FA_INST_0[0].FA_INST_1[91].FA_  ( .A(A[91]), .B(B[91]), .CI(C[91]), 
        .S(S[91]), .CO(C[92]) );
  FA_1956 \FA_INST_0[0].FA_INST_1[92].FA_  ( .A(A[92]), .B(B[92]), .CI(C[92]), 
        .S(S[92]), .CO(C[93]) );
  FA_1955 \FA_INST_0[0].FA_INST_1[93].FA_  ( .A(A[93]), .B(B[93]), .CI(C[93]), 
        .S(S[93]), .CO(C[94]) );
  FA_1954 \FA_INST_0[0].FA_INST_1[94].FA_  ( .A(A[94]), .B(B[94]), .CI(C[94]), 
        .S(S[94]), .CO(C[95]) );
  FA_1953 \FA_INST_0[0].FA_INST_1[95].FA_  ( .A(A[95]), .B(B[95]), .CI(C[95]), 
        .S(S[95]), .CO(C[96]) );
  FA_1952 \FA_INST_0[0].FA_INST_1[96].FA_  ( .A(A[96]), .B(B[96]), .CI(C[96]), 
        .S(S[96]), .CO(C[97]) );
  FA_1951 \FA_INST_0[0].FA_INST_1[97].FA_  ( .A(A[97]), .B(B[97]), .CI(C[97]), 
        .S(S[97]), .CO(C[98]) );
  FA_1950 \FA_INST_0[0].FA_INST_1[98].FA_  ( .A(A[98]), .B(B[98]), .CI(C[98]), 
        .S(S[98]), .CO(C[99]) );
  FA_1949 \FA_INST_0[0].FA_INST_1[99].FA_  ( .A(A[99]), .B(B[99]), .CI(C[99]), 
        .S(S[99]), .CO(C[100]) );
  FA_1948 \FA_INST_0[0].FA_INST_1[100].FA_  ( .A(A[100]), .B(B[100]), .CI(
        C[100]), .S(S[100]), .CO(C[101]) );
  FA_1947 \FA_INST_0[0].FA_INST_1[101].FA_  ( .A(A[101]), .B(B[101]), .CI(
        C[101]), .S(S[101]), .CO(C[102]) );
  FA_1946 \FA_INST_0[0].FA_INST_1[102].FA_  ( .A(A[102]), .B(B[102]), .CI(
        C[102]), .S(S[102]), .CO(C[103]) );
  FA_1945 \FA_INST_0[0].FA_INST_1[103].FA_  ( .A(A[103]), .B(B[103]), .CI(
        C[103]), .S(S[103]), .CO(C[104]) );
  FA_1944 \FA_INST_0[0].FA_INST_1[104].FA_  ( .A(A[104]), .B(B[104]), .CI(
        C[104]), .S(S[104]), .CO(C[105]) );
  FA_1943 \FA_INST_0[0].FA_INST_1[105].FA_  ( .A(A[105]), .B(B[105]), .CI(
        C[105]), .S(S[105]), .CO(C[106]) );
  FA_1942 \FA_INST_0[0].FA_INST_1[106].FA_  ( .A(A[106]), .B(B[106]), .CI(
        C[106]), .S(S[106]), .CO(C[107]) );
  FA_1941 \FA_INST_0[0].FA_INST_1[107].FA_  ( .A(A[107]), .B(B[107]), .CI(
        C[107]), .S(S[107]), .CO(C[108]) );
  FA_1940 \FA_INST_0[0].FA_INST_1[108].FA_  ( .A(A[108]), .B(B[108]), .CI(
        C[108]), .S(S[108]), .CO(C[109]) );
  FA_1939 \FA_INST_0[0].FA_INST_1[109].FA_  ( .A(A[109]), .B(B[109]), .CI(
        C[109]), .S(S[109]), .CO(C[110]) );
  FA_1938 \FA_INST_0[0].FA_INST_1[110].FA_  ( .A(A[110]), .B(B[110]), .CI(
        C[110]), .S(S[110]), .CO(C[111]) );
  FA_1937 \FA_INST_0[0].FA_INST_1[111].FA_  ( .A(A[111]), .B(B[111]), .CI(
        C[111]), .S(S[111]), .CO(C[112]) );
  FA_1936 \FA_INST_0[0].FA_INST_1[112].FA_  ( .A(A[112]), .B(B[112]), .CI(
        C[112]), .S(S[112]), .CO(C[113]) );
  FA_1935 \FA_INST_0[0].FA_INST_1[113].FA_  ( .A(A[113]), .B(B[113]), .CI(
        C[113]), .S(S[113]), .CO(C[114]) );
  FA_1934 \FA_INST_0[0].FA_INST_1[114].FA_  ( .A(A[114]), .B(B[114]), .CI(
        C[114]), .S(S[114]), .CO(C[115]) );
  FA_1933 \FA_INST_0[0].FA_INST_1[115].FA_  ( .A(A[115]), .B(B[115]), .CI(
        C[115]), .S(S[115]), .CO(C[116]) );
  FA_1932 \FA_INST_0[0].FA_INST_1[116].FA_  ( .A(A[116]), .B(B[116]), .CI(
        C[116]), .S(S[116]), .CO(C[117]) );
  FA_1931 \FA_INST_0[0].FA_INST_1[117].FA_  ( .A(A[117]), .B(B[117]), .CI(
        C[117]), .S(S[117]), .CO(C[118]) );
  FA_1930 \FA_INST_0[0].FA_INST_1[118].FA_  ( .A(A[118]), .B(B[118]), .CI(
        C[118]), .S(S[118]), .CO(C[119]) );
  FA_1929 \FA_INST_0[0].FA_INST_1[119].FA_  ( .A(A[119]), .B(B[119]), .CI(
        C[119]), .S(S[119]), .CO(C[120]) );
  FA_1928 \FA_INST_0[0].FA_INST_1[120].FA_  ( .A(A[120]), .B(B[120]), .CI(
        C[120]), .S(S[120]), .CO(C[121]) );
  FA_1927 \FA_INST_0[0].FA_INST_1[121].FA_  ( .A(A[121]), .B(B[121]), .CI(
        C[121]), .S(S[121]), .CO(C[122]) );
  FA_1926 \FA_INST_0[0].FA_INST_1[122].FA_  ( .A(A[122]), .B(B[122]), .CI(
        C[122]), .S(S[122]), .CO(C[123]) );
  FA_1925 \FA_INST_0[0].FA_INST_1[123].FA_  ( .A(A[123]), .B(B[123]), .CI(
        C[123]), .S(S[123]), .CO(C[124]) );
  FA_1924 \FA_INST_0[0].FA_INST_1[124].FA_  ( .A(A[124]), .B(B[124]), .CI(
        C[124]), .S(S[124]), .CO(C[125]) );
  FA_1923 \FA_INST_0[0].FA_INST_1[125].FA_  ( .A(A[125]), .B(B[125]), .CI(
        C[125]), .S(S[125]), .CO(C[126]) );
  FA_1922 \FA_INST_0[0].FA_INST_1[126].FA_  ( .A(A[126]), .B(B[126]), .CI(
        C[126]), .S(S[126]), .CO(C[127]) );
  FA_1921 \FA_INST_0[0].FA_INST_1[127].FA_  ( .A(A[127]), .B(B[127]), .CI(
        C[127]), .S(S[127]), .CO(C[128]) );
  FA_1920 \FA_INST_0[0].FA_INST_1[128].FA_  ( .A(A[128]), .B(B[128]), .CI(
        C[128]), .S(S[128]), .CO(C[129]) );
  FA_1919 \FA_INST_0[0].FA_INST_1[129].FA_  ( .A(A[129]), .B(B[129]), .CI(
        C[129]), .S(S[129]), .CO(C[130]) );
  FA_1918 \FA_INST_0[0].FA_INST_1[130].FA_  ( .A(A[130]), .B(B[130]), .CI(
        C[130]), .S(S[130]), .CO(C[131]) );
  FA_1917 \FA_INST_0[0].FA_INST_1[131].FA_  ( .A(A[131]), .B(B[131]), .CI(
        C[131]), .S(S[131]), .CO(C[132]) );
  FA_1916 \FA_INST_0[0].FA_INST_1[132].FA_  ( .A(A[132]), .B(B[132]), .CI(
        C[132]), .S(S[132]), .CO(C[133]) );
  FA_1915 \FA_INST_0[0].FA_INST_1[133].FA_  ( .A(A[133]), .B(B[133]), .CI(
        C[133]), .S(S[133]), .CO(C[134]) );
  FA_1914 \FA_INST_0[0].FA_INST_1[134].FA_  ( .A(A[134]), .B(B[134]), .CI(
        C[134]), .S(S[134]), .CO(C[135]) );
  FA_1913 \FA_INST_0[0].FA_INST_1[135].FA_  ( .A(A[135]), .B(B[135]), .CI(
        C[135]), .S(S[135]), .CO(C[136]) );
  FA_1912 \FA_INST_0[0].FA_INST_1[136].FA_  ( .A(A[136]), .B(B[136]), .CI(
        C[136]), .S(S[136]), .CO(C[137]) );
  FA_1911 \FA_INST_0[0].FA_INST_1[137].FA_  ( .A(A[137]), .B(B[137]), .CI(
        C[137]), .S(S[137]), .CO(C[138]) );
  FA_1910 \FA_INST_0[0].FA_INST_1[138].FA_  ( .A(A[138]), .B(B[138]), .CI(
        C[138]), .S(S[138]), .CO(C[139]) );
  FA_1909 \FA_INST_0[0].FA_INST_1[139].FA_  ( .A(A[139]), .B(B[139]), .CI(
        C[139]), .S(S[139]), .CO(C[140]) );
  FA_1908 \FA_INST_0[0].FA_INST_1[140].FA_  ( .A(A[140]), .B(B[140]), .CI(
        C[140]), .S(S[140]), .CO(C[141]) );
  FA_1907 \FA_INST_0[0].FA_INST_1[141].FA_  ( .A(A[141]), .B(B[141]), .CI(
        C[141]), .S(S[141]), .CO(C[142]) );
  FA_1906 \FA_INST_0[0].FA_INST_1[142].FA_  ( .A(A[142]), .B(B[142]), .CI(
        C[142]), .S(S[142]), .CO(C[143]) );
  FA_1905 \FA_INST_0[0].FA_INST_1[143].FA_  ( .A(A[143]), .B(B[143]), .CI(
        C[143]), .S(S[143]), .CO(C[144]) );
  FA_1904 \FA_INST_0[0].FA_INST_1[144].FA_  ( .A(A[144]), .B(B[144]), .CI(
        C[144]), .S(S[144]), .CO(C[145]) );
  FA_1903 \FA_INST_0[0].FA_INST_1[145].FA_  ( .A(A[145]), .B(B[145]), .CI(
        C[145]), .S(S[145]), .CO(C[146]) );
  FA_1902 \FA_INST_0[0].FA_INST_1[146].FA_  ( .A(A[146]), .B(B[146]), .CI(
        C[146]), .S(S[146]), .CO(C[147]) );
  FA_1901 \FA_INST_0[0].FA_INST_1[147].FA_  ( .A(A[147]), .B(B[147]), .CI(
        C[147]), .S(S[147]), .CO(C[148]) );
  FA_1900 \FA_INST_0[0].FA_INST_1[148].FA_  ( .A(A[148]), .B(B[148]), .CI(
        C[148]), .S(S[148]), .CO(C[149]) );
  FA_1899 \FA_INST_0[0].FA_INST_1[149].FA_  ( .A(A[149]), .B(B[149]), .CI(
        C[149]), .S(S[149]), .CO(C[150]) );
  FA_1898 \FA_INST_0[0].FA_INST_1[150].FA_  ( .A(A[150]), .B(B[150]), .CI(
        C[150]), .S(S[150]), .CO(C[151]) );
  FA_1897 \FA_INST_0[0].FA_INST_1[151].FA_  ( .A(A[151]), .B(B[151]), .CI(
        C[151]), .S(S[151]), .CO(C[152]) );
  FA_1896 \FA_INST_0[0].FA_INST_1[152].FA_  ( .A(A[152]), .B(B[152]), .CI(
        C[152]), .S(S[152]), .CO(C[153]) );
  FA_1895 \FA_INST_0[0].FA_INST_1[153].FA_  ( .A(A[153]), .B(B[153]), .CI(
        C[153]), .S(S[153]), .CO(C[154]) );
  FA_1894 \FA_INST_0[0].FA_INST_1[154].FA_  ( .A(A[154]), .B(B[154]), .CI(
        C[154]), .S(S[154]), .CO(C[155]) );
  FA_1893 \FA_INST_0[0].FA_INST_1[155].FA_  ( .A(A[155]), .B(B[155]), .CI(
        C[155]), .S(S[155]), .CO(C[156]) );
  FA_1892 \FA_INST_0[0].FA_INST_1[156].FA_  ( .A(A[156]), .B(B[156]), .CI(
        C[156]), .S(S[156]), .CO(C[157]) );
  FA_1891 \FA_INST_0[0].FA_INST_1[157].FA_  ( .A(A[157]), .B(B[157]), .CI(
        C[157]), .S(S[157]), .CO(C[158]) );
  FA_1890 \FA_INST_0[0].FA_INST_1[158].FA_  ( .A(A[158]), .B(B[158]), .CI(
        C[158]), .S(S[158]), .CO(C[159]) );
  FA_1889 \FA_INST_0[0].FA_INST_1[159].FA_  ( .A(A[159]), .B(B[159]), .CI(
        C[159]), .S(S[159]), .CO(C[160]) );
  FA_1888 \FA_INST_0[0].FA_INST_1[160].FA_  ( .A(A[160]), .B(B[160]), .CI(
        C[160]), .S(S[160]), .CO(C[161]) );
  FA_1887 \FA_INST_0[0].FA_INST_1[161].FA_  ( .A(A[161]), .B(B[161]), .CI(
        C[161]), .S(S[161]), .CO(C[162]) );
  FA_1886 \FA_INST_0[0].FA_INST_1[162].FA_  ( .A(A[162]), .B(B[162]), .CI(
        C[162]), .S(S[162]), .CO(C[163]) );
  FA_1885 \FA_INST_0[0].FA_INST_1[163].FA_  ( .A(A[163]), .B(B[163]), .CI(
        C[163]), .S(S[163]), .CO(C[164]) );
  FA_1884 \FA_INST_0[0].FA_INST_1[164].FA_  ( .A(A[164]), .B(B[164]), .CI(
        C[164]), .S(S[164]), .CO(C[165]) );
  FA_1883 \FA_INST_0[0].FA_INST_1[165].FA_  ( .A(A[165]), .B(B[165]), .CI(
        C[165]), .S(S[165]), .CO(C[166]) );
  FA_1882 \FA_INST_0[0].FA_INST_1[166].FA_  ( .A(A[166]), .B(B[166]), .CI(
        C[166]), .S(S[166]), .CO(C[167]) );
  FA_1881 \FA_INST_0[0].FA_INST_1[167].FA_  ( .A(A[167]), .B(B[167]), .CI(
        C[167]), .S(S[167]), .CO(C[168]) );
  FA_1880 \FA_INST_0[0].FA_INST_1[168].FA_  ( .A(A[168]), .B(B[168]), .CI(
        C[168]), .S(S[168]), .CO(C[169]) );
  FA_1879 \FA_INST_0[0].FA_INST_1[169].FA_  ( .A(A[169]), .B(B[169]), .CI(
        C[169]), .S(S[169]), .CO(C[170]) );
  FA_1878 \FA_INST_0[0].FA_INST_1[170].FA_  ( .A(A[170]), .B(B[170]), .CI(
        C[170]), .S(S[170]), .CO(C[171]) );
  FA_1877 \FA_INST_0[0].FA_INST_1[171].FA_  ( .A(A[171]), .B(B[171]), .CI(
        C[171]), .S(S[171]), .CO(C[172]) );
  FA_1876 \FA_INST_0[0].FA_INST_1[172].FA_  ( .A(A[172]), .B(B[172]), .CI(
        C[172]), .S(S[172]), .CO(C[173]) );
  FA_1875 \FA_INST_0[0].FA_INST_1[173].FA_  ( .A(A[173]), .B(B[173]), .CI(
        C[173]), .S(S[173]), .CO(C[174]) );
  FA_1874 \FA_INST_0[0].FA_INST_1[174].FA_  ( .A(A[174]), .B(B[174]), .CI(
        C[174]), .S(S[174]), .CO(C[175]) );
  FA_1873 \FA_INST_0[0].FA_INST_1[175].FA_  ( .A(A[175]), .B(B[175]), .CI(
        C[175]), .S(S[175]), .CO(C[176]) );
  FA_1872 \FA_INST_0[0].FA_INST_1[176].FA_  ( .A(A[176]), .B(B[176]), .CI(
        C[176]), .S(S[176]), .CO(C[177]) );
  FA_1871 \FA_INST_0[0].FA_INST_1[177].FA_  ( .A(A[177]), .B(B[177]), .CI(
        C[177]), .S(S[177]), .CO(C[178]) );
  FA_1870 \FA_INST_0[0].FA_INST_1[178].FA_  ( .A(A[178]), .B(B[178]), .CI(
        C[178]), .S(S[178]), .CO(C[179]) );
  FA_1869 \FA_INST_0[0].FA_INST_1[179].FA_  ( .A(A[179]), .B(B[179]), .CI(
        C[179]), .S(S[179]), .CO(C[180]) );
  FA_1868 \FA_INST_0[0].FA_INST_1[180].FA_  ( .A(A[180]), .B(B[180]), .CI(
        C[180]), .S(S[180]), .CO(C[181]) );
  FA_1867 \FA_INST_0[0].FA_INST_1[181].FA_  ( .A(A[181]), .B(B[181]), .CI(
        C[181]), .S(S[181]), .CO(C[182]) );
  FA_1866 \FA_INST_0[0].FA_INST_1[182].FA_  ( .A(A[182]), .B(B[182]), .CI(
        C[182]), .S(S[182]), .CO(C[183]) );
  FA_1865 \FA_INST_0[0].FA_INST_1[183].FA_  ( .A(A[183]), .B(B[183]), .CI(
        C[183]), .S(S[183]), .CO(C[184]) );
  FA_1864 \FA_INST_0[0].FA_INST_1[184].FA_  ( .A(A[184]), .B(B[184]), .CI(
        C[184]), .S(S[184]), .CO(C[185]) );
  FA_1863 \FA_INST_0[0].FA_INST_1[185].FA_  ( .A(A[185]), .B(B[185]), .CI(
        C[185]), .S(S[185]), .CO(C[186]) );
  FA_1862 \FA_INST_0[0].FA_INST_1[186].FA_  ( .A(A[186]), .B(B[186]), .CI(
        C[186]), .S(S[186]), .CO(C[187]) );
  FA_1861 \FA_INST_0[0].FA_INST_1[187].FA_  ( .A(A[187]), .B(B[187]), .CI(
        C[187]), .S(S[187]), .CO(C[188]) );
  FA_1860 \FA_INST_0[0].FA_INST_1[188].FA_  ( .A(A[188]), .B(B[188]), .CI(
        C[188]), .S(S[188]), .CO(C[189]) );
  FA_1859 \FA_INST_0[0].FA_INST_1[189].FA_  ( .A(A[189]), .B(B[189]), .CI(
        C[189]), .S(S[189]), .CO(C[190]) );
  FA_1858 \FA_INST_0[0].FA_INST_1[190].FA_  ( .A(A[190]), .B(B[190]), .CI(
        C[190]), .S(S[190]), .CO(C[191]) );
  FA_1857 \FA_INST_0[0].FA_INST_1[191].FA_  ( .A(A[191]), .B(B[191]), .CI(
        C[191]), .S(S[191]), .CO(C[192]) );
  FA_1856 \FA_INST_0[0].FA_INST_1[192].FA_  ( .A(A[192]), .B(B[192]), .CI(
        C[192]), .S(S[192]), .CO(C[193]) );
  FA_1855 \FA_INST_0[0].FA_INST_1[193].FA_  ( .A(A[193]), .B(B[193]), .CI(
        C[193]), .S(S[193]), .CO(C[194]) );
  FA_1854 \FA_INST_0[0].FA_INST_1[194].FA_  ( .A(A[194]), .B(B[194]), .CI(
        C[194]), .S(S[194]), .CO(C[195]) );
  FA_1853 \FA_INST_0[0].FA_INST_1[195].FA_  ( .A(A[195]), .B(B[195]), .CI(
        C[195]), .S(S[195]), .CO(C[196]) );
  FA_1852 \FA_INST_0[0].FA_INST_1[196].FA_  ( .A(A[196]), .B(B[196]), .CI(
        C[196]), .S(S[196]), .CO(C[197]) );
  FA_1851 \FA_INST_0[0].FA_INST_1[197].FA_  ( .A(A[197]), .B(B[197]), .CI(
        C[197]), .S(S[197]), .CO(C[198]) );
  FA_1850 \FA_INST_0[0].FA_INST_1[198].FA_  ( .A(A[198]), .B(B[198]), .CI(
        C[198]), .S(S[198]), .CO(C[199]) );
  FA_1849 \FA_INST_0[0].FA_INST_1[199].FA_  ( .A(A[199]), .B(B[199]), .CI(
        C[199]), .S(S[199]), .CO(C[200]) );
  FA_1848 \FA_INST_0[0].FA_INST_1[200].FA_  ( .A(A[200]), .B(B[200]), .CI(
        C[200]), .S(S[200]), .CO(C[201]) );
  FA_1847 \FA_INST_0[0].FA_INST_1[201].FA_  ( .A(A[201]), .B(B[201]), .CI(
        C[201]), .S(S[201]), .CO(C[202]) );
  FA_1846 \FA_INST_0[0].FA_INST_1[202].FA_  ( .A(A[202]), .B(B[202]), .CI(
        C[202]), .S(S[202]), .CO(C[203]) );
  FA_1845 \FA_INST_0[0].FA_INST_1[203].FA_  ( .A(A[203]), .B(B[203]), .CI(
        C[203]), .S(S[203]), .CO(C[204]) );
  FA_1844 \FA_INST_0[0].FA_INST_1[204].FA_  ( .A(A[204]), .B(B[204]), .CI(
        C[204]), .S(S[204]), .CO(C[205]) );
  FA_1843 \FA_INST_0[0].FA_INST_1[205].FA_  ( .A(A[205]), .B(B[205]), .CI(
        C[205]), .S(S[205]), .CO(C[206]) );
  FA_1842 \FA_INST_0[0].FA_INST_1[206].FA_  ( .A(A[206]), .B(B[206]), .CI(
        C[206]), .S(S[206]), .CO(C[207]) );
  FA_1841 \FA_INST_0[0].FA_INST_1[207].FA_  ( .A(A[207]), .B(B[207]), .CI(
        C[207]), .S(S[207]), .CO(C[208]) );
  FA_1840 \FA_INST_0[0].FA_INST_1[208].FA_  ( .A(A[208]), .B(B[208]), .CI(
        C[208]), .S(S[208]), .CO(C[209]) );
  FA_1839 \FA_INST_0[0].FA_INST_1[209].FA_  ( .A(A[209]), .B(B[209]), .CI(
        C[209]), .S(S[209]), .CO(C[210]) );
  FA_1838 \FA_INST_0[0].FA_INST_1[210].FA_  ( .A(A[210]), .B(B[210]), .CI(
        C[210]), .S(S[210]), .CO(C[211]) );
  FA_1837 \FA_INST_0[0].FA_INST_1[211].FA_  ( .A(A[211]), .B(B[211]), .CI(
        C[211]), .S(S[211]), .CO(C[212]) );
  FA_1836 \FA_INST_0[0].FA_INST_1[212].FA_  ( .A(A[212]), .B(B[212]), .CI(
        C[212]), .S(S[212]), .CO(C[213]) );
  FA_1835 \FA_INST_0[0].FA_INST_1[213].FA_  ( .A(A[213]), .B(B[213]), .CI(
        C[213]), .S(S[213]), .CO(C[214]) );
  FA_1834 \FA_INST_0[0].FA_INST_1[214].FA_  ( .A(A[214]), .B(B[214]), .CI(
        C[214]), .S(S[214]), .CO(C[215]) );
  FA_1833 \FA_INST_0[0].FA_INST_1[215].FA_  ( .A(A[215]), .B(B[215]), .CI(
        C[215]), .S(S[215]), .CO(C[216]) );
  FA_1832 \FA_INST_0[0].FA_INST_1[216].FA_  ( .A(A[216]), .B(B[216]), .CI(
        C[216]), .S(S[216]), .CO(C[217]) );
  FA_1831 \FA_INST_0[0].FA_INST_1[217].FA_  ( .A(A[217]), .B(B[217]), .CI(
        C[217]), .S(S[217]), .CO(C[218]) );
  FA_1830 \FA_INST_0[0].FA_INST_1[218].FA_  ( .A(A[218]), .B(B[218]), .CI(
        C[218]), .S(S[218]), .CO(C[219]) );
  FA_1829 \FA_INST_0[0].FA_INST_1[219].FA_  ( .A(A[219]), .B(B[219]), .CI(
        C[219]), .S(S[219]), .CO(C[220]) );
  FA_1828 \FA_INST_0[0].FA_INST_1[220].FA_  ( .A(A[220]), .B(B[220]), .CI(
        C[220]), .S(S[220]), .CO(C[221]) );
  FA_1827 \FA_INST_0[0].FA_INST_1[221].FA_  ( .A(A[221]), .B(B[221]), .CI(
        C[221]), .S(S[221]), .CO(C[222]) );
  FA_1826 \FA_INST_0[0].FA_INST_1[222].FA_  ( .A(A[222]), .B(B[222]), .CI(
        C[222]), .S(S[222]), .CO(C[223]) );
  FA_1825 \FA_INST_0[0].FA_INST_1[223].FA_  ( .A(A[223]), .B(B[223]), .CI(
        C[223]), .S(S[223]), .CO(C[224]) );
  FA_1824 \FA_INST_0[0].FA_INST_1[224].FA_  ( .A(A[224]), .B(B[224]), .CI(
        C[224]), .S(S[224]), .CO(C[225]) );
  FA_1823 \FA_INST_0[0].FA_INST_1[225].FA_  ( .A(A[225]), .B(B[225]), .CI(
        C[225]), .S(S[225]), .CO(C[226]) );
  FA_1822 \FA_INST_0[0].FA_INST_1[226].FA_  ( .A(A[226]), .B(B[226]), .CI(
        C[226]), .S(S[226]), .CO(C[227]) );
  FA_1821 \FA_INST_0[0].FA_INST_1[227].FA_  ( .A(A[227]), .B(B[227]), .CI(
        C[227]), .S(S[227]), .CO(C[228]) );
  FA_1820 \FA_INST_0[0].FA_INST_1[228].FA_  ( .A(A[228]), .B(B[228]), .CI(
        C[228]), .S(S[228]), .CO(C[229]) );
  FA_1819 \FA_INST_0[0].FA_INST_1[229].FA_  ( .A(A[229]), .B(B[229]), .CI(
        C[229]), .S(S[229]), .CO(C[230]) );
  FA_1818 \FA_INST_0[0].FA_INST_1[230].FA_  ( .A(A[230]), .B(B[230]), .CI(
        C[230]), .S(S[230]), .CO(C[231]) );
  FA_1817 \FA_INST_0[0].FA_INST_1[231].FA_  ( .A(A[231]), .B(B[231]), .CI(
        C[231]), .S(S[231]), .CO(C[232]) );
  FA_1816 \FA_INST_0[0].FA_INST_1[232].FA_  ( .A(A[232]), .B(B[232]), .CI(
        C[232]), .S(S[232]), .CO(C[233]) );
  FA_1815 \FA_INST_0[0].FA_INST_1[233].FA_  ( .A(A[233]), .B(B[233]), .CI(
        C[233]), .S(S[233]), .CO(C[234]) );
  FA_1814 \FA_INST_0[0].FA_INST_1[234].FA_  ( .A(A[234]), .B(B[234]), .CI(
        C[234]), .S(S[234]), .CO(C[235]) );
  FA_1813 \FA_INST_0[0].FA_INST_1[235].FA_  ( .A(A[235]), .B(B[235]), .CI(
        C[235]), .S(S[235]), .CO(C[236]) );
  FA_1812 \FA_INST_0[0].FA_INST_1[236].FA_  ( .A(A[236]), .B(B[236]), .CI(
        C[236]), .S(S[236]), .CO(C[237]) );
  FA_1811 \FA_INST_0[0].FA_INST_1[237].FA_  ( .A(A[237]), .B(B[237]), .CI(
        C[237]), .S(S[237]), .CO(C[238]) );
  FA_1810 \FA_INST_0[0].FA_INST_1[238].FA_  ( .A(A[238]), .B(B[238]), .CI(
        C[238]), .S(S[238]), .CO(C[239]) );
  FA_1809 \FA_INST_0[0].FA_INST_1[239].FA_  ( .A(A[239]), .B(B[239]), .CI(
        C[239]), .S(S[239]), .CO(C[240]) );
  FA_1808 \FA_INST_0[0].FA_INST_1[240].FA_  ( .A(A[240]), .B(B[240]), .CI(
        C[240]), .S(S[240]), .CO(C[241]) );
  FA_1807 \FA_INST_0[0].FA_INST_1[241].FA_  ( .A(A[241]), .B(B[241]), .CI(
        C[241]), .S(S[241]), .CO(C[242]) );
  FA_1806 \FA_INST_0[0].FA_INST_1[242].FA_  ( .A(A[242]), .B(B[242]), .CI(
        C[242]), .S(S[242]), .CO(C[243]) );
  FA_1805 \FA_INST_0[0].FA_INST_1[243].FA_  ( .A(A[243]), .B(B[243]), .CI(
        C[243]), .S(S[243]), .CO(C[244]) );
  FA_1804 \FA_INST_0[0].FA_INST_1[244].FA_  ( .A(A[244]), .B(B[244]), .CI(
        C[244]), .S(S[244]), .CO(C[245]) );
  FA_1803 \FA_INST_0[0].FA_INST_1[245].FA_  ( .A(A[245]), .B(B[245]), .CI(
        C[245]), .S(S[245]), .CO(C[246]) );
  FA_1802 \FA_INST_0[0].FA_INST_1[246].FA_  ( .A(A[246]), .B(B[246]), .CI(
        C[246]), .S(S[246]), .CO(C[247]) );
  FA_1801 \FA_INST_0[0].FA_INST_1[247].FA_  ( .A(A[247]), .B(B[247]), .CI(
        C[247]), .S(S[247]), .CO(C[248]) );
  FA_1800 \FA_INST_0[0].FA_INST_1[248].FA_  ( .A(A[248]), .B(B[248]), .CI(
        C[248]), .S(S[248]), .CO(C[249]) );
  FA_1799 \FA_INST_0[0].FA_INST_1[249].FA_  ( .A(A[249]), .B(B[249]), .CI(
        C[249]), .S(S[249]), .CO(C[250]) );
  FA_1798 \FA_INST_0[0].FA_INST_1[250].FA_  ( .A(A[250]), .B(B[250]), .CI(
        C[250]), .S(S[250]), .CO(C[251]) );
  FA_1797 \FA_INST_0[0].FA_INST_1[251].FA_  ( .A(A[251]), .B(B[251]), .CI(
        C[251]), .S(S[251]), .CO(C[252]) );
  FA_1796 \FA_INST_0[0].FA_INST_1[252].FA_  ( .A(A[252]), .B(B[252]), .CI(
        C[252]), .S(S[252]), .CO(C[253]) );
  FA_1795 \FA_INST_0[0].FA_INST_1[253].FA_  ( .A(A[253]), .B(B[253]), .CI(
        C[253]), .S(S[253]), .CO(C[254]) );
  FA_1794 \FA_INST_0[0].FA_INST_1[254].FA_  ( .A(A[254]), .B(B[254]), .CI(
        C[254]), .S(S[254]), .CO(C[255]) );
  FA_1793 \FA_INST_0[0].FA_INST_1[255].FA_  ( .A(A[255]), .B(B[255]), .CI(
        C[255]), .S(S[255]), .CO(C[256]) );
  FA_1792 \FA_INST_0[0].FA_INST_1[256].FA_  ( .A(A[256]), .B(B[256]), .CI(
        C[256]), .S(S[256]), .CO(C[257]) );
  FA_1791 \FA_INST_0[0].FA_INST_1[257].FA_  ( .A(A[257]), .B(B[257]), .CI(
        C[257]), .S(S[257]), .CO(C[258]) );
  FA_1790 \FA_INST_0[0].FA_INST_1[258].FA_  ( .A(A[258]), .B(B[258]), .CI(
        C[258]), .S(S[258]), .CO(C[259]) );
  FA_1789 \FA_INST_0[0].FA_INST_1[259].FA_  ( .A(A[259]), .B(B[259]), .CI(
        C[259]), .S(S[259]), .CO(C[260]) );
  FA_1788 \FA_INST_0[0].FA_INST_1[260].FA_  ( .A(A[260]), .B(B[260]), .CI(
        C[260]), .S(S[260]), .CO(C[261]) );
  FA_1787 \FA_INST_0[0].FA_INST_1[261].FA_  ( .A(A[261]), .B(B[261]), .CI(
        C[261]), .S(S[261]), .CO(C[262]) );
  FA_1786 \FA_INST_0[0].FA_INST_1[262].FA_  ( .A(A[262]), .B(B[262]), .CI(
        C[262]), .S(S[262]), .CO(C[263]) );
  FA_1785 \FA_INST_0[0].FA_INST_1[263].FA_  ( .A(A[263]), .B(B[263]), .CI(
        C[263]), .S(S[263]), .CO(C[264]) );
  FA_1784 \FA_INST_0[0].FA_INST_1[264].FA_  ( .A(A[264]), .B(B[264]), .CI(
        C[264]), .S(S[264]), .CO(C[265]) );
  FA_1783 \FA_INST_0[0].FA_INST_1[265].FA_  ( .A(A[265]), .B(B[265]), .CI(
        C[265]), .S(S[265]), .CO(C[266]) );
  FA_1782 \FA_INST_0[0].FA_INST_1[266].FA_  ( .A(A[266]), .B(B[266]), .CI(
        C[266]), .S(S[266]), .CO(C[267]) );
  FA_1781 \FA_INST_0[0].FA_INST_1[267].FA_  ( .A(A[267]), .B(B[267]), .CI(
        C[267]), .S(S[267]), .CO(C[268]) );
  FA_1780 \FA_INST_0[0].FA_INST_1[268].FA_  ( .A(A[268]), .B(B[268]), .CI(
        C[268]), .S(S[268]), .CO(C[269]) );
  FA_1779 \FA_INST_0[0].FA_INST_1[269].FA_  ( .A(A[269]), .B(B[269]), .CI(
        C[269]), .S(S[269]), .CO(C[270]) );
  FA_1778 \FA_INST_0[0].FA_INST_1[270].FA_  ( .A(A[270]), .B(B[270]), .CI(
        C[270]), .S(S[270]), .CO(C[271]) );
  FA_1777 \FA_INST_0[0].FA_INST_1[271].FA_  ( .A(A[271]), .B(B[271]), .CI(
        C[271]), .S(S[271]), .CO(C[272]) );
  FA_1776 \FA_INST_0[0].FA_INST_1[272].FA_  ( .A(A[272]), .B(B[272]), .CI(
        C[272]), .S(S[272]), .CO(C[273]) );
  FA_1775 \FA_INST_0[0].FA_INST_1[273].FA_  ( .A(A[273]), .B(B[273]), .CI(
        C[273]), .S(S[273]), .CO(C[274]) );
  FA_1774 \FA_INST_0[0].FA_INST_1[274].FA_  ( .A(A[274]), .B(B[274]), .CI(
        C[274]), .S(S[274]), .CO(C[275]) );
  FA_1773 \FA_INST_0[0].FA_INST_1[275].FA_  ( .A(A[275]), .B(B[275]), .CI(
        C[275]), .S(S[275]), .CO(C[276]) );
  FA_1772 \FA_INST_0[0].FA_INST_1[276].FA_  ( .A(A[276]), .B(B[276]), .CI(
        C[276]), .S(S[276]), .CO(C[277]) );
  FA_1771 \FA_INST_0[0].FA_INST_1[277].FA_  ( .A(A[277]), .B(B[277]), .CI(
        C[277]), .S(S[277]), .CO(C[278]) );
  FA_1770 \FA_INST_0[0].FA_INST_1[278].FA_  ( .A(A[278]), .B(B[278]), .CI(
        C[278]), .S(S[278]), .CO(C[279]) );
  FA_1769 \FA_INST_0[0].FA_INST_1[279].FA_  ( .A(A[279]), .B(B[279]), .CI(
        C[279]), .S(S[279]), .CO(C[280]) );
  FA_1768 \FA_INST_0[0].FA_INST_1[280].FA_  ( .A(A[280]), .B(B[280]), .CI(
        C[280]), .S(S[280]), .CO(C[281]) );
  FA_1767 \FA_INST_0[0].FA_INST_1[281].FA_  ( .A(A[281]), .B(B[281]), .CI(
        C[281]), .S(S[281]), .CO(C[282]) );
  FA_1766 \FA_INST_0[0].FA_INST_1[282].FA_  ( .A(A[282]), .B(B[282]), .CI(
        C[282]), .S(S[282]), .CO(C[283]) );
  FA_1765 \FA_INST_0[0].FA_INST_1[283].FA_  ( .A(A[283]), .B(B[283]), .CI(
        C[283]), .S(S[283]), .CO(C[284]) );
  FA_1764 \FA_INST_0[0].FA_INST_1[284].FA_  ( .A(A[284]), .B(B[284]), .CI(
        C[284]), .S(S[284]), .CO(C[285]) );
  FA_1763 \FA_INST_0[0].FA_INST_1[285].FA_  ( .A(A[285]), .B(B[285]), .CI(
        C[285]), .S(S[285]), .CO(C[286]) );
  FA_1762 \FA_INST_0[0].FA_INST_1[286].FA_  ( .A(A[286]), .B(B[286]), .CI(
        C[286]), .S(S[286]), .CO(C[287]) );
  FA_1761 \FA_INST_0[0].FA_INST_1[287].FA_  ( .A(A[287]), .B(B[287]), .CI(
        C[287]), .S(S[287]), .CO(C[288]) );
  FA_1760 \FA_INST_0[0].FA_INST_1[288].FA_  ( .A(A[288]), .B(B[288]), .CI(
        C[288]), .S(S[288]), .CO(C[289]) );
  FA_1759 \FA_INST_0[0].FA_INST_1[289].FA_  ( .A(A[289]), .B(B[289]), .CI(
        C[289]), .S(S[289]), .CO(C[290]) );
  FA_1758 \FA_INST_0[0].FA_INST_1[290].FA_  ( .A(A[290]), .B(B[290]), .CI(
        C[290]), .S(S[290]), .CO(C[291]) );
  FA_1757 \FA_INST_0[0].FA_INST_1[291].FA_  ( .A(A[291]), .B(B[291]), .CI(
        C[291]), .S(S[291]), .CO(C[292]) );
  FA_1756 \FA_INST_0[0].FA_INST_1[292].FA_  ( .A(A[292]), .B(B[292]), .CI(
        C[292]), .S(S[292]), .CO(C[293]) );
  FA_1755 \FA_INST_0[0].FA_INST_1[293].FA_  ( .A(A[293]), .B(B[293]), .CI(
        C[293]), .S(S[293]), .CO(C[294]) );
  FA_1754 \FA_INST_0[0].FA_INST_1[294].FA_  ( .A(A[294]), .B(B[294]), .CI(
        C[294]), .S(S[294]), .CO(C[295]) );
  FA_1753 \FA_INST_0[0].FA_INST_1[295].FA_  ( .A(A[295]), .B(B[295]), .CI(
        C[295]), .S(S[295]), .CO(C[296]) );
  FA_1752 \FA_INST_0[0].FA_INST_1[296].FA_  ( .A(A[296]), .B(B[296]), .CI(
        C[296]), .S(S[296]), .CO(C[297]) );
  FA_1751 \FA_INST_0[0].FA_INST_1[297].FA_  ( .A(A[297]), .B(B[297]), .CI(
        C[297]), .S(S[297]), .CO(C[298]) );
  FA_1750 \FA_INST_0[0].FA_INST_1[298].FA_  ( .A(A[298]), .B(B[298]), .CI(
        C[298]), .S(S[298]), .CO(C[299]) );
  FA_1749 \FA_INST_0[0].FA_INST_1[299].FA_  ( .A(A[299]), .B(B[299]), .CI(
        C[299]), .S(S[299]), .CO(C[300]) );
  FA_1748 \FA_INST_0[0].FA_INST_1[300].FA_  ( .A(A[300]), .B(B[300]), .CI(
        C[300]), .S(S[300]), .CO(C[301]) );
  FA_1747 \FA_INST_0[0].FA_INST_1[301].FA_  ( .A(A[301]), .B(B[301]), .CI(
        C[301]), .S(S[301]), .CO(C[302]) );
  FA_1746 \FA_INST_0[0].FA_INST_1[302].FA_  ( .A(A[302]), .B(B[302]), .CI(
        C[302]), .S(S[302]), .CO(C[303]) );
  FA_1745 \FA_INST_0[0].FA_INST_1[303].FA_  ( .A(A[303]), .B(B[303]), .CI(
        C[303]), .S(S[303]), .CO(C[304]) );
  FA_1744 \FA_INST_0[0].FA_INST_1[304].FA_  ( .A(A[304]), .B(B[304]), .CI(
        C[304]), .S(S[304]), .CO(C[305]) );
  FA_1743 \FA_INST_0[0].FA_INST_1[305].FA_  ( .A(A[305]), .B(B[305]), .CI(
        C[305]), .S(S[305]), .CO(C[306]) );
  FA_1742 \FA_INST_0[0].FA_INST_1[306].FA_  ( .A(A[306]), .B(B[306]), .CI(
        C[306]), .S(S[306]), .CO(C[307]) );
  FA_1741 \FA_INST_0[0].FA_INST_1[307].FA_  ( .A(A[307]), .B(B[307]), .CI(
        C[307]), .S(S[307]), .CO(C[308]) );
  FA_1740 \FA_INST_0[0].FA_INST_1[308].FA_  ( .A(A[308]), .B(B[308]), .CI(
        C[308]), .S(S[308]), .CO(C[309]) );
  FA_1739 \FA_INST_0[0].FA_INST_1[309].FA_  ( .A(A[309]), .B(B[309]), .CI(
        C[309]), .S(S[309]), .CO(C[310]) );
  FA_1738 \FA_INST_0[0].FA_INST_1[310].FA_  ( .A(A[310]), .B(B[310]), .CI(
        C[310]), .S(S[310]), .CO(C[311]) );
  FA_1737 \FA_INST_0[0].FA_INST_1[311].FA_  ( .A(A[311]), .B(B[311]), .CI(
        C[311]), .S(S[311]), .CO(C[312]) );
  FA_1736 \FA_INST_0[0].FA_INST_1[312].FA_  ( .A(A[312]), .B(B[312]), .CI(
        C[312]), .S(S[312]), .CO(C[313]) );
  FA_1735 \FA_INST_0[0].FA_INST_1[313].FA_  ( .A(A[313]), .B(B[313]), .CI(
        C[313]), .S(S[313]), .CO(C[314]) );
  FA_1734 \FA_INST_0[0].FA_INST_1[314].FA_  ( .A(A[314]), .B(B[314]), .CI(
        C[314]), .S(S[314]), .CO(C[315]) );
  FA_1733 \FA_INST_0[0].FA_INST_1[315].FA_  ( .A(A[315]), .B(B[315]), .CI(
        C[315]), .S(S[315]), .CO(C[316]) );
  FA_1732 \FA_INST_0[0].FA_INST_1[316].FA_  ( .A(A[316]), .B(B[316]), .CI(
        C[316]), .S(S[316]), .CO(C[317]) );
  FA_1731 \FA_INST_0[0].FA_INST_1[317].FA_  ( .A(A[317]), .B(B[317]), .CI(
        C[317]), .S(S[317]), .CO(C[318]) );
  FA_1730 \FA_INST_0[0].FA_INST_1[318].FA_  ( .A(A[318]), .B(B[318]), .CI(
        C[318]), .S(S[318]), .CO(C[319]) );
  FA_1729 \FA_INST_0[0].FA_INST_1[319].FA_  ( .A(A[319]), .B(B[319]), .CI(
        C[319]), .S(S[319]), .CO(C[320]) );
  FA_1728 \FA_INST_0[0].FA_INST_1[320].FA_  ( .A(A[320]), .B(B[320]), .CI(
        C[320]), .S(S[320]), .CO(C[321]) );
  FA_1727 \FA_INST_0[0].FA_INST_1[321].FA_  ( .A(A[321]), .B(B[321]), .CI(
        C[321]), .S(S[321]), .CO(C[322]) );
  FA_1726 \FA_INST_0[0].FA_INST_1[322].FA_  ( .A(A[322]), .B(B[322]), .CI(
        C[322]), .S(S[322]), .CO(C[323]) );
  FA_1725 \FA_INST_0[0].FA_INST_1[323].FA_  ( .A(A[323]), .B(B[323]), .CI(
        C[323]), .S(S[323]), .CO(C[324]) );
  FA_1724 \FA_INST_0[0].FA_INST_1[324].FA_  ( .A(A[324]), .B(B[324]), .CI(
        C[324]), .S(S[324]), .CO(C[325]) );
  FA_1723 \FA_INST_0[0].FA_INST_1[325].FA_  ( .A(A[325]), .B(B[325]), .CI(
        C[325]), .S(S[325]), .CO(C[326]) );
  FA_1722 \FA_INST_0[0].FA_INST_1[326].FA_  ( .A(A[326]), .B(B[326]), .CI(
        C[326]), .S(S[326]), .CO(C[327]) );
  FA_1721 \FA_INST_0[0].FA_INST_1[327].FA_  ( .A(A[327]), .B(B[327]), .CI(
        C[327]), .S(S[327]), .CO(C[328]) );
  FA_1720 \FA_INST_0[0].FA_INST_1[328].FA_  ( .A(A[328]), .B(B[328]), .CI(
        C[328]), .S(S[328]), .CO(C[329]) );
  FA_1719 \FA_INST_0[0].FA_INST_1[329].FA_  ( .A(A[329]), .B(B[329]), .CI(
        C[329]), .S(S[329]), .CO(C[330]) );
  FA_1718 \FA_INST_0[0].FA_INST_1[330].FA_  ( .A(A[330]), .B(B[330]), .CI(
        C[330]), .S(S[330]), .CO(C[331]) );
  FA_1717 \FA_INST_0[0].FA_INST_1[331].FA_  ( .A(A[331]), .B(B[331]), .CI(
        C[331]), .S(S[331]), .CO(C[332]) );
  FA_1716 \FA_INST_0[0].FA_INST_1[332].FA_  ( .A(A[332]), .B(B[332]), .CI(
        C[332]), .S(S[332]), .CO(C[333]) );
  FA_1715 \FA_INST_0[0].FA_INST_1[333].FA_  ( .A(A[333]), .B(B[333]), .CI(
        C[333]), .S(S[333]), .CO(C[334]) );
  FA_1714 \FA_INST_0[0].FA_INST_1[334].FA_  ( .A(A[334]), .B(B[334]), .CI(
        C[334]), .S(S[334]), .CO(C[335]) );
  FA_1713 \FA_INST_0[0].FA_INST_1[335].FA_  ( .A(A[335]), .B(B[335]), .CI(
        C[335]), .S(S[335]), .CO(C[336]) );
  FA_1712 \FA_INST_0[0].FA_INST_1[336].FA_  ( .A(A[336]), .B(B[336]), .CI(
        C[336]), .S(S[336]), .CO(C[337]) );
  FA_1711 \FA_INST_0[0].FA_INST_1[337].FA_  ( .A(A[337]), .B(B[337]), .CI(
        C[337]), .S(S[337]), .CO(C[338]) );
  FA_1710 \FA_INST_0[0].FA_INST_1[338].FA_  ( .A(A[338]), .B(B[338]), .CI(
        C[338]), .S(S[338]), .CO(C[339]) );
  FA_1709 \FA_INST_0[0].FA_INST_1[339].FA_  ( .A(A[339]), .B(B[339]), .CI(
        C[339]), .S(S[339]), .CO(C[340]) );
  FA_1708 \FA_INST_0[0].FA_INST_1[340].FA_  ( .A(A[340]), .B(B[340]), .CI(
        C[340]), .S(S[340]), .CO(C[341]) );
  FA_1707 \FA_INST_0[0].FA_INST_1[341].FA_  ( .A(A[341]), .B(B[341]), .CI(
        C[341]), .S(S[341]), .CO(C[342]) );
  FA_1706 \FA_INST_0[0].FA_INST_1[342].FA_  ( .A(A[342]), .B(B[342]), .CI(
        C[342]), .S(S[342]), .CO(C[343]) );
  FA_1705 \FA_INST_0[0].FA_INST_1[343].FA_  ( .A(A[343]), .B(B[343]), .CI(
        C[343]), .S(S[343]), .CO(C[344]) );
  FA_1704 \FA_INST_0[0].FA_INST_1[344].FA_  ( .A(A[344]), .B(B[344]), .CI(
        C[344]), .S(S[344]), .CO(C[345]) );
  FA_1703 \FA_INST_0[0].FA_INST_1[345].FA_  ( .A(A[345]), .B(B[345]), .CI(
        C[345]), .S(S[345]), .CO(C[346]) );
  FA_1702 \FA_INST_0[0].FA_INST_1[346].FA_  ( .A(A[346]), .B(B[346]), .CI(
        C[346]), .S(S[346]), .CO(C[347]) );
  FA_1701 \FA_INST_0[0].FA_INST_1[347].FA_  ( .A(A[347]), .B(B[347]), .CI(
        C[347]), .S(S[347]), .CO(C[348]) );
  FA_1700 \FA_INST_0[0].FA_INST_1[348].FA_  ( .A(A[348]), .B(B[348]), .CI(
        C[348]), .S(S[348]), .CO(C[349]) );
  FA_1699 \FA_INST_0[0].FA_INST_1[349].FA_  ( .A(A[349]), .B(B[349]), .CI(
        C[349]), .S(S[349]), .CO(C[350]) );
  FA_1698 \FA_INST_0[0].FA_INST_1[350].FA_  ( .A(A[350]), .B(B[350]), .CI(
        C[350]), .S(S[350]), .CO(C[351]) );
  FA_1697 \FA_INST_0[0].FA_INST_1[351].FA_  ( .A(A[351]), .B(B[351]), .CI(
        C[351]), .S(S[351]), .CO(C[352]) );
  FA_1696 \FA_INST_0[0].FA_INST_1[352].FA_  ( .A(A[352]), .B(B[352]), .CI(
        C[352]), .S(S[352]), .CO(C[353]) );
  FA_1695 \FA_INST_0[0].FA_INST_1[353].FA_  ( .A(A[353]), .B(B[353]), .CI(
        C[353]), .S(S[353]), .CO(C[354]) );
  FA_1694 \FA_INST_0[0].FA_INST_1[354].FA_  ( .A(A[354]), .B(B[354]), .CI(
        C[354]), .S(S[354]), .CO(C[355]) );
  FA_1693 \FA_INST_0[0].FA_INST_1[355].FA_  ( .A(A[355]), .B(B[355]), .CI(
        C[355]), .S(S[355]), .CO(C[356]) );
  FA_1692 \FA_INST_0[0].FA_INST_1[356].FA_  ( .A(A[356]), .B(B[356]), .CI(
        C[356]), .S(S[356]), .CO(C[357]) );
  FA_1691 \FA_INST_0[0].FA_INST_1[357].FA_  ( .A(A[357]), .B(B[357]), .CI(
        C[357]), .S(S[357]), .CO(C[358]) );
  FA_1690 \FA_INST_0[0].FA_INST_1[358].FA_  ( .A(A[358]), .B(B[358]), .CI(
        C[358]), .S(S[358]), .CO(C[359]) );
  FA_1689 \FA_INST_0[0].FA_INST_1[359].FA_  ( .A(A[359]), .B(B[359]), .CI(
        C[359]), .S(S[359]), .CO(C[360]) );
  FA_1688 \FA_INST_0[0].FA_INST_1[360].FA_  ( .A(A[360]), .B(B[360]), .CI(
        C[360]), .S(S[360]), .CO(C[361]) );
  FA_1687 \FA_INST_0[0].FA_INST_1[361].FA_  ( .A(A[361]), .B(B[361]), .CI(
        C[361]), .S(S[361]), .CO(C[362]) );
  FA_1686 \FA_INST_0[0].FA_INST_1[362].FA_  ( .A(A[362]), .B(B[362]), .CI(
        C[362]), .S(S[362]), .CO(C[363]) );
  FA_1685 \FA_INST_0[0].FA_INST_1[363].FA_  ( .A(A[363]), .B(B[363]), .CI(
        C[363]), .S(S[363]), .CO(C[364]) );
  FA_1684 \FA_INST_0[0].FA_INST_1[364].FA_  ( .A(A[364]), .B(B[364]), .CI(
        C[364]), .S(S[364]), .CO(C[365]) );
  FA_1683 \FA_INST_0[0].FA_INST_1[365].FA_  ( .A(A[365]), .B(B[365]), .CI(
        C[365]), .S(S[365]), .CO(C[366]) );
  FA_1682 \FA_INST_0[0].FA_INST_1[366].FA_  ( .A(A[366]), .B(B[366]), .CI(
        C[366]), .S(S[366]), .CO(C[367]) );
  FA_1681 \FA_INST_0[0].FA_INST_1[367].FA_  ( .A(A[367]), .B(B[367]), .CI(
        C[367]), .S(S[367]), .CO(C[368]) );
  FA_1680 \FA_INST_0[0].FA_INST_1[368].FA_  ( .A(A[368]), .B(B[368]), .CI(
        C[368]), .S(S[368]), .CO(C[369]) );
  FA_1679 \FA_INST_0[0].FA_INST_1[369].FA_  ( .A(A[369]), .B(B[369]), .CI(
        C[369]), .S(S[369]), .CO(C[370]) );
  FA_1678 \FA_INST_0[0].FA_INST_1[370].FA_  ( .A(A[370]), .B(B[370]), .CI(
        C[370]), .S(S[370]), .CO(C[371]) );
  FA_1677 \FA_INST_0[0].FA_INST_1[371].FA_  ( .A(A[371]), .B(B[371]), .CI(
        C[371]), .S(S[371]), .CO(C[372]) );
  FA_1676 \FA_INST_0[0].FA_INST_1[372].FA_  ( .A(A[372]), .B(B[372]), .CI(
        C[372]), .S(S[372]), .CO(C[373]) );
  FA_1675 \FA_INST_0[0].FA_INST_1[373].FA_  ( .A(A[373]), .B(B[373]), .CI(
        C[373]), .S(S[373]), .CO(C[374]) );
  FA_1674 \FA_INST_0[0].FA_INST_1[374].FA_  ( .A(A[374]), .B(B[374]), .CI(
        C[374]), .S(S[374]), .CO(C[375]) );
  FA_1673 \FA_INST_0[0].FA_INST_1[375].FA_  ( .A(A[375]), .B(B[375]), .CI(
        C[375]), .S(S[375]), .CO(C[376]) );
  FA_1672 \FA_INST_0[0].FA_INST_1[376].FA_  ( .A(A[376]), .B(B[376]), .CI(
        C[376]), .S(S[376]), .CO(C[377]) );
  FA_1671 \FA_INST_0[0].FA_INST_1[377].FA_  ( .A(A[377]), .B(B[377]), .CI(
        C[377]), .S(S[377]), .CO(C[378]) );
  FA_1670 \FA_INST_0[0].FA_INST_1[378].FA_  ( .A(A[378]), .B(B[378]), .CI(
        C[378]), .S(S[378]), .CO(C[379]) );
  FA_1669 \FA_INST_0[0].FA_INST_1[379].FA_  ( .A(A[379]), .B(B[379]), .CI(
        C[379]), .S(S[379]), .CO(C[380]) );
  FA_1668 \FA_INST_0[0].FA_INST_1[380].FA_  ( .A(A[380]), .B(B[380]), .CI(
        C[380]), .S(S[380]), .CO(C[381]) );
  FA_1667 \FA_INST_0[0].FA_INST_1[381].FA_  ( .A(A[381]), .B(B[381]), .CI(
        C[381]), .S(S[381]), .CO(C[382]) );
  FA_1666 \FA_INST_0[0].FA_INST_1[382].FA_  ( .A(A[382]), .B(B[382]), .CI(
        C[382]), .S(S[382]), .CO(C[383]) );
  FA_1665 \FA_INST_0[0].FA_INST_1[383].FA_  ( .A(A[383]), .B(B[383]), .CI(
        C[383]), .S(S[383]), .CO(C[384]) );
  FA_1664 \FA_INST_0[0].FA_INST_1[384].FA_  ( .A(A[384]), .B(B[384]), .CI(
        C[384]), .S(S[384]), .CO(C[385]) );
  FA_1663 \FA_INST_0[0].FA_INST_1[385].FA_  ( .A(A[385]), .B(B[385]), .CI(
        C[385]), .S(S[385]), .CO(C[386]) );
  FA_1662 \FA_INST_0[0].FA_INST_1[386].FA_  ( .A(A[386]), .B(B[386]), .CI(
        C[386]), .S(S[386]), .CO(C[387]) );
  FA_1661 \FA_INST_0[0].FA_INST_1[387].FA_  ( .A(A[387]), .B(B[387]), .CI(
        C[387]), .S(S[387]), .CO(C[388]) );
  FA_1660 \FA_INST_0[0].FA_INST_1[388].FA_  ( .A(A[388]), .B(B[388]), .CI(
        C[388]), .S(S[388]), .CO(C[389]) );
  FA_1659 \FA_INST_0[0].FA_INST_1[389].FA_  ( .A(A[389]), .B(B[389]), .CI(
        C[389]), .S(S[389]), .CO(C[390]) );
  FA_1658 \FA_INST_0[0].FA_INST_1[390].FA_  ( .A(A[390]), .B(B[390]), .CI(
        C[390]), .S(S[390]), .CO(C[391]) );
  FA_1657 \FA_INST_0[0].FA_INST_1[391].FA_  ( .A(A[391]), .B(B[391]), .CI(
        C[391]), .S(S[391]), .CO(C[392]) );
  FA_1656 \FA_INST_0[0].FA_INST_1[392].FA_  ( .A(A[392]), .B(B[392]), .CI(
        C[392]), .S(S[392]), .CO(C[393]) );
  FA_1655 \FA_INST_0[0].FA_INST_1[393].FA_  ( .A(A[393]), .B(B[393]), .CI(
        C[393]), .S(S[393]), .CO(C[394]) );
  FA_1654 \FA_INST_0[0].FA_INST_1[394].FA_  ( .A(A[394]), .B(B[394]), .CI(
        C[394]), .S(S[394]), .CO(C[395]) );
  FA_1653 \FA_INST_0[0].FA_INST_1[395].FA_  ( .A(A[395]), .B(B[395]), .CI(
        C[395]), .S(S[395]), .CO(C[396]) );
  FA_1652 \FA_INST_0[0].FA_INST_1[396].FA_  ( .A(A[396]), .B(B[396]), .CI(
        C[396]), .S(S[396]), .CO(C[397]) );
  FA_1651 \FA_INST_0[0].FA_INST_1[397].FA_  ( .A(A[397]), .B(B[397]), .CI(
        C[397]), .S(S[397]), .CO(C[398]) );
  FA_1650 \FA_INST_0[0].FA_INST_1[398].FA_  ( .A(A[398]), .B(B[398]), .CI(
        C[398]), .S(S[398]), .CO(C[399]) );
  FA_1649 \FA_INST_0[0].FA_INST_1[399].FA_  ( .A(A[399]), .B(B[399]), .CI(
        C[399]), .S(S[399]), .CO(C[400]) );
  FA_1648 \FA_INST_0[0].FA_INST_1[400].FA_  ( .A(A[400]), .B(B[400]), .CI(
        C[400]), .S(S[400]), .CO(C[401]) );
  FA_1647 \FA_INST_0[0].FA_INST_1[401].FA_  ( .A(A[401]), .B(B[401]), .CI(
        C[401]), .S(S[401]), .CO(C[402]) );
  FA_1646 \FA_INST_0[0].FA_INST_1[402].FA_  ( .A(A[402]), .B(B[402]), .CI(
        C[402]), .S(S[402]), .CO(C[403]) );
  FA_1645 \FA_INST_0[0].FA_INST_1[403].FA_  ( .A(A[403]), .B(B[403]), .CI(
        C[403]), .S(S[403]), .CO(C[404]) );
  FA_1644 \FA_INST_0[0].FA_INST_1[404].FA_  ( .A(A[404]), .B(B[404]), .CI(
        C[404]), .S(S[404]), .CO(C[405]) );
  FA_1643 \FA_INST_0[0].FA_INST_1[405].FA_  ( .A(A[405]), .B(B[405]), .CI(
        C[405]), .S(S[405]), .CO(C[406]) );
  FA_1642 \FA_INST_0[0].FA_INST_1[406].FA_  ( .A(A[406]), .B(B[406]), .CI(
        C[406]), .S(S[406]), .CO(C[407]) );
  FA_1641 \FA_INST_0[0].FA_INST_1[407].FA_  ( .A(A[407]), .B(B[407]), .CI(
        C[407]), .S(S[407]), .CO(C[408]) );
  FA_1640 \FA_INST_0[0].FA_INST_1[408].FA_  ( .A(A[408]), .B(B[408]), .CI(
        C[408]), .S(S[408]), .CO(C[409]) );
  FA_1639 \FA_INST_0[0].FA_INST_1[409].FA_  ( .A(A[409]), .B(B[409]), .CI(
        C[409]), .S(S[409]), .CO(C[410]) );
  FA_1638 \FA_INST_0[0].FA_INST_1[410].FA_  ( .A(A[410]), .B(B[410]), .CI(
        C[410]), .S(S[410]), .CO(C[411]) );
  FA_1637 \FA_INST_0[0].FA_INST_1[411].FA_  ( .A(A[411]), .B(B[411]), .CI(
        C[411]), .S(S[411]), .CO(C[412]) );
  FA_1636 \FA_INST_0[0].FA_INST_1[412].FA_  ( .A(A[412]), .B(B[412]), .CI(
        C[412]), .S(S[412]), .CO(C[413]) );
  FA_1635 \FA_INST_0[0].FA_INST_1[413].FA_  ( .A(A[413]), .B(B[413]), .CI(
        C[413]), .S(S[413]), .CO(C[414]) );
  FA_1634 \FA_INST_0[0].FA_INST_1[414].FA_  ( .A(A[414]), .B(B[414]), .CI(
        C[414]), .S(S[414]), .CO(C[415]) );
  FA_1633 \FA_INST_0[0].FA_INST_1[415].FA_  ( .A(A[415]), .B(B[415]), .CI(
        C[415]), .S(S[415]), .CO(C[416]) );
  FA_1632 \FA_INST_0[0].FA_INST_1[416].FA_  ( .A(A[416]), .B(B[416]), .CI(
        C[416]), .S(S[416]), .CO(C[417]) );
  FA_1631 \FA_INST_0[0].FA_INST_1[417].FA_  ( .A(A[417]), .B(B[417]), .CI(
        C[417]), .S(S[417]), .CO(C[418]) );
  FA_1630 \FA_INST_0[0].FA_INST_1[418].FA_  ( .A(A[418]), .B(B[418]), .CI(
        C[418]), .S(S[418]), .CO(C[419]) );
  FA_1629 \FA_INST_0[0].FA_INST_1[419].FA_  ( .A(A[419]), .B(B[419]), .CI(
        C[419]), .S(S[419]), .CO(C[420]) );
  FA_1628 \FA_INST_0[0].FA_INST_1[420].FA_  ( .A(A[420]), .B(B[420]), .CI(
        C[420]), .S(S[420]), .CO(C[421]) );
  FA_1627 \FA_INST_0[0].FA_INST_1[421].FA_  ( .A(A[421]), .B(B[421]), .CI(
        C[421]), .S(S[421]), .CO(C[422]) );
  FA_1626 \FA_INST_0[0].FA_INST_1[422].FA_  ( .A(A[422]), .B(B[422]), .CI(
        C[422]), .S(S[422]), .CO(C[423]) );
  FA_1625 \FA_INST_0[0].FA_INST_1[423].FA_  ( .A(A[423]), .B(B[423]), .CI(
        C[423]), .S(S[423]), .CO(C[424]) );
  FA_1624 \FA_INST_0[0].FA_INST_1[424].FA_  ( .A(A[424]), .B(B[424]), .CI(
        C[424]), .S(S[424]), .CO(C[425]) );
  FA_1623 \FA_INST_0[0].FA_INST_1[425].FA_  ( .A(A[425]), .B(B[425]), .CI(
        C[425]), .S(S[425]), .CO(C[426]) );
  FA_1622 \FA_INST_0[0].FA_INST_1[426].FA_  ( .A(A[426]), .B(B[426]), .CI(
        C[426]), .S(S[426]), .CO(C[427]) );
  FA_1621 \FA_INST_0[0].FA_INST_1[427].FA_  ( .A(A[427]), .B(B[427]), .CI(
        C[427]), .S(S[427]), .CO(C[428]) );
  FA_1620 \FA_INST_0[0].FA_INST_1[428].FA_  ( .A(A[428]), .B(B[428]), .CI(
        C[428]), .S(S[428]), .CO(C[429]) );
  FA_1619 \FA_INST_0[0].FA_INST_1[429].FA_  ( .A(A[429]), .B(B[429]), .CI(
        C[429]), .S(S[429]), .CO(C[430]) );
  FA_1618 \FA_INST_0[0].FA_INST_1[430].FA_  ( .A(A[430]), .B(B[430]), .CI(
        C[430]), .S(S[430]), .CO(C[431]) );
  FA_1617 \FA_INST_0[0].FA_INST_1[431].FA_  ( .A(A[431]), .B(B[431]), .CI(
        C[431]), .S(S[431]), .CO(C[432]) );
  FA_1616 \FA_INST_0[0].FA_INST_1[432].FA_  ( .A(A[432]), .B(B[432]), .CI(
        C[432]), .S(S[432]), .CO(C[433]) );
  FA_1615 \FA_INST_0[0].FA_INST_1[433].FA_  ( .A(A[433]), .B(B[433]), .CI(
        C[433]), .S(S[433]), .CO(C[434]) );
  FA_1614 \FA_INST_0[0].FA_INST_1[434].FA_  ( .A(A[434]), .B(B[434]), .CI(
        C[434]), .S(S[434]), .CO(C[435]) );
  FA_1613 \FA_INST_0[0].FA_INST_1[435].FA_  ( .A(A[435]), .B(B[435]), .CI(
        C[435]), .S(S[435]), .CO(C[436]) );
  FA_1612 \FA_INST_0[0].FA_INST_1[436].FA_  ( .A(A[436]), .B(B[436]), .CI(
        C[436]), .S(S[436]), .CO(C[437]) );
  FA_1611 \FA_INST_0[0].FA_INST_1[437].FA_  ( .A(A[437]), .B(B[437]), .CI(
        C[437]), .S(S[437]), .CO(C[438]) );
  FA_1610 \FA_INST_0[0].FA_INST_1[438].FA_  ( .A(A[438]), .B(B[438]), .CI(
        C[438]), .S(S[438]), .CO(C[439]) );
  FA_1609 \FA_INST_0[0].FA_INST_1[439].FA_  ( .A(A[439]), .B(B[439]), .CI(
        C[439]), .S(S[439]), .CO(C[440]) );
  FA_1608 \FA_INST_0[0].FA_INST_1[440].FA_  ( .A(A[440]), .B(B[440]), .CI(
        C[440]), .S(S[440]), .CO(C[441]) );
  FA_1607 \FA_INST_0[0].FA_INST_1[441].FA_  ( .A(A[441]), .B(B[441]), .CI(
        C[441]), .S(S[441]), .CO(C[442]) );
  FA_1606 \FA_INST_0[0].FA_INST_1[442].FA_  ( .A(A[442]), .B(B[442]), .CI(
        C[442]), .S(S[442]), .CO(C[443]) );
  FA_1605 \FA_INST_0[0].FA_INST_1[443].FA_  ( .A(A[443]), .B(B[443]), .CI(
        C[443]), .S(S[443]), .CO(C[444]) );
  FA_1604 \FA_INST_0[0].FA_INST_1[444].FA_  ( .A(A[444]), .B(B[444]), .CI(
        C[444]), .S(S[444]), .CO(C[445]) );
  FA_1603 \FA_INST_0[0].FA_INST_1[445].FA_  ( .A(A[445]), .B(B[445]), .CI(
        C[445]), .S(S[445]), .CO(C[446]) );
  FA_1602 \FA_INST_0[0].FA_INST_1[446].FA_  ( .A(A[446]), .B(B[446]), .CI(
        C[446]), .S(S[446]), .CO(C[447]) );
  FA_1601 \FA_INST_0[0].FA_INST_1[447].FA_  ( .A(A[447]), .B(B[447]), .CI(
        C[447]), .S(S[447]), .CO(C[448]) );
  FA_1600 \FA_INST_0[0].FA_INST_1[448].FA_  ( .A(A[448]), .B(B[448]), .CI(
        C[448]), .S(S[448]), .CO(C[449]) );
  FA_1599 \FA_INST_0[0].FA_INST_1[449].FA_  ( .A(A[449]), .B(B[449]), .CI(
        C[449]), .S(S[449]), .CO(C[450]) );
  FA_1598 \FA_INST_0[0].FA_INST_1[450].FA_  ( .A(A[450]), .B(B[450]), .CI(
        C[450]), .S(S[450]), .CO(C[451]) );
  FA_1597 \FA_INST_0[0].FA_INST_1[451].FA_  ( .A(A[451]), .B(B[451]), .CI(
        C[451]), .S(S[451]), .CO(C[452]) );
  FA_1596 \FA_INST_0[0].FA_INST_1[452].FA_  ( .A(A[452]), .B(B[452]), .CI(
        C[452]), .S(S[452]), .CO(C[453]) );
  FA_1595 \FA_INST_0[0].FA_INST_1[453].FA_  ( .A(A[453]), .B(B[453]), .CI(
        C[453]), .S(S[453]), .CO(C[454]) );
  FA_1594 \FA_INST_0[0].FA_INST_1[454].FA_  ( .A(A[454]), .B(B[454]), .CI(
        C[454]), .S(S[454]), .CO(C[455]) );
  FA_1593 \FA_INST_0[0].FA_INST_1[455].FA_  ( .A(A[455]), .B(B[455]), .CI(
        C[455]), .S(S[455]), .CO(C[456]) );
  FA_1592 \FA_INST_0[0].FA_INST_1[456].FA_  ( .A(A[456]), .B(B[456]), .CI(
        C[456]), .S(S[456]), .CO(C[457]) );
  FA_1591 \FA_INST_0[0].FA_INST_1[457].FA_  ( .A(A[457]), .B(B[457]), .CI(
        C[457]), .S(S[457]), .CO(C[458]) );
  FA_1590 \FA_INST_0[0].FA_INST_1[458].FA_  ( .A(A[458]), .B(B[458]), .CI(
        C[458]), .S(S[458]), .CO(C[459]) );
  FA_1589 \FA_INST_0[0].FA_INST_1[459].FA_  ( .A(A[459]), .B(B[459]), .CI(
        C[459]), .S(S[459]), .CO(C[460]) );
  FA_1588 \FA_INST_0[0].FA_INST_1[460].FA_  ( .A(A[460]), .B(B[460]), .CI(
        C[460]), .S(S[460]), .CO(C[461]) );
  FA_1587 \FA_INST_0[0].FA_INST_1[461].FA_  ( .A(A[461]), .B(B[461]), .CI(
        C[461]), .S(S[461]), .CO(C[462]) );
  FA_1586 \FA_INST_0[0].FA_INST_1[462].FA_  ( .A(A[462]), .B(B[462]), .CI(
        C[462]), .S(S[462]), .CO(C[463]) );
  FA_1585 \FA_INST_0[0].FA_INST_1[463].FA_  ( .A(A[463]), .B(B[463]), .CI(
        C[463]), .S(S[463]), .CO(C[464]) );
  FA_1584 \FA_INST_0[0].FA_INST_1[464].FA_  ( .A(A[464]), .B(B[464]), .CI(
        C[464]), .S(S[464]), .CO(C[465]) );
  FA_1583 \FA_INST_0[0].FA_INST_1[465].FA_  ( .A(A[465]), .B(B[465]), .CI(
        C[465]), .S(S[465]), .CO(C[466]) );
  FA_1582 \FA_INST_0[0].FA_INST_1[466].FA_  ( .A(A[466]), .B(B[466]), .CI(
        C[466]), .S(S[466]), .CO(C[467]) );
  FA_1581 \FA_INST_0[0].FA_INST_1[467].FA_  ( .A(A[467]), .B(B[467]), .CI(
        C[467]), .S(S[467]), .CO(C[468]) );
  FA_1580 \FA_INST_0[0].FA_INST_1[468].FA_  ( .A(A[468]), .B(B[468]), .CI(
        C[468]), .S(S[468]), .CO(C[469]) );
  FA_1579 \FA_INST_0[0].FA_INST_1[469].FA_  ( .A(A[469]), .B(B[469]), .CI(
        C[469]), .S(S[469]), .CO(C[470]) );
  FA_1578 \FA_INST_0[0].FA_INST_1[470].FA_  ( .A(A[470]), .B(B[470]), .CI(
        C[470]), .S(S[470]), .CO(C[471]) );
  FA_1577 \FA_INST_0[0].FA_INST_1[471].FA_  ( .A(A[471]), .B(B[471]), .CI(
        C[471]), .S(S[471]), .CO(C[472]) );
  FA_1576 \FA_INST_0[0].FA_INST_1[472].FA_  ( .A(A[472]), .B(B[472]), .CI(
        C[472]), .S(S[472]), .CO(C[473]) );
  FA_1575 \FA_INST_0[0].FA_INST_1[473].FA_  ( .A(A[473]), .B(B[473]), .CI(
        C[473]), .S(S[473]), .CO(C[474]) );
  FA_1574 \FA_INST_0[0].FA_INST_1[474].FA_  ( .A(A[474]), .B(B[474]), .CI(
        C[474]), .S(S[474]), .CO(C[475]) );
  FA_1573 \FA_INST_0[0].FA_INST_1[475].FA_  ( .A(A[475]), .B(B[475]), .CI(
        C[475]), .S(S[475]), .CO(C[476]) );
  FA_1572 \FA_INST_0[0].FA_INST_1[476].FA_  ( .A(A[476]), .B(B[476]), .CI(
        C[476]), .S(S[476]), .CO(C[477]) );
  FA_1571 \FA_INST_0[0].FA_INST_1[477].FA_  ( .A(A[477]), .B(B[477]), .CI(
        C[477]), .S(S[477]), .CO(C[478]) );
  FA_1570 \FA_INST_0[0].FA_INST_1[478].FA_  ( .A(A[478]), .B(B[478]), .CI(
        C[478]), .S(S[478]), .CO(C[479]) );
  FA_1569 \FA_INST_0[0].FA_INST_1[479].FA_  ( .A(A[479]), .B(B[479]), .CI(
        C[479]), .S(S[479]), .CO(C[480]) );
  FA_1568 \FA_INST_0[0].FA_INST_1[480].FA_  ( .A(A[480]), .B(B[480]), .CI(
        C[480]), .S(S[480]), .CO(C[481]) );
  FA_1567 \FA_INST_0[0].FA_INST_1[481].FA_  ( .A(A[481]), .B(B[481]), .CI(
        C[481]), .S(S[481]), .CO(C[482]) );
  FA_1566 \FA_INST_0[0].FA_INST_1[482].FA_  ( .A(A[482]), .B(B[482]), .CI(
        C[482]), .S(S[482]), .CO(C[483]) );
  FA_1565 \FA_INST_0[0].FA_INST_1[483].FA_  ( .A(A[483]), .B(B[483]), .CI(
        C[483]), .S(S[483]), .CO(C[484]) );
  FA_1564 \FA_INST_0[0].FA_INST_1[484].FA_  ( .A(A[484]), .B(B[484]), .CI(
        C[484]), .S(S[484]), .CO(C[485]) );
  FA_1563 \FA_INST_0[0].FA_INST_1[485].FA_  ( .A(A[485]), .B(B[485]), .CI(
        C[485]), .S(S[485]), .CO(C[486]) );
  FA_1562 \FA_INST_0[0].FA_INST_1[486].FA_  ( .A(A[486]), .B(B[486]), .CI(
        C[486]), .S(S[486]), .CO(C[487]) );
  FA_1561 \FA_INST_0[0].FA_INST_1[487].FA_  ( .A(A[487]), .B(B[487]), .CI(
        C[487]), .S(S[487]), .CO(C[488]) );
  FA_1560 \FA_INST_0[0].FA_INST_1[488].FA_  ( .A(A[488]), .B(B[488]), .CI(
        C[488]), .S(S[488]), .CO(C[489]) );
  FA_1559 \FA_INST_0[0].FA_INST_1[489].FA_  ( .A(A[489]), .B(B[489]), .CI(
        C[489]), .S(S[489]), .CO(C[490]) );
  FA_1558 \FA_INST_0[0].FA_INST_1[490].FA_  ( .A(A[490]), .B(B[490]), .CI(
        C[490]), .S(S[490]), .CO(C[491]) );
  FA_1557 \FA_INST_0[0].FA_INST_1[491].FA_  ( .A(A[491]), .B(B[491]), .CI(
        C[491]), .S(S[491]), .CO(C[492]) );
  FA_1556 \FA_INST_0[0].FA_INST_1[492].FA_  ( .A(A[492]), .B(B[492]), .CI(
        C[492]), .S(S[492]), .CO(C[493]) );
  FA_1555 \FA_INST_0[0].FA_INST_1[493].FA_  ( .A(A[493]), .B(B[493]), .CI(
        C[493]), .S(S[493]), .CO(C[494]) );
  FA_1554 \FA_INST_0[0].FA_INST_1[494].FA_  ( .A(A[494]), .B(B[494]), .CI(
        C[494]), .S(S[494]), .CO(C[495]) );
  FA_1553 \FA_INST_0[0].FA_INST_1[495].FA_  ( .A(A[495]), .B(B[495]), .CI(
        C[495]), .S(S[495]), .CO(C[496]) );
  FA_1552 \FA_INST_0[0].FA_INST_1[496].FA_  ( .A(A[496]), .B(B[496]), .CI(
        C[496]), .S(S[496]), .CO(C[497]) );
  FA_1551 \FA_INST_0[0].FA_INST_1[497].FA_  ( .A(A[497]), .B(B[497]), .CI(
        C[497]), .S(S[497]), .CO(C[498]) );
  FA_1550 \FA_INST_0[0].FA_INST_1[498].FA_  ( .A(A[498]), .B(B[498]), .CI(
        C[498]), .S(S[498]), .CO(C[499]) );
  FA_1549 \FA_INST_0[0].FA_INST_1[499].FA_  ( .A(A[499]), .B(B[499]), .CI(
        C[499]), .S(S[499]), .CO(C[500]) );
  FA_1548 \FA_INST_0[0].FA_INST_1[500].FA_  ( .A(A[500]), .B(B[500]), .CI(
        C[500]), .S(S[500]), .CO(C[501]) );
  FA_1547 \FA_INST_0[0].FA_INST_1[501].FA_  ( .A(A[501]), .B(B[501]), .CI(
        C[501]), .S(S[501]), .CO(C[502]) );
  FA_1546 \FA_INST_0[0].FA_INST_1[502].FA_  ( .A(A[502]), .B(B[502]), .CI(
        C[502]), .S(S[502]), .CO(C[503]) );
  FA_1545 \FA_INST_0[0].FA_INST_1[503].FA_  ( .A(A[503]), .B(B[503]), .CI(
        C[503]), .S(S[503]), .CO(C[504]) );
  FA_1544 \FA_INST_0[0].FA_INST_1[504].FA_  ( .A(A[504]), .B(B[504]), .CI(
        C[504]), .S(S[504]), .CO(C[505]) );
  FA_1543 \FA_INST_0[0].FA_INST_1[505].FA_  ( .A(A[505]), .B(B[505]), .CI(
        C[505]), .S(S[505]), .CO(C[506]) );
  FA_1542 \FA_INST_0[0].FA_INST_1[506].FA_  ( .A(A[506]), .B(B[506]), .CI(
        C[506]), .S(S[506]), .CO(C[507]) );
  FA_1541 \FA_INST_0[0].FA_INST_1[507].FA_  ( .A(A[507]), .B(B[507]), .CI(
        C[507]), .S(S[507]), .CO(C[508]) );
  FA_1540 \FA_INST_0[0].FA_INST_1[508].FA_  ( .A(A[508]), .B(B[508]), .CI(
        C[508]), .S(S[508]), .CO(C[509]) );
  FA_1539 \FA_INST_0[0].FA_INST_1[509].FA_  ( .A(A[509]), .B(B[509]), .CI(
        C[509]), .S(S[509]), .CO(C[510]) );
  FA_1538 \FA_INST_0[0].FA_INST_1[510].FA_  ( .A(A[510]), .B(B[510]), .CI(
        C[510]), .S(S[510]), .CO(C[511]) );
  FA_1537 \FA_INST_0[0].FA_INST_1[511].FA_  ( .A(A[511]), .B(B[511]), .CI(
        C[511]), .S(S[511]), .CO(C[512]) );
  FA_1536 \FA_INST_0[1].FA_INST_1[0].FA_  ( .A(A[512]), .B(B[512]), .CI(C[512]), .S(S[512]), .CO(C[513]) );
  FA_1535 \FA_INST_0[1].FA_INST_1[1].FA_  ( .A(A[513]), .B(B[513]), .CI(C[513]), .S(S[513]), .CO(C[514]) );
  FA_1534 \FA_INST_0[1].FA_INST_1[2].FA_  ( .A(A[514]), .B(B[514]), .CI(C[514]), .S(S[514]), .CO(C[515]) );
  FA_1533 \FA_INST_0[1].FA_INST_1[3].FA_  ( .A(A[515]), .B(B[515]), .CI(C[515]), .S(S[515]), .CO(C[516]) );
  FA_1532 \FA_INST_0[1].FA_INST_1[4].FA_  ( .A(A[516]), .B(B[516]), .CI(C[516]), .S(S[516]), .CO(C[517]) );
  FA_1531 \FA_INST_0[1].FA_INST_1[5].FA_  ( .A(A[517]), .B(B[517]), .CI(C[517]), .S(S[517]), .CO(C[518]) );
  FA_1530 \FA_INST_0[1].FA_INST_1[6].FA_  ( .A(A[518]), .B(B[518]), .CI(C[518]), .S(S[518]), .CO(C[519]) );
  FA_1529 \FA_INST_0[1].FA_INST_1[7].FA_  ( .A(A[519]), .B(B[519]), .CI(C[519]), .S(S[519]), .CO(C[520]) );
  FA_1528 \FA_INST_0[1].FA_INST_1[8].FA_  ( .A(A[520]), .B(B[520]), .CI(C[520]), .S(S[520]), .CO(C[521]) );
  FA_1527 \FA_INST_0[1].FA_INST_1[9].FA_  ( .A(A[521]), .B(B[521]), .CI(C[521]), .S(S[521]), .CO(C[522]) );
  FA_1526 \FA_INST_0[1].FA_INST_1[10].FA_  ( .A(A[522]), .B(B[522]), .CI(
        C[522]), .S(S[522]), .CO(C[523]) );
  FA_1525 \FA_INST_0[1].FA_INST_1[11].FA_  ( .A(A[523]), .B(B[523]), .CI(
        C[523]), .S(S[523]), .CO(C[524]) );
  FA_1524 \FA_INST_0[1].FA_INST_1[12].FA_  ( .A(A[524]), .B(B[524]), .CI(
        C[524]), .S(S[524]), .CO(C[525]) );
  FA_1523 \FA_INST_0[1].FA_INST_1[13].FA_  ( .A(A[525]), .B(B[525]), .CI(
        C[525]), .S(S[525]), .CO(C[526]) );
  FA_1522 \FA_INST_0[1].FA_INST_1[14].FA_  ( .A(A[526]), .B(B[526]), .CI(
        C[526]), .S(S[526]), .CO(C[527]) );
  FA_1521 \FA_INST_0[1].FA_INST_1[15].FA_  ( .A(A[527]), .B(B[527]), .CI(
        C[527]), .S(S[527]), .CO(C[528]) );
  FA_1520 \FA_INST_0[1].FA_INST_1[16].FA_  ( .A(A[528]), .B(B[528]), .CI(
        C[528]), .S(S[528]), .CO(C[529]) );
  FA_1519 \FA_INST_0[1].FA_INST_1[17].FA_  ( .A(A[529]), .B(B[529]), .CI(
        C[529]), .S(S[529]), .CO(C[530]) );
  FA_1518 \FA_INST_0[1].FA_INST_1[18].FA_  ( .A(A[530]), .B(B[530]), .CI(
        C[530]), .S(S[530]), .CO(C[531]) );
  FA_1517 \FA_INST_0[1].FA_INST_1[19].FA_  ( .A(A[531]), .B(B[531]), .CI(
        C[531]), .S(S[531]), .CO(C[532]) );
  FA_1516 \FA_INST_0[1].FA_INST_1[20].FA_  ( .A(A[532]), .B(B[532]), .CI(
        C[532]), .S(S[532]), .CO(C[533]) );
  FA_1515 \FA_INST_0[1].FA_INST_1[21].FA_  ( .A(A[533]), .B(B[533]), .CI(
        C[533]), .S(S[533]), .CO(C[534]) );
  FA_1514 \FA_INST_0[1].FA_INST_1[22].FA_  ( .A(A[534]), .B(B[534]), .CI(
        C[534]), .S(S[534]), .CO(C[535]) );
  FA_1513 \FA_INST_0[1].FA_INST_1[23].FA_  ( .A(A[535]), .B(B[535]), .CI(
        C[535]), .S(S[535]), .CO(C[536]) );
  FA_1512 \FA_INST_0[1].FA_INST_1[24].FA_  ( .A(A[536]), .B(B[536]), .CI(
        C[536]), .S(S[536]), .CO(C[537]) );
  FA_1511 \FA_INST_0[1].FA_INST_1[25].FA_  ( .A(A[537]), .B(B[537]), .CI(
        C[537]), .S(S[537]), .CO(C[538]) );
  FA_1510 \FA_INST_0[1].FA_INST_1[26].FA_  ( .A(A[538]), .B(B[538]), .CI(
        C[538]), .S(S[538]), .CO(C[539]) );
  FA_1509 \FA_INST_0[1].FA_INST_1[27].FA_  ( .A(A[539]), .B(B[539]), .CI(
        C[539]), .S(S[539]), .CO(C[540]) );
  FA_1508 \FA_INST_0[1].FA_INST_1[28].FA_  ( .A(A[540]), .B(B[540]), .CI(
        C[540]), .S(S[540]), .CO(C[541]) );
  FA_1507 \FA_INST_0[1].FA_INST_1[29].FA_  ( .A(A[541]), .B(B[541]), .CI(
        C[541]), .S(S[541]), .CO(C[542]) );
  FA_1506 \FA_INST_0[1].FA_INST_1[30].FA_  ( .A(A[542]), .B(B[542]), .CI(
        C[542]), .S(S[542]), .CO(C[543]) );
  FA_1505 \FA_INST_0[1].FA_INST_1[31].FA_  ( .A(A[543]), .B(B[543]), .CI(
        C[543]), .S(S[543]), .CO(C[544]) );
  FA_1504 \FA_INST_0[1].FA_INST_1[32].FA_  ( .A(A[544]), .B(B[544]), .CI(
        C[544]), .S(S[544]), .CO(C[545]) );
  FA_1503 \FA_INST_0[1].FA_INST_1[33].FA_  ( .A(A[545]), .B(B[545]), .CI(
        C[545]), .S(S[545]), .CO(C[546]) );
  FA_1502 \FA_INST_0[1].FA_INST_1[34].FA_  ( .A(A[546]), .B(B[546]), .CI(
        C[546]), .S(S[546]), .CO(C[547]) );
  FA_1501 \FA_INST_0[1].FA_INST_1[35].FA_  ( .A(A[547]), .B(B[547]), .CI(
        C[547]), .S(S[547]), .CO(C[548]) );
  FA_1500 \FA_INST_0[1].FA_INST_1[36].FA_  ( .A(A[548]), .B(B[548]), .CI(
        C[548]), .S(S[548]), .CO(C[549]) );
  FA_1499 \FA_INST_0[1].FA_INST_1[37].FA_  ( .A(A[549]), .B(B[549]), .CI(
        C[549]), .S(S[549]), .CO(C[550]) );
  FA_1498 \FA_INST_0[1].FA_INST_1[38].FA_  ( .A(A[550]), .B(B[550]), .CI(
        C[550]), .S(S[550]), .CO(C[551]) );
  FA_1497 \FA_INST_0[1].FA_INST_1[39].FA_  ( .A(A[551]), .B(B[551]), .CI(
        C[551]), .S(S[551]), .CO(C[552]) );
  FA_1496 \FA_INST_0[1].FA_INST_1[40].FA_  ( .A(A[552]), .B(B[552]), .CI(
        C[552]), .S(S[552]), .CO(C[553]) );
  FA_1495 \FA_INST_0[1].FA_INST_1[41].FA_  ( .A(A[553]), .B(B[553]), .CI(
        C[553]), .S(S[553]), .CO(C[554]) );
  FA_1494 \FA_INST_0[1].FA_INST_1[42].FA_  ( .A(A[554]), .B(B[554]), .CI(
        C[554]), .S(S[554]), .CO(C[555]) );
  FA_1493 \FA_INST_0[1].FA_INST_1[43].FA_  ( .A(A[555]), .B(B[555]), .CI(
        C[555]), .S(S[555]), .CO(C[556]) );
  FA_1492 \FA_INST_0[1].FA_INST_1[44].FA_  ( .A(A[556]), .B(B[556]), .CI(
        C[556]), .S(S[556]), .CO(C[557]) );
  FA_1491 \FA_INST_0[1].FA_INST_1[45].FA_  ( .A(A[557]), .B(B[557]), .CI(
        C[557]), .S(S[557]), .CO(C[558]) );
  FA_1490 \FA_INST_0[1].FA_INST_1[46].FA_  ( .A(A[558]), .B(B[558]), .CI(
        C[558]), .S(S[558]), .CO(C[559]) );
  FA_1489 \FA_INST_0[1].FA_INST_1[47].FA_  ( .A(A[559]), .B(B[559]), .CI(
        C[559]), .S(S[559]), .CO(C[560]) );
  FA_1488 \FA_INST_0[1].FA_INST_1[48].FA_  ( .A(A[560]), .B(B[560]), .CI(
        C[560]), .S(S[560]), .CO(C[561]) );
  FA_1487 \FA_INST_0[1].FA_INST_1[49].FA_  ( .A(A[561]), .B(B[561]), .CI(
        C[561]), .S(S[561]), .CO(C[562]) );
  FA_1486 \FA_INST_0[1].FA_INST_1[50].FA_  ( .A(A[562]), .B(B[562]), .CI(
        C[562]), .S(S[562]), .CO(C[563]) );
  FA_1485 \FA_INST_0[1].FA_INST_1[51].FA_  ( .A(A[563]), .B(B[563]), .CI(
        C[563]), .S(S[563]), .CO(C[564]) );
  FA_1484 \FA_INST_0[1].FA_INST_1[52].FA_  ( .A(A[564]), .B(B[564]), .CI(
        C[564]), .S(S[564]), .CO(C[565]) );
  FA_1483 \FA_INST_0[1].FA_INST_1[53].FA_  ( .A(A[565]), .B(B[565]), .CI(
        C[565]), .S(S[565]), .CO(C[566]) );
  FA_1482 \FA_INST_0[1].FA_INST_1[54].FA_  ( .A(A[566]), .B(B[566]), .CI(
        C[566]), .S(S[566]), .CO(C[567]) );
  FA_1481 \FA_INST_0[1].FA_INST_1[55].FA_  ( .A(A[567]), .B(B[567]), .CI(
        C[567]), .S(S[567]), .CO(C[568]) );
  FA_1480 \FA_INST_0[1].FA_INST_1[56].FA_  ( .A(A[568]), .B(B[568]), .CI(
        C[568]), .S(S[568]), .CO(C[569]) );
  FA_1479 \FA_INST_0[1].FA_INST_1[57].FA_  ( .A(A[569]), .B(B[569]), .CI(
        C[569]), .S(S[569]), .CO(C[570]) );
  FA_1478 \FA_INST_0[1].FA_INST_1[58].FA_  ( .A(A[570]), .B(B[570]), .CI(
        C[570]), .S(S[570]), .CO(C[571]) );
  FA_1477 \FA_INST_0[1].FA_INST_1[59].FA_  ( .A(A[571]), .B(B[571]), .CI(
        C[571]), .S(S[571]), .CO(C[572]) );
  FA_1476 \FA_INST_0[1].FA_INST_1[60].FA_  ( .A(A[572]), .B(B[572]), .CI(
        C[572]), .S(S[572]), .CO(C[573]) );
  FA_1475 \FA_INST_0[1].FA_INST_1[61].FA_  ( .A(A[573]), .B(B[573]), .CI(
        C[573]), .S(S[573]), .CO(C[574]) );
  FA_1474 \FA_INST_0[1].FA_INST_1[62].FA_  ( .A(A[574]), .B(B[574]), .CI(
        C[574]), .S(S[574]), .CO(C[575]) );
  FA_1473 \FA_INST_0[1].FA_INST_1[63].FA_  ( .A(A[575]), .B(B[575]), .CI(
        C[575]), .S(S[575]), .CO(C[576]) );
  FA_1472 \FA_INST_0[1].FA_INST_1[64].FA_  ( .A(A[576]), .B(B[576]), .CI(
        C[576]), .S(S[576]), .CO(C[577]) );
  FA_1471 \FA_INST_0[1].FA_INST_1[65].FA_  ( .A(A[577]), .B(B[577]), .CI(
        C[577]), .S(S[577]), .CO(C[578]) );
  FA_1470 \FA_INST_0[1].FA_INST_1[66].FA_  ( .A(A[578]), .B(B[578]), .CI(
        C[578]), .S(S[578]), .CO(C[579]) );
  FA_1469 \FA_INST_0[1].FA_INST_1[67].FA_  ( .A(A[579]), .B(B[579]), .CI(
        C[579]), .S(S[579]), .CO(C[580]) );
  FA_1468 \FA_INST_0[1].FA_INST_1[68].FA_  ( .A(A[580]), .B(B[580]), .CI(
        C[580]), .S(S[580]), .CO(C[581]) );
  FA_1467 \FA_INST_0[1].FA_INST_1[69].FA_  ( .A(A[581]), .B(B[581]), .CI(
        C[581]), .S(S[581]), .CO(C[582]) );
  FA_1466 \FA_INST_0[1].FA_INST_1[70].FA_  ( .A(A[582]), .B(B[582]), .CI(
        C[582]), .S(S[582]), .CO(C[583]) );
  FA_1465 \FA_INST_0[1].FA_INST_1[71].FA_  ( .A(A[583]), .B(B[583]), .CI(
        C[583]), .S(S[583]), .CO(C[584]) );
  FA_1464 \FA_INST_0[1].FA_INST_1[72].FA_  ( .A(A[584]), .B(B[584]), .CI(
        C[584]), .S(S[584]), .CO(C[585]) );
  FA_1463 \FA_INST_0[1].FA_INST_1[73].FA_  ( .A(A[585]), .B(B[585]), .CI(
        C[585]), .S(S[585]), .CO(C[586]) );
  FA_1462 \FA_INST_0[1].FA_INST_1[74].FA_  ( .A(A[586]), .B(B[586]), .CI(
        C[586]), .S(S[586]), .CO(C[587]) );
  FA_1461 \FA_INST_0[1].FA_INST_1[75].FA_  ( .A(A[587]), .B(B[587]), .CI(
        C[587]), .S(S[587]), .CO(C[588]) );
  FA_1460 \FA_INST_0[1].FA_INST_1[76].FA_  ( .A(A[588]), .B(B[588]), .CI(
        C[588]), .S(S[588]), .CO(C[589]) );
  FA_1459 \FA_INST_0[1].FA_INST_1[77].FA_  ( .A(A[589]), .B(B[589]), .CI(
        C[589]), .S(S[589]), .CO(C[590]) );
  FA_1458 \FA_INST_0[1].FA_INST_1[78].FA_  ( .A(A[590]), .B(B[590]), .CI(
        C[590]), .S(S[590]), .CO(C[591]) );
  FA_1457 \FA_INST_0[1].FA_INST_1[79].FA_  ( .A(A[591]), .B(B[591]), .CI(
        C[591]), .S(S[591]), .CO(C[592]) );
  FA_1456 \FA_INST_0[1].FA_INST_1[80].FA_  ( .A(A[592]), .B(B[592]), .CI(
        C[592]), .S(S[592]), .CO(C[593]) );
  FA_1455 \FA_INST_0[1].FA_INST_1[81].FA_  ( .A(A[593]), .B(B[593]), .CI(
        C[593]), .S(S[593]), .CO(C[594]) );
  FA_1454 \FA_INST_0[1].FA_INST_1[82].FA_  ( .A(A[594]), .B(B[594]), .CI(
        C[594]), .S(S[594]), .CO(C[595]) );
  FA_1453 \FA_INST_0[1].FA_INST_1[83].FA_  ( .A(A[595]), .B(B[595]), .CI(
        C[595]), .S(S[595]), .CO(C[596]) );
  FA_1452 \FA_INST_0[1].FA_INST_1[84].FA_  ( .A(A[596]), .B(B[596]), .CI(
        C[596]), .S(S[596]), .CO(C[597]) );
  FA_1451 \FA_INST_0[1].FA_INST_1[85].FA_  ( .A(A[597]), .B(B[597]), .CI(
        C[597]), .S(S[597]), .CO(C[598]) );
  FA_1450 \FA_INST_0[1].FA_INST_1[86].FA_  ( .A(A[598]), .B(B[598]), .CI(
        C[598]), .S(S[598]), .CO(C[599]) );
  FA_1449 \FA_INST_0[1].FA_INST_1[87].FA_  ( .A(A[599]), .B(B[599]), .CI(
        C[599]), .S(S[599]), .CO(C[600]) );
  FA_1448 \FA_INST_0[1].FA_INST_1[88].FA_  ( .A(A[600]), .B(B[600]), .CI(
        C[600]), .S(S[600]), .CO(C[601]) );
  FA_1447 \FA_INST_0[1].FA_INST_1[89].FA_  ( .A(A[601]), .B(B[601]), .CI(
        C[601]), .S(S[601]), .CO(C[602]) );
  FA_1446 \FA_INST_0[1].FA_INST_1[90].FA_  ( .A(A[602]), .B(B[602]), .CI(
        C[602]), .S(S[602]), .CO(C[603]) );
  FA_1445 \FA_INST_0[1].FA_INST_1[91].FA_  ( .A(A[603]), .B(B[603]), .CI(
        C[603]), .S(S[603]), .CO(C[604]) );
  FA_1444 \FA_INST_0[1].FA_INST_1[92].FA_  ( .A(A[604]), .B(B[604]), .CI(
        C[604]), .S(S[604]), .CO(C[605]) );
  FA_1443 \FA_INST_0[1].FA_INST_1[93].FA_  ( .A(A[605]), .B(B[605]), .CI(
        C[605]), .S(S[605]), .CO(C[606]) );
  FA_1442 \FA_INST_0[1].FA_INST_1[94].FA_  ( .A(A[606]), .B(B[606]), .CI(
        C[606]), .S(S[606]), .CO(C[607]) );
  FA_1441 \FA_INST_0[1].FA_INST_1[95].FA_  ( .A(A[607]), .B(B[607]), .CI(
        C[607]), .S(S[607]), .CO(C[608]) );
  FA_1440 \FA_INST_0[1].FA_INST_1[96].FA_  ( .A(A[608]), .B(B[608]), .CI(
        C[608]), .S(S[608]), .CO(C[609]) );
  FA_1439 \FA_INST_0[1].FA_INST_1[97].FA_  ( .A(A[609]), .B(B[609]), .CI(
        C[609]), .S(S[609]), .CO(C[610]) );
  FA_1438 \FA_INST_0[1].FA_INST_1[98].FA_  ( .A(A[610]), .B(B[610]), .CI(
        C[610]), .S(S[610]), .CO(C[611]) );
  FA_1437 \FA_INST_0[1].FA_INST_1[99].FA_  ( .A(A[611]), .B(B[611]), .CI(
        C[611]), .S(S[611]), .CO(C[612]) );
  FA_1436 \FA_INST_0[1].FA_INST_1[100].FA_  ( .A(A[612]), .B(B[612]), .CI(
        C[612]), .S(S[612]), .CO(C[613]) );
  FA_1435 \FA_INST_0[1].FA_INST_1[101].FA_  ( .A(A[613]), .B(B[613]), .CI(
        C[613]), .S(S[613]), .CO(C[614]) );
  FA_1434 \FA_INST_0[1].FA_INST_1[102].FA_  ( .A(A[614]), .B(B[614]), .CI(
        C[614]), .S(S[614]), .CO(C[615]) );
  FA_1433 \FA_INST_0[1].FA_INST_1[103].FA_  ( .A(A[615]), .B(B[615]), .CI(
        C[615]), .S(S[615]), .CO(C[616]) );
  FA_1432 \FA_INST_0[1].FA_INST_1[104].FA_  ( .A(A[616]), .B(B[616]), .CI(
        C[616]), .S(S[616]), .CO(C[617]) );
  FA_1431 \FA_INST_0[1].FA_INST_1[105].FA_  ( .A(A[617]), .B(B[617]), .CI(
        C[617]), .S(S[617]), .CO(C[618]) );
  FA_1430 \FA_INST_0[1].FA_INST_1[106].FA_  ( .A(A[618]), .B(B[618]), .CI(
        C[618]), .S(S[618]), .CO(C[619]) );
  FA_1429 \FA_INST_0[1].FA_INST_1[107].FA_  ( .A(A[619]), .B(B[619]), .CI(
        C[619]), .S(S[619]), .CO(C[620]) );
  FA_1428 \FA_INST_0[1].FA_INST_1[108].FA_  ( .A(A[620]), .B(B[620]), .CI(
        C[620]), .S(S[620]), .CO(C[621]) );
  FA_1427 \FA_INST_0[1].FA_INST_1[109].FA_  ( .A(A[621]), .B(B[621]), .CI(
        C[621]), .S(S[621]), .CO(C[622]) );
  FA_1426 \FA_INST_0[1].FA_INST_1[110].FA_  ( .A(A[622]), .B(B[622]), .CI(
        C[622]), .S(S[622]), .CO(C[623]) );
  FA_1425 \FA_INST_0[1].FA_INST_1[111].FA_  ( .A(A[623]), .B(B[623]), .CI(
        C[623]), .S(S[623]), .CO(C[624]) );
  FA_1424 \FA_INST_0[1].FA_INST_1[112].FA_  ( .A(A[624]), .B(B[624]), .CI(
        C[624]), .S(S[624]), .CO(C[625]) );
  FA_1423 \FA_INST_0[1].FA_INST_1[113].FA_  ( .A(A[625]), .B(B[625]), .CI(
        C[625]), .S(S[625]), .CO(C[626]) );
  FA_1422 \FA_INST_0[1].FA_INST_1[114].FA_  ( .A(A[626]), .B(B[626]), .CI(
        C[626]), .S(S[626]), .CO(C[627]) );
  FA_1421 \FA_INST_0[1].FA_INST_1[115].FA_  ( .A(A[627]), .B(B[627]), .CI(
        C[627]), .S(S[627]), .CO(C[628]) );
  FA_1420 \FA_INST_0[1].FA_INST_1[116].FA_  ( .A(A[628]), .B(B[628]), .CI(
        C[628]), .S(S[628]), .CO(C[629]) );
  FA_1419 \FA_INST_0[1].FA_INST_1[117].FA_  ( .A(A[629]), .B(B[629]), .CI(
        C[629]), .S(S[629]), .CO(C[630]) );
  FA_1418 \FA_INST_0[1].FA_INST_1[118].FA_  ( .A(A[630]), .B(B[630]), .CI(
        C[630]), .S(S[630]), .CO(C[631]) );
  FA_1417 \FA_INST_0[1].FA_INST_1[119].FA_  ( .A(A[631]), .B(B[631]), .CI(
        C[631]), .S(S[631]), .CO(C[632]) );
  FA_1416 \FA_INST_0[1].FA_INST_1[120].FA_  ( .A(A[632]), .B(B[632]), .CI(
        C[632]), .S(S[632]), .CO(C[633]) );
  FA_1415 \FA_INST_0[1].FA_INST_1[121].FA_  ( .A(A[633]), .B(B[633]), .CI(
        C[633]), .S(S[633]), .CO(C[634]) );
  FA_1414 \FA_INST_0[1].FA_INST_1[122].FA_  ( .A(A[634]), .B(B[634]), .CI(
        C[634]), .S(S[634]), .CO(C[635]) );
  FA_1413 \FA_INST_0[1].FA_INST_1[123].FA_  ( .A(A[635]), .B(B[635]), .CI(
        C[635]), .S(S[635]), .CO(C[636]) );
  FA_1412 \FA_INST_0[1].FA_INST_1[124].FA_  ( .A(A[636]), .B(B[636]), .CI(
        C[636]), .S(S[636]), .CO(C[637]) );
  FA_1411 \FA_INST_0[1].FA_INST_1[125].FA_  ( .A(A[637]), .B(B[637]), .CI(
        C[637]), .S(S[637]), .CO(C[638]) );
  FA_1410 \FA_INST_0[1].FA_INST_1[126].FA_  ( .A(A[638]), .B(B[638]), .CI(
        C[638]), .S(S[638]), .CO(C[639]) );
  FA_1409 \FA_INST_0[1].FA_INST_1[127].FA_  ( .A(A[639]), .B(B[639]), .CI(
        C[639]), .S(S[639]), .CO(C[640]) );
  FA_1408 \FA_INST_0[1].FA_INST_1[128].FA_  ( .A(A[640]), .B(B[640]), .CI(
        C[640]), .S(S[640]), .CO(C[641]) );
  FA_1407 \FA_INST_0[1].FA_INST_1[129].FA_  ( .A(A[641]), .B(B[641]), .CI(
        C[641]), .S(S[641]), .CO(C[642]) );
  FA_1406 \FA_INST_0[1].FA_INST_1[130].FA_  ( .A(A[642]), .B(B[642]), .CI(
        C[642]), .S(S[642]), .CO(C[643]) );
  FA_1405 \FA_INST_0[1].FA_INST_1[131].FA_  ( .A(A[643]), .B(B[643]), .CI(
        C[643]), .S(S[643]), .CO(C[644]) );
  FA_1404 \FA_INST_0[1].FA_INST_1[132].FA_  ( .A(A[644]), .B(B[644]), .CI(
        C[644]), .S(S[644]), .CO(C[645]) );
  FA_1403 \FA_INST_0[1].FA_INST_1[133].FA_  ( .A(A[645]), .B(B[645]), .CI(
        C[645]), .S(S[645]), .CO(C[646]) );
  FA_1402 \FA_INST_0[1].FA_INST_1[134].FA_  ( .A(A[646]), .B(B[646]), .CI(
        C[646]), .S(S[646]), .CO(C[647]) );
  FA_1401 \FA_INST_0[1].FA_INST_1[135].FA_  ( .A(A[647]), .B(B[647]), .CI(
        C[647]), .S(S[647]), .CO(C[648]) );
  FA_1400 \FA_INST_0[1].FA_INST_1[136].FA_  ( .A(A[648]), .B(B[648]), .CI(
        C[648]), .S(S[648]), .CO(C[649]) );
  FA_1399 \FA_INST_0[1].FA_INST_1[137].FA_  ( .A(A[649]), .B(B[649]), .CI(
        C[649]), .S(S[649]), .CO(C[650]) );
  FA_1398 \FA_INST_0[1].FA_INST_1[138].FA_  ( .A(A[650]), .B(B[650]), .CI(
        C[650]), .S(S[650]), .CO(C[651]) );
  FA_1397 \FA_INST_0[1].FA_INST_1[139].FA_  ( .A(A[651]), .B(B[651]), .CI(
        C[651]), .S(S[651]), .CO(C[652]) );
  FA_1396 \FA_INST_0[1].FA_INST_1[140].FA_  ( .A(A[652]), .B(B[652]), .CI(
        C[652]), .S(S[652]), .CO(C[653]) );
  FA_1395 \FA_INST_0[1].FA_INST_1[141].FA_  ( .A(A[653]), .B(B[653]), .CI(
        C[653]), .S(S[653]), .CO(C[654]) );
  FA_1394 \FA_INST_0[1].FA_INST_1[142].FA_  ( .A(A[654]), .B(B[654]), .CI(
        C[654]), .S(S[654]), .CO(C[655]) );
  FA_1393 \FA_INST_0[1].FA_INST_1[143].FA_  ( .A(A[655]), .B(B[655]), .CI(
        C[655]), .S(S[655]), .CO(C[656]) );
  FA_1392 \FA_INST_0[1].FA_INST_1[144].FA_  ( .A(A[656]), .B(B[656]), .CI(
        C[656]), .S(S[656]), .CO(C[657]) );
  FA_1391 \FA_INST_0[1].FA_INST_1[145].FA_  ( .A(A[657]), .B(B[657]), .CI(
        C[657]), .S(S[657]), .CO(C[658]) );
  FA_1390 \FA_INST_0[1].FA_INST_1[146].FA_  ( .A(A[658]), .B(B[658]), .CI(
        C[658]), .S(S[658]), .CO(C[659]) );
  FA_1389 \FA_INST_0[1].FA_INST_1[147].FA_  ( .A(A[659]), .B(B[659]), .CI(
        C[659]), .S(S[659]), .CO(C[660]) );
  FA_1388 \FA_INST_0[1].FA_INST_1[148].FA_  ( .A(A[660]), .B(B[660]), .CI(
        C[660]), .S(S[660]), .CO(C[661]) );
  FA_1387 \FA_INST_0[1].FA_INST_1[149].FA_  ( .A(A[661]), .B(B[661]), .CI(
        C[661]), .S(S[661]), .CO(C[662]) );
  FA_1386 \FA_INST_0[1].FA_INST_1[150].FA_  ( .A(A[662]), .B(B[662]), .CI(
        C[662]), .S(S[662]), .CO(C[663]) );
  FA_1385 \FA_INST_0[1].FA_INST_1[151].FA_  ( .A(A[663]), .B(B[663]), .CI(
        C[663]), .S(S[663]), .CO(C[664]) );
  FA_1384 \FA_INST_0[1].FA_INST_1[152].FA_  ( .A(A[664]), .B(B[664]), .CI(
        C[664]), .S(S[664]), .CO(C[665]) );
  FA_1383 \FA_INST_0[1].FA_INST_1[153].FA_  ( .A(A[665]), .B(B[665]), .CI(
        C[665]), .S(S[665]), .CO(C[666]) );
  FA_1382 \FA_INST_0[1].FA_INST_1[154].FA_  ( .A(A[666]), .B(B[666]), .CI(
        C[666]), .S(S[666]), .CO(C[667]) );
  FA_1381 \FA_INST_0[1].FA_INST_1[155].FA_  ( .A(A[667]), .B(B[667]), .CI(
        C[667]), .S(S[667]), .CO(C[668]) );
  FA_1380 \FA_INST_0[1].FA_INST_1[156].FA_  ( .A(A[668]), .B(B[668]), .CI(
        C[668]), .S(S[668]), .CO(C[669]) );
  FA_1379 \FA_INST_0[1].FA_INST_1[157].FA_  ( .A(A[669]), .B(B[669]), .CI(
        C[669]), .S(S[669]), .CO(C[670]) );
  FA_1378 \FA_INST_0[1].FA_INST_1[158].FA_  ( .A(A[670]), .B(B[670]), .CI(
        C[670]), .S(S[670]), .CO(C[671]) );
  FA_1377 \FA_INST_0[1].FA_INST_1[159].FA_  ( .A(A[671]), .B(B[671]), .CI(
        C[671]), .S(S[671]), .CO(C[672]) );
  FA_1376 \FA_INST_0[1].FA_INST_1[160].FA_  ( .A(A[672]), .B(B[672]), .CI(
        C[672]), .S(S[672]), .CO(C[673]) );
  FA_1375 \FA_INST_0[1].FA_INST_1[161].FA_  ( .A(A[673]), .B(B[673]), .CI(
        C[673]), .S(S[673]), .CO(C[674]) );
  FA_1374 \FA_INST_0[1].FA_INST_1[162].FA_  ( .A(A[674]), .B(B[674]), .CI(
        C[674]), .S(S[674]), .CO(C[675]) );
  FA_1373 \FA_INST_0[1].FA_INST_1[163].FA_  ( .A(A[675]), .B(B[675]), .CI(
        C[675]), .S(S[675]), .CO(C[676]) );
  FA_1372 \FA_INST_0[1].FA_INST_1[164].FA_  ( .A(A[676]), .B(B[676]), .CI(
        C[676]), .S(S[676]), .CO(C[677]) );
  FA_1371 \FA_INST_0[1].FA_INST_1[165].FA_  ( .A(A[677]), .B(B[677]), .CI(
        C[677]), .S(S[677]), .CO(C[678]) );
  FA_1370 \FA_INST_0[1].FA_INST_1[166].FA_  ( .A(A[678]), .B(B[678]), .CI(
        C[678]), .S(S[678]), .CO(C[679]) );
  FA_1369 \FA_INST_0[1].FA_INST_1[167].FA_  ( .A(A[679]), .B(B[679]), .CI(
        C[679]), .S(S[679]), .CO(C[680]) );
  FA_1368 \FA_INST_0[1].FA_INST_1[168].FA_  ( .A(A[680]), .B(B[680]), .CI(
        C[680]), .S(S[680]), .CO(C[681]) );
  FA_1367 \FA_INST_0[1].FA_INST_1[169].FA_  ( .A(A[681]), .B(B[681]), .CI(
        C[681]), .S(S[681]), .CO(C[682]) );
  FA_1366 \FA_INST_0[1].FA_INST_1[170].FA_  ( .A(A[682]), .B(B[682]), .CI(
        C[682]), .S(S[682]), .CO(C[683]) );
  FA_1365 \FA_INST_0[1].FA_INST_1[171].FA_  ( .A(A[683]), .B(B[683]), .CI(
        C[683]), .S(S[683]), .CO(C[684]) );
  FA_1364 \FA_INST_0[1].FA_INST_1[172].FA_  ( .A(A[684]), .B(B[684]), .CI(
        C[684]), .S(S[684]), .CO(C[685]) );
  FA_1363 \FA_INST_0[1].FA_INST_1[173].FA_  ( .A(A[685]), .B(B[685]), .CI(
        C[685]), .S(S[685]), .CO(C[686]) );
  FA_1362 \FA_INST_0[1].FA_INST_1[174].FA_  ( .A(A[686]), .B(B[686]), .CI(
        C[686]), .S(S[686]), .CO(C[687]) );
  FA_1361 \FA_INST_0[1].FA_INST_1[175].FA_  ( .A(A[687]), .B(B[687]), .CI(
        C[687]), .S(S[687]), .CO(C[688]) );
  FA_1360 \FA_INST_0[1].FA_INST_1[176].FA_  ( .A(A[688]), .B(B[688]), .CI(
        C[688]), .S(S[688]), .CO(C[689]) );
  FA_1359 \FA_INST_0[1].FA_INST_1[177].FA_  ( .A(A[689]), .B(B[689]), .CI(
        C[689]), .S(S[689]), .CO(C[690]) );
  FA_1358 \FA_INST_0[1].FA_INST_1[178].FA_  ( .A(A[690]), .B(B[690]), .CI(
        C[690]), .S(S[690]), .CO(C[691]) );
  FA_1357 \FA_INST_0[1].FA_INST_1[179].FA_  ( .A(A[691]), .B(B[691]), .CI(
        C[691]), .S(S[691]), .CO(C[692]) );
  FA_1356 \FA_INST_0[1].FA_INST_1[180].FA_  ( .A(A[692]), .B(B[692]), .CI(
        C[692]), .S(S[692]), .CO(C[693]) );
  FA_1355 \FA_INST_0[1].FA_INST_1[181].FA_  ( .A(A[693]), .B(B[693]), .CI(
        C[693]), .S(S[693]), .CO(C[694]) );
  FA_1354 \FA_INST_0[1].FA_INST_1[182].FA_  ( .A(A[694]), .B(B[694]), .CI(
        C[694]), .S(S[694]), .CO(C[695]) );
  FA_1353 \FA_INST_0[1].FA_INST_1[183].FA_  ( .A(A[695]), .B(B[695]), .CI(
        C[695]), .S(S[695]), .CO(C[696]) );
  FA_1352 \FA_INST_0[1].FA_INST_1[184].FA_  ( .A(A[696]), .B(B[696]), .CI(
        C[696]), .S(S[696]), .CO(C[697]) );
  FA_1351 \FA_INST_0[1].FA_INST_1[185].FA_  ( .A(A[697]), .B(B[697]), .CI(
        C[697]), .S(S[697]), .CO(C[698]) );
  FA_1350 \FA_INST_0[1].FA_INST_1[186].FA_  ( .A(A[698]), .B(B[698]), .CI(
        C[698]), .S(S[698]), .CO(C[699]) );
  FA_1349 \FA_INST_0[1].FA_INST_1[187].FA_  ( .A(A[699]), .B(B[699]), .CI(
        C[699]), .S(S[699]), .CO(C[700]) );
  FA_1348 \FA_INST_0[1].FA_INST_1[188].FA_  ( .A(A[700]), .B(B[700]), .CI(
        C[700]), .S(S[700]), .CO(C[701]) );
  FA_1347 \FA_INST_0[1].FA_INST_1[189].FA_  ( .A(A[701]), .B(B[701]), .CI(
        C[701]), .S(S[701]), .CO(C[702]) );
  FA_1346 \FA_INST_0[1].FA_INST_1[190].FA_  ( .A(A[702]), .B(B[702]), .CI(
        C[702]), .S(S[702]), .CO(C[703]) );
  FA_1345 \FA_INST_0[1].FA_INST_1[191].FA_  ( .A(A[703]), .B(B[703]), .CI(
        C[703]), .S(S[703]), .CO(C[704]) );
  FA_1344 \FA_INST_0[1].FA_INST_1[192].FA_  ( .A(A[704]), .B(B[704]), .CI(
        C[704]), .S(S[704]), .CO(C[705]) );
  FA_1343 \FA_INST_0[1].FA_INST_1[193].FA_  ( .A(A[705]), .B(B[705]), .CI(
        C[705]), .S(S[705]), .CO(C[706]) );
  FA_1342 \FA_INST_0[1].FA_INST_1[194].FA_  ( .A(A[706]), .B(B[706]), .CI(
        C[706]), .S(S[706]), .CO(C[707]) );
  FA_1341 \FA_INST_0[1].FA_INST_1[195].FA_  ( .A(A[707]), .B(B[707]), .CI(
        C[707]), .S(S[707]), .CO(C[708]) );
  FA_1340 \FA_INST_0[1].FA_INST_1[196].FA_  ( .A(A[708]), .B(B[708]), .CI(
        C[708]), .S(S[708]), .CO(C[709]) );
  FA_1339 \FA_INST_0[1].FA_INST_1[197].FA_  ( .A(A[709]), .B(B[709]), .CI(
        C[709]), .S(S[709]), .CO(C[710]) );
  FA_1338 \FA_INST_0[1].FA_INST_1[198].FA_  ( .A(A[710]), .B(B[710]), .CI(
        C[710]), .S(S[710]), .CO(C[711]) );
  FA_1337 \FA_INST_0[1].FA_INST_1[199].FA_  ( .A(A[711]), .B(B[711]), .CI(
        C[711]), .S(S[711]), .CO(C[712]) );
  FA_1336 \FA_INST_0[1].FA_INST_1[200].FA_  ( .A(A[712]), .B(B[712]), .CI(
        C[712]), .S(S[712]), .CO(C[713]) );
  FA_1335 \FA_INST_0[1].FA_INST_1[201].FA_  ( .A(A[713]), .B(B[713]), .CI(
        C[713]), .S(S[713]), .CO(C[714]) );
  FA_1334 \FA_INST_0[1].FA_INST_1[202].FA_  ( .A(A[714]), .B(B[714]), .CI(
        C[714]), .S(S[714]), .CO(C[715]) );
  FA_1333 \FA_INST_0[1].FA_INST_1[203].FA_  ( .A(A[715]), .B(B[715]), .CI(
        C[715]), .S(S[715]), .CO(C[716]) );
  FA_1332 \FA_INST_0[1].FA_INST_1[204].FA_  ( .A(A[716]), .B(B[716]), .CI(
        C[716]), .S(S[716]), .CO(C[717]) );
  FA_1331 \FA_INST_0[1].FA_INST_1[205].FA_  ( .A(A[717]), .B(B[717]), .CI(
        C[717]), .S(S[717]), .CO(C[718]) );
  FA_1330 \FA_INST_0[1].FA_INST_1[206].FA_  ( .A(A[718]), .B(B[718]), .CI(
        C[718]), .S(S[718]), .CO(C[719]) );
  FA_1329 \FA_INST_0[1].FA_INST_1[207].FA_  ( .A(A[719]), .B(B[719]), .CI(
        C[719]), .S(S[719]), .CO(C[720]) );
  FA_1328 \FA_INST_0[1].FA_INST_1[208].FA_  ( .A(A[720]), .B(B[720]), .CI(
        C[720]), .S(S[720]), .CO(C[721]) );
  FA_1327 \FA_INST_0[1].FA_INST_1[209].FA_  ( .A(A[721]), .B(B[721]), .CI(
        C[721]), .S(S[721]), .CO(C[722]) );
  FA_1326 \FA_INST_0[1].FA_INST_1[210].FA_  ( .A(A[722]), .B(B[722]), .CI(
        C[722]), .S(S[722]), .CO(C[723]) );
  FA_1325 \FA_INST_0[1].FA_INST_1[211].FA_  ( .A(A[723]), .B(B[723]), .CI(
        C[723]), .S(S[723]), .CO(C[724]) );
  FA_1324 \FA_INST_0[1].FA_INST_1[212].FA_  ( .A(A[724]), .B(B[724]), .CI(
        C[724]), .S(S[724]), .CO(C[725]) );
  FA_1323 \FA_INST_0[1].FA_INST_1[213].FA_  ( .A(A[725]), .B(B[725]), .CI(
        C[725]), .S(S[725]), .CO(C[726]) );
  FA_1322 \FA_INST_0[1].FA_INST_1[214].FA_  ( .A(A[726]), .B(B[726]), .CI(
        C[726]), .S(S[726]), .CO(C[727]) );
  FA_1321 \FA_INST_0[1].FA_INST_1[215].FA_  ( .A(A[727]), .B(B[727]), .CI(
        C[727]), .S(S[727]), .CO(C[728]) );
  FA_1320 \FA_INST_0[1].FA_INST_1[216].FA_  ( .A(A[728]), .B(B[728]), .CI(
        C[728]), .S(S[728]), .CO(C[729]) );
  FA_1319 \FA_INST_0[1].FA_INST_1[217].FA_  ( .A(A[729]), .B(B[729]), .CI(
        C[729]), .S(S[729]), .CO(C[730]) );
  FA_1318 \FA_INST_0[1].FA_INST_1[218].FA_  ( .A(A[730]), .B(B[730]), .CI(
        C[730]), .S(S[730]), .CO(C[731]) );
  FA_1317 \FA_INST_0[1].FA_INST_1[219].FA_  ( .A(A[731]), .B(B[731]), .CI(
        C[731]), .S(S[731]), .CO(C[732]) );
  FA_1316 \FA_INST_0[1].FA_INST_1[220].FA_  ( .A(A[732]), .B(B[732]), .CI(
        C[732]), .S(S[732]), .CO(C[733]) );
  FA_1315 \FA_INST_0[1].FA_INST_1[221].FA_  ( .A(A[733]), .B(B[733]), .CI(
        C[733]), .S(S[733]), .CO(C[734]) );
  FA_1314 \FA_INST_0[1].FA_INST_1[222].FA_  ( .A(A[734]), .B(B[734]), .CI(
        C[734]), .S(S[734]), .CO(C[735]) );
  FA_1313 \FA_INST_0[1].FA_INST_1[223].FA_  ( .A(A[735]), .B(B[735]), .CI(
        C[735]), .S(S[735]), .CO(C[736]) );
  FA_1312 \FA_INST_0[1].FA_INST_1[224].FA_  ( .A(A[736]), .B(B[736]), .CI(
        C[736]), .S(S[736]), .CO(C[737]) );
  FA_1311 \FA_INST_0[1].FA_INST_1[225].FA_  ( .A(A[737]), .B(B[737]), .CI(
        C[737]), .S(S[737]), .CO(C[738]) );
  FA_1310 \FA_INST_0[1].FA_INST_1[226].FA_  ( .A(A[738]), .B(B[738]), .CI(
        C[738]), .S(S[738]), .CO(C[739]) );
  FA_1309 \FA_INST_0[1].FA_INST_1[227].FA_  ( .A(A[739]), .B(B[739]), .CI(
        C[739]), .S(S[739]), .CO(C[740]) );
  FA_1308 \FA_INST_0[1].FA_INST_1[228].FA_  ( .A(A[740]), .B(B[740]), .CI(
        C[740]), .S(S[740]), .CO(C[741]) );
  FA_1307 \FA_INST_0[1].FA_INST_1[229].FA_  ( .A(A[741]), .B(B[741]), .CI(
        C[741]), .S(S[741]), .CO(C[742]) );
  FA_1306 \FA_INST_0[1].FA_INST_1[230].FA_  ( .A(A[742]), .B(B[742]), .CI(
        C[742]), .S(S[742]), .CO(C[743]) );
  FA_1305 \FA_INST_0[1].FA_INST_1[231].FA_  ( .A(A[743]), .B(B[743]), .CI(
        C[743]), .S(S[743]), .CO(C[744]) );
  FA_1304 \FA_INST_0[1].FA_INST_1[232].FA_  ( .A(A[744]), .B(B[744]), .CI(
        C[744]), .S(S[744]), .CO(C[745]) );
  FA_1303 \FA_INST_0[1].FA_INST_1[233].FA_  ( .A(A[745]), .B(B[745]), .CI(
        C[745]), .S(S[745]), .CO(C[746]) );
  FA_1302 \FA_INST_0[1].FA_INST_1[234].FA_  ( .A(A[746]), .B(B[746]), .CI(
        C[746]), .S(S[746]), .CO(C[747]) );
  FA_1301 \FA_INST_0[1].FA_INST_1[235].FA_  ( .A(A[747]), .B(B[747]), .CI(
        C[747]), .S(S[747]), .CO(C[748]) );
  FA_1300 \FA_INST_0[1].FA_INST_1[236].FA_  ( .A(A[748]), .B(B[748]), .CI(
        C[748]), .S(S[748]), .CO(C[749]) );
  FA_1299 \FA_INST_0[1].FA_INST_1[237].FA_  ( .A(A[749]), .B(B[749]), .CI(
        C[749]), .S(S[749]), .CO(C[750]) );
  FA_1298 \FA_INST_0[1].FA_INST_1[238].FA_  ( .A(A[750]), .B(B[750]), .CI(
        C[750]), .S(S[750]), .CO(C[751]) );
  FA_1297 \FA_INST_0[1].FA_INST_1[239].FA_  ( .A(A[751]), .B(B[751]), .CI(
        C[751]), .S(S[751]), .CO(C[752]) );
  FA_1296 \FA_INST_0[1].FA_INST_1[240].FA_  ( .A(A[752]), .B(B[752]), .CI(
        C[752]), .S(S[752]), .CO(C[753]) );
  FA_1295 \FA_INST_0[1].FA_INST_1[241].FA_  ( .A(A[753]), .B(B[753]), .CI(
        C[753]), .S(S[753]), .CO(C[754]) );
  FA_1294 \FA_INST_0[1].FA_INST_1[242].FA_  ( .A(A[754]), .B(B[754]), .CI(
        C[754]), .S(S[754]), .CO(C[755]) );
  FA_1293 \FA_INST_0[1].FA_INST_1[243].FA_  ( .A(A[755]), .B(B[755]), .CI(
        C[755]), .S(S[755]), .CO(C[756]) );
  FA_1292 \FA_INST_0[1].FA_INST_1[244].FA_  ( .A(A[756]), .B(B[756]), .CI(
        C[756]), .S(S[756]), .CO(C[757]) );
  FA_1291 \FA_INST_0[1].FA_INST_1[245].FA_  ( .A(A[757]), .B(B[757]), .CI(
        C[757]), .S(S[757]), .CO(C[758]) );
  FA_1290 \FA_INST_0[1].FA_INST_1[246].FA_  ( .A(A[758]), .B(B[758]), .CI(
        C[758]), .S(S[758]), .CO(C[759]) );
  FA_1289 \FA_INST_0[1].FA_INST_1[247].FA_  ( .A(A[759]), .B(B[759]), .CI(
        C[759]), .S(S[759]), .CO(C[760]) );
  FA_1288 \FA_INST_0[1].FA_INST_1[248].FA_  ( .A(A[760]), .B(B[760]), .CI(
        C[760]), .S(S[760]), .CO(C[761]) );
  FA_1287 \FA_INST_0[1].FA_INST_1[249].FA_  ( .A(A[761]), .B(B[761]), .CI(
        C[761]), .S(S[761]), .CO(C[762]) );
  FA_1286 \FA_INST_0[1].FA_INST_1[250].FA_  ( .A(A[762]), .B(B[762]), .CI(
        C[762]), .S(S[762]), .CO(C[763]) );
  FA_1285 \FA_INST_0[1].FA_INST_1[251].FA_  ( .A(A[763]), .B(B[763]), .CI(
        C[763]), .S(S[763]), .CO(C[764]) );
  FA_1284 \FA_INST_0[1].FA_INST_1[252].FA_  ( .A(A[764]), .B(B[764]), .CI(
        C[764]), .S(S[764]), .CO(C[765]) );
  FA_1283 \FA_INST_0[1].FA_INST_1[253].FA_  ( .A(A[765]), .B(B[765]), .CI(
        C[765]), .S(S[765]), .CO(C[766]) );
  FA_1282 \FA_INST_0[1].FA_INST_1[254].FA_  ( .A(A[766]), .B(B[766]), .CI(
        C[766]), .S(S[766]), .CO(C[767]) );
  FA_1281 \FA_INST_0[1].FA_INST_1[255].FA_  ( .A(A[767]), .B(B[767]), .CI(
        C[767]), .S(S[767]), .CO(C[768]) );
  FA_1280 \FA_INST_0[1].FA_INST_1[256].FA_  ( .A(A[768]), .B(B[768]), .CI(
        C[768]), .S(S[768]), .CO(C[769]) );
  FA_1279 \FA_INST_0[1].FA_INST_1[257].FA_  ( .A(A[769]), .B(B[769]), .CI(
        C[769]), .S(S[769]), .CO(C[770]) );
  FA_1278 \FA_INST_0[1].FA_INST_1[258].FA_  ( .A(A[770]), .B(B[770]), .CI(
        C[770]), .S(S[770]), .CO(C[771]) );
  FA_1277 \FA_INST_0[1].FA_INST_1[259].FA_  ( .A(A[771]), .B(B[771]), .CI(
        C[771]), .S(S[771]), .CO(C[772]) );
  FA_1276 \FA_INST_0[1].FA_INST_1[260].FA_  ( .A(A[772]), .B(B[772]), .CI(
        C[772]), .S(S[772]), .CO(C[773]) );
  FA_1275 \FA_INST_0[1].FA_INST_1[261].FA_  ( .A(A[773]), .B(B[773]), .CI(
        C[773]), .S(S[773]), .CO(C[774]) );
  FA_1274 \FA_INST_0[1].FA_INST_1[262].FA_  ( .A(A[774]), .B(B[774]), .CI(
        C[774]), .S(S[774]), .CO(C[775]) );
  FA_1273 \FA_INST_0[1].FA_INST_1[263].FA_  ( .A(A[775]), .B(B[775]), .CI(
        C[775]), .S(S[775]), .CO(C[776]) );
  FA_1272 \FA_INST_0[1].FA_INST_1[264].FA_  ( .A(A[776]), .B(B[776]), .CI(
        C[776]), .S(S[776]), .CO(C[777]) );
  FA_1271 \FA_INST_0[1].FA_INST_1[265].FA_  ( .A(A[777]), .B(B[777]), .CI(
        C[777]), .S(S[777]), .CO(C[778]) );
  FA_1270 \FA_INST_0[1].FA_INST_1[266].FA_  ( .A(A[778]), .B(B[778]), .CI(
        C[778]), .S(S[778]), .CO(C[779]) );
  FA_1269 \FA_INST_0[1].FA_INST_1[267].FA_  ( .A(A[779]), .B(B[779]), .CI(
        C[779]), .S(S[779]), .CO(C[780]) );
  FA_1268 \FA_INST_0[1].FA_INST_1[268].FA_  ( .A(A[780]), .B(B[780]), .CI(
        C[780]), .S(S[780]), .CO(C[781]) );
  FA_1267 \FA_INST_0[1].FA_INST_1[269].FA_  ( .A(A[781]), .B(B[781]), .CI(
        C[781]), .S(S[781]), .CO(C[782]) );
  FA_1266 \FA_INST_0[1].FA_INST_1[270].FA_  ( .A(A[782]), .B(B[782]), .CI(
        C[782]), .S(S[782]), .CO(C[783]) );
  FA_1265 \FA_INST_0[1].FA_INST_1[271].FA_  ( .A(A[783]), .B(B[783]), .CI(
        C[783]), .S(S[783]), .CO(C[784]) );
  FA_1264 \FA_INST_0[1].FA_INST_1[272].FA_  ( .A(A[784]), .B(B[784]), .CI(
        C[784]), .S(S[784]), .CO(C[785]) );
  FA_1263 \FA_INST_0[1].FA_INST_1[273].FA_  ( .A(A[785]), .B(B[785]), .CI(
        C[785]), .S(S[785]), .CO(C[786]) );
  FA_1262 \FA_INST_0[1].FA_INST_1[274].FA_  ( .A(A[786]), .B(B[786]), .CI(
        C[786]), .S(S[786]), .CO(C[787]) );
  FA_1261 \FA_INST_0[1].FA_INST_1[275].FA_  ( .A(A[787]), .B(B[787]), .CI(
        C[787]), .S(S[787]), .CO(C[788]) );
  FA_1260 \FA_INST_0[1].FA_INST_1[276].FA_  ( .A(A[788]), .B(B[788]), .CI(
        C[788]), .S(S[788]), .CO(C[789]) );
  FA_1259 \FA_INST_0[1].FA_INST_1[277].FA_  ( .A(A[789]), .B(B[789]), .CI(
        C[789]), .S(S[789]), .CO(C[790]) );
  FA_1258 \FA_INST_0[1].FA_INST_1[278].FA_  ( .A(A[790]), .B(B[790]), .CI(
        C[790]), .S(S[790]), .CO(C[791]) );
  FA_1257 \FA_INST_0[1].FA_INST_1[279].FA_  ( .A(A[791]), .B(B[791]), .CI(
        C[791]), .S(S[791]), .CO(C[792]) );
  FA_1256 \FA_INST_0[1].FA_INST_1[280].FA_  ( .A(A[792]), .B(B[792]), .CI(
        C[792]), .S(S[792]), .CO(C[793]) );
  FA_1255 \FA_INST_0[1].FA_INST_1[281].FA_  ( .A(A[793]), .B(B[793]), .CI(
        C[793]), .S(S[793]), .CO(C[794]) );
  FA_1254 \FA_INST_0[1].FA_INST_1[282].FA_  ( .A(A[794]), .B(B[794]), .CI(
        C[794]), .S(S[794]), .CO(C[795]) );
  FA_1253 \FA_INST_0[1].FA_INST_1[283].FA_  ( .A(A[795]), .B(B[795]), .CI(
        C[795]), .S(S[795]), .CO(C[796]) );
  FA_1252 \FA_INST_0[1].FA_INST_1[284].FA_  ( .A(A[796]), .B(B[796]), .CI(
        C[796]), .S(S[796]), .CO(C[797]) );
  FA_1251 \FA_INST_0[1].FA_INST_1[285].FA_  ( .A(A[797]), .B(B[797]), .CI(
        C[797]), .S(S[797]), .CO(C[798]) );
  FA_1250 \FA_INST_0[1].FA_INST_1[286].FA_  ( .A(A[798]), .B(B[798]), .CI(
        C[798]), .S(S[798]), .CO(C[799]) );
  FA_1249 \FA_INST_0[1].FA_INST_1[287].FA_  ( .A(A[799]), .B(B[799]), .CI(
        C[799]), .S(S[799]), .CO(C[800]) );
  FA_1248 \FA_INST_0[1].FA_INST_1[288].FA_  ( .A(A[800]), .B(B[800]), .CI(
        C[800]), .S(S[800]), .CO(C[801]) );
  FA_1247 \FA_INST_0[1].FA_INST_1[289].FA_  ( .A(A[801]), .B(B[801]), .CI(
        C[801]), .S(S[801]), .CO(C[802]) );
  FA_1246 \FA_INST_0[1].FA_INST_1[290].FA_  ( .A(A[802]), .B(B[802]), .CI(
        C[802]), .S(S[802]), .CO(C[803]) );
  FA_1245 \FA_INST_0[1].FA_INST_1[291].FA_  ( .A(A[803]), .B(B[803]), .CI(
        C[803]), .S(S[803]), .CO(C[804]) );
  FA_1244 \FA_INST_0[1].FA_INST_1[292].FA_  ( .A(A[804]), .B(B[804]), .CI(
        C[804]), .S(S[804]), .CO(C[805]) );
  FA_1243 \FA_INST_0[1].FA_INST_1[293].FA_  ( .A(A[805]), .B(B[805]), .CI(
        C[805]), .S(S[805]), .CO(C[806]) );
  FA_1242 \FA_INST_0[1].FA_INST_1[294].FA_  ( .A(A[806]), .B(B[806]), .CI(
        C[806]), .S(S[806]), .CO(C[807]) );
  FA_1241 \FA_INST_0[1].FA_INST_1[295].FA_  ( .A(A[807]), .B(B[807]), .CI(
        C[807]), .S(S[807]), .CO(C[808]) );
  FA_1240 \FA_INST_0[1].FA_INST_1[296].FA_  ( .A(A[808]), .B(B[808]), .CI(
        C[808]), .S(S[808]), .CO(C[809]) );
  FA_1239 \FA_INST_0[1].FA_INST_1[297].FA_  ( .A(A[809]), .B(B[809]), .CI(
        C[809]), .S(S[809]), .CO(C[810]) );
  FA_1238 \FA_INST_0[1].FA_INST_1[298].FA_  ( .A(A[810]), .B(B[810]), .CI(
        C[810]), .S(S[810]), .CO(C[811]) );
  FA_1237 \FA_INST_0[1].FA_INST_1[299].FA_  ( .A(A[811]), .B(B[811]), .CI(
        C[811]), .S(S[811]), .CO(C[812]) );
  FA_1236 \FA_INST_0[1].FA_INST_1[300].FA_  ( .A(A[812]), .B(B[812]), .CI(
        C[812]), .S(S[812]), .CO(C[813]) );
  FA_1235 \FA_INST_0[1].FA_INST_1[301].FA_  ( .A(A[813]), .B(B[813]), .CI(
        C[813]), .S(S[813]), .CO(C[814]) );
  FA_1234 \FA_INST_0[1].FA_INST_1[302].FA_  ( .A(A[814]), .B(B[814]), .CI(
        C[814]), .S(S[814]), .CO(C[815]) );
  FA_1233 \FA_INST_0[1].FA_INST_1[303].FA_  ( .A(A[815]), .B(B[815]), .CI(
        C[815]), .S(S[815]), .CO(C[816]) );
  FA_1232 \FA_INST_0[1].FA_INST_1[304].FA_  ( .A(A[816]), .B(B[816]), .CI(
        C[816]), .S(S[816]), .CO(C[817]) );
  FA_1231 \FA_INST_0[1].FA_INST_1[305].FA_  ( .A(A[817]), .B(B[817]), .CI(
        C[817]), .S(S[817]), .CO(C[818]) );
  FA_1230 \FA_INST_0[1].FA_INST_1[306].FA_  ( .A(A[818]), .B(B[818]), .CI(
        C[818]), .S(S[818]), .CO(C[819]) );
  FA_1229 \FA_INST_0[1].FA_INST_1[307].FA_  ( .A(A[819]), .B(B[819]), .CI(
        C[819]), .S(S[819]), .CO(C[820]) );
  FA_1228 \FA_INST_0[1].FA_INST_1[308].FA_  ( .A(A[820]), .B(B[820]), .CI(
        C[820]), .S(S[820]), .CO(C[821]) );
  FA_1227 \FA_INST_0[1].FA_INST_1[309].FA_  ( .A(A[821]), .B(B[821]), .CI(
        C[821]), .S(S[821]), .CO(C[822]) );
  FA_1226 \FA_INST_0[1].FA_INST_1[310].FA_  ( .A(A[822]), .B(B[822]), .CI(
        C[822]), .S(S[822]), .CO(C[823]) );
  FA_1225 \FA_INST_0[1].FA_INST_1[311].FA_  ( .A(A[823]), .B(B[823]), .CI(
        C[823]), .S(S[823]), .CO(C[824]) );
  FA_1224 \FA_INST_0[1].FA_INST_1[312].FA_  ( .A(A[824]), .B(B[824]), .CI(
        C[824]), .S(S[824]), .CO(C[825]) );
  FA_1223 \FA_INST_0[1].FA_INST_1[313].FA_  ( .A(A[825]), .B(B[825]), .CI(
        C[825]), .S(S[825]), .CO(C[826]) );
  FA_1222 \FA_INST_0[1].FA_INST_1[314].FA_  ( .A(A[826]), .B(B[826]), .CI(
        C[826]), .S(S[826]), .CO(C[827]) );
  FA_1221 \FA_INST_0[1].FA_INST_1[315].FA_  ( .A(A[827]), .B(B[827]), .CI(
        C[827]), .S(S[827]), .CO(C[828]) );
  FA_1220 \FA_INST_0[1].FA_INST_1[316].FA_  ( .A(A[828]), .B(B[828]), .CI(
        C[828]), .S(S[828]), .CO(C[829]) );
  FA_1219 \FA_INST_0[1].FA_INST_1[317].FA_  ( .A(A[829]), .B(B[829]), .CI(
        C[829]), .S(S[829]), .CO(C[830]) );
  FA_1218 \FA_INST_0[1].FA_INST_1[318].FA_  ( .A(A[830]), .B(B[830]), .CI(
        C[830]), .S(S[830]), .CO(C[831]) );
  FA_1217 \FA_INST_0[1].FA_INST_1[319].FA_  ( .A(A[831]), .B(B[831]), .CI(
        C[831]), .S(S[831]), .CO(C[832]) );
  FA_1216 \FA_INST_0[1].FA_INST_1[320].FA_  ( .A(A[832]), .B(B[832]), .CI(
        C[832]), .S(S[832]), .CO(C[833]) );
  FA_1215 \FA_INST_0[1].FA_INST_1[321].FA_  ( .A(A[833]), .B(B[833]), .CI(
        C[833]), .S(S[833]), .CO(C[834]) );
  FA_1214 \FA_INST_0[1].FA_INST_1[322].FA_  ( .A(A[834]), .B(B[834]), .CI(
        C[834]), .S(S[834]), .CO(C[835]) );
  FA_1213 \FA_INST_0[1].FA_INST_1[323].FA_  ( .A(A[835]), .B(B[835]), .CI(
        C[835]), .S(S[835]), .CO(C[836]) );
  FA_1212 \FA_INST_0[1].FA_INST_1[324].FA_  ( .A(A[836]), .B(B[836]), .CI(
        C[836]), .S(S[836]), .CO(C[837]) );
  FA_1211 \FA_INST_0[1].FA_INST_1[325].FA_  ( .A(A[837]), .B(B[837]), .CI(
        C[837]), .S(S[837]), .CO(C[838]) );
  FA_1210 \FA_INST_0[1].FA_INST_1[326].FA_  ( .A(A[838]), .B(B[838]), .CI(
        C[838]), .S(S[838]), .CO(C[839]) );
  FA_1209 \FA_INST_0[1].FA_INST_1[327].FA_  ( .A(A[839]), .B(B[839]), .CI(
        C[839]), .S(S[839]), .CO(C[840]) );
  FA_1208 \FA_INST_0[1].FA_INST_1[328].FA_  ( .A(A[840]), .B(B[840]), .CI(
        C[840]), .S(S[840]), .CO(C[841]) );
  FA_1207 \FA_INST_0[1].FA_INST_1[329].FA_  ( .A(A[841]), .B(B[841]), .CI(
        C[841]), .S(S[841]), .CO(C[842]) );
  FA_1206 \FA_INST_0[1].FA_INST_1[330].FA_  ( .A(A[842]), .B(B[842]), .CI(
        C[842]), .S(S[842]), .CO(C[843]) );
  FA_1205 \FA_INST_0[1].FA_INST_1[331].FA_  ( .A(A[843]), .B(B[843]), .CI(
        C[843]), .S(S[843]), .CO(C[844]) );
  FA_1204 \FA_INST_0[1].FA_INST_1[332].FA_  ( .A(A[844]), .B(B[844]), .CI(
        C[844]), .S(S[844]), .CO(C[845]) );
  FA_1203 \FA_INST_0[1].FA_INST_1[333].FA_  ( .A(A[845]), .B(B[845]), .CI(
        C[845]), .S(S[845]), .CO(C[846]) );
  FA_1202 \FA_INST_0[1].FA_INST_1[334].FA_  ( .A(A[846]), .B(B[846]), .CI(
        C[846]), .S(S[846]), .CO(C[847]) );
  FA_1201 \FA_INST_0[1].FA_INST_1[335].FA_  ( .A(A[847]), .B(B[847]), .CI(
        C[847]), .S(S[847]), .CO(C[848]) );
  FA_1200 \FA_INST_0[1].FA_INST_1[336].FA_  ( .A(A[848]), .B(B[848]), .CI(
        C[848]), .S(S[848]), .CO(C[849]) );
  FA_1199 \FA_INST_0[1].FA_INST_1[337].FA_  ( .A(A[849]), .B(B[849]), .CI(
        C[849]), .S(S[849]), .CO(C[850]) );
  FA_1198 \FA_INST_0[1].FA_INST_1[338].FA_  ( .A(A[850]), .B(B[850]), .CI(
        C[850]), .S(S[850]), .CO(C[851]) );
  FA_1197 \FA_INST_0[1].FA_INST_1[339].FA_  ( .A(A[851]), .B(B[851]), .CI(
        C[851]), .S(S[851]), .CO(C[852]) );
  FA_1196 \FA_INST_0[1].FA_INST_1[340].FA_  ( .A(A[852]), .B(B[852]), .CI(
        C[852]), .S(S[852]), .CO(C[853]) );
  FA_1195 \FA_INST_0[1].FA_INST_1[341].FA_  ( .A(A[853]), .B(B[853]), .CI(
        C[853]), .S(S[853]), .CO(C[854]) );
  FA_1194 \FA_INST_0[1].FA_INST_1[342].FA_  ( .A(A[854]), .B(B[854]), .CI(
        C[854]), .S(S[854]), .CO(C[855]) );
  FA_1193 \FA_INST_0[1].FA_INST_1[343].FA_  ( .A(A[855]), .B(B[855]), .CI(
        C[855]), .S(S[855]), .CO(C[856]) );
  FA_1192 \FA_INST_0[1].FA_INST_1[344].FA_  ( .A(A[856]), .B(B[856]), .CI(
        C[856]), .S(S[856]), .CO(C[857]) );
  FA_1191 \FA_INST_0[1].FA_INST_1[345].FA_  ( .A(A[857]), .B(B[857]), .CI(
        C[857]), .S(S[857]), .CO(C[858]) );
  FA_1190 \FA_INST_0[1].FA_INST_1[346].FA_  ( .A(A[858]), .B(B[858]), .CI(
        C[858]), .S(S[858]), .CO(C[859]) );
  FA_1189 \FA_INST_0[1].FA_INST_1[347].FA_  ( .A(A[859]), .B(B[859]), .CI(
        C[859]), .S(S[859]), .CO(C[860]) );
  FA_1188 \FA_INST_0[1].FA_INST_1[348].FA_  ( .A(A[860]), .B(B[860]), .CI(
        C[860]), .S(S[860]), .CO(C[861]) );
  FA_1187 \FA_INST_0[1].FA_INST_1[349].FA_  ( .A(A[861]), .B(B[861]), .CI(
        C[861]), .S(S[861]), .CO(C[862]) );
  FA_1186 \FA_INST_0[1].FA_INST_1[350].FA_  ( .A(A[862]), .B(B[862]), .CI(
        C[862]), .S(S[862]), .CO(C[863]) );
  FA_1185 \FA_INST_0[1].FA_INST_1[351].FA_  ( .A(A[863]), .B(B[863]), .CI(
        C[863]), .S(S[863]), .CO(C[864]) );
  FA_1184 \FA_INST_0[1].FA_INST_1[352].FA_  ( .A(A[864]), .B(B[864]), .CI(
        C[864]), .S(S[864]), .CO(C[865]) );
  FA_1183 \FA_INST_0[1].FA_INST_1[353].FA_  ( .A(A[865]), .B(B[865]), .CI(
        C[865]), .S(S[865]), .CO(C[866]) );
  FA_1182 \FA_INST_0[1].FA_INST_1[354].FA_  ( .A(A[866]), .B(B[866]), .CI(
        C[866]), .S(S[866]), .CO(C[867]) );
  FA_1181 \FA_INST_0[1].FA_INST_1[355].FA_  ( .A(A[867]), .B(B[867]), .CI(
        C[867]), .S(S[867]), .CO(C[868]) );
  FA_1180 \FA_INST_0[1].FA_INST_1[356].FA_  ( .A(A[868]), .B(B[868]), .CI(
        C[868]), .S(S[868]), .CO(C[869]) );
  FA_1179 \FA_INST_0[1].FA_INST_1[357].FA_  ( .A(A[869]), .B(B[869]), .CI(
        C[869]), .S(S[869]), .CO(C[870]) );
  FA_1178 \FA_INST_0[1].FA_INST_1[358].FA_  ( .A(A[870]), .B(B[870]), .CI(
        C[870]), .S(S[870]), .CO(C[871]) );
  FA_1177 \FA_INST_0[1].FA_INST_1[359].FA_  ( .A(A[871]), .B(B[871]), .CI(
        C[871]), .S(S[871]), .CO(C[872]) );
  FA_1176 \FA_INST_0[1].FA_INST_1[360].FA_  ( .A(A[872]), .B(B[872]), .CI(
        C[872]), .S(S[872]), .CO(C[873]) );
  FA_1175 \FA_INST_0[1].FA_INST_1[361].FA_  ( .A(A[873]), .B(B[873]), .CI(
        C[873]), .S(S[873]), .CO(C[874]) );
  FA_1174 \FA_INST_0[1].FA_INST_1[362].FA_  ( .A(A[874]), .B(B[874]), .CI(
        C[874]), .S(S[874]), .CO(C[875]) );
  FA_1173 \FA_INST_0[1].FA_INST_1[363].FA_  ( .A(A[875]), .B(B[875]), .CI(
        C[875]), .S(S[875]), .CO(C[876]) );
  FA_1172 \FA_INST_0[1].FA_INST_1[364].FA_  ( .A(A[876]), .B(B[876]), .CI(
        C[876]), .S(S[876]), .CO(C[877]) );
  FA_1171 \FA_INST_0[1].FA_INST_1[365].FA_  ( .A(A[877]), .B(B[877]), .CI(
        C[877]), .S(S[877]), .CO(C[878]) );
  FA_1170 \FA_INST_0[1].FA_INST_1[366].FA_  ( .A(A[878]), .B(B[878]), .CI(
        C[878]), .S(S[878]), .CO(C[879]) );
  FA_1169 \FA_INST_0[1].FA_INST_1[367].FA_  ( .A(A[879]), .B(B[879]), .CI(
        C[879]), .S(S[879]), .CO(C[880]) );
  FA_1168 \FA_INST_0[1].FA_INST_1[368].FA_  ( .A(A[880]), .B(B[880]), .CI(
        C[880]), .S(S[880]), .CO(C[881]) );
  FA_1167 \FA_INST_0[1].FA_INST_1[369].FA_  ( .A(A[881]), .B(B[881]), .CI(
        C[881]), .S(S[881]), .CO(C[882]) );
  FA_1166 \FA_INST_0[1].FA_INST_1[370].FA_  ( .A(A[882]), .B(B[882]), .CI(
        C[882]), .S(S[882]), .CO(C[883]) );
  FA_1165 \FA_INST_0[1].FA_INST_1[371].FA_  ( .A(A[883]), .B(B[883]), .CI(
        C[883]), .S(S[883]), .CO(C[884]) );
  FA_1164 \FA_INST_0[1].FA_INST_1[372].FA_  ( .A(A[884]), .B(B[884]), .CI(
        C[884]), .S(S[884]), .CO(C[885]) );
  FA_1163 \FA_INST_0[1].FA_INST_1[373].FA_  ( .A(A[885]), .B(B[885]), .CI(
        C[885]), .S(S[885]), .CO(C[886]) );
  FA_1162 \FA_INST_0[1].FA_INST_1[374].FA_  ( .A(A[886]), .B(B[886]), .CI(
        C[886]), .S(S[886]), .CO(C[887]) );
  FA_1161 \FA_INST_0[1].FA_INST_1[375].FA_  ( .A(A[887]), .B(B[887]), .CI(
        C[887]), .S(S[887]), .CO(C[888]) );
  FA_1160 \FA_INST_0[1].FA_INST_1[376].FA_  ( .A(A[888]), .B(B[888]), .CI(
        C[888]), .S(S[888]), .CO(C[889]) );
  FA_1159 \FA_INST_0[1].FA_INST_1[377].FA_  ( .A(A[889]), .B(B[889]), .CI(
        C[889]), .S(S[889]), .CO(C[890]) );
  FA_1158 \FA_INST_0[1].FA_INST_1[378].FA_  ( .A(A[890]), .B(B[890]), .CI(
        C[890]), .S(S[890]), .CO(C[891]) );
  FA_1157 \FA_INST_0[1].FA_INST_1[379].FA_  ( .A(A[891]), .B(B[891]), .CI(
        C[891]), .S(S[891]), .CO(C[892]) );
  FA_1156 \FA_INST_0[1].FA_INST_1[380].FA_  ( .A(A[892]), .B(B[892]), .CI(
        C[892]), .S(S[892]), .CO(C[893]) );
  FA_1155 \FA_INST_0[1].FA_INST_1[381].FA_  ( .A(A[893]), .B(B[893]), .CI(
        C[893]), .S(S[893]), .CO(C[894]) );
  FA_1154 \FA_INST_0[1].FA_INST_1[382].FA_  ( .A(A[894]), .B(B[894]), .CI(
        C[894]), .S(S[894]), .CO(C[895]) );
  FA_1153 \FA_INST_0[1].FA_INST_1[383].FA_  ( .A(A[895]), .B(B[895]), .CI(
        C[895]), .S(S[895]), .CO(C[896]) );
  FA_1152 \FA_INST_0[1].FA_INST_1[384].FA_  ( .A(A[896]), .B(B[896]), .CI(
        C[896]), .S(S[896]), .CO(C[897]) );
  FA_1151 \FA_INST_0[1].FA_INST_1[385].FA_  ( .A(A[897]), .B(B[897]), .CI(
        C[897]), .S(S[897]), .CO(C[898]) );
  FA_1150 \FA_INST_0[1].FA_INST_1[386].FA_  ( .A(A[898]), .B(B[898]), .CI(
        C[898]), .S(S[898]), .CO(C[899]) );
  FA_1149 \FA_INST_0[1].FA_INST_1[387].FA_  ( .A(A[899]), .B(B[899]), .CI(
        C[899]), .S(S[899]), .CO(C[900]) );
  FA_1148 \FA_INST_0[1].FA_INST_1[388].FA_  ( .A(A[900]), .B(B[900]), .CI(
        C[900]), .S(S[900]), .CO(C[901]) );
  FA_1147 \FA_INST_0[1].FA_INST_1[389].FA_  ( .A(A[901]), .B(B[901]), .CI(
        C[901]), .S(S[901]), .CO(C[902]) );
  FA_1146 \FA_INST_0[1].FA_INST_1[390].FA_  ( .A(A[902]), .B(B[902]), .CI(
        C[902]), .S(S[902]), .CO(C[903]) );
  FA_1145 \FA_INST_0[1].FA_INST_1[391].FA_  ( .A(A[903]), .B(B[903]), .CI(
        C[903]), .S(S[903]), .CO(C[904]) );
  FA_1144 \FA_INST_0[1].FA_INST_1[392].FA_  ( .A(A[904]), .B(B[904]), .CI(
        C[904]), .S(S[904]), .CO(C[905]) );
  FA_1143 \FA_INST_0[1].FA_INST_1[393].FA_  ( .A(A[905]), .B(B[905]), .CI(
        C[905]), .S(S[905]), .CO(C[906]) );
  FA_1142 \FA_INST_0[1].FA_INST_1[394].FA_  ( .A(A[906]), .B(B[906]), .CI(
        C[906]), .S(S[906]), .CO(C[907]) );
  FA_1141 \FA_INST_0[1].FA_INST_1[395].FA_  ( .A(A[907]), .B(B[907]), .CI(
        C[907]), .S(S[907]), .CO(C[908]) );
  FA_1140 \FA_INST_0[1].FA_INST_1[396].FA_  ( .A(A[908]), .B(B[908]), .CI(
        C[908]), .S(S[908]), .CO(C[909]) );
  FA_1139 \FA_INST_0[1].FA_INST_1[397].FA_  ( .A(A[909]), .B(B[909]), .CI(
        C[909]), .S(S[909]), .CO(C[910]) );
  FA_1138 \FA_INST_0[1].FA_INST_1[398].FA_  ( .A(A[910]), .B(B[910]), .CI(
        C[910]), .S(S[910]), .CO(C[911]) );
  FA_1137 \FA_INST_0[1].FA_INST_1[399].FA_  ( .A(A[911]), .B(B[911]), .CI(
        C[911]), .S(S[911]), .CO(C[912]) );
  FA_1136 \FA_INST_0[1].FA_INST_1[400].FA_  ( .A(A[912]), .B(B[912]), .CI(
        C[912]), .S(S[912]), .CO(C[913]) );
  FA_1135 \FA_INST_0[1].FA_INST_1[401].FA_  ( .A(A[913]), .B(B[913]), .CI(
        C[913]), .S(S[913]), .CO(C[914]) );
  FA_1134 \FA_INST_0[1].FA_INST_1[402].FA_  ( .A(A[914]), .B(B[914]), .CI(
        C[914]), .S(S[914]), .CO(C[915]) );
  FA_1133 \FA_INST_0[1].FA_INST_1[403].FA_  ( .A(A[915]), .B(B[915]), .CI(
        C[915]), .S(S[915]), .CO(C[916]) );
  FA_1132 \FA_INST_0[1].FA_INST_1[404].FA_  ( .A(A[916]), .B(B[916]), .CI(
        C[916]), .S(S[916]), .CO(C[917]) );
  FA_1131 \FA_INST_0[1].FA_INST_1[405].FA_  ( .A(A[917]), .B(B[917]), .CI(
        C[917]), .S(S[917]), .CO(C[918]) );
  FA_1130 \FA_INST_0[1].FA_INST_1[406].FA_  ( .A(A[918]), .B(B[918]), .CI(
        C[918]), .S(S[918]), .CO(C[919]) );
  FA_1129 \FA_INST_0[1].FA_INST_1[407].FA_  ( .A(A[919]), .B(B[919]), .CI(
        C[919]), .S(S[919]), .CO(C[920]) );
  FA_1128 \FA_INST_0[1].FA_INST_1[408].FA_  ( .A(A[920]), .B(B[920]), .CI(
        C[920]), .S(S[920]), .CO(C[921]) );
  FA_1127 \FA_INST_0[1].FA_INST_1[409].FA_  ( .A(A[921]), .B(B[921]), .CI(
        C[921]), .S(S[921]), .CO(C[922]) );
  FA_1126 \FA_INST_0[1].FA_INST_1[410].FA_  ( .A(A[922]), .B(B[922]), .CI(
        C[922]), .S(S[922]), .CO(C[923]) );
  FA_1125 \FA_INST_0[1].FA_INST_1[411].FA_  ( .A(A[923]), .B(B[923]), .CI(
        C[923]), .S(S[923]), .CO(C[924]) );
  FA_1124 \FA_INST_0[1].FA_INST_1[412].FA_  ( .A(A[924]), .B(B[924]), .CI(
        C[924]), .S(S[924]), .CO(C[925]) );
  FA_1123 \FA_INST_0[1].FA_INST_1[413].FA_  ( .A(A[925]), .B(B[925]), .CI(
        C[925]), .S(S[925]), .CO(C[926]) );
  FA_1122 \FA_INST_0[1].FA_INST_1[414].FA_  ( .A(A[926]), .B(B[926]), .CI(
        C[926]), .S(S[926]), .CO(C[927]) );
  FA_1121 \FA_INST_0[1].FA_INST_1[415].FA_  ( .A(A[927]), .B(B[927]), .CI(
        C[927]), .S(S[927]), .CO(C[928]) );
  FA_1120 \FA_INST_0[1].FA_INST_1[416].FA_  ( .A(A[928]), .B(B[928]), .CI(
        C[928]), .S(S[928]), .CO(C[929]) );
  FA_1119 \FA_INST_0[1].FA_INST_1[417].FA_  ( .A(A[929]), .B(B[929]), .CI(
        C[929]), .S(S[929]), .CO(C[930]) );
  FA_1118 \FA_INST_0[1].FA_INST_1[418].FA_  ( .A(A[930]), .B(B[930]), .CI(
        C[930]), .S(S[930]), .CO(C[931]) );
  FA_1117 \FA_INST_0[1].FA_INST_1[419].FA_  ( .A(A[931]), .B(B[931]), .CI(
        C[931]), .S(S[931]), .CO(C[932]) );
  FA_1116 \FA_INST_0[1].FA_INST_1[420].FA_  ( .A(A[932]), .B(B[932]), .CI(
        C[932]), .S(S[932]), .CO(C[933]) );
  FA_1115 \FA_INST_0[1].FA_INST_1[421].FA_  ( .A(A[933]), .B(B[933]), .CI(
        C[933]), .S(S[933]), .CO(C[934]) );
  FA_1114 \FA_INST_0[1].FA_INST_1[422].FA_  ( .A(A[934]), .B(B[934]), .CI(
        C[934]), .S(S[934]), .CO(C[935]) );
  FA_1113 \FA_INST_0[1].FA_INST_1[423].FA_  ( .A(A[935]), .B(B[935]), .CI(
        C[935]), .S(S[935]), .CO(C[936]) );
  FA_1112 \FA_INST_0[1].FA_INST_1[424].FA_  ( .A(A[936]), .B(B[936]), .CI(
        C[936]), .S(S[936]), .CO(C[937]) );
  FA_1111 \FA_INST_0[1].FA_INST_1[425].FA_  ( .A(A[937]), .B(B[937]), .CI(
        C[937]), .S(S[937]), .CO(C[938]) );
  FA_1110 \FA_INST_0[1].FA_INST_1[426].FA_  ( .A(A[938]), .B(B[938]), .CI(
        C[938]), .S(S[938]), .CO(C[939]) );
  FA_1109 \FA_INST_0[1].FA_INST_1[427].FA_  ( .A(A[939]), .B(B[939]), .CI(
        C[939]), .S(S[939]), .CO(C[940]) );
  FA_1108 \FA_INST_0[1].FA_INST_1[428].FA_  ( .A(A[940]), .B(B[940]), .CI(
        C[940]), .S(S[940]), .CO(C[941]) );
  FA_1107 \FA_INST_0[1].FA_INST_1[429].FA_  ( .A(A[941]), .B(B[941]), .CI(
        C[941]), .S(S[941]), .CO(C[942]) );
  FA_1106 \FA_INST_0[1].FA_INST_1[430].FA_  ( .A(A[942]), .B(B[942]), .CI(
        C[942]), .S(S[942]), .CO(C[943]) );
  FA_1105 \FA_INST_0[1].FA_INST_1[431].FA_  ( .A(A[943]), .B(B[943]), .CI(
        C[943]), .S(S[943]), .CO(C[944]) );
  FA_1104 \FA_INST_0[1].FA_INST_1[432].FA_  ( .A(A[944]), .B(B[944]), .CI(
        C[944]), .S(S[944]), .CO(C[945]) );
  FA_1103 \FA_INST_0[1].FA_INST_1[433].FA_  ( .A(A[945]), .B(B[945]), .CI(
        C[945]), .S(S[945]), .CO(C[946]) );
  FA_1102 \FA_INST_0[1].FA_INST_1[434].FA_  ( .A(A[946]), .B(B[946]), .CI(
        C[946]), .S(S[946]), .CO(C[947]) );
  FA_1101 \FA_INST_0[1].FA_INST_1[435].FA_  ( .A(A[947]), .B(B[947]), .CI(
        C[947]), .S(S[947]), .CO(C[948]) );
  FA_1100 \FA_INST_0[1].FA_INST_1[436].FA_  ( .A(A[948]), .B(B[948]), .CI(
        C[948]), .S(S[948]), .CO(C[949]) );
  FA_1099 \FA_INST_0[1].FA_INST_1[437].FA_  ( .A(A[949]), .B(B[949]), .CI(
        C[949]), .S(S[949]), .CO(C[950]) );
  FA_1098 \FA_INST_0[1].FA_INST_1[438].FA_  ( .A(A[950]), .B(B[950]), .CI(
        C[950]), .S(S[950]), .CO(C[951]) );
  FA_1097 \FA_INST_0[1].FA_INST_1[439].FA_  ( .A(A[951]), .B(B[951]), .CI(
        C[951]), .S(S[951]), .CO(C[952]) );
  FA_1096 \FA_INST_0[1].FA_INST_1[440].FA_  ( .A(A[952]), .B(B[952]), .CI(
        C[952]), .S(S[952]), .CO(C[953]) );
  FA_1095 \FA_INST_0[1].FA_INST_1[441].FA_  ( .A(A[953]), .B(B[953]), .CI(
        C[953]), .S(S[953]), .CO(C[954]) );
  FA_1094 \FA_INST_0[1].FA_INST_1[442].FA_  ( .A(A[954]), .B(B[954]), .CI(
        C[954]), .S(S[954]), .CO(C[955]) );
  FA_1093 \FA_INST_0[1].FA_INST_1[443].FA_  ( .A(A[955]), .B(B[955]), .CI(
        C[955]), .S(S[955]), .CO(C[956]) );
  FA_1092 \FA_INST_0[1].FA_INST_1[444].FA_  ( .A(A[956]), .B(B[956]), .CI(
        C[956]), .S(S[956]), .CO(C[957]) );
  FA_1091 \FA_INST_0[1].FA_INST_1[445].FA_  ( .A(A[957]), .B(B[957]), .CI(
        C[957]), .S(S[957]), .CO(C[958]) );
  FA_1090 \FA_INST_0[1].FA_INST_1[446].FA_  ( .A(A[958]), .B(B[958]), .CI(
        C[958]), .S(S[958]), .CO(C[959]) );
  FA_1089 \FA_INST_0[1].FA_INST_1[447].FA_  ( .A(A[959]), .B(B[959]), .CI(
        C[959]), .S(S[959]), .CO(C[960]) );
  FA_1088 \FA_INST_0[1].FA_INST_1[448].FA_  ( .A(A[960]), .B(B[960]), .CI(
        C[960]), .S(S[960]), .CO(C[961]) );
  FA_1087 \FA_INST_0[1].FA_INST_1[449].FA_  ( .A(A[961]), .B(B[961]), .CI(
        C[961]), .S(S[961]), .CO(C[962]) );
  FA_1086 \FA_INST_0[1].FA_INST_1[450].FA_  ( .A(A[962]), .B(B[962]), .CI(
        C[962]), .S(S[962]), .CO(C[963]) );
  FA_1085 \FA_INST_0[1].FA_INST_1[451].FA_  ( .A(A[963]), .B(B[963]), .CI(
        C[963]), .S(S[963]), .CO(C[964]) );
  FA_1084 \FA_INST_0[1].FA_INST_1[452].FA_  ( .A(A[964]), .B(B[964]), .CI(
        C[964]), .S(S[964]), .CO(C[965]) );
  FA_1083 \FA_INST_0[1].FA_INST_1[453].FA_  ( .A(A[965]), .B(B[965]), .CI(
        C[965]), .S(S[965]), .CO(C[966]) );
  FA_1082 \FA_INST_0[1].FA_INST_1[454].FA_  ( .A(A[966]), .B(B[966]), .CI(
        C[966]), .S(S[966]), .CO(C[967]) );
  FA_1081 \FA_INST_0[1].FA_INST_1[455].FA_  ( .A(A[967]), .B(B[967]), .CI(
        C[967]), .S(S[967]), .CO(C[968]) );
  FA_1080 \FA_INST_0[1].FA_INST_1[456].FA_  ( .A(A[968]), .B(B[968]), .CI(
        C[968]), .S(S[968]), .CO(C[969]) );
  FA_1079 \FA_INST_0[1].FA_INST_1[457].FA_  ( .A(A[969]), .B(B[969]), .CI(
        C[969]), .S(S[969]), .CO(C[970]) );
  FA_1078 \FA_INST_0[1].FA_INST_1[458].FA_  ( .A(A[970]), .B(B[970]), .CI(
        C[970]), .S(S[970]), .CO(C[971]) );
  FA_1077 \FA_INST_0[1].FA_INST_1[459].FA_  ( .A(A[971]), .B(B[971]), .CI(
        C[971]), .S(S[971]), .CO(C[972]) );
  FA_1076 \FA_INST_0[1].FA_INST_1[460].FA_  ( .A(A[972]), .B(B[972]), .CI(
        C[972]), .S(S[972]), .CO(C[973]) );
  FA_1075 \FA_INST_0[1].FA_INST_1[461].FA_  ( .A(A[973]), .B(B[973]), .CI(
        C[973]), .S(S[973]), .CO(C[974]) );
  FA_1074 \FA_INST_0[1].FA_INST_1[462].FA_  ( .A(A[974]), .B(B[974]), .CI(
        C[974]), .S(S[974]), .CO(C[975]) );
  FA_1073 \FA_INST_0[1].FA_INST_1[463].FA_  ( .A(A[975]), .B(B[975]), .CI(
        C[975]), .S(S[975]), .CO(C[976]) );
  FA_1072 \FA_INST_0[1].FA_INST_1[464].FA_  ( .A(A[976]), .B(B[976]), .CI(
        C[976]), .S(S[976]), .CO(C[977]) );
  FA_1071 \FA_INST_0[1].FA_INST_1[465].FA_  ( .A(A[977]), .B(B[977]), .CI(
        C[977]), .S(S[977]), .CO(C[978]) );
  FA_1070 \FA_INST_0[1].FA_INST_1[466].FA_  ( .A(A[978]), .B(B[978]), .CI(
        C[978]), .S(S[978]), .CO(C[979]) );
  FA_1069 \FA_INST_0[1].FA_INST_1[467].FA_  ( .A(A[979]), .B(B[979]), .CI(
        C[979]), .S(S[979]), .CO(C[980]) );
  FA_1068 \FA_INST_0[1].FA_INST_1[468].FA_  ( .A(A[980]), .B(B[980]), .CI(
        C[980]), .S(S[980]), .CO(C[981]) );
  FA_1067 \FA_INST_0[1].FA_INST_1[469].FA_  ( .A(A[981]), .B(B[981]), .CI(
        C[981]), .S(S[981]), .CO(C[982]) );
  FA_1066 \FA_INST_0[1].FA_INST_1[470].FA_  ( .A(A[982]), .B(B[982]), .CI(
        C[982]), .S(S[982]), .CO(C[983]) );
  FA_1065 \FA_INST_0[1].FA_INST_1[471].FA_  ( .A(A[983]), .B(B[983]), .CI(
        C[983]), .S(S[983]), .CO(C[984]) );
  FA_1064 \FA_INST_0[1].FA_INST_1[472].FA_  ( .A(A[984]), .B(B[984]), .CI(
        C[984]), .S(S[984]), .CO(C[985]) );
  FA_1063 \FA_INST_0[1].FA_INST_1[473].FA_  ( .A(A[985]), .B(B[985]), .CI(
        C[985]), .S(S[985]), .CO(C[986]) );
  FA_1062 \FA_INST_0[1].FA_INST_1[474].FA_  ( .A(A[986]), .B(B[986]), .CI(
        C[986]), .S(S[986]), .CO(C[987]) );
  FA_1061 \FA_INST_0[1].FA_INST_1[475].FA_  ( .A(A[987]), .B(B[987]), .CI(
        C[987]), .S(S[987]), .CO(C[988]) );
  FA_1060 \FA_INST_0[1].FA_INST_1[476].FA_  ( .A(A[988]), .B(B[988]), .CI(
        C[988]), .S(S[988]), .CO(C[989]) );
  FA_1059 \FA_INST_0[1].FA_INST_1[477].FA_  ( .A(A[989]), .B(B[989]), .CI(
        C[989]), .S(S[989]), .CO(C[990]) );
  FA_1058 \FA_INST_0[1].FA_INST_1[478].FA_  ( .A(A[990]), .B(B[990]), .CI(
        C[990]), .S(S[990]), .CO(C[991]) );
  FA_1057 \FA_INST_0[1].FA_INST_1[479].FA_  ( .A(A[991]), .B(B[991]), .CI(
        C[991]), .S(S[991]), .CO(C[992]) );
  FA_1056 \FA_INST_0[1].FA_INST_1[480].FA_  ( .A(A[992]), .B(B[992]), .CI(
        C[992]), .S(S[992]), .CO(C[993]) );
  FA_1055 \FA_INST_0[1].FA_INST_1[481].FA_  ( .A(A[993]), .B(B[993]), .CI(
        C[993]), .S(S[993]), .CO(C[994]) );
  FA_1054 \FA_INST_0[1].FA_INST_1[482].FA_  ( .A(A[994]), .B(B[994]), .CI(
        C[994]), .S(S[994]), .CO(C[995]) );
  FA_1053 \FA_INST_0[1].FA_INST_1[483].FA_  ( .A(A[995]), .B(B[995]), .CI(
        C[995]), .S(S[995]), .CO(C[996]) );
  FA_1052 \FA_INST_0[1].FA_INST_1[484].FA_  ( .A(A[996]), .B(B[996]), .CI(
        C[996]), .S(S[996]), .CO(C[997]) );
  FA_1051 \FA_INST_0[1].FA_INST_1[485].FA_  ( .A(A[997]), .B(B[997]), .CI(
        C[997]), .S(S[997]), .CO(C[998]) );
  FA_1050 \FA_INST_0[1].FA_INST_1[486].FA_  ( .A(A[998]), .B(B[998]), .CI(
        C[998]), .S(S[998]), .CO(C[999]) );
  FA_1049 \FA_INST_0[1].FA_INST_1[487].FA_  ( .A(A[999]), .B(B[999]), .CI(
        C[999]), .S(S[999]), .CO(C[1000]) );
  FA_1048 \FA_INST_0[1].FA_INST_1[488].FA_  ( .A(A[1000]), .B(B[1000]), .CI(
        C[1000]), .S(S[1000]), .CO(C[1001]) );
  FA_1047 \FA_INST_0[1].FA_INST_1[489].FA_  ( .A(A[1001]), .B(B[1001]), .CI(
        C[1001]), .S(S[1001]), .CO(C[1002]) );
  FA_1046 \FA_INST_0[1].FA_INST_1[490].FA_  ( .A(A[1002]), .B(B[1002]), .CI(
        C[1002]), .S(S[1002]), .CO(C[1003]) );
  FA_1045 \FA_INST_0[1].FA_INST_1[491].FA_  ( .A(A[1003]), .B(B[1003]), .CI(
        C[1003]), .S(S[1003]), .CO(C[1004]) );
  FA_1044 \FA_INST_0[1].FA_INST_1[492].FA_  ( .A(A[1004]), .B(B[1004]), .CI(
        C[1004]), .S(S[1004]), .CO(C[1005]) );
  FA_1043 \FA_INST_0[1].FA_INST_1[493].FA_  ( .A(A[1005]), .B(B[1005]), .CI(
        C[1005]), .S(S[1005]), .CO(C[1006]) );
  FA_1042 \FA_INST_0[1].FA_INST_1[494].FA_  ( .A(A[1006]), .B(B[1006]), .CI(
        C[1006]), .S(S[1006]), .CO(C[1007]) );
  FA_1041 \FA_INST_0[1].FA_INST_1[495].FA_  ( .A(A[1007]), .B(B[1007]), .CI(
        C[1007]), .S(S[1007]), .CO(C[1008]) );
  FA_1040 \FA_INST_0[1].FA_INST_1[496].FA_  ( .A(A[1008]), .B(B[1008]), .CI(
        C[1008]), .S(S[1008]), .CO(C[1009]) );
  FA_1039 \FA_INST_0[1].FA_INST_1[497].FA_  ( .A(A[1009]), .B(B[1009]), .CI(
        C[1009]), .S(S[1009]), .CO(C[1010]) );
  FA_1038 \FA_INST_0[1].FA_INST_1[498].FA_  ( .A(A[1010]), .B(B[1010]), .CI(
        C[1010]), .S(S[1010]), .CO(C[1011]) );
  FA_1037 \FA_INST_0[1].FA_INST_1[499].FA_  ( .A(A[1011]), .B(B[1011]), .CI(
        C[1011]), .S(S[1011]), .CO(C[1012]) );
  FA_1036 \FA_INST_0[1].FA_INST_1[500].FA_  ( .A(A[1012]), .B(B[1012]), .CI(
        C[1012]), .S(S[1012]), .CO(C[1013]) );
  FA_1035 \FA_INST_0[1].FA_INST_1[501].FA_  ( .A(A[1013]), .B(B[1013]), .CI(
        C[1013]), .S(S[1013]), .CO(C[1014]) );
  FA_1034 \FA_INST_0[1].FA_INST_1[502].FA_  ( .A(A[1014]), .B(B[1014]), .CI(
        C[1014]), .S(S[1014]), .CO(C[1015]) );
  FA_1033 \FA_INST_0[1].FA_INST_1[503].FA_  ( .A(A[1015]), .B(B[1015]), .CI(
        C[1015]), .S(S[1015]), .CO(C[1016]) );
  FA_1032 \FA_INST_0[1].FA_INST_1[504].FA_  ( .A(A[1016]), .B(B[1016]), .CI(
        C[1016]), .S(S[1016]), .CO(C[1017]) );
  FA_1031 \FA_INST_0[1].FA_INST_1[505].FA_  ( .A(A[1017]), .B(B[1017]), .CI(
        C[1017]), .S(S[1017]), .CO(C[1018]) );
  FA_1030 \FA_INST_0[1].FA_INST_1[506].FA_  ( .A(A[1018]), .B(B[1018]), .CI(
        C[1018]), .S(S[1018]), .CO(C[1019]) );
  FA_1029 \FA_INST_0[1].FA_INST_1[507].FA_  ( .A(A[1019]), .B(B[1019]), .CI(
        C[1019]), .S(S[1019]), .CO(C[1020]) );
  FA_1028 \FA_INST_0[1].FA_INST_1[508].FA_  ( .A(A[1020]), .B(B[1020]), .CI(
        C[1020]), .S(S[1020]), .CO(C[1021]) );
  FA_1027 \FA_INST_0[1].FA_INST_1[509].FA_  ( .A(A[1021]), .B(B[1021]), .CI(
        C[1021]), .S(S[1021]), .CO(C[1022]) );
  FA_1026 \FA_INST_0[1].FA_INST_1[510].FA_  ( .A(1'b0), .B(B[1022]), .CI(
        C[1022]), .S(S[1022]) );
  FA_1025 \FA_INST_0[1].FA_INST_1[511].FA_  ( .A(1'b0), .B(B[1023]), .CI(1'b0), 
        .S(S[1023]) );
endmodule


module mult_N1024_CC512_DW01_add_0 ( A, B, CI, SUM, CO );
  input [1023:0] A;
  input [1023:0] B;
  output [1023:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905;

  NAND U2 ( .A(n27), .B(n30), .Z(n31) );
  XOR U3 ( .A(n1), .B(n2), .Z(SUM[9]) );
  NANDN U4 ( .A(n3), .B(n4), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[99]) );
  NANDN U6 ( .A(n7), .B(n8), .Z(n6) );
  ANDN U7 ( .B(n9), .A(n10), .Z(n5) );
  NAND U8 ( .A(n11), .B(n12), .Z(n9) );
  XOR U9 ( .A(n13), .B(n14), .Z(SUM[999]) );
  NANDN U10 ( .A(n15), .B(n16), .Z(n14) );
  ANDN U11 ( .B(n17), .A(n18), .Z(n13) );
  NAND U12 ( .A(n19), .B(n20), .Z(n17) );
  XNOR U13 ( .A(n19), .B(n21), .Z(SUM[998]) );
  NANDN U14 ( .A(n18), .B(n20), .Z(n21) );
  NANDN U15 ( .A(n22), .B(n23), .Z(n19) );
  NAND U16 ( .A(n24), .B(n25), .Z(n23) );
  XNOR U17 ( .A(n24), .B(n26), .Z(SUM[997]) );
  NANDN U18 ( .A(n22), .B(n25), .Z(n26) );
  NAND U19 ( .A(n27), .B(n28), .Z(n24) );
  NANDN U20 ( .A(n29), .B(n30), .Z(n28) );
  XOR U21 ( .A(n29), .B(n31), .Z(SUM[996]) );
  XOR U22 ( .A(n32), .B(n33), .Z(SUM[995]) );
  NANDN U23 ( .A(n34), .B(n35), .Z(n33) );
  ANDN U24 ( .B(n36), .A(n37), .Z(n32) );
  NAND U25 ( .A(n38), .B(n39), .Z(n36) );
  XNOR U26 ( .A(n38), .B(n40), .Z(SUM[994]) );
  NANDN U27 ( .A(n37), .B(n39), .Z(n40) );
  NANDN U28 ( .A(n41), .B(n42), .Z(n38) );
  NAND U29 ( .A(n43), .B(n44), .Z(n42) );
  XNOR U30 ( .A(n43), .B(n45), .Z(SUM[993]) );
  NANDN U31 ( .A(n41), .B(n44), .Z(n45) );
  NANDN U32 ( .A(n46), .B(n47), .Z(n43) );
  OR U33 ( .A(n48), .B(n49), .Z(n47) );
  XOR U34 ( .A(n48), .B(n50), .Z(SUM[992]) );
  OR U35 ( .A(n49), .B(n46), .Z(n50) );
  XOR U36 ( .A(n51), .B(n52), .Z(SUM[991]) );
  OR U37 ( .A(n53), .B(n54), .Z(n52) );
  ANDN U38 ( .B(n55), .A(n56), .Z(n51) );
  NANDN U39 ( .A(n57), .B(n58), .Z(n55) );
  XNOR U40 ( .A(n58), .B(n59), .Z(SUM[990]) );
  OR U41 ( .A(n57), .B(n56), .Z(n59) );
  NANDN U42 ( .A(n60), .B(n61), .Z(n58) );
  NANDN U43 ( .A(n62), .B(n63), .Z(n61) );
  XNOR U44 ( .A(n11), .B(n64), .Z(SUM[98]) );
  NANDN U45 ( .A(n10), .B(n12), .Z(n64) );
  NANDN U46 ( .A(n65), .B(n66), .Z(n11) );
  NAND U47 ( .A(n67), .B(n68), .Z(n66) );
  XNOR U48 ( .A(n63), .B(n69), .Z(SUM[989]) );
  OR U49 ( .A(n62), .B(n60), .Z(n69) );
  NANDN U50 ( .A(n70), .B(n71), .Z(n63) );
  NANDN U51 ( .A(n72), .B(n73), .Z(n71) );
  XNOR U52 ( .A(n73), .B(n74), .Z(SUM[988]) );
  OR U53 ( .A(n72), .B(n70), .Z(n74) );
  NANDN U54 ( .A(n75), .B(n76), .Z(n73) );
  NANDN U55 ( .A(n77), .B(n78), .Z(n76) );
  XOR U56 ( .A(n79), .B(n80), .Z(SUM[987]) );
  NANDN U57 ( .A(n81), .B(n82), .Z(n80) );
  ANDN U58 ( .B(n83), .A(n84), .Z(n79) );
  NAND U59 ( .A(n85), .B(n86), .Z(n83) );
  XNOR U60 ( .A(n85), .B(n87), .Z(SUM[986]) );
  NANDN U61 ( .A(n84), .B(n86), .Z(n87) );
  NANDN U62 ( .A(n88), .B(n89), .Z(n85) );
  NAND U63 ( .A(n90), .B(n91), .Z(n89) );
  XNOR U64 ( .A(n90), .B(n92), .Z(SUM[985]) );
  NANDN U65 ( .A(n88), .B(n91), .Z(n92) );
  NANDN U66 ( .A(n93), .B(n94), .Z(n90) );
  NAND U67 ( .A(n78), .B(n95), .Z(n94) );
  XNOR U68 ( .A(n78), .B(n96), .Z(SUM[984]) );
  NANDN U69 ( .A(n93), .B(n95), .Z(n96) );
  NANDN U70 ( .A(n97), .B(n98), .Z(n78) );
  OR U71 ( .A(n99), .B(n100), .Z(n98) );
  XOR U72 ( .A(n101), .B(n102), .Z(SUM[983]) );
  NANDN U73 ( .A(n103), .B(n104), .Z(n102) );
  ANDN U74 ( .B(n105), .A(n106), .Z(n101) );
  NAND U75 ( .A(n107), .B(n108), .Z(n105) );
  XNOR U76 ( .A(n107), .B(n109), .Z(SUM[982]) );
  NANDN U77 ( .A(n106), .B(n108), .Z(n109) );
  NANDN U78 ( .A(n110), .B(n111), .Z(n107) );
  NAND U79 ( .A(n112), .B(n113), .Z(n111) );
  XNOR U80 ( .A(n112), .B(n114), .Z(SUM[981]) );
  NANDN U81 ( .A(n110), .B(n113), .Z(n114) );
  NANDN U82 ( .A(n115), .B(n116), .Z(n112) );
  NANDN U83 ( .A(n100), .B(n117), .Z(n116) );
  XOR U84 ( .A(n100), .B(n118), .Z(SUM[980]) );
  NANDN U85 ( .A(n115), .B(n117), .Z(n118) );
  NOR U86 ( .A(n119), .B(n120), .Z(n100) );
  XNOR U87 ( .A(n67), .B(n121), .Z(SUM[97]) );
  NANDN U88 ( .A(n65), .B(n68), .Z(n121) );
  NANDN U89 ( .A(n122), .B(n123), .Z(n67) );
  OR U90 ( .A(n124), .B(n125), .Z(n123) );
  XOR U91 ( .A(n126), .B(n127), .Z(SUM[979]) );
  NANDN U92 ( .A(n128), .B(n129), .Z(n127) );
  ANDN U93 ( .B(n130), .A(n131), .Z(n126) );
  NAND U94 ( .A(n132), .B(n133), .Z(n130) );
  XNOR U95 ( .A(n132), .B(n134), .Z(SUM[978]) );
  NANDN U96 ( .A(n131), .B(n133), .Z(n134) );
  NANDN U97 ( .A(n135), .B(n136), .Z(n132) );
  NAND U98 ( .A(n137), .B(n138), .Z(n136) );
  XNOR U99 ( .A(n137), .B(n139), .Z(SUM[977]) );
  NANDN U100 ( .A(n135), .B(n138), .Z(n139) );
  NANDN U101 ( .A(n140), .B(n141), .Z(n137) );
  OR U102 ( .A(n142), .B(n143), .Z(n141) );
  XOR U103 ( .A(n142), .B(n144), .Z(SUM[976]) );
  OR U104 ( .A(n143), .B(n140), .Z(n144) );
  XOR U105 ( .A(n145), .B(n146), .Z(SUM[975]) );
  OR U106 ( .A(n147), .B(n148), .Z(n146) );
  ANDN U107 ( .B(n149), .A(n150), .Z(n145) );
  NANDN U108 ( .A(n151), .B(n152), .Z(n149) );
  XNOR U109 ( .A(n152), .B(n153), .Z(SUM[974]) );
  OR U110 ( .A(n151), .B(n150), .Z(n153) );
  NANDN U111 ( .A(n154), .B(n155), .Z(n152) );
  NANDN U112 ( .A(n156), .B(n157), .Z(n155) );
  XNOR U113 ( .A(n157), .B(n158), .Z(SUM[973]) );
  OR U114 ( .A(n156), .B(n154), .Z(n158) );
  NANDN U115 ( .A(n159), .B(n160), .Z(n157) );
  NANDN U116 ( .A(n161), .B(n162), .Z(n160) );
  XNOR U117 ( .A(n162), .B(n163), .Z(SUM[972]) );
  OR U118 ( .A(n161), .B(n159), .Z(n163) );
  NANDN U119 ( .A(n164), .B(n165), .Z(n162) );
  NANDN U120 ( .A(n166), .B(n167), .Z(n165) );
  XOR U121 ( .A(n168), .B(n169), .Z(SUM[971]) );
  NANDN U122 ( .A(n170), .B(n171), .Z(n169) );
  ANDN U123 ( .B(n172), .A(n173), .Z(n168) );
  NAND U124 ( .A(n174), .B(n175), .Z(n172) );
  XNOR U125 ( .A(n174), .B(n176), .Z(SUM[970]) );
  NANDN U126 ( .A(n173), .B(n175), .Z(n176) );
  NANDN U127 ( .A(n177), .B(n178), .Z(n174) );
  NAND U128 ( .A(n179), .B(n180), .Z(n178) );
  XOR U129 ( .A(n125), .B(n181), .Z(SUM[96]) );
  OR U130 ( .A(n124), .B(n122), .Z(n181) );
  XNOR U131 ( .A(n179), .B(n182), .Z(SUM[969]) );
  NANDN U132 ( .A(n177), .B(n180), .Z(n182) );
  NANDN U133 ( .A(n183), .B(n184), .Z(n179) );
  NAND U134 ( .A(n167), .B(n185), .Z(n184) );
  XNOR U135 ( .A(n167), .B(n186), .Z(SUM[968]) );
  NANDN U136 ( .A(n183), .B(n185), .Z(n186) );
  NANDN U137 ( .A(n187), .B(n188), .Z(n167) );
  OR U138 ( .A(n189), .B(n190), .Z(n188) );
  XOR U139 ( .A(n191), .B(n192), .Z(SUM[967]) );
  NANDN U140 ( .A(n193), .B(n194), .Z(n192) );
  ANDN U141 ( .B(n195), .A(n196), .Z(n191) );
  NAND U142 ( .A(n197), .B(n198), .Z(n195) );
  XNOR U143 ( .A(n197), .B(n199), .Z(SUM[966]) );
  NANDN U144 ( .A(n196), .B(n198), .Z(n199) );
  NANDN U145 ( .A(n200), .B(n201), .Z(n197) );
  NAND U146 ( .A(n202), .B(n203), .Z(n201) );
  XNOR U147 ( .A(n202), .B(n204), .Z(SUM[965]) );
  NANDN U148 ( .A(n200), .B(n203), .Z(n204) );
  NANDN U149 ( .A(n205), .B(n206), .Z(n202) );
  NANDN U150 ( .A(n190), .B(n207), .Z(n206) );
  XOR U151 ( .A(n190), .B(n208), .Z(SUM[964]) );
  NANDN U152 ( .A(n205), .B(n207), .Z(n208) );
  NOR U153 ( .A(n209), .B(n210), .Z(n190) );
  XOR U154 ( .A(n211), .B(n212), .Z(SUM[963]) );
  NANDN U155 ( .A(n213), .B(n214), .Z(n212) );
  ANDN U156 ( .B(n215), .A(n216), .Z(n211) );
  NAND U157 ( .A(n217), .B(n218), .Z(n215) );
  XNOR U158 ( .A(n217), .B(n219), .Z(SUM[962]) );
  NANDN U159 ( .A(n216), .B(n218), .Z(n219) );
  NANDN U160 ( .A(n220), .B(n221), .Z(n217) );
  NAND U161 ( .A(n222), .B(n223), .Z(n221) );
  XNOR U162 ( .A(n222), .B(n224), .Z(SUM[961]) );
  NANDN U163 ( .A(n220), .B(n223), .Z(n224) );
  NANDN U164 ( .A(n225), .B(n226), .Z(n222) );
  OR U165 ( .A(n227), .B(n228), .Z(n226) );
  XOR U166 ( .A(n227), .B(n229), .Z(SUM[960]) );
  OR U167 ( .A(n228), .B(n225), .Z(n229) );
  XOR U168 ( .A(n230), .B(n231), .Z(SUM[95]) );
  NANDN U169 ( .A(n232), .B(n233), .Z(n231) );
  ANDN U170 ( .B(n234), .A(n235), .Z(n230) );
  NANDN U171 ( .A(n236), .B(n237), .Z(n234) );
  XOR U172 ( .A(n238), .B(n239), .Z(SUM[959]) );
  OR U173 ( .A(n240), .B(n241), .Z(n239) );
  ANDN U174 ( .B(n242), .A(n243), .Z(n238) );
  NANDN U175 ( .A(n244), .B(n245), .Z(n242) );
  XNOR U176 ( .A(n245), .B(n246), .Z(SUM[958]) );
  OR U177 ( .A(n244), .B(n243), .Z(n246) );
  NANDN U178 ( .A(n247), .B(n248), .Z(n245) );
  NANDN U179 ( .A(n249), .B(n250), .Z(n248) );
  XNOR U180 ( .A(n250), .B(n251), .Z(SUM[957]) );
  OR U181 ( .A(n249), .B(n247), .Z(n251) );
  NANDN U182 ( .A(n252), .B(n253), .Z(n250) );
  NAND U183 ( .A(n254), .B(n255), .Z(n253) );
  XNOR U184 ( .A(n254), .B(n256), .Z(SUM[956]) );
  NANDN U185 ( .A(n252), .B(n255), .Z(n256) );
  NANDN U186 ( .A(n257), .B(n258), .Z(n254) );
  NANDN U187 ( .A(n259), .B(n260), .Z(n258) );
  XOR U188 ( .A(n261), .B(n262), .Z(SUM[955]) );
  NANDN U189 ( .A(n263), .B(n264), .Z(n262) );
  ANDN U190 ( .B(n265), .A(n266), .Z(n261) );
  NAND U191 ( .A(n267), .B(n268), .Z(n265) );
  XNOR U192 ( .A(n267), .B(n269), .Z(SUM[954]) );
  NANDN U193 ( .A(n266), .B(n268), .Z(n269) );
  NANDN U194 ( .A(n270), .B(n271), .Z(n267) );
  NAND U195 ( .A(n272), .B(n273), .Z(n271) );
  XNOR U196 ( .A(n272), .B(n274), .Z(SUM[953]) );
  NANDN U197 ( .A(n270), .B(n273), .Z(n274) );
  NANDN U198 ( .A(n275), .B(n276), .Z(n272) );
  NAND U199 ( .A(n260), .B(n277), .Z(n276) );
  XNOR U200 ( .A(n260), .B(n278), .Z(SUM[952]) );
  NANDN U201 ( .A(n275), .B(n277), .Z(n278) );
  NANDN U202 ( .A(n279), .B(n280), .Z(n260) );
  NANDN U203 ( .A(n281), .B(n282), .Z(n280) );
  XOR U204 ( .A(n283), .B(n284), .Z(SUM[951]) );
  NANDN U205 ( .A(n285), .B(n286), .Z(n284) );
  ANDN U206 ( .B(n287), .A(n288), .Z(n283) );
  NAND U207 ( .A(n289), .B(n290), .Z(n287) );
  XNOR U208 ( .A(n289), .B(n291), .Z(SUM[950]) );
  NANDN U209 ( .A(n288), .B(n290), .Z(n291) );
  NANDN U210 ( .A(n292), .B(n293), .Z(n289) );
  NAND U211 ( .A(n294), .B(n295), .Z(n293) );
  XNOR U212 ( .A(n237), .B(n296), .Z(SUM[94]) );
  OR U213 ( .A(n236), .B(n235), .Z(n296) );
  NANDN U214 ( .A(n297), .B(n298), .Z(n237) );
  NAND U215 ( .A(n299), .B(n300), .Z(n298) );
  XNOR U216 ( .A(n294), .B(n301), .Z(SUM[949]) );
  NANDN U217 ( .A(n292), .B(n295), .Z(n301) );
  NANDN U218 ( .A(n302), .B(n303), .Z(n294) );
  NANDN U219 ( .A(n281), .B(n304), .Z(n303) );
  XOR U220 ( .A(n281), .B(n305), .Z(SUM[948]) );
  NANDN U221 ( .A(n302), .B(n304), .Z(n305) );
  ANDN U222 ( .B(n306), .A(n307), .Z(n281) );
  OR U223 ( .A(n308), .B(n309), .Z(n306) );
  XOR U224 ( .A(n310), .B(n311), .Z(SUM[947]) );
  NANDN U225 ( .A(n312), .B(n313), .Z(n311) );
  ANDN U226 ( .B(n314), .A(n315), .Z(n310) );
  NANDN U227 ( .A(n316), .B(n317), .Z(n314) );
  XNOR U228 ( .A(n317), .B(n318), .Z(SUM[946]) );
  OR U229 ( .A(n316), .B(n315), .Z(n318) );
  NANDN U230 ( .A(n319), .B(n320), .Z(n317) );
  NAND U231 ( .A(n321), .B(n322), .Z(n320) );
  XNOR U232 ( .A(n321), .B(n323), .Z(SUM[945]) );
  NANDN U233 ( .A(n319), .B(n322), .Z(n323) );
  NANDN U234 ( .A(n324), .B(n325), .Z(n321) );
  NANDN U235 ( .A(n309), .B(n326), .Z(n325) );
  XOR U236 ( .A(n309), .B(n327), .Z(SUM[944]) );
  NANDN U237 ( .A(n324), .B(n326), .Z(n327) );
  XOR U238 ( .A(n328), .B(n329), .Z(SUM[943]) );
  OR U239 ( .A(n330), .B(n331), .Z(n329) );
  ANDN U240 ( .B(n332), .A(n333), .Z(n328) );
  NANDN U241 ( .A(n334), .B(n335), .Z(n332) );
  XNOR U242 ( .A(n335), .B(n336), .Z(SUM[942]) );
  OR U243 ( .A(n334), .B(n333), .Z(n336) );
  NANDN U244 ( .A(n337), .B(n338), .Z(n335) );
  NANDN U245 ( .A(n339), .B(n340), .Z(n338) );
  XNOR U246 ( .A(n340), .B(n341), .Z(SUM[941]) );
  OR U247 ( .A(n339), .B(n337), .Z(n341) );
  NANDN U248 ( .A(n342), .B(n343), .Z(n340) );
  NAND U249 ( .A(n344), .B(n345), .Z(n343) );
  XNOR U250 ( .A(n344), .B(n346), .Z(SUM[940]) );
  NANDN U251 ( .A(n342), .B(n345), .Z(n346) );
  NANDN U252 ( .A(n347), .B(n348), .Z(n344) );
  NANDN U253 ( .A(n349), .B(n350), .Z(n348) );
  XNOR U254 ( .A(n299), .B(n351), .Z(SUM[93]) );
  NANDN U255 ( .A(n297), .B(n300), .Z(n351) );
  NANDN U256 ( .A(n352), .B(n353), .Z(n299) );
  NANDN U257 ( .A(n354), .B(n355), .Z(n353) );
  XOR U258 ( .A(n356), .B(n357), .Z(SUM[939]) );
  NANDN U259 ( .A(n358), .B(n359), .Z(n357) );
  ANDN U260 ( .B(n360), .A(n361), .Z(n356) );
  NAND U261 ( .A(n362), .B(n363), .Z(n360) );
  XNOR U262 ( .A(n362), .B(n364), .Z(SUM[938]) );
  NANDN U263 ( .A(n361), .B(n363), .Z(n364) );
  NANDN U264 ( .A(n365), .B(n366), .Z(n362) );
  NAND U265 ( .A(n367), .B(n368), .Z(n366) );
  XNOR U266 ( .A(n367), .B(n369), .Z(SUM[937]) );
  NANDN U267 ( .A(n365), .B(n368), .Z(n369) );
  NANDN U268 ( .A(n370), .B(n371), .Z(n367) );
  NAND U269 ( .A(n350), .B(n372), .Z(n371) );
  XNOR U270 ( .A(n350), .B(n373), .Z(SUM[936]) );
  NANDN U271 ( .A(n370), .B(n372), .Z(n373) );
  NANDN U272 ( .A(n374), .B(n375), .Z(n350) );
  NANDN U273 ( .A(n376), .B(n377), .Z(n375) );
  XOR U274 ( .A(n378), .B(n379), .Z(SUM[935]) );
  NANDN U275 ( .A(n380), .B(n381), .Z(n379) );
  ANDN U276 ( .B(n382), .A(n383), .Z(n378) );
  NAND U277 ( .A(n384), .B(n385), .Z(n382) );
  XNOR U278 ( .A(n384), .B(n386), .Z(SUM[934]) );
  NANDN U279 ( .A(n383), .B(n385), .Z(n386) );
  NANDN U280 ( .A(n387), .B(n388), .Z(n384) );
  NAND U281 ( .A(n389), .B(n390), .Z(n388) );
  XNOR U282 ( .A(n389), .B(n391), .Z(SUM[933]) );
  NANDN U283 ( .A(n387), .B(n390), .Z(n391) );
  NANDN U284 ( .A(n392), .B(n393), .Z(n389) );
  NANDN U285 ( .A(n376), .B(n394), .Z(n393) );
  XOR U286 ( .A(n376), .B(n395), .Z(SUM[932]) );
  NANDN U287 ( .A(n392), .B(n394), .Z(n395) );
  ANDN U288 ( .B(n396), .A(n397), .Z(n376) );
  OR U289 ( .A(n398), .B(n399), .Z(n396) );
  XOR U290 ( .A(n400), .B(n401), .Z(SUM[931]) );
  NANDN U291 ( .A(n402), .B(n403), .Z(n401) );
  ANDN U292 ( .B(n404), .A(n405), .Z(n400) );
  NANDN U293 ( .A(n406), .B(n407), .Z(n404) );
  XNOR U294 ( .A(n407), .B(n408), .Z(SUM[930]) );
  OR U295 ( .A(n406), .B(n405), .Z(n408) );
  NANDN U296 ( .A(n409), .B(n410), .Z(n407) );
  NAND U297 ( .A(n411), .B(n412), .Z(n410) );
  XNOR U298 ( .A(n355), .B(n413), .Z(SUM[92]) );
  OR U299 ( .A(n354), .B(n352), .Z(n413) );
  NANDN U300 ( .A(n414), .B(n415), .Z(n355) );
  NANDN U301 ( .A(n416), .B(n417), .Z(n415) );
  XNOR U302 ( .A(n411), .B(n418), .Z(SUM[929]) );
  NANDN U303 ( .A(n409), .B(n412), .Z(n418) );
  NANDN U304 ( .A(n419), .B(n420), .Z(n411) );
  NANDN U305 ( .A(n399), .B(n421), .Z(n420) );
  XOR U306 ( .A(n399), .B(n422), .Z(SUM[928]) );
  NANDN U307 ( .A(n419), .B(n421), .Z(n422) );
  XOR U308 ( .A(n423), .B(n424), .Z(SUM[927]) );
  OR U309 ( .A(n425), .B(n426), .Z(n424) );
  ANDN U310 ( .B(n427), .A(n428), .Z(n423) );
  NANDN U311 ( .A(n429), .B(n430), .Z(n427) );
  XNOR U312 ( .A(n430), .B(n431), .Z(SUM[926]) );
  OR U313 ( .A(n429), .B(n428), .Z(n431) );
  NANDN U314 ( .A(n432), .B(n433), .Z(n430) );
  NANDN U315 ( .A(n434), .B(n435), .Z(n433) );
  XNOR U316 ( .A(n435), .B(n436), .Z(SUM[925]) );
  OR U317 ( .A(n434), .B(n432), .Z(n436) );
  NANDN U318 ( .A(n437), .B(n438), .Z(n435) );
  NAND U319 ( .A(n439), .B(n440), .Z(n438) );
  XNOR U320 ( .A(n439), .B(n441), .Z(SUM[924]) );
  NANDN U321 ( .A(n437), .B(n440), .Z(n441) );
  NANDN U322 ( .A(n442), .B(n443), .Z(n439) );
  NANDN U323 ( .A(n444), .B(n445), .Z(n443) );
  XOR U324 ( .A(n446), .B(n447), .Z(SUM[923]) );
  NANDN U325 ( .A(n448), .B(n449), .Z(n447) );
  ANDN U326 ( .B(n450), .A(n451), .Z(n446) );
  NAND U327 ( .A(n452), .B(n453), .Z(n450) );
  XNOR U328 ( .A(n452), .B(n454), .Z(SUM[922]) );
  NANDN U329 ( .A(n451), .B(n453), .Z(n454) );
  NANDN U330 ( .A(n455), .B(n456), .Z(n452) );
  NAND U331 ( .A(n457), .B(n458), .Z(n456) );
  XNOR U332 ( .A(n457), .B(n459), .Z(SUM[921]) );
  NANDN U333 ( .A(n455), .B(n458), .Z(n459) );
  NANDN U334 ( .A(n460), .B(n461), .Z(n457) );
  NAND U335 ( .A(n445), .B(n462), .Z(n461) );
  XNOR U336 ( .A(n445), .B(n463), .Z(SUM[920]) );
  NANDN U337 ( .A(n460), .B(n462), .Z(n463) );
  NANDN U338 ( .A(n464), .B(n465), .Z(n445) );
  NANDN U339 ( .A(n466), .B(n467), .Z(n465) );
  XOR U340 ( .A(n468), .B(n469), .Z(SUM[91]) );
  NANDN U341 ( .A(n470), .B(n471), .Z(n469) );
  ANDN U342 ( .B(n472), .A(n473), .Z(n468) );
  NAND U343 ( .A(n474), .B(n475), .Z(n472) );
  XOR U344 ( .A(n476), .B(n477), .Z(SUM[919]) );
  NANDN U345 ( .A(n478), .B(n479), .Z(n477) );
  ANDN U346 ( .B(n480), .A(n481), .Z(n476) );
  NAND U347 ( .A(n482), .B(n483), .Z(n480) );
  XNOR U348 ( .A(n482), .B(n484), .Z(SUM[918]) );
  NANDN U349 ( .A(n481), .B(n483), .Z(n484) );
  NANDN U350 ( .A(n485), .B(n486), .Z(n482) );
  NAND U351 ( .A(n487), .B(n488), .Z(n486) );
  XNOR U352 ( .A(n487), .B(n489), .Z(SUM[917]) );
  NANDN U353 ( .A(n485), .B(n488), .Z(n489) );
  NANDN U354 ( .A(n490), .B(n491), .Z(n487) );
  NANDN U355 ( .A(n466), .B(n492), .Z(n491) );
  XOR U356 ( .A(n466), .B(n493), .Z(SUM[916]) );
  NANDN U357 ( .A(n490), .B(n492), .Z(n493) );
  ANDN U358 ( .B(n494), .A(n495), .Z(n466) );
  OR U359 ( .A(n496), .B(n497), .Z(n494) );
  XOR U360 ( .A(n498), .B(n499), .Z(SUM[915]) );
  NANDN U361 ( .A(n500), .B(n501), .Z(n499) );
  ANDN U362 ( .B(n502), .A(n503), .Z(n498) );
  NANDN U363 ( .A(n504), .B(n505), .Z(n502) );
  XNOR U364 ( .A(n505), .B(n506), .Z(SUM[914]) );
  OR U365 ( .A(n504), .B(n503), .Z(n506) );
  NANDN U366 ( .A(n507), .B(n508), .Z(n505) );
  NAND U367 ( .A(n509), .B(n510), .Z(n508) );
  XNOR U368 ( .A(n509), .B(n511), .Z(SUM[913]) );
  NANDN U369 ( .A(n507), .B(n510), .Z(n511) );
  NANDN U370 ( .A(n512), .B(n513), .Z(n509) );
  NANDN U371 ( .A(n497), .B(n514), .Z(n513) );
  XOR U372 ( .A(n497), .B(n515), .Z(SUM[912]) );
  NANDN U373 ( .A(n512), .B(n514), .Z(n515) );
  XOR U374 ( .A(n516), .B(n517), .Z(SUM[911]) );
  OR U375 ( .A(n518), .B(n519), .Z(n517) );
  ANDN U376 ( .B(n520), .A(n521), .Z(n516) );
  NANDN U377 ( .A(n522), .B(n523), .Z(n520) );
  XNOR U378 ( .A(n523), .B(n524), .Z(SUM[910]) );
  OR U379 ( .A(n522), .B(n521), .Z(n524) );
  NANDN U380 ( .A(n525), .B(n526), .Z(n523) );
  NANDN U381 ( .A(n527), .B(n528), .Z(n526) );
  XNOR U382 ( .A(n474), .B(n529), .Z(SUM[90]) );
  NANDN U383 ( .A(n473), .B(n475), .Z(n529) );
  NANDN U384 ( .A(n530), .B(n531), .Z(n474) );
  NAND U385 ( .A(n532), .B(n533), .Z(n531) );
  XNOR U386 ( .A(n528), .B(n534), .Z(SUM[909]) );
  OR U387 ( .A(n527), .B(n525), .Z(n534) );
  NANDN U388 ( .A(n535), .B(n536), .Z(n528) );
  NAND U389 ( .A(n537), .B(n538), .Z(n536) );
  XNOR U390 ( .A(n537), .B(n539), .Z(SUM[908]) );
  NANDN U391 ( .A(n535), .B(n538), .Z(n539) );
  NANDN U392 ( .A(n540), .B(n541), .Z(n537) );
  NANDN U393 ( .A(n542), .B(n543), .Z(n541) );
  XOR U394 ( .A(n544), .B(n545), .Z(SUM[907]) );
  NANDN U395 ( .A(n546), .B(n547), .Z(n545) );
  ANDN U396 ( .B(n548), .A(n549), .Z(n544) );
  NAND U397 ( .A(n550), .B(n551), .Z(n548) );
  XNOR U398 ( .A(n550), .B(n552), .Z(SUM[906]) );
  NANDN U399 ( .A(n549), .B(n551), .Z(n552) );
  NANDN U400 ( .A(n553), .B(n554), .Z(n550) );
  NAND U401 ( .A(n555), .B(n556), .Z(n554) );
  XNOR U402 ( .A(n555), .B(n557), .Z(SUM[905]) );
  NANDN U403 ( .A(n553), .B(n556), .Z(n557) );
  NANDN U404 ( .A(n558), .B(n559), .Z(n555) );
  NAND U405 ( .A(n543), .B(n560), .Z(n559) );
  XNOR U406 ( .A(n543), .B(n561), .Z(SUM[904]) );
  NANDN U407 ( .A(n558), .B(n560), .Z(n561) );
  NANDN U408 ( .A(n562), .B(n563), .Z(n543) );
  NANDN U409 ( .A(n564), .B(n565), .Z(n563) );
  XOR U410 ( .A(n566), .B(n567), .Z(SUM[903]) );
  NANDN U411 ( .A(n568), .B(n569), .Z(n567) );
  ANDN U412 ( .B(n570), .A(n571), .Z(n566) );
  NAND U413 ( .A(n572), .B(n573), .Z(n570) );
  XNOR U414 ( .A(n572), .B(n574), .Z(SUM[902]) );
  NANDN U415 ( .A(n571), .B(n573), .Z(n574) );
  NANDN U416 ( .A(n575), .B(n576), .Z(n572) );
  NAND U417 ( .A(n577), .B(n578), .Z(n576) );
  XNOR U418 ( .A(n577), .B(n579), .Z(SUM[901]) );
  NANDN U419 ( .A(n575), .B(n578), .Z(n579) );
  NANDN U420 ( .A(n580), .B(n581), .Z(n577) );
  NANDN U421 ( .A(n564), .B(n582), .Z(n581) );
  XOR U422 ( .A(n564), .B(n583), .Z(SUM[900]) );
  NANDN U423 ( .A(n580), .B(n582), .Z(n583) );
  ANDN U424 ( .B(n584), .A(n585), .Z(n564) );
  OR U425 ( .A(n586), .B(n587), .Z(n584) );
  XOR U426 ( .A(n588), .B(n589), .Z(SUM[8]) );
  OR U427 ( .A(n590), .B(n591), .Z(n589) );
  XNOR U428 ( .A(n532), .B(n592), .Z(SUM[89]) );
  NANDN U429 ( .A(n530), .B(n533), .Z(n592) );
  NANDN U430 ( .A(n593), .B(n594), .Z(n532) );
  NAND U431 ( .A(n417), .B(n595), .Z(n594) );
  XOR U432 ( .A(n596), .B(n597), .Z(SUM[899]) );
  NANDN U433 ( .A(n598), .B(n599), .Z(n597) );
  ANDN U434 ( .B(n600), .A(n601), .Z(n596) );
  NANDN U435 ( .A(n602), .B(n603), .Z(n600) );
  XNOR U436 ( .A(n603), .B(n604), .Z(SUM[898]) );
  OR U437 ( .A(n602), .B(n601), .Z(n604) );
  NANDN U438 ( .A(n605), .B(n606), .Z(n603) );
  NAND U439 ( .A(n607), .B(n608), .Z(n606) );
  XNOR U440 ( .A(n607), .B(n609), .Z(SUM[897]) );
  NANDN U441 ( .A(n605), .B(n608), .Z(n609) );
  NANDN U442 ( .A(n610), .B(n611), .Z(n607) );
  NANDN U443 ( .A(n587), .B(n612), .Z(n611) );
  XOR U444 ( .A(n587), .B(n613), .Z(SUM[896]) );
  NANDN U445 ( .A(n610), .B(n612), .Z(n613) );
  XOR U446 ( .A(n614), .B(n615), .Z(SUM[895]) );
  OR U447 ( .A(n616), .B(n617), .Z(n615) );
  ANDN U448 ( .B(n618), .A(n619), .Z(n614) );
  NANDN U449 ( .A(n620), .B(n621), .Z(n618) );
  XNOR U450 ( .A(n621), .B(n622), .Z(SUM[894]) );
  OR U451 ( .A(n620), .B(n619), .Z(n622) );
  NANDN U452 ( .A(n623), .B(n624), .Z(n621) );
  NANDN U453 ( .A(n625), .B(n626), .Z(n624) );
  XNOR U454 ( .A(n626), .B(n627), .Z(SUM[893]) );
  OR U455 ( .A(n625), .B(n623), .Z(n627) );
  NANDN U456 ( .A(n628), .B(n629), .Z(n626) );
  NAND U457 ( .A(n630), .B(n631), .Z(n629) );
  XNOR U458 ( .A(n630), .B(n632), .Z(SUM[892]) );
  NANDN U459 ( .A(n628), .B(n631), .Z(n632) );
  NANDN U460 ( .A(n633), .B(n634), .Z(n630) );
  NANDN U461 ( .A(n635), .B(n636), .Z(n634) );
  XOR U462 ( .A(n637), .B(n638), .Z(SUM[891]) );
  NANDN U463 ( .A(n639), .B(n640), .Z(n638) );
  ANDN U464 ( .B(n641), .A(n642), .Z(n637) );
  NAND U465 ( .A(n643), .B(n644), .Z(n641) );
  XNOR U466 ( .A(n643), .B(n645), .Z(SUM[890]) );
  NANDN U467 ( .A(n642), .B(n644), .Z(n645) );
  NANDN U468 ( .A(n646), .B(n647), .Z(n643) );
  NAND U469 ( .A(n648), .B(n649), .Z(n647) );
  XNOR U470 ( .A(n417), .B(n650), .Z(SUM[88]) );
  NANDN U471 ( .A(n593), .B(n595), .Z(n650) );
  NANDN U472 ( .A(n651), .B(n652), .Z(n417) );
  NANDN U473 ( .A(n653), .B(n654), .Z(n652) );
  XNOR U474 ( .A(n648), .B(n655), .Z(SUM[889]) );
  NANDN U475 ( .A(n646), .B(n649), .Z(n655) );
  NANDN U476 ( .A(n656), .B(n657), .Z(n648) );
  NAND U477 ( .A(n636), .B(n658), .Z(n657) );
  XNOR U478 ( .A(n636), .B(n659), .Z(SUM[888]) );
  NANDN U479 ( .A(n656), .B(n658), .Z(n659) );
  NANDN U480 ( .A(n660), .B(n661), .Z(n636) );
  NANDN U481 ( .A(n662), .B(n663), .Z(n661) );
  XOR U482 ( .A(n664), .B(n665), .Z(SUM[887]) );
  NANDN U483 ( .A(n666), .B(n667), .Z(n665) );
  ANDN U484 ( .B(n668), .A(n669), .Z(n664) );
  NAND U485 ( .A(n670), .B(n671), .Z(n668) );
  XNOR U486 ( .A(n670), .B(n672), .Z(SUM[886]) );
  NANDN U487 ( .A(n669), .B(n671), .Z(n672) );
  NANDN U488 ( .A(n673), .B(n674), .Z(n670) );
  NAND U489 ( .A(n675), .B(n676), .Z(n674) );
  XNOR U490 ( .A(n675), .B(n677), .Z(SUM[885]) );
  NANDN U491 ( .A(n673), .B(n676), .Z(n677) );
  NANDN U492 ( .A(n678), .B(n679), .Z(n675) );
  NANDN U493 ( .A(n662), .B(n680), .Z(n679) );
  XOR U494 ( .A(n662), .B(n681), .Z(SUM[884]) );
  NANDN U495 ( .A(n678), .B(n680), .Z(n681) );
  ANDN U496 ( .B(n682), .A(n683), .Z(n662) );
  OR U497 ( .A(n684), .B(n685), .Z(n682) );
  XOR U498 ( .A(n686), .B(n687), .Z(SUM[883]) );
  NANDN U499 ( .A(n688), .B(n689), .Z(n687) );
  ANDN U500 ( .B(n690), .A(n691), .Z(n686) );
  NANDN U501 ( .A(n692), .B(n693), .Z(n690) );
  XNOR U502 ( .A(n693), .B(n694), .Z(SUM[882]) );
  OR U503 ( .A(n692), .B(n691), .Z(n694) );
  NANDN U504 ( .A(n695), .B(n696), .Z(n693) );
  NAND U505 ( .A(n697), .B(n698), .Z(n696) );
  XNOR U506 ( .A(n697), .B(n699), .Z(SUM[881]) );
  NANDN U507 ( .A(n695), .B(n698), .Z(n699) );
  NANDN U508 ( .A(n700), .B(n701), .Z(n697) );
  NANDN U509 ( .A(n685), .B(n702), .Z(n701) );
  XOR U510 ( .A(n685), .B(n703), .Z(SUM[880]) );
  NANDN U511 ( .A(n700), .B(n702), .Z(n703) );
  XOR U512 ( .A(n704), .B(n705), .Z(SUM[87]) );
  NANDN U513 ( .A(n706), .B(n707), .Z(n705) );
  ANDN U514 ( .B(n708), .A(n709), .Z(n704) );
  NAND U515 ( .A(n710), .B(n711), .Z(n708) );
  XOR U516 ( .A(n712), .B(n713), .Z(SUM[879]) );
  OR U517 ( .A(n714), .B(n715), .Z(n713) );
  ANDN U518 ( .B(n716), .A(n717), .Z(n712) );
  NANDN U519 ( .A(n718), .B(n719), .Z(n716) );
  XNOR U520 ( .A(n719), .B(n720), .Z(SUM[878]) );
  OR U521 ( .A(n718), .B(n717), .Z(n720) );
  NANDN U522 ( .A(n721), .B(n722), .Z(n719) );
  NANDN U523 ( .A(n723), .B(n724), .Z(n722) );
  XNOR U524 ( .A(n724), .B(n725), .Z(SUM[877]) );
  OR U525 ( .A(n723), .B(n721), .Z(n725) );
  NANDN U526 ( .A(n726), .B(n727), .Z(n724) );
  NAND U527 ( .A(n728), .B(n729), .Z(n727) );
  XNOR U528 ( .A(n728), .B(n730), .Z(SUM[876]) );
  NANDN U529 ( .A(n726), .B(n729), .Z(n730) );
  NANDN U530 ( .A(n731), .B(n732), .Z(n728) );
  NANDN U531 ( .A(n733), .B(n734), .Z(n732) );
  XOR U532 ( .A(n735), .B(n736), .Z(SUM[875]) );
  NANDN U533 ( .A(n737), .B(n738), .Z(n736) );
  ANDN U534 ( .B(n739), .A(n740), .Z(n735) );
  NAND U535 ( .A(n741), .B(n742), .Z(n739) );
  XNOR U536 ( .A(n741), .B(n743), .Z(SUM[874]) );
  NANDN U537 ( .A(n740), .B(n742), .Z(n743) );
  NANDN U538 ( .A(n744), .B(n745), .Z(n741) );
  NAND U539 ( .A(n746), .B(n747), .Z(n745) );
  XNOR U540 ( .A(n746), .B(n748), .Z(SUM[873]) );
  NANDN U541 ( .A(n744), .B(n747), .Z(n748) );
  NANDN U542 ( .A(n749), .B(n750), .Z(n746) );
  NAND U543 ( .A(n734), .B(n751), .Z(n750) );
  XNOR U544 ( .A(n734), .B(n752), .Z(SUM[872]) );
  NANDN U545 ( .A(n749), .B(n751), .Z(n752) );
  NANDN U546 ( .A(n753), .B(n754), .Z(n734) );
  NANDN U547 ( .A(n755), .B(n756), .Z(n754) );
  XOR U548 ( .A(n757), .B(n758), .Z(SUM[871]) );
  NANDN U549 ( .A(n759), .B(n760), .Z(n758) );
  ANDN U550 ( .B(n761), .A(n762), .Z(n757) );
  NAND U551 ( .A(n763), .B(n764), .Z(n761) );
  XNOR U552 ( .A(n763), .B(n765), .Z(SUM[870]) );
  NANDN U553 ( .A(n762), .B(n764), .Z(n765) );
  NANDN U554 ( .A(n766), .B(n767), .Z(n763) );
  NAND U555 ( .A(n768), .B(n769), .Z(n767) );
  XNOR U556 ( .A(n710), .B(n770), .Z(SUM[86]) );
  NANDN U557 ( .A(n709), .B(n711), .Z(n770) );
  NANDN U558 ( .A(n771), .B(n772), .Z(n710) );
  NAND U559 ( .A(n773), .B(n774), .Z(n772) );
  XNOR U560 ( .A(n768), .B(n775), .Z(SUM[869]) );
  NANDN U561 ( .A(n766), .B(n769), .Z(n775) );
  NANDN U562 ( .A(n776), .B(n777), .Z(n768) );
  NANDN U563 ( .A(n755), .B(n778), .Z(n777) );
  XOR U564 ( .A(n755), .B(n779), .Z(SUM[868]) );
  NANDN U565 ( .A(n776), .B(n778), .Z(n779) );
  ANDN U566 ( .B(n780), .A(n781), .Z(n755) );
  OR U567 ( .A(n782), .B(n783), .Z(n780) );
  XOR U568 ( .A(n784), .B(n785), .Z(SUM[867]) );
  NANDN U569 ( .A(n786), .B(n787), .Z(n785) );
  ANDN U570 ( .B(n788), .A(n789), .Z(n784) );
  NANDN U571 ( .A(n790), .B(n791), .Z(n788) );
  XNOR U572 ( .A(n791), .B(n792), .Z(SUM[866]) );
  OR U573 ( .A(n790), .B(n789), .Z(n792) );
  NANDN U574 ( .A(n793), .B(n794), .Z(n791) );
  NAND U575 ( .A(n795), .B(n796), .Z(n794) );
  XNOR U576 ( .A(n795), .B(n797), .Z(SUM[865]) );
  NANDN U577 ( .A(n793), .B(n796), .Z(n797) );
  NANDN U578 ( .A(n798), .B(n799), .Z(n795) );
  NANDN U579 ( .A(n783), .B(n800), .Z(n799) );
  XOR U580 ( .A(n783), .B(n801), .Z(SUM[864]) );
  NANDN U581 ( .A(n798), .B(n800), .Z(n801) );
  XOR U582 ( .A(n802), .B(n803), .Z(SUM[863]) );
  OR U583 ( .A(n804), .B(n805), .Z(n803) );
  ANDN U584 ( .B(n806), .A(n807), .Z(n802) );
  NANDN U585 ( .A(n808), .B(n809), .Z(n806) );
  XNOR U586 ( .A(n809), .B(n810), .Z(SUM[862]) );
  OR U587 ( .A(n808), .B(n807), .Z(n810) );
  NANDN U588 ( .A(n811), .B(n812), .Z(n809) );
  NANDN U589 ( .A(n813), .B(n814), .Z(n812) );
  XNOR U590 ( .A(n814), .B(n815), .Z(SUM[861]) );
  OR U591 ( .A(n813), .B(n811), .Z(n815) );
  NANDN U592 ( .A(n816), .B(n817), .Z(n814) );
  NAND U593 ( .A(n818), .B(n819), .Z(n817) );
  XNOR U594 ( .A(n818), .B(n820), .Z(SUM[860]) );
  NANDN U595 ( .A(n816), .B(n819), .Z(n820) );
  NANDN U596 ( .A(n821), .B(n822), .Z(n818) );
  NANDN U597 ( .A(n823), .B(n824), .Z(n822) );
  XNOR U598 ( .A(n773), .B(n825), .Z(SUM[85]) );
  NANDN U599 ( .A(n771), .B(n774), .Z(n825) );
  NANDN U600 ( .A(n826), .B(n827), .Z(n773) );
  NANDN U601 ( .A(n653), .B(n828), .Z(n827) );
  XOR U602 ( .A(n829), .B(n830), .Z(SUM[859]) );
  NANDN U603 ( .A(n831), .B(n832), .Z(n830) );
  ANDN U604 ( .B(n833), .A(n834), .Z(n829) );
  NAND U605 ( .A(n835), .B(n836), .Z(n833) );
  XNOR U606 ( .A(n835), .B(n837), .Z(SUM[858]) );
  NANDN U607 ( .A(n834), .B(n836), .Z(n837) );
  NANDN U608 ( .A(n838), .B(n839), .Z(n835) );
  NAND U609 ( .A(n840), .B(n841), .Z(n839) );
  XNOR U610 ( .A(n840), .B(n842), .Z(SUM[857]) );
  NANDN U611 ( .A(n838), .B(n841), .Z(n842) );
  NANDN U612 ( .A(n843), .B(n844), .Z(n840) );
  NAND U613 ( .A(n824), .B(n845), .Z(n844) );
  XNOR U614 ( .A(n824), .B(n846), .Z(SUM[856]) );
  NANDN U615 ( .A(n843), .B(n845), .Z(n846) );
  NANDN U616 ( .A(n847), .B(n848), .Z(n824) );
  NANDN U617 ( .A(n849), .B(n850), .Z(n848) );
  XOR U618 ( .A(n851), .B(n852), .Z(SUM[855]) );
  NANDN U619 ( .A(n853), .B(n854), .Z(n852) );
  ANDN U620 ( .B(n855), .A(n856), .Z(n851) );
  NAND U621 ( .A(n857), .B(n858), .Z(n855) );
  XNOR U622 ( .A(n857), .B(n859), .Z(SUM[854]) );
  NANDN U623 ( .A(n856), .B(n858), .Z(n859) );
  NANDN U624 ( .A(n860), .B(n861), .Z(n857) );
  NAND U625 ( .A(n862), .B(n863), .Z(n861) );
  XNOR U626 ( .A(n862), .B(n864), .Z(SUM[853]) );
  NANDN U627 ( .A(n860), .B(n863), .Z(n864) );
  NANDN U628 ( .A(n865), .B(n866), .Z(n862) );
  NANDN U629 ( .A(n849), .B(n867), .Z(n866) );
  XOR U630 ( .A(n849), .B(n868), .Z(SUM[852]) );
  NANDN U631 ( .A(n865), .B(n867), .Z(n868) );
  ANDN U632 ( .B(n869), .A(n870), .Z(n849) );
  OR U633 ( .A(n871), .B(n872), .Z(n869) );
  XOR U634 ( .A(n873), .B(n874), .Z(SUM[851]) );
  NANDN U635 ( .A(n875), .B(n876), .Z(n874) );
  ANDN U636 ( .B(n877), .A(n878), .Z(n873) );
  NANDN U637 ( .A(n879), .B(n880), .Z(n877) );
  XNOR U638 ( .A(n880), .B(n881), .Z(SUM[850]) );
  OR U639 ( .A(n879), .B(n878), .Z(n881) );
  NANDN U640 ( .A(n882), .B(n883), .Z(n880) );
  NAND U641 ( .A(n884), .B(n885), .Z(n883) );
  XOR U642 ( .A(n653), .B(n886), .Z(SUM[84]) );
  NANDN U643 ( .A(n826), .B(n828), .Z(n886) );
  ANDN U644 ( .B(n887), .A(n888), .Z(n653) );
  OR U645 ( .A(n889), .B(n890), .Z(n887) );
  XNOR U646 ( .A(n884), .B(n891), .Z(SUM[849]) );
  NANDN U647 ( .A(n882), .B(n885), .Z(n891) );
  NANDN U648 ( .A(n892), .B(n893), .Z(n884) );
  NANDN U649 ( .A(n872), .B(n894), .Z(n893) );
  XOR U650 ( .A(n872), .B(n895), .Z(SUM[848]) );
  NANDN U651 ( .A(n892), .B(n894), .Z(n895) );
  XOR U652 ( .A(n896), .B(n897), .Z(SUM[847]) );
  OR U653 ( .A(n898), .B(n899), .Z(n897) );
  ANDN U654 ( .B(n900), .A(n901), .Z(n896) );
  NANDN U655 ( .A(n902), .B(n903), .Z(n900) );
  XNOR U656 ( .A(n903), .B(n904), .Z(SUM[846]) );
  OR U657 ( .A(n902), .B(n901), .Z(n904) );
  NANDN U658 ( .A(n905), .B(n906), .Z(n903) );
  NANDN U659 ( .A(n907), .B(n908), .Z(n906) );
  XNOR U660 ( .A(n908), .B(n909), .Z(SUM[845]) );
  OR U661 ( .A(n907), .B(n905), .Z(n909) );
  NANDN U662 ( .A(n910), .B(n911), .Z(n908) );
  NAND U663 ( .A(n912), .B(n913), .Z(n911) );
  XNOR U664 ( .A(n912), .B(n914), .Z(SUM[844]) );
  NANDN U665 ( .A(n910), .B(n913), .Z(n914) );
  NANDN U666 ( .A(n915), .B(n916), .Z(n912) );
  NANDN U667 ( .A(n917), .B(n918), .Z(n916) );
  XOR U668 ( .A(n919), .B(n920), .Z(SUM[843]) );
  NANDN U669 ( .A(n921), .B(n922), .Z(n920) );
  ANDN U670 ( .B(n923), .A(n924), .Z(n919) );
  NAND U671 ( .A(n925), .B(n926), .Z(n923) );
  XNOR U672 ( .A(n925), .B(n927), .Z(SUM[842]) );
  NANDN U673 ( .A(n924), .B(n926), .Z(n927) );
  NANDN U674 ( .A(n928), .B(n929), .Z(n925) );
  NAND U675 ( .A(n930), .B(n931), .Z(n929) );
  XNOR U676 ( .A(n930), .B(n932), .Z(SUM[841]) );
  NANDN U677 ( .A(n928), .B(n931), .Z(n932) );
  NANDN U678 ( .A(n933), .B(n934), .Z(n930) );
  NAND U679 ( .A(n918), .B(n935), .Z(n934) );
  XNOR U680 ( .A(n918), .B(n936), .Z(SUM[840]) );
  NANDN U681 ( .A(n933), .B(n935), .Z(n936) );
  NANDN U682 ( .A(n937), .B(n938), .Z(n918) );
  NANDN U683 ( .A(n939), .B(n940), .Z(n938) );
  XOR U684 ( .A(n941), .B(n942), .Z(SUM[83]) );
  NANDN U685 ( .A(n943), .B(n944), .Z(n942) );
  ANDN U686 ( .B(n945), .A(n946), .Z(n941) );
  NANDN U687 ( .A(n947), .B(n948), .Z(n945) );
  XOR U688 ( .A(n949), .B(n950), .Z(SUM[839]) );
  NANDN U689 ( .A(n951), .B(n952), .Z(n950) );
  ANDN U690 ( .B(n953), .A(n954), .Z(n949) );
  NAND U691 ( .A(n955), .B(n956), .Z(n953) );
  XNOR U692 ( .A(n955), .B(n957), .Z(SUM[838]) );
  NANDN U693 ( .A(n954), .B(n956), .Z(n957) );
  NANDN U694 ( .A(n958), .B(n959), .Z(n955) );
  NAND U695 ( .A(n960), .B(n961), .Z(n959) );
  XNOR U696 ( .A(n960), .B(n962), .Z(SUM[837]) );
  NANDN U697 ( .A(n958), .B(n961), .Z(n962) );
  NANDN U698 ( .A(n963), .B(n964), .Z(n960) );
  NANDN U699 ( .A(n939), .B(n965), .Z(n964) );
  XOR U700 ( .A(n939), .B(n966), .Z(SUM[836]) );
  NANDN U701 ( .A(n963), .B(n965), .Z(n966) );
  ANDN U702 ( .B(n967), .A(n968), .Z(n939) );
  OR U703 ( .A(n969), .B(n970), .Z(n967) );
  XOR U704 ( .A(n971), .B(n972), .Z(SUM[835]) );
  NANDN U705 ( .A(n973), .B(n974), .Z(n972) );
  ANDN U706 ( .B(n975), .A(n976), .Z(n971) );
  NANDN U707 ( .A(n977), .B(n978), .Z(n975) );
  XNOR U708 ( .A(n978), .B(n979), .Z(SUM[834]) );
  OR U709 ( .A(n977), .B(n976), .Z(n979) );
  NANDN U710 ( .A(n980), .B(n981), .Z(n978) );
  NAND U711 ( .A(n982), .B(n983), .Z(n981) );
  XNOR U712 ( .A(n982), .B(n984), .Z(SUM[833]) );
  NANDN U713 ( .A(n980), .B(n983), .Z(n984) );
  NANDN U714 ( .A(n985), .B(n986), .Z(n982) );
  NANDN U715 ( .A(n970), .B(n987), .Z(n986) );
  XOR U716 ( .A(n970), .B(n988), .Z(SUM[832]) );
  NANDN U717 ( .A(n985), .B(n987), .Z(n988) );
  XOR U718 ( .A(n989), .B(n990), .Z(SUM[831]) );
  OR U719 ( .A(n991), .B(n992), .Z(n990) );
  ANDN U720 ( .B(n993), .A(n994), .Z(n989) );
  NANDN U721 ( .A(n995), .B(n996), .Z(n993) );
  XNOR U722 ( .A(n996), .B(n997), .Z(SUM[830]) );
  OR U723 ( .A(n995), .B(n994), .Z(n997) );
  NANDN U724 ( .A(n998), .B(n999), .Z(n996) );
  NANDN U725 ( .A(n1000), .B(n1001), .Z(n999) );
  XNOR U726 ( .A(n948), .B(n1002), .Z(SUM[82]) );
  OR U727 ( .A(n947), .B(n946), .Z(n1002) );
  NANDN U728 ( .A(n1003), .B(n1004), .Z(n948) );
  NAND U729 ( .A(n1005), .B(n1006), .Z(n1004) );
  XNOR U730 ( .A(n1001), .B(n1007), .Z(SUM[829]) );
  OR U731 ( .A(n1000), .B(n998), .Z(n1007) );
  NANDN U732 ( .A(n1008), .B(n1009), .Z(n1001) );
  NAND U733 ( .A(n1010), .B(n1011), .Z(n1009) );
  XNOR U734 ( .A(n1010), .B(n1012), .Z(SUM[828]) );
  NANDN U735 ( .A(n1008), .B(n1011), .Z(n1012) );
  NANDN U736 ( .A(n1013), .B(n1014), .Z(n1010) );
  NANDN U737 ( .A(n1015), .B(n1016), .Z(n1014) );
  XOR U738 ( .A(n1017), .B(n1018), .Z(SUM[827]) );
  NANDN U739 ( .A(n1019), .B(n1020), .Z(n1018) );
  ANDN U740 ( .B(n1021), .A(n1022), .Z(n1017) );
  NAND U741 ( .A(n1023), .B(n1024), .Z(n1021) );
  XNOR U742 ( .A(n1023), .B(n1025), .Z(SUM[826]) );
  NANDN U743 ( .A(n1022), .B(n1024), .Z(n1025) );
  NANDN U744 ( .A(n1026), .B(n1027), .Z(n1023) );
  NAND U745 ( .A(n1028), .B(n1029), .Z(n1027) );
  XNOR U746 ( .A(n1028), .B(n1030), .Z(SUM[825]) );
  NANDN U747 ( .A(n1026), .B(n1029), .Z(n1030) );
  NANDN U748 ( .A(n1031), .B(n1032), .Z(n1028) );
  NAND U749 ( .A(n1016), .B(n1033), .Z(n1032) );
  XNOR U750 ( .A(n1016), .B(n1034), .Z(SUM[824]) );
  NANDN U751 ( .A(n1031), .B(n1033), .Z(n1034) );
  NANDN U752 ( .A(n1035), .B(n1036), .Z(n1016) );
  NANDN U753 ( .A(n1037), .B(n1038), .Z(n1036) );
  XOR U754 ( .A(n1039), .B(n1040), .Z(SUM[823]) );
  NANDN U755 ( .A(n1041), .B(n1042), .Z(n1040) );
  ANDN U756 ( .B(n1043), .A(n1044), .Z(n1039) );
  NAND U757 ( .A(n1045), .B(n1046), .Z(n1043) );
  XNOR U758 ( .A(n1045), .B(n1047), .Z(SUM[822]) );
  NANDN U759 ( .A(n1044), .B(n1046), .Z(n1047) );
  NANDN U760 ( .A(n1048), .B(n1049), .Z(n1045) );
  NAND U761 ( .A(n1050), .B(n1051), .Z(n1049) );
  XNOR U762 ( .A(n1050), .B(n1052), .Z(SUM[821]) );
  NANDN U763 ( .A(n1048), .B(n1051), .Z(n1052) );
  NANDN U764 ( .A(n1053), .B(n1054), .Z(n1050) );
  NANDN U765 ( .A(n1037), .B(n1055), .Z(n1054) );
  XOR U766 ( .A(n1037), .B(n1056), .Z(SUM[820]) );
  NANDN U767 ( .A(n1053), .B(n1055), .Z(n1056) );
  ANDN U768 ( .B(n1057), .A(n1058), .Z(n1037) );
  OR U769 ( .A(n1059), .B(n1060), .Z(n1057) );
  XNOR U770 ( .A(n1005), .B(n1061), .Z(SUM[81]) );
  NANDN U771 ( .A(n1003), .B(n1006), .Z(n1061) );
  NANDN U772 ( .A(n1062), .B(n1063), .Z(n1005) );
  NANDN U773 ( .A(n890), .B(n1064), .Z(n1063) );
  XOR U774 ( .A(n1065), .B(n1066), .Z(SUM[819]) );
  NANDN U775 ( .A(n1067), .B(n1068), .Z(n1066) );
  ANDN U776 ( .B(n1069), .A(n1070), .Z(n1065) );
  NANDN U777 ( .A(n1071), .B(n1072), .Z(n1069) );
  XNOR U778 ( .A(n1072), .B(n1073), .Z(SUM[818]) );
  OR U779 ( .A(n1071), .B(n1070), .Z(n1073) );
  NANDN U780 ( .A(n1074), .B(n1075), .Z(n1072) );
  NAND U781 ( .A(n1076), .B(n1077), .Z(n1075) );
  XNOR U782 ( .A(n1076), .B(n1078), .Z(SUM[817]) );
  NANDN U783 ( .A(n1074), .B(n1077), .Z(n1078) );
  NANDN U784 ( .A(n1079), .B(n1080), .Z(n1076) );
  NANDN U785 ( .A(n1060), .B(n1081), .Z(n1080) );
  XOR U786 ( .A(n1060), .B(n1082), .Z(SUM[816]) );
  NANDN U787 ( .A(n1079), .B(n1081), .Z(n1082) );
  XOR U788 ( .A(n1083), .B(n1084), .Z(SUM[815]) );
  OR U789 ( .A(n1085), .B(n1086), .Z(n1084) );
  ANDN U790 ( .B(n1087), .A(n1088), .Z(n1083) );
  NANDN U791 ( .A(n1089), .B(n1090), .Z(n1087) );
  XNOR U792 ( .A(n1090), .B(n1091), .Z(SUM[814]) );
  OR U793 ( .A(n1089), .B(n1088), .Z(n1091) );
  NANDN U794 ( .A(n1092), .B(n1093), .Z(n1090) );
  NANDN U795 ( .A(n1094), .B(n1095), .Z(n1093) );
  XNOR U796 ( .A(n1095), .B(n1096), .Z(SUM[813]) );
  OR U797 ( .A(n1094), .B(n1092), .Z(n1096) );
  NANDN U798 ( .A(n1097), .B(n1098), .Z(n1095) );
  NAND U799 ( .A(n1099), .B(n1100), .Z(n1098) );
  XNOR U800 ( .A(n1099), .B(n1101), .Z(SUM[812]) );
  NANDN U801 ( .A(n1097), .B(n1100), .Z(n1101) );
  NANDN U802 ( .A(n1102), .B(n1103), .Z(n1099) );
  NANDN U803 ( .A(n1104), .B(n1105), .Z(n1103) );
  XOR U804 ( .A(n1106), .B(n1107), .Z(SUM[811]) );
  NANDN U805 ( .A(n1108), .B(n1109), .Z(n1107) );
  ANDN U806 ( .B(n1110), .A(n1111), .Z(n1106) );
  NAND U807 ( .A(n1112), .B(n1113), .Z(n1110) );
  XNOR U808 ( .A(n1112), .B(n1114), .Z(SUM[810]) );
  NANDN U809 ( .A(n1111), .B(n1113), .Z(n1114) );
  NANDN U810 ( .A(n1115), .B(n1116), .Z(n1112) );
  NAND U811 ( .A(n1117), .B(n1118), .Z(n1116) );
  XOR U812 ( .A(n890), .B(n1119), .Z(SUM[80]) );
  NANDN U813 ( .A(n1062), .B(n1064), .Z(n1119) );
  XNOR U814 ( .A(n1117), .B(n1120), .Z(SUM[809]) );
  NANDN U815 ( .A(n1115), .B(n1118), .Z(n1120) );
  NANDN U816 ( .A(n1121), .B(n1122), .Z(n1117) );
  NAND U817 ( .A(n1105), .B(n1123), .Z(n1122) );
  XNOR U818 ( .A(n1105), .B(n1124), .Z(SUM[808]) );
  NANDN U819 ( .A(n1121), .B(n1123), .Z(n1124) );
  NANDN U820 ( .A(n1125), .B(n1126), .Z(n1105) );
  NANDN U821 ( .A(n1127), .B(n1128), .Z(n1126) );
  XOR U822 ( .A(n1129), .B(n1130), .Z(SUM[807]) );
  NANDN U823 ( .A(n1131), .B(n1132), .Z(n1130) );
  ANDN U824 ( .B(n1133), .A(n1134), .Z(n1129) );
  NAND U825 ( .A(n1135), .B(n1136), .Z(n1133) );
  XNOR U826 ( .A(n1135), .B(n1137), .Z(SUM[806]) );
  NANDN U827 ( .A(n1134), .B(n1136), .Z(n1137) );
  NANDN U828 ( .A(n1138), .B(n1139), .Z(n1135) );
  NAND U829 ( .A(n1140), .B(n1141), .Z(n1139) );
  XNOR U830 ( .A(n1140), .B(n1142), .Z(SUM[805]) );
  NANDN U831 ( .A(n1138), .B(n1141), .Z(n1142) );
  NANDN U832 ( .A(n1143), .B(n1144), .Z(n1140) );
  NANDN U833 ( .A(n1127), .B(n1145), .Z(n1144) );
  XOR U834 ( .A(n1127), .B(n1146), .Z(SUM[804]) );
  NANDN U835 ( .A(n1143), .B(n1145), .Z(n1146) );
  ANDN U836 ( .B(n1147), .A(n1148), .Z(n1127) );
  OR U837 ( .A(n1149), .B(n1150), .Z(n1147) );
  XOR U838 ( .A(n1151), .B(n1152), .Z(SUM[803]) );
  NANDN U839 ( .A(n1153), .B(n1154), .Z(n1152) );
  ANDN U840 ( .B(n1155), .A(n1156), .Z(n1151) );
  NANDN U841 ( .A(n1157), .B(n1158), .Z(n1155) );
  XNOR U842 ( .A(n1158), .B(n1159), .Z(SUM[802]) );
  OR U843 ( .A(n1157), .B(n1156), .Z(n1159) );
  NANDN U844 ( .A(n1160), .B(n1161), .Z(n1158) );
  NAND U845 ( .A(n1162), .B(n1163), .Z(n1161) );
  XNOR U846 ( .A(n1162), .B(n1164), .Z(SUM[801]) );
  NANDN U847 ( .A(n1160), .B(n1163), .Z(n1164) );
  NANDN U848 ( .A(n1165), .B(n1166), .Z(n1162) );
  NANDN U849 ( .A(n1150), .B(n1167), .Z(n1166) );
  XOR U850 ( .A(n1150), .B(n1168), .Z(SUM[800]) );
  NANDN U851 ( .A(n1165), .B(n1167), .Z(n1168) );
  XOR U852 ( .A(n1169), .B(n1170), .Z(SUM[7]) );
  OR U853 ( .A(n1171), .B(n1172), .Z(n1170) );
  ANDN U854 ( .B(n1173), .A(n1174), .Z(n1169) );
  XOR U855 ( .A(n1175), .B(n1176), .Z(SUM[79]) );
  NANDN U856 ( .A(n1177), .B(n1178), .Z(n1176) );
  ANDN U857 ( .B(n1179), .A(n1180), .Z(n1175) );
  NANDN U858 ( .A(n1181), .B(n1182), .Z(n1179) );
  XOR U859 ( .A(n1183), .B(n1184), .Z(SUM[799]) );
  OR U860 ( .A(n1185), .B(n1186), .Z(n1184) );
  ANDN U861 ( .B(n1187), .A(n1188), .Z(n1183) );
  NANDN U862 ( .A(n1189), .B(n1190), .Z(n1187) );
  XNOR U863 ( .A(n1190), .B(n1191), .Z(SUM[798]) );
  OR U864 ( .A(n1189), .B(n1188), .Z(n1191) );
  NANDN U865 ( .A(n1192), .B(n1193), .Z(n1190) );
  NANDN U866 ( .A(n1194), .B(n1195), .Z(n1193) );
  XNOR U867 ( .A(n1195), .B(n1196), .Z(SUM[797]) );
  OR U868 ( .A(n1194), .B(n1192), .Z(n1196) );
  NANDN U869 ( .A(n1197), .B(n1198), .Z(n1195) );
  NAND U870 ( .A(n1199), .B(n1200), .Z(n1198) );
  XNOR U871 ( .A(n1199), .B(n1201), .Z(SUM[796]) );
  NANDN U872 ( .A(n1197), .B(n1200), .Z(n1201) );
  NANDN U873 ( .A(n1202), .B(n1203), .Z(n1199) );
  NANDN U874 ( .A(n1204), .B(n1205), .Z(n1203) );
  XOR U875 ( .A(n1206), .B(n1207), .Z(SUM[795]) );
  NANDN U876 ( .A(n1208), .B(n1209), .Z(n1207) );
  ANDN U877 ( .B(n1210), .A(n1211), .Z(n1206) );
  NAND U878 ( .A(n1212), .B(n1213), .Z(n1210) );
  XNOR U879 ( .A(n1212), .B(n1214), .Z(SUM[794]) );
  NANDN U880 ( .A(n1211), .B(n1213), .Z(n1214) );
  NANDN U881 ( .A(n1215), .B(n1216), .Z(n1212) );
  NAND U882 ( .A(n1217), .B(n1218), .Z(n1216) );
  XNOR U883 ( .A(n1217), .B(n1219), .Z(SUM[793]) );
  NANDN U884 ( .A(n1215), .B(n1218), .Z(n1219) );
  NANDN U885 ( .A(n1220), .B(n1221), .Z(n1217) );
  NAND U886 ( .A(n1205), .B(n1222), .Z(n1221) );
  XNOR U887 ( .A(n1205), .B(n1223), .Z(SUM[792]) );
  NANDN U888 ( .A(n1220), .B(n1222), .Z(n1223) );
  NANDN U889 ( .A(n1224), .B(n1225), .Z(n1205) );
  NANDN U890 ( .A(n1226), .B(n1227), .Z(n1225) );
  XOR U891 ( .A(n1228), .B(n1229), .Z(SUM[791]) );
  NANDN U892 ( .A(n1230), .B(n1231), .Z(n1229) );
  ANDN U893 ( .B(n1232), .A(n1233), .Z(n1228) );
  NAND U894 ( .A(n1234), .B(n1235), .Z(n1232) );
  XNOR U895 ( .A(n1234), .B(n1236), .Z(SUM[790]) );
  NANDN U896 ( .A(n1233), .B(n1235), .Z(n1236) );
  NANDN U897 ( .A(n1237), .B(n1238), .Z(n1234) );
  NAND U898 ( .A(n1239), .B(n1240), .Z(n1238) );
  XNOR U899 ( .A(n1182), .B(n1241), .Z(SUM[78]) );
  OR U900 ( .A(n1181), .B(n1180), .Z(n1241) );
  NANDN U901 ( .A(n1242), .B(n1243), .Z(n1182) );
  NAND U902 ( .A(n1244), .B(n1245), .Z(n1243) );
  XNOR U903 ( .A(n1239), .B(n1246), .Z(SUM[789]) );
  NANDN U904 ( .A(n1237), .B(n1240), .Z(n1246) );
  NANDN U905 ( .A(n1247), .B(n1248), .Z(n1239) );
  NANDN U906 ( .A(n1226), .B(n1249), .Z(n1248) );
  XOR U907 ( .A(n1226), .B(n1250), .Z(SUM[788]) );
  NANDN U908 ( .A(n1247), .B(n1249), .Z(n1250) );
  ANDN U909 ( .B(n1251), .A(n1252), .Z(n1226) );
  OR U910 ( .A(n1253), .B(n1254), .Z(n1251) );
  XOR U911 ( .A(n1255), .B(n1256), .Z(SUM[787]) );
  NANDN U912 ( .A(n1257), .B(n1258), .Z(n1256) );
  ANDN U913 ( .B(n1259), .A(n1260), .Z(n1255) );
  NANDN U914 ( .A(n1261), .B(n1262), .Z(n1259) );
  XNOR U915 ( .A(n1262), .B(n1263), .Z(SUM[786]) );
  OR U916 ( .A(n1261), .B(n1260), .Z(n1263) );
  NANDN U917 ( .A(n1264), .B(n1265), .Z(n1262) );
  NAND U918 ( .A(n1266), .B(n1267), .Z(n1265) );
  XNOR U919 ( .A(n1266), .B(n1268), .Z(SUM[785]) );
  NANDN U920 ( .A(n1264), .B(n1267), .Z(n1268) );
  NANDN U921 ( .A(n1269), .B(n1270), .Z(n1266) );
  NANDN U922 ( .A(n1254), .B(n1271), .Z(n1270) );
  XOR U923 ( .A(n1254), .B(n1272), .Z(SUM[784]) );
  NANDN U924 ( .A(n1269), .B(n1271), .Z(n1272) );
  XOR U925 ( .A(n1273), .B(n1274), .Z(SUM[783]) );
  OR U926 ( .A(n1275), .B(n1276), .Z(n1274) );
  ANDN U927 ( .B(n1277), .A(n1278), .Z(n1273) );
  NANDN U928 ( .A(n1279), .B(n1280), .Z(n1277) );
  XNOR U929 ( .A(n1280), .B(n1281), .Z(SUM[782]) );
  OR U930 ( .A(n1279), .B(n1278), .Z(n1281) );
  NANDN U931 ( .A(n1282), .B(n1283), .Z(n1280) );
  NANDN U932 ( .A(n1284), .B(n1285), .Z(n1283) );
  XNOR U933 ( .A(n1285), .B(n1286), .Z(SUM[781]) );
  OR U934 ( .A(n1284), .B(n1282), .Z(n1286) );
  NANDN U935 ( .A(n1287), .B(n1288), .Z(n1285) );
  NAND U936 ( .A(n1289), .B(n1290), .Z(n1288) );
  XNOR U937 ( .A(n1289), .B(n1291), .Z(SUM[780]) );
  NANDN U938 ( .A(n1287), .B(n1290), .Z(n1291) );
  NANDN U939 ( .A(n1292), .B(n1293), .Z(n1289) );
  NANDN U940 ( .A(n1294), .B(n1295), .Z(n1293) );
  XNOR U941 ( .A(n1244), .B(n1296), .Z(SUM[77]) );
  NANDN U942 ( .A(n1242), .B(n1245), .Z(n1296) );
  NANDN U943 ( .A(n1297), .B(n1298), .Z(n1244) );
  NANDN U944 ( .A(n1299), .B(n1300), .Z(n1298) );
  XOR U945 ( .A(n1301), .B(n1302), .Z(SUM[779]) );
  NANDN U946 ( .A(n1303), .B(n1304), .Z(n1302) );
  ANDN U947 ( .B(n1305), .A(n1306), .Z(n1301) );
  NAND U948 ( .A(n1307), .B(n1308), .Z(n1305) );
  XNOR U949 ( .A(n1307), .B(n1309), .Z(SUM[778]) );
  NANDN U950 ( .A(n1306), .B(n1308), .Z(n1309) );
  NANDN U951 ( .A(n1310), .B(n1311), .Z(n1307) );
  NAND U952 ( .A(n1312), .B(n1313), .Z(n1311) );
  XNOR U953 ( .A(n1312), .B(n1314), .Z(SUM[777]) );
  NANDN U954 ( .A(n1310), .B(n1313), .Z(n1314) );
  NANDN U955 ( .A(n1315), .B(n1316), .Z(n1312) );
  NAND U956 ( .A(n1295), .B(n1317), .Z(n1316) );
  XNOR U957 ( .A(n1295), .B(n1318), .Z(SUM[776]) );
  NANDN U958 ( .A(n1315), .B(n1317), .Z(n1318) );
  NANDN U959 ( .A(n1319), .B(n1320), .Z(n1295) );
  NANDN U960 ( .A(n1321), .B(n1322), .Z(n1320) );
  XOR U961 ( .A(n1323), .B(n1324), .Z(SUM[775]) );
  NANDN U962 ( .A(n1325), .B(n1326), .Z(n1324) );
  ANDN U963 ( .B(n1327), .A(n1328), .Z(n1323) );
  NAND U964 ( .A(n1329), .B(n1330), .Z(n1327) );
  XNOR U965 ( .A(n1329), .B(n1331), .Z(SUM[774]) );
  NANDN U966 ( .A(n1328), .B(n1330), .Z(n1331) );
  NANDN U967 ( .A(n1332), .B(n1333), .Z(n1329) );
  NAND U968 ( .A(n1334), .B(n1335), .Z(n1333) );
  XNOR U969 ( .A(n1334), .B(n1336), .Z(SUM[773]) );
  NANDN U970 ( .A(n1332), .B(n1335), .Z(n1336) );
  NANDN U971 ( .A(n1337), .B(n1338), .Z(n1334) );
  NANDN U972 ( .A(n1321), .B(n1339), .Z(n1338) );
  XOR U973 ( .A(n1321), .B(n1340), .Z(SUM[772]) );
  NANDN U974 ( .A(n1337), .B(n1339), .Z(n1340) );
  ANDN U975 ( .B(n1341), .A(n1342), .Z(n1321) );
  OR U976 ( .A(n1343), .B(n1344), .Z(n1341) );
  XOR U977 ( .A(n1345), .B(n1346), .Z(SUM[771]) );
  NANDN U978 ( .A(n1347), .B(n1348), .Z(n1346) );
  ANDN U979 ( .B(n1349), .A(n1350), .Z(n1345) );
  NANDN U980 ( .A(n1351), .B(n1352), .Z(n1349) );
  XNOR U981 ( .A(n1352), .B(n1353), .Z(SUM[770]) );
  OR U982 ( .A(n1351), .B(n1350), .Z(n1353) );
  NANDN U983 ( .A(n1354), .B(n1355), .Z(n1352) );
  NAND U984 ( .A(n1356), .B(n1357), .Z(n1355) );
  XNOR U985 ( .A(n1300), .B(n1358), .Z(SUM[76]) );
  OR U986 ( .A(n1299), .B(n1297), .Z(n1358) );
  NANDN U987 ( .A(n1359), .B(n1360), .Z(n1300) );
  NANDN U988 ( .A(n1361), .B(n1362), .Z(n1360) );
  XNOR U989 ( .A(n1356), .B(n1363), .Z(SUM[769]) );
  NANDN U990 ( .A(n1354), .B(n1357), .Z(n1363) );
  NANDN U991 ( .A(n1364), .B(n1365), .Z(n1356) );
  NANDN U992 ( .A(n1344), .B(n1366), .Z(n1365) );
  XOR U993 ( .A(n1344), .B(n1367), .Z(SUM[768]) );
  NANDN U994 ( .A(n1364), .B(n1366), .Z(n1367) );
  XOR U995 ( .A(n1368), .B(n1369), .Z(SUM[767]) );
  OR U996 ( .A(n1370), .B(n1371), .Z(n1369) );
  ANDN U997 ( .B(n1372), .A(n1373), .Z(n1368) );
  NAND U998 ( .A(n1374), .B(n1375), .Z(n1372) );
  XNOR U999 ( .A(n1374), .B(n1376), .Z(SUM[766]) );
  NANDN U1000 ( .A(n1373), .B(n1375), .Z(n1376) );
  NANDN U1001 ( .A(n1377), .B(n1378), .Z(n1374) );
  NAND U1002 ( .A(n1379), .B(n1380), .Z(n1378) );
  XNOR U1003 ( .A(n1379), .B(n1381), .Z(SUM[765]) );
  NANDN U1004 ( .A(n1377), .B(n1380), .Z(n1381) );
  NANDN U1005 ( .A(n1382), .B(n1383), .Z(n1379) );
  NANDN U1006 ( .A(n1384), .B(n1385), .Z(n1383) );
  XNOR U1007 ( .A(n1385), .B(n1386), .Z(SUM[764]) );
  OR U1008 ( .A(n1384), .B(n1382), .Z(n1386) );
  NANDN U1009 ( .A(n1387), .B(n1388), .Z(n1385) );
  NANDN U1010 ( .A(n1389), .B(n1390), .Z(n1388) );
  XOR U1011 ( .A(n1391), .B(n1392), .Z(SUM[763]) );
  NANDN U1012 ( .A(n1393), .B(n1394), .Z(n1392) );
  ANDN U1013 ( .B(n1395), .A(n1396), .Z(n1391) );
  NAND U1014 ( .A(n1397), .B(n1398), .Z(n1395) );
  XNOR U1015 ( .A(n1397), .B(n1399), .Z(SUM[762]) );
  NANDN U1016 ( .A(n1396), .B(n1398), .Z(n1399) );
  NANDN U1017 ( .A(n1400), .B(n1401), .Z(n1397) );
  NAND U1018 ( .A(n1402), .B(n1403), .Z(n1401) );
  XNOR U1019 ( .A(n1402), .B(n1404), .Z(SUM[761]) );
  NANDN U1020 ( .A(n1400), .B(n1403), .Z(n1404) );
  NANDN U1021 ( .A(n1405), .B(n1406), .Z(n1402) );
  NAND U1022 ( .A(n1390), .B(n1407), .Z(n1406) );
  XNOR U1023 ( .A(n1390), .B(n1408), .Z(SUM[760]) );
  NANDN U1024 ( .A(n1405), .B(n1407), .Z(n1408) );
  NANDN U1025 ( .A(n1409), .B(n1410), .Z(n1390) );
  NANDN U1026 ( .A(n1411), .B(n1412), .Z(n1410) );
  XOR U1027 ( .A(n1413), .B(n1414), .Z(SUM[75]) );
  NANDN U1028 ( .A(n1415), .B(n1416), .Z(n1414) );
  ANDN U1029 ( .B(n1417), .A(n1418), .Z(n1413) );
  NAND U1030 ( .A(n1419), .B(n1420), .Z(n1417) );
  XOR U1031 ( .A(n1421), .B(n1422), .Z(SUM[759]) );
  NANDN U1032 ( .A(n1423), .B(n1424), .Z(n1422) );
  ANDN U1033 ( .B(n1425), .A(n1426), .Z(n1421) );
  NAND U1034 ( .A(n1427), .B(n1428), .Z(n1425) );
  XNOR U1035 ( .A(n1427), .B(n1429), .Z(SUM[758]) );
  NANDN U1036 ( .A(n1426), .B(n1428), .Z(n1429) );
  NANDN U1037 ( .A(n1430), .B(n1431), .Z(n1427) );
  NAND U1038 ( .A(n1432), .B(n1433), .Z(n1431) );
  XNOR U1039 ( .A(n1432), .B(n1434), .Z(SUM[757]) );
  NANDN U1040 ( .A(n1430), .B(n1433), .Z(n1434) );
  NANDN U1041 ( .A(n1435), .B(n1436), .Z(n1432) );
  NANDN U1042 ( .A(n1411), .B(n1437), .Z(n1436) );
  XOR U1043 ( .A(n1411), .B(n1438), .Z(SUM[756]) );
  NANDN U1044 ( .A(n1435), .B(n1437), .Z(n1438) );
  ANDN U1045 ( .B(n1439), .A(n1440), .Z(n1411) );
  NANDN U1046 ( .A(n1441), .B(n1442), .Z(n1439) );
  XOR U1047 ( .A(n1443), .B(n1444), .Z(SUM[755]) );
  NANDN U1048 ( .A(n1445), .B(n1446), .Z(n1444) );
  ANDN U1049 ( .B(n1447), .A(n1448), .Z(n1443) );
  NANDN U1050 ( .A(n1449), .B(n1450), .Z(n1447) );
  XNOR U1051 ( .A(n1450), .B(n1451), .Z(SUM[754]) );
  OR U1052 ( .A(n1449), .B(n1448), .Z(n1451) );
  NANDN U1053 ( .A(n1452), .B(n1453), .Z(n1450) );
  NAND U1054 ( .A(n1454), .B(n1455), .Z(n1453) );
  XNOR U1055 ( .A(n1454), .B(n1456), .Z(SUM[753]) );
  NANDN U1056 ( .A(n1452), .B(n1455), .Z(n1456) );
  NANDN U1057 ( .A(n1457), .B(n1458), .Z(n1454) );
  NAND U1058 ( .A(n1442), .B(n1459), .Z(n1458) );
  XNOR U1059 ( .A(n1442), .B(n1460), .Z(SUM[752]) );
  NANDN U1060 ( .A(n1457), .B(n1459), .Z(n1460) );
  NANDN U1061 ( .A(n1461), .B(n1462), .Z(n1442) );
  NANDN U1062 ( .A(n1463), .B(n1464), .Z(n1462) );
  XOR U1063 ( .A(n1465), .B(n1466), .Z(SUM[751]) );
  NANDN U1064 ( .A(n1467), .B(n1468), .Z(n1466) );
  ANDN U1065 ( .B(n1469), .A(n1470), .Z(n1465) );
  NAND U1066 ( .A(n1471), .B(n1472), .Z(n1469) );
  XNOR U1067 ( .A(n1471), .B(n1473), .Z(SUM[750]) );
  NANDN U1068 ( .A(n1470), .B(n1472), .Z(n1473) );
  NANDN U1069 ( .A(n1474), .B(n1475), .Z(n1471) );
  NAND U1070 ( .A(n1476), .B(n1477), .Z(n1475) );
  XNOR U1071 ( .A(n1419), .B(n1478), .Z(SUM[74]) );
  NANDN U1072 ( .A(n1418), .B(n1420), .Z(n1478) );
  NANDN U1073 ( .A(n1479), .B(n1480), .Z(n1419) );
  NAND U1074 ( .A(n1481), .B(n1482), .Z(n1480) );
  XNOR U1075 ( .A(n1476), .B(n1483), .Z(SUM[749]) );
  NANDN U1076 ( .A(n1474), .B(n1477), .Z(n1483) );
  NANDN U1077 ( .A(n1484), .B(n1485), .Z(n1476) );
  NAND U1078 ( .A(n1486), .B(n1487), .Z(n1485) );
  XNOR U1079 ( .A(n1486), .B(n1488), .Z(SUM[748]) );
  NANDN U1080 ( .A(n1484), .B(n1487), .Z(n1488) );
  NANDN U1081 ( .A(n1489), .B(n1490), .Z(n1486) );
  NAND U1082 ( .A(n1491), .B(n1492), .Z(n1490) );
  XOR U1083 ( .A(n1493), .B(n1494), .Z(SUM[747]) );
  NANDN U1084 ( .A(n1495), .B(n1496), .Z(n1494) );
  ANDN U1085 ( .B(n1497), .A(n1498), .Z(n1493) );
  NAND U1086 ( .A(n1499), .B(n1500), .Z(n1497) );
  XNOR U1087 ( .A(n1499), .B(n1501), .Z(SUM[746]) );
  NANDN U1088 ( .A(n1498), .B(n1500), .Z(n1501) );
  NANDN U1089 ( .A(n1502), .B(n1503), .Z(n1499) );
  NAND U1090 ( .A(n1504), .B(n1505), .Z(n1503) );
  XNOR U1091 ( .A(n1504), .B(n1506), .Z(SUM[745]) );
  NANDN U1092 ( .A(n1502), .B(n1505), .Z(n1506) );
  NANDN U1093 ( .A(n1507), .B(n1508), .Z(n1504) );
  NAND U1094 ( .A(n1492), .B(n1509), .Z(n1508) );
  XNOR U1095 ( .A(n1492), .B(n1510), .Z(SUM[744]) );
  NANDN U1096 ( .A(n1507), .B(n1509), .Z(n1510) );
  NANDN U1097 ( .A(n1511), .B(n1512), .Z(n1492) );
  OR U1098 ( .A(n1513), .B(n1514), .Z(n1512) );
  XOR U1099 ( .A(n1515), .B(n1516), .Z(SUM[743]) );
  NANDN U1100 ( .A(n1517), .B(n1518), .Z(n1516) );
  ANDN U1101 ( .B(n1519), .A(n1520), .Z(n1515) );
  NAND U1102 ( .A(n1521), .B(n1522), .Z(n1519) );
  XNOR U1103 ( .A(n1521), .B(n1523), .Z(SUM[742]) );
  NANDN U1104 ( .A(n1520), .B(n1522), .Z(n1523) );
  NANDN U1105 ( .A(n1524), .B(n1525), .Z(n1521) );
  NAND U1106 ( .A(n1526), .B(n1527), .Z(n1525) );
  XNOR U1107 ( .A(n1526), .B(n1528), .Z(SUM[741]) );
  NANDN U1108 ( .A(n1524), .B(n1527), .Z(n1528) );
  NANDN U1109 ( .A(n1529), .B(n1530), .Z(n1526) );
  NANDN U1110 ( .A(n1514), .B(n1531), .Z(n1530) );
  XOR U1111 ( .A(n1514), .B(n1532), .Z(SUM[740]) );
  NANDN U1112 ( .A(n1529), .B(n1531), .Z(n1532) );
  ANDN U1113 ( .B(n1533), .A(n1534), .Z(n1514) );
  NANDN U1114 ( .A(n1535), .B(n1464), .Z(n1533) );
  XNOR U1115 ( .A(n1481), .B(n1536), .Z(SUM[73]) );
  NANDN U1116 ( .A(n1479), .B(n1482), .Z(n1536) );
  NANDN U1117 ( .A(n1537), .B(n1538), .Z(n1481) );
  NAND U1118 ( .A(n1362), .B(n1539), .Z(n1538) );
  XOR U1119 ( .A(n1540), .B(n1541), .Z(SUM[739]) );
  NANDN U1120 ( .A(n1542), .B(n1543), .Z(n1541) );
  ANDN U1121 ( .B(n1544), .A(n1545), .Z(n1540) );
  NAND U1122 ( .A(n1546), .B(n1547), .Z(n1544) );
  XNOR U1123 ( .A(n1546), .B(n1548), .Z(SUM[738]) );
  NANDN U1124 ( .A(n1545), .B(n1547), .Z(n1548) );
  NANDN U1125 ( .A(n1549), .B(n1550), .Z(n1546) );
  NAND U1126 ( .A(n1551), .B(n1552), .Z(n1550) );
  XNOR U1127 ( .A(n1551), .B(n1553), .Z(SUM[737]) );
  NANDN U1128 ( .A(n1549), .B(n1552), .Z(n1553) );
  NANDN U1129 ( .A(n1554), .B(n1555), .Z(n1551) );
  NAND U1130 ( .A(n1464), .B(n1556), .Z(n1555) );
  XNOR U1131 ( .A(n1464), .B(n1557), .Z(SUM[736]) );
  NANDN U1132 ( .A(n1554), .B(n1556), .Z(n1557) );
  NANDN U1133 ( .A(n1558), .B(n1559), .Z(n1464) );
  NANDN U1134 ( .A(n1560), .B(n1561), .Z(n1559) );
  XOR U1135 ( .A(n1562), .B(n1563), .Z(SUM[735]) );
  NANDN U1136 ( .A(n1564), .B(n1565), .Z(n1563) );
  ANDN U1137 ( .B(n1566), .A(n1567), .Z(n1562) );
  NAND U1138 ( .A(n1568), .B(n1569), .Z(n1566) );
  XNOR U1139 ( .A(n1568), .B(n1570), .Z(SUM[734]) );
  NANDN U1140 ( .A(n1567), .B(n1569), .Z(n1570) );
  NANDN U1141 ( .A(n1571), .B(n1572), .Z(n1568) );
  NAND U1142 ( .A(n1573), .B(n1574), .Z(n1572) );
  XNOR U1143 ( .A(n1573), .B(n1575), .Z(SUM[733]) );
  NANDN U1144 ( .A(n1571), .B(n1574), .Z(n1575) );
  NANDN U1145 ( .A(n1576), .B(n1577), .Z(n1573) );
  NAND U1146 ( .A(n1578), .B(n1579), .Z(n1577) );
  XNOR U1147 ( .A(n1578), .B(n1580), .Z(SUM[732]) );
  NANDN U1148 ( .A(n1576), .B(n1579), .Z(n1580) );
  NANDN U1149 ( .A(n1581), .B(n1582), .Z(n1578) );
  NAND U1150 ( .A(n1583), .B(n1584), .Z(n1582) );
  XOR U1151 ( .A(n1585), .B(n1586), .Z(SUM[731]) );
  NANDN U1152 ( .A(n1587), .B(n1588), .Z(n1586) );
  ANDN U1153 ( .B(n1589), .A(n1590), .Z(n1585) );
  NAND U1154 ( .A(n1591), .B(n1592), .Z(n1589) );
  XNOR U1155 ( .A(n1591), .B(n1593), .Z(SUM[730]) );
  NANDN U1156 ( .A(n1590), .B(n1592), .Z(n1593) );
  NANDN U1157 ( .A(n1594), .B(n1595), .Z(n1591) );
  NAND U1158 ( .A(n1596), .B(n1597), .Z(n1595) );
  XNOR U1159 ( .A(n1362), .B(n1598), .Z(SUM[72]) );
  NANDN U1160 ( .A(n1537), .B(n1539), .Z(n1598) );
  NANDN U1161 ( .A(n1599), .B(n1600), .Z(n1362) );
  NANDN U1162 ( .A(n1601), .B(n1602), .Z(n1600) );
  XNOR U1163 ( .A(n1596), .B(n1603), .Z(SUM[729]) );
  NANDN U1164 ( .A(n1594), .B(n1597), .Z(n1603) );
  NANDN U1165 ( .A(n1604), .B(n1605), .Z(n1596) );
  NAND U1166 ( .A(n1584), .B(n1606), .Z(n1605) );
  XNOR U1167 ( .A(n1584), .B(n1607), .Z(SUM[728]) );
  NANDN U1168 ( .A(n1604), .B(n1606), .Z(n1607) );
  NANDN U1169 ( .A(n1608), .B(n1609), .Z(n1584) );
  OR U1170 ( .A(n1610), .B(n1611), .Z(n1609) );
  XOR U1171 ( .A(n1612), .B(n1613), .Z(SUM[727]) );
  NANDN U1172 ( .A(n1614), .B(n1615), .Z(n1613) );
  ANDN U1173 ( .B(n1616), .A(n1617), .Z(n1612) );
  NAND U1174 ( .A(n1618), .B(n1619), .Z(n1616) );
  XNOR U1175 ( .A(n1618), .B(n1620), .Z(SUM[726]) );
  NANDN U1176 ( .A(n1617), .B(n1619), .Z(n1620) );
  NANDN U1177 ( .A(n1621), .B(n1622), .Z(n1618) );
  NAND U1178 ( .A(n1623), .B(n1624), .Z(n1622) );
  XNOR U1179 ( .A(n1623), .B(n1625), .Z(SUM[725]) );
  NANDN U1180 ( .A(n1621), .B(n1624), .Z(n1625) );
  NANDN U1181 ( .A(n1626), .B(n1627), .Z(n1623) );
  NANDN U1182 ( .A(n1611), .B(n1628), .Z(n1627) );
  XOR U1183 ( .A(n1611), .B(n1629), .Z(SUM[724]) );
  NANDN U1184 ( .A(n1626), .B(n1628), .Z(n1629) );
  ANDN U1185 ( .B(n1630), .A(n1631), .Z(n1611) );
  NANDN U1186 ( .A(n1632), .B(n1561), .Z(n1630) );
  XOR U1187 ( .A(n1633), .B(n1634), .Z(SUM[723]) );
  NANDN U1188 ( .A(n1635), .B(n1636), .Z(n1634) );
  ANDN U1189 ( .B(n1637), .A(n1638), .Z(n1633) );
  NAND U1190 ( .A(n1639), .B(n1640), .Z(n1637) );
  XNOR U1191 ( .A(n1639), .B(n1641), .Z(SUM[722]) );
  NANDN U1192 ( .A(n1638), .B(n1640), .Z(n1641) );
  NANDN U1193 ( .A(n1642), .B(n1643), .Z(n1639) );
  NAND U1194 ( .A(n1644), .B(n1645), .Z(n1643) );
  XNOR U1195 ( .A(n1644), .B(n1646), .Z(SUM[721]) );
  NANDN U1196 ( .A(n1642), .B(n1645), .Z(n1646) );
  NANDN U1197 ( .A(n1647), .B(n1648), .Z(n1644) );
  NAND U1198 ( .A(n1561), .B(n1649), .Z(n1648) );
  XNOR U1199 ( .A(n1561), .B(n1650), .Z(SUM[720]) );
  NANDN U1200 ( .A(n1647), .B(n1649), .Z(n1650) );
  NANDN U1201 ( .A(n1651), .B(n1652), .Z(n1561) );
  NANDN U1202 ( .A(n1653), .B(n1654), .Z(n1652) );
  XOR U1203 ( .A(n1655), .B(n1656), .Z(SUM[71]) );
  NANDN U1204 ( .A(n1657), .B(n1658), .Z(n1656) );
  ANDN U1205 ( .B(n1659), .A(n1660), .Z(n1655) );
  NAND U1206 ( .A(n1661), .B(n1662), .Z(n1659) );
  XOR U1207 ( .A(n1663), .B(n1664), .Z(SUM[719]) );
  NANDN U1208 ( .A(n1665), .B(n1666), .Z(n1664) );
  ANDN U1209 ( .B(n1667), .A(n1668), .Z(n1663) );
  NAND U1210 ( .A(n1669), .B(n1670), .Z(n1667) );
  XNOR U1211 ( .A(n1669), .B(n1671), .Z(SUM[718]) );
  NANDN U1212 ( .A(n1668), .B(n1670), .Z(n1671) );
  NANDN U1213 ( .A(n1672), .B(n1673), .Z(n1669) );
  NAND U1214 ( .A(n1674), .B(n1675), .Z(n1673) );
  XNOR U1215 ( .A(n1674), .B(n1676), .Z(SUM[717]) );
  NANDN U1216 ( .A(n1672), .B(n1675), .Z(n1676) );
  NANDN U1217 ( .A(n1677), .B(n1678), .Z(n1674) );
  NAND U1218 ( .A(n1679), .B(n1680), .Z(n1678) );
  XNOR U1219 ( .A(n1679), .B(n1681), .Z(SUM[716]) );
  NANDN U1220 ( .A(n1677), .B(n1680), .Z(n1681) );
  NANDN U1221 ( .A(n1682), .B(n1683), .Z(n1679) );
  NAND U1222 ( .A(n1684), .B(n1685), .Z(n1683) );
  XOR U1223 ( .A(n1686), .B(n1687), .Z(SUM[715]) );
  NANDN U1224 ( .A(n1688), .B(n1689), .Z(n1687) );
  ANDN U1225 ( .B(n1690), .A(n1691), .Z(n1686) );
  NAND U1226 ( .A(n1692), .B(n1693), .Z(n1690) );
  XNOR U1227 ( .A(n1692), .B(n1694), .Z(SUM[714]) );
  NANDN U1228 ( .A(n1691), .B(n1693), .Z(n1694) );
  NANDN U1229 ( .A(n1695), .B(n1696), .Z(n1692) );
  NAND U1230 ( .A(n1697), .B(n1698), .Z(n1696) );
  XNOR U1231 ( .A(n1697), .B(n1699), .Z(SUM[713]) );
  NANDN U1232 ( .A(n1695), .B(n1698), .Z(n1699) );
  NANDN U1233 ( .A(n1700), .B(n1701), .Z(n1697) );
  NAND U1234 ( .A(n1685), .B(n1702), .Z(n1701) );
  XNOR U1235 ( .A(n1685), .B(n1703), .Z(SUM[712]) );
  NANDN U1236 ( .A(n1700), .B(n1702), .Z(n1703) );
  NANDN U1237 ( .A(n1704), .B(n1705), .Z(n1685) );
  OR U1238 ( .A(n1706), .B(n1707), .Z(n1705) );
  XOR U1239 ( .A(n1708), .B(n1709), .Z(SUM[711]) );
  NANDN U1240 ( .A(n1710), .B(n1711), .Z(n1709) );
  ANDN U1241 ( .B(n1712), .A(n1713), .Z(n1708) );
  NAND U1242 ( .A(n1714), .B(n1715), .Z(n1712) );
  XNOR U1243 ( .A(n1714), .B(n1716), .Z(SUM[710]) );
  NANDN U1244 ( .A(n1713), .B(n1715), .Z(n1716) );
  NANDN U1245 ( .A(n1717), .B(n1718), .Z(n1714) );
  NAND U1246 ( .A(n1719), .B(n1720), .Z(n1718) );
  XNOR U1247 ( .A(n1661), .B(n1721), .Z(SUM[70]) );
  NANDN U1248 ( .A(n1660), .B(n1662), .Z(n1721) );
  NANDN U1249 ( .A(n1722), .B(n1723), .Z(n1661) );
  NAND U1250 ( .A(n1724), .B(n1725), .Z(n1723) );
  XNOR U1251 ( .A(n1719), .B(n1726), .Z(SUM[709]) );
  NANDN U1252 ( .A(n1717), .B(n1720), .Z(n1726) );
  NANDN U1253 ( .A(n1727), .B(n1728), .Z(n1719) );
  NANDN U1254 ( .A(n1707), .B(n1729), .Z(n1728) );
  XOR U1255 ( .A(n1707), .B(n1730), .Z(SUM[708]) );
  NANDN U1256 ( .A(n1727), .B(n1729), .Z(n1730) );
  ANDN U1257 ( .B(n1731), .A(n1732), .Z(n1707) );
  NANDN U1258 ( .A(n1733), .B(n1654), .Z(n1731) );
  XOR U1259 ( .A(n1734), .B(n1735), .Z(SUM[707]) );
  NANDN U1260 ( .A(n1736), .B(n1737), .Z(n1735) );
  ANDN U1261 ( .B(n1738), .A(n1739), .Z(n1734) );
  NAND U1262 ( .A(n1740), .B(n1741), .Z(n1738) );
  XNOR U1263 ( .A(n1740), .B(n1742), .Z(SUM[706]) );
  NANDN U1264 ( .A(n1739), .B(n1741), .Z(n1742) );
  NANDN U1265 ( .A(n1743), .B(n1744), .Z(n1740) );
  NAND U1266 ( .A(n1745), .B(n1746), .Z(n1744) );
  XNOR U1267 ( .A(n1745), .B(n1747), .Z(SUM[705]) );
  NANDN U1268 ( .A(n1743), .B(n1746), .Z(n1747) );
  NANDN U1269 ( .A(n1748), .B(n1749), .Z(n1745) );
  NAND U1270 ( .A(n1654), .B(n1750), .Z(n1749) );
  XNOR U1271 ( .A(n1654), .B(n1751), .Z(SUM[704]) );
  NANDN U1272 ( .A(n1748), .B(n1750), .Z(n1751) );
  NANDN U1273 ( .A(n1752), .B(n1753), .Z(n1654) );
  NANDN U1274 ( .A(n1754), .B(n1755), .Z(n1753) );
  XOR U1275 ( .A(n1756), .B(n1757), .Z(SUM[703]) );
  NANDN U1276 ( .A(n1758), .B(n1759), .Z(n1757) );
  ANDN U1277 ( .B(n1760), .A(n1761), .Z(n1756) );
  NAND U1278 ( .A(n1762), .B(n1763), .Z(n1760) );
  XNOR U1279 ( .A(n1762), .B(n1764), .Z(SUM[702]) );
  NANDN U1280 ( .A(n1761), .B(n1763), .Z(n1764) );
  NANDN U1281 ( .A(n1765), .B(n1766), .Z(n1762) );
  NAND U1282 ( .A(n1767), .B(n1768), .Z(n1766) );
  XNOR U1283 ( .A(n1767), .B(n1769), .Z(SUM[701]) );
  NANDN U1284 ( .A(n1765), .B(n1768), .Z(n1769) );
  NANDN U1285 ( .A(n1770), .B(n1771), .Z(n1767) );
  NAND U1286 ( .A(n1772), .B(n1773), .Z(n1771) );
  XNOR U1287 ( .A(n1772), .B(n1774), .Z(SUM[700]) );
  NANDN U1288 ( .A(n1770), .B(n1773), .Z(n1774) );
  NANDN U1289 ( .A(n1775), .B(n1776), .Z(n1772) );
  NANDN U1290 ( .A(n1777), .B(n1778), .Z(n1776) );
  XNOR U1291 ( .A(n1779), .B(n1780), .Z(SUM[6]) );
  OR U1292 ( .A(n1781), .B(n1174), .Z(n1780) );
  XNOR U1293 ( .A(n1724), .B(n1782), .Z(SUM[69]) );
  NANDN U1294 ( .A(n1722), .B(n1725), .Z(n1782) );
  NANDN U1295 ( .A(n1783), .B(n1784), .Z(n1724) );
  NANDN U1296 ( .A(n1601), .B(n1785), .Z(n1784) );
  XOR U1297 ( .A(n1786), .B(n1787), .Z(SUM[699]) );
  NANDN U1298 ( .A(n1788), .B(n1789), .Z(n1787) );
  ANDN U1299 ( .B(n1790), .A(n1791), .Z(n1786) );
  NAND U1300 ( .A(n1792), .B(n1793), .Z(n1790) );
  XNOR U1301 ( .A(n1792), .B(n1794), .Z(SUM[698]) );
  NANDN U1302 ( .A(n1791), .B(n1793), .Z(n1794) );
  NANDN U1303 ( .A(n1795), .B(n1796), .Z(n1792) );
  NAND U1304 ( .A(n1797), .B(n1798), .Z(n1796) );
  XNOR U1305 ( .A(n1797), .B(n1799), .Z(SUM[697]) );
  NANDN U1306 ( .A(n1795), .B(n1798), .Z(n1799) );
  NANDN U1307 ( .A(n1800), .B(n1801), .Z(n1797) );
  NAND U1308 ( .A(n1778), .B(n1802), .Z(n1801) );
  XNOR U1309 ( .A(n1778), .B(n1803), .Z(SUM[696]) );
  NANDN U1310 ( .A(n1800), .B(n1802), .Z(n1803) );
  NANDN U1311 ( .A(n1804), .B(n1805), .Z(n1778) );
  OR U1312 ( .A(n1806), .B(n1807), .Z(n1805) );
  XOR U1313 ( .A(n1808), .B(n1809), .Z(SUM[695]) );
  NANDN U1314 ( .A(n1810), .B(n1811), .Z(n1809) );
  ANDN U1315 ( .B(n1812), .A(n1813), .Z(n1808) );
  NAND U1316 ( .A(n1814), .B(n1815), .Z(n1812) );
  XNOR U1317 ( .A(n1814), .B(n1816), .Z(SUM[694]) );
  NANDN U1318 ( .A(n1813), .B(n1815), .Z(n1816) );
  NANDN U1319 ( .A(n1817), .B(n1818), .Z(n1814) );
  NAND U1320 ( .A(n1819), .B(n1820), .Z(n1818) );
  XNOR U1321 ( .A(n1819), .B(n1821), .Z(SUM[693]) );
  NANDN U1322 ( .A(n1817), .B(n1820), .Z(n1821) );
  NANDN U1323 ( .A(n1822), .B(n1823), .Z(n1819) );
  NANDN U1324 ( .A(n1807), .B(n1824), .Z(n1823) );
  XOR U1325 ( .A(n1807), .B(n1825), .Z(SUM[692]) );
  NANDN U1326 ( .A(n1822), .B(n1824), .Z(n1825) );
  ANDN U1327 ( .B(n1826), .A(n1827), .Z(n1807) );
  NANDN U1328 ( .A(n1828), .B(n1829), .Z(n1826) );
  XOR U1329 ( .A(n1830), .B(n1831), .Z(SUM[691]) );
  NANDN U1330 ( .A(n1832), .B(n1833), .Z(n1831) );
  ANDN U1331 ( .B(n1834), .A(n1835), .Z(n1830) );
  NAND U1332 ( .A(n1836), .B(n1837), .Z(n1834) );
  XNOR U1333 ( .A(n1836), .B(n1838), .Z(SUM[690]) );
  NANDN U1334 ( .A(n1835), .B(n1837), .Z(n1838) );
  NANDN U1335 ( .A(n1839), .B(n1840), .Z(n1836) );
  NAND U1336 ( .A(n1841), .B(n1842), .Z(n1840) );
  XOR U1337 ( .A(n1601), .B(n1843), .Z(SUM[68]) );
  NANDN U1338 ( .A(n1783), .B(n1785), .Z(n1843) );
  ANDN U1339 ( .B(n1844), .A(n1845), .Z(n1601) );
  OR U1340 ( .A(n1846), .B(n1847), .Z(n1844) );
  XNOR U1341 ( .A(n1841), .B(n1848), .Z(SUM[689]) );
  NANDN U1342 ( .A(n1839), .B(n1842), .Z(n1848) );
  NANDN U1343 ( .A(n1849), .B(n1850), .Z(n1841) );
  NAND U1344 ( .A(n1829), .B(n1851), .Z(n1850) );
  XNOR U1345 ( .A(n1829), .B(n1852), .Z(SUM[688]) );
  NANDN U1346 ( .A(n1849), .B(n1851), .Z(n1852) );
  NANDN U1347 ( .A(n1853), .B(n1854), .Z(n1829) );
  NAND U1348 ( .A(n1855), .B(n1856), .Z(n1854) );
  XOR U1349 ( .A(n1857), .B(n1858), .Z(SUM[687]) );
  NANDN U1350 ( .A(n1859), .B(n1860), .Z(n1858) );
  ANDN U1351 ( .B(n1861), .A(n1862), .Z(n1857) );
  NAND U1352 ( .A(n1863), .B(n1864), .Z(n1861) );
  XNOR U1353 ( .A(n1863), .B(n1865), .Z(SUM[686]) );
  NANDN U1354 ( .A(n1862), .B(n1864), .Z(n1865) );
  NANDN U1355 ( .A(n1866), .B(n1867), .Z(n1863) );
  NAND U1356 ( .A(n1868), .B(n1869), .Z(n1867) );
  XNOR U1357 ( .A(n1868), .B(n1870), .Z(SUM[685]) );
  NANDN U1358 ( .A(n1866), .B(n1869), .Z(n1870) );
  NANDN U1359 ( .A(n1871), .B(n1872), .Z(n1868) );
  NAND U1360 ( .A(n1873), .B(n1874), .Z(n1872) );
  XNOR U1361 ( .A(n1873), .B(n1875), .Z(SUM[684]) );
  NANDN U1362 ( .A(n1871), .B(n1874), .Z(n1875) );
  NANDN U1363 ( .A(n1876), .B(n1877), .Z(n1873) );
  NAND U1364 ( .A(n1878), .B(n1879), .Z(n1877) );
  XOR U1365 ( .A(n1880), .B(n1881), .Z(SUM[683]) );
  NANDN U1366 ( .A(n1882), .B(n1883), .Z(n1881) );
  ANDN U1367 ( .B(n1884), .A(n1885), .Z(n1880) );
  NAND U1368 ( .A(n1886), .B(n1887), .Z(n1884) );
  XNOR U1369 ( .A(n1886), .B(n1888), .Z(SUM[682]) );
  NANDN U1370 ( .A(n1885), .B(n1887), .Z(n1888) );
  NANDN U1371 ( .A(n1889), .B(n1890), .Z(n1886) );
  NAND U1372 ( .A(n1891), .B(n1892), .Z(n1890) );
  XNOR U1373 ( .A(n1891), .B(n1893), .Z(SUM[681]) );
  NANDN U1374 ( .A(n1889), .B(n1892), .Z(n1893) );
  NANDN U1375 ( .A(n1894), .B(n1895), .Z(n1891) );
  NAND U1376 ( .A(n1879), .B(n1896), .Z(n1895) );
  XNOR U1377 ( .A(n1879), .B(n1897), .Z(SUM[680]) );
  NANDN U1378 ( .A(n1894), .B(n1896), .Z(n1897) );
  NANDN U1379 ( .A(n1898), .B(n1899), .Z(n1879) );
  OR U1380 ( .A(n1900), .B(n1901), .Z(n1899) );
  XOR U1381 ( .A(n1902), .B(n1903), .Z(SUM[67]) );
  NANDN U1382 ( .A(n1904), .B(n1905), .Z(n1903) );
  ANDN U1383 ( .B(n1906), .A(n1907), .Z(n1902) );
  NANDN U1384 ( .A(n1908), .B(n1909), .Z(n1906) );
  XOR U1385 ( .A(n1910), .B(n1911), .Z(SUM[679]) );
  NANDN U1386 ( .A(n1912), .B(n1913), .Z(n1911) );
  ANDN U1387 ( .B(n1914), .A(n1915), .Z(n1910) );
  NAND U1388 ( .A(n1916), .B(n1917), .Z(n1914) );
  XNOR U1389 ( .A(n1916), .B(n1918), .Z(SUM[678]) );
  NANDN U1390 ( .A(n1915), .B(n1917), .Z(n1918) );
  NANDN U1391 ( .A(n1919), .B(n1920), .Z(n1916) );
  NAND U1392 ( .A(n1921), .B(n1922), .Z(n1920) );
  XNOR U1393 ( .A(n1921), .B(n1923), .Z(SUM[677]) );
  NANDN U1394 ( .A(n1919), .B(n1922), .Z(n1923) );
  NANDN U1395 ( .A(n1924), .B(n1925), .Z(n1921) );
  NANDN U1396 ( .A(n1901), .B(n1926), .Z(n1925) );
  XOR U1397 ( .A(n1901), .B(n1927), .Z(SUM[676]) );
  NANDN U1398 ( .A(n1924), .B(n1926), .Z(n1927) );
  ANDN U1399 ( .B(n1928), .A(n1929), .Z(n1901) );
  NANDN U1400 ( .A(n1930), .B(n1856), .Z(n1928) );
  XOR U1401 ( .A(n1931), .B(n1932), .Z(SUM[675]) );
  NANDN U1402 ( .A(n1933), .B(n1934), .Z(n1932) );
  ANDN U1403 ( .B(n1935), .A(n1936), .Z(n1931) );
  NAND U1404 ( .A(n1937), .B(n1938), .Z(n1935) );
  XNOR U1405 ( .A(n1937), .B(n1939), .Z(SUM[674]) );
  NANDN U1406 ( .A(n1936), .B(n1938), .Z(n1939) );
  NANDN U1407 ( .A(n1940), .B(n1941), .Z(n1937) );
  NAND U1408 ( .A(n1942), .B(n1943), .Z(n1941) );
  XNOR U1409 ( .A(n1942), .B(n1944), .Z(SUM[673]) );
  NANDN U1410 ( .A(n1940), .B(n1943), .Z(n1944) );
  NANDN U1411 ( .A(n1945), .B(n1946), .Z(n1942) );
  NAND U1412 ( .A(n1856), .B(n1947), .Z(n1946) );
  XNOR U1413 ( .A(n1856), .B(n1948), .Z(SUM[672]) );
  NANDN U1414 ( .A(n1945), .B(n1947), .Z(n1948) );
  NANDN U1415 ( .A(n1949), .B(n1950), .Z(n1856) );
  OR U1416 ( .A(n1951), .B(n1952), .Z(n1950) );
  XOR U1417 ( .A(n1953), .B(n1954), .Z(SUM[671]) );
  NANDN U1418 ( .A(n1955), .B(n1956), .Z(n1954) );
  ANDN U1419 ( .B(n1957), .A(n1958), .Z(n1953) );
  NAND U1420 ( .A(n1959), .B(n1960), .Z(n1957) );
  XNOR U1421 ( .A(n1959), .B(n1961), .Z(SUM[670]) );
  NANDN U1422 ( .A(n1958), .B(n1960), .Z(n1961) );
  NANDN U1423 ( .A(n1962), .B(n1963), .Z(n1959) );
  NAND U1424 ( .A(n1964), .B(n1965), .Z(n1963) );
  XNOR U1425 ( .A(n1909), .B(n1966), .Z(SUM[66]) );
  OR U1426 ( .A(n1908), .B(n1907), .Z(n1966) );
  NANDN U1427 ( .A(n1967), .B(n1968), .Z(n1909) );
  NAND U1428 ( .A(n1969), .B(n1970), .Z(n1968) );
  XNOR U1429 ( .A(n1964), .B(n1971), .Z(SUM[669]) );
  NANDN U1430 ( .A(n1962), .B(n1965), .Z(n1971) );
  NANDN U1431 ( .A(n1972), .B(n1973), .Z(n1964) );
  NAND U1432 ( .A(n1974), .B(n1975), .Z(n1973) );
  XNOR U1433 ( .A(n1974), .B(n1976), .Z(SUM[668]) );
  NANDN U1434 ( .A(n1972), .B(n1975), .Z(n1976) );
  NANDN U1435 ( .A(n1977), .B(n1978), .Z(n1974) );
  NAND U1436 ( .A(n1979), .B(n1980), .Z(n1978) );
  XOR U1437 ( .A(n1981), .B(n1982), .Z(SUM[667]) );
  NANDN U1438 ( .A(n1983), .B(n1984), .Z(n1982) );
  ANDN U1439 ( .B(n1985), .A(n1986), .Z(n1981) );
  NAND U1440 ( .A(n1987), .B(n1988), .Z(n1985) );
  XNOR U1441 ( .A(n1987), .B(n1989), .Z(SUM[666]) );
  NANDN U1442 ( .A(n1986), .B(n1988), .Z(n1989) );
  NANDN U1443 ( .A(n1990), .B(n1991), .Z(n1987) );
  NAND U1444 ( .A(n1992), .B(n1993), .Z(n1991) );
  XNOR U1445 ( .A(n1992), .B(n1994), .Z(SUM[665]) );
  NANDN U1446 ( .A(n1990), .B(n1993), .Z(n1994) );
  NANDN U1447 ( .A(n1995), .B(n1996), .Z(n1992) );
  NAND U1448 ( .A(n1980), .B(n1997), .Z(n1996) );
  XNOR U1449 ( .A(n1980), .B(n1998), .Z(SUM[664]) );
  NANDN U1450 ( .A(n1995), .B(n1997), .Z(n1998) );
  NANDN U1451 ( .A(n1999), .B(n2000), .Z(n1980) );
  OR U1452 ( .A(n2001), .B(n2002), .Z(n2000) );
  XOR U1453 ( .A(n2003), .B(n2004), .Z(SUM[663]) );
  NANDN U1454 ( .A(n2005), .B(n2006), .Z(n2004) );
  ANDN U1455 ( .B(n2007), .A(n2008), .Z(n2003) );
  NAND U1456 ( .A(n2009), .B(n2010), .Z(n2007) );
  XNOR U1457 ( .A(n2009), .B(n2011), .Z(SUM[662]) );
  NANDN U1458 ( .A(n2008), .B(n2010), .Z(n2011) );
  NANDN U1459 ( .A(n2012), .B(n2013), .Z(n2009) );
  NAND U1460 ( .A(n2014), .B(n2015), .Z(n2013) );
  XNOR U1461 ( .A(n2014), .B(n2016), .Z(SUM[661]) );
  NANDN U1462 ( .A(n2012), .B(n2015), .Z(n2016) );
  NANDN U1463 ( .A(n2017), .B(n2018), .Z(n2014) );
  NANDN U1464 ( .A(n2002), .B(n2019), .Z(n2018) );
  XOR U1465 ( .A(n2002), .B(n2020), .Z(SUM[660]) );
  NANDN U1466 ( .A(n2017), .B(n2019), .Z(n2020) );
  ANDN U1467 ( .B(n2021), .A(n2022), .Z(n2002) );
  OR U1468 ( .A(n2023), .B(n1952), .Z(n2021) );
  XNOR U1469 ( .A(n1969), .B(n2024), .Z(SUM[65]) );
  NANDN U1470 ( .A(n1967), .B(n1970), .Z(n2024) );
  NANDN U1471 ( .A(n2025), .B(n2026), .Z(n1969) );
  NANDN U1472 ( .A(n1847), .B(n2027), .Z(n2026) );
  XOR U1473 ( .A(n2028), .B(n2029), .Z(SUM[659]) );
  NANDN U1474 ( .A(n2030), .B(n2031), .Z(n2029) );
  ANDN U1475 ( .B(n2032), .A(n2033), .Z(n2028) );
  NAND U1476 ( .A(n2034), .B(n2035), .Z(n2032) );
  XNOR U1477 ( .A(n2034), .B(n2036), .Z(SUM[658]) );
  NANDN U1478 ( .A(n2033), .B(n2035), .Z(n2036) );
  NANDN U1479 ( .A(n2037), .B(n2038), .Z(n2034) );
  NAND U1480 ( .A(n2039), .B(n2040), .Z(n2038) );
  XNOR U1481 ( .A(n2039), .B(n2041), .Z(SUM[657]) );
  NANDN U1482 ( .A(n2037), .B(n2040), .Z(n2041) );
  NANDN U1483 ( .A(n2042), .B(n2043), .Z(n2039) );
  NANDN U1484 ( .A(n1952), .B(n2044), .Z(n2043) );
  XOR U1485 ( .A(n1952), .B(n2045), .Z(SUM[656]) );
  NANDN U1486 ( .A(n2042), .B(n2044), .Z(n2045) );
  ANDN U1487 ( .B(n2046), .A(n2047), .Z(n1952) );
  NANDN U1488 ( .A(n2048), .B(n1755), .Z(n2046) );
  XOR U1489 ( .A(n2049), .B(n2050), .Z(SUM[655]) );
  NANDN U1490 ( .A(n2051), .B(n2052), .Z(n2050) );
  ANDN U1491 ( .B(n2053), .A(n2054), .Z(n2049) );
  NAND U1492 ( .A(n2055), .B(n2056), .Z(n2053) );
  XNOR U1493 ( .A(n2055), .B(n2057), .Z(SUM[654]) );
  NANDN U1494 ( .A(n2054), .B(n2056), .Z(n2057) );
  NANDN U1495 ( .A(n2058), .B(n2059), .Z(n2055) );
  NAND U1496 ( .A(n2060), .B(n2061), .Z(n2059) );
  XNOR U1497 ( .A(n2060), .B(n2062), .Z(SUM[653]) );
  NANDN U1498 ( .A(n2058), .B(n2061), .Z(n2062) );
  NANDN U1499 ( .A(n2063), .B(n2064), .Z(n2060) );
  NAND U1500 ( .A(n2065), .B(n2066), .Z(n2064) );
  XNOR U1501 ( .A(n2065), .B(n2067), .Z(SUM[652]) );
  NANDN U1502 ( .A(n2063), .B(n2066), .Z(n2067) );
  NANDN U1503 ( .A(n2068), .B(n2069), .Z(n2065) );
  NAND U1504 ( .A(n2070), .B(n2071), .Z(n2069) );
  XOR U1505 ( .A(n2072), .B(n2073), .Z(SUM[651]) );
  NANDN U1506 ( .A(n2074), .B(n2075), .Z(n2073) );
  ANDN U1507 ( .B(n2076), .A(n2077), .Z(n2072) );
  NAND U1508 ( .A(n2078), .B(n2079), .Z(n2076) );
  XNOR U1509 ( .A(n2078), .B(n2080), .Z(SUM[650]) );
  NANDN U1510 ( .A(n2077), .B(n2079), .Z(n2080) );
  NANDN U1511 ( .A(n2081), .B(n2082), .Z(n2078) );
  NAND U1512 ( .A(n2083), .B(n2084), .Z(n2082) );
  XOR U1513 ( .A(n1847), .B(n2085), .Z(SUM[64]) );
  NANDN U1514 ( .A(n2025), .B(n2027), .Z(n2085) );
  XNOR U1515 ( .A(n2083), .B(n2086), .Z(SUM[649]) );
  NANDN U1516 ( .A(n2081), .B(n2084), .Z(n2086) );
  NANDN U1517 ( .A(n2087), .B(n2088), .Z(n2083) );
  NAND U1518 ( .A(n2071), .B(n2089), .Z(n2088) );
  XNOR U1519 ( .A(n2071), .B(n2090), .Z(SUM[648]) );
  NANDN U1520 ( .A(n2087), .B(n2089), .Z(n2090) );
  NANDN U1521 ( .A(n2091), .B(n2092), .Z(n2071) );
  OR U1522 ( .A(n2093), .B(n2094), .Z(n2092) );
  XOR U1523 ( .A(n2095), .B(n2096), .Z(SUM[647]) );
  NANDN U1524 ( .A(n2097), .B(n2098), .Z(n2096) );
  ANDN U1525 ( .B(n2099), .A(n2100), .Z(n2095) );
  NAND U1526 ( .A(n2101), .B(n2102), .Z(n2099) );
  XNOR U1527 ( .A(n2101), .B(n2103), .Z(SUM[646]) );
  NANDN U1528 ( .A(n2100), .B(n2102), .Z(n2103) );
  NANDN U1529 ( .A(n2104), .B(n2105), .Z(n2101) );
  NAND U1530 ( .A(n2106), .B(n2107), .Z(n2105) );
  XNOR U1531 ( .A(n2106), .B(n2108), .Z(SUM[645]) );
  NANDN U1532 ( .A(n2104), .B(n2107), .Z(n2108) );
  NANDN U1533 ( .A(n2109), .B(n2110), .Z(n2106) );
  NANDN U1534 ( .A(n2094), .B(n2111), .Z(n2110) );
  XOR U1535 ( .A(n2094), .B(n2112), .Z(SUM[644]) );
  NANDN U1536 ( .A(n2109), .B(n2111), .Z(n2112) );
  ANDN U1537 ( .B(n2113), .A(n2114), .Z(n2094) );
  NANDN U1538 ( .A(n2115), .B(n1755), .Z(n2113) );
  XOR U1539 ( .A(n2116), .B(n2117), .Z(SUM[643]) );
  NANDN U1540 ( .A(n2118), .B(n2119), .Z(n2117) );
  ANDN U1541 ( .B(n2120), .A(n2121), .Z(n2116) );
  NAND U1542 ( .A(n2122), .B(n2123), .Z(n2120) );
  XNOR U1543 ( .A(n2122), .B(n2124), .Z(SUM[642]) );
  NANDN U1544 ( .A(n2121), .B(n2123), .Z(n2124) );
  NANDN U1545 ( .A(n2125), .B(n2126), .Z(n2122) );
  NAND U1546 ( .A(n2127), .B(n2128), .Z(n2126) );
  XNOR U1547 ( .A(n2127), .B(n2129), .Z(SUM[641]) );
  NANDN U1548 ( .A(n2125), .B(n2128), .Z(n2129) );
  NANDN U1549 ( .A(n2130), .B(n2131), .Z(n2127) );
  NAND U1550 ( .A(n1755), .B(n2132), .Z(n2131) );
  XNOR U1551 ( .A(n1755), .B(n2133), .Z(SUM[640]) );
  NANDN U1552 ( .A(n2130), .B(n2132), .Z(n2133) );
  NANDN U1553 ( .A(n2134), .B(n2135), .Z(n1755) );
  OR U1554 ( .A(n2136), .B(n2137), .Z(n2135) );
  XOR U1555 ( .A(n2138), .B(n2139), .Z(SUM[63]) );
  OR U1556 ( .A(n2140), .B(n2141), .Z(n2139) );
  ANDN U1557 ( .B(n2142), .A(n2143), .Z(n2138) );
  NANDN U1558 ( .A(n2144), .B(n2145), .Z(n2142) );
  XOR U1559 ( .A(n2146), .B(n2147), .Z(SUM[639]) );
  NANDN U1560 ( .A(n2148), .B(n2149), .Z(n2147) );
  ANDN U1561 ( .B(n2150), .A(n2151), .Z(n2146) );
  NAND U1562 ( .A(n2152), .B(n2153), .Z(n2150) );
  XNOR U1563 ( .A(n2152), .B(n2154), .Z(SUM[638]) );
  NANDN U1564 ( .A(n2151), .B(n2153), .Z(n2154) );
  NANDN U1565 ( .A(n2155), .B(n2156), .Z(n2152) );
  NAND U1566 ( .A(n2157), .B(n2158), .Z(n2156) );
  XNOR U1567 ( .A(n2157), .B(n2159), .Z(SUM[637]) );
  NANDN U1568 ( .A(n2155), .B(n2158), .Z(n2159) );
  NANDN U1569 ( .A(n2160), .B(n2161), .Z(n2157) );
  NAND U1570 ( .A(n2162), .B(n2163), .Z(n2161) );
  XNOR U1571 ( .A(n2162), .B(n2164), .Z(SUM[636]) );
  NANDN U1572 ( .A(n2160), .B(n2163), .Z(n2164) );
  NANDN U1573 ( .A(n2165), .B(n2166), .Z(n2162) );
  NANDN U1574 ( .A(n2167), .B(n2168), .Z(n2166) );
  XOR U1575 ( .A(n2169), .B(n2170), .Z(SUM[635]) );
  NANDN U1576 ( .A(n2171), .B(n2172), .Z(n2170) );
  ANDN U1577 ( .B(n2173), .A(n2174), .Z(n2169) );
  NAND U1578 ( .A(n2175), .B(n2176), .Z(n2173) );
  XNOR U1579 ( .A(n2175), .B(n2177), .Z(SUM[634]) );
  NANDN U1580 ( .A(n2174), .B(n2176), .Z(n2177) );
  NANDN U1581 ( .A(n2178), .B(n2179), .Z(n2175) );
  NAND U1582 ( .A(n2180), .B(n2181), .Z(n2179) );
  XNOR U1583 ( .A(n2180), .B(n2182), .Z(SUM[633]) );
  NANDN U1584 ( .A(n2178), .B(n2181), .Z(n2182) );
  NANDN U1585 ( .A(n2183), .B(n2184), .Z(n2180) );
  NAND U1586 ( .A(n2168), .B(n2185), .Z(n2184) );
  XNOR U1587 ( .A(n2168), .B(n2186), .Z(SUM[632]) );
  NANDN U1588 ( .A(n2183), .B(n2185), .Z(n2186) );
  NANDN U1589 ( .A(n2187), .B(n2188), .Z(n2168) );
  OR U1590 ( .A(n2189), .B(n2190), .Z(n2188) );
  XOR U1591 ( .A(n2191), .B(n2192), .Z(SUM[631]) );
  NANDN U1592 ( .A(n2193), .B(n2194), .Z(n2192) );
  ANDN U1593 ( .B(n2195), .A(n2196), .Z(n2191) );
  NAND U1594 ( .A(n2197), .B(n2198), .Z(n2195) );
  XNOR U1595 ( .A(n2197), .B(n2199), .Z(SUM[630]) );
  NANDN U1596 ( .A(n2196), .B(n2198), .Z(n2199) );
  NANDN U1597 ( .A(n2200), .B(n2201), .Z(n2197) );
  NAND U1598 ( .A(n2202), .B(n2203), .Z(n2201) );
  XNOR U1599 ( .A(n2145), .B(n2204), .Z(SUM[62]) );
  OR U1600 ( .A(n2144), .B(n2143), .Z(n2204) );
  NANDN U1601 ( .A(n2205), .B(n2206), .Z(n2145) );
  NANDN U1602 ( .A(n2207), .B(n2208), .Z(n2206) );
  XNOR U1603 ( .A(n2202), .B(n2209), .Z(SUM[629]) );
  NANDN U1604 ( .A(n2200), .B(n2203), .Z(n2209) );
  NANDN U1605 ( .A(n2210), .B(n2211), .Z(n2202) );
  NANDN U1606 ( .A(n2190), .B(n2212), .Z(n2211) );
  XOR U1607 ( .A(n2190), .B(n2213), .Z(SUM[628]) );
  NANDN U1608 ( .A(n2210), .B(n2212), .Z(n2213) );
  ANDN U1609 ( .B(n2214), .A(n2215), .Z(n2190) );
  NANDN U1610 ( .A(n2216), .B(n2217), .Z(n2214) );
  XOR U1611 ( .A(n2218), .B(n2219), .Z(SUM[627]) );
  NANDN U1612 ( .A(n2220), .B(n2221), .Z(n2219) );
  ANDN U1613 ( .B(n2222), .A(n2223), .Z(n2218) );
  NAND U1614 ( .A(n2224), .B(n2225), .Z(n2222) );
  XNOR U1615 ( .A(n2224), .B(n2226), .Z(SUM[626]) );
  NANDN U1616 ( .A(n2223), .B(n2225), .Z(n2226) );
  NANDN U1617 ( .A(n2227), .B(n2228), .Z(n2224) );
  NAND U1618 ( .A(n2229), .B(n2230), .Z(n2228) );
  XNOR U1619 ( .A(n2229), .B(n2231), .Z(SUM[625]) );
  NANDN U1620 ( .A(n2227), .B(n2230), .Z(n2231) );
  NANDN U1621 ( .A(n2232), .B(n2233), .Z(n2229) );
  NAND U1622 ( .A(n2217), .B(n2234), .Z(n2233) );
  XNOR U1623 ( .A(n2217), .B(n2235), .Z(SUM[624]) );
  NANDN U1624 ( .A(n2232), .B(n2234), .Z(n2235) );
  NANDN U1625 ( .A(n2236), .B(n2237), .Z(n2217) );
  NANDN U1626 ( .A(n2238), .B(n2239), .Z(n2237) );
  XOR U1627 ( .A(n2240), .B(n2241), .Z(SUM[623]) );
  NANDN U1628 ( .A(n2242), .B(n2243), .Z(n2241) );
  ANDN U1629 ( .B(n2244), .A(n2245), .Z(n2240) );
  NAND U1630 ( .A(n2246), .B(n2247), .Z(n2244) );
  XNOR U1631 ( .A(n2246), .B(n2248), .Z(SUM[622]) );
  NANDN U1632 ( .A(n2245), .B(n2247), .Z(n2248) );
  NANDN U1633 ( .A(n2249), .B(n2250), .Z(n2246) );
  NAND U1634 ( .A(n2251), .B(n2252), .Z(n2250) );
  XNOR U1635 ( .A(n2251), .B(n2253), .Z(SUM[621]) );
  NANDN U1636 ( .A(n2249), .B(n2252), .Z(n2253) );
  NANDN U1637 ( .A(n2254), .B(n2255), .Z(n2251) );
  NAND U1638 ( .A(n2256), .B(n2257), .Z(n2255) );
  XNOR U1639 ( .A(n2256), .B(n2258), .Z(SUM[620]) );
  NANDN U1640 ( .A(n2254), .B(n2257), .Z(n2258) );
  NANDN U1641 ( .A(n2259), .B(n2260), .Z(n2256) );
  NANDN U1642 ( .A(n2261), .B(n2262), .Z(n2260) );
  XNOR U1643 ( .A(n2208), .B(n2263), .Z(SUM[61]) );
  OR U1644 ( .A(n2207), .B(n2205), .Z(n2263) );
  NANDN U1645 ( .A(n2264), .B(n2265), .Z(n2208) );
  NANDN U1646 ( .A(n2266), .B(n2267), .Z(n2265) );
  XOR U1647 ( .A(n2268), .B(n2269), .Z(SUM[619]) );
  NANDN U1648 ( .A(n2270), .B(n2271), .Z(n2269) );
  ANDN U1649 ( .B(n2272), .A(n2273), .Z(n2268) );
  NAND U1650 ( .A(n2274), .B(n2275), .Z(n2272) );
  XNOR U1651 ( .A(n2274), .B(n2276), .Z(SUM[618]) );
  NANDN U1652 ( .A(n2273), .B(n2275), .Z(n2276) );
  NANDN U1653 ( .A(n2277), .B(n2278), .Z(n2274) );
  NAND U1654 ( .A(n2279), .B(n2280), .Z(n2278) );
  XNOR U1655 ( .A(n2279), .B(n2281), .Z(SUM[617]) );
  NANDN U1656 ( .A(n2277), .B(n2280), .Z(n2281) );
  NANDN U1657 ( .A(n2282), .B(n2283), .Z(n2279) );
  NAND U1658 ( .A(n2262), .B(n2284), .Z(n2283) );
  XNOR U1659 ( .A(n2262), .B(n2285), .Z(SUM[616]) );
  NANDN U1660 ( .A(n2282), .B(n2284), .Z(n2285) );
  NANDN U1661 ( .A(n2286), .B(n2287), .Z(n2262) );
  OR U1662 ( .A(n2288), .B(n2289), .Z(n2287) );
  XOR U1663 ( .A(n2290), .B(n2291), .Z(SUM[615]) );
  NANDN U1664 ( .A(n2292), .B(n2293), .Z(n2291) );
  ANDN U1665 ( .B(n2294), .A(n2295), .Z(n2290) );
  NAND U1666 ( .A(n2296), .B(n2297), .Z(n2294) );
  XNOR U1667 ( .A(n2296), .B(n2298), .Z(SUM[614]) );
  NANDN U1668 ( .A(n2295), .B(n2297), .Z(n2298) );
  NANDN U1669 ( .A(n2299), .B(n2300), .Z(n2296) );
  NAND U1670 ( .A(n2301), .B(n2302), .Z(n2300) );
  XNOR U1671 ( .A(n2301), .B(n2303), .Z(SUM[613]) );
  NANDN U1672 ( .A(n2299), .B(n2302), .Z(n2303) );
  NANDN U1673 ( .A(n2304), .B(n2305), .Z(n2301) );
  NANDN U1674 ( .A(n2289), .B(n2306), .Z(n2305) );
  XOR U1675 ( .A(n2289), .B(n2307), .Z(SUM[612]) );
  NANDN U1676 ( .A(n2304), .B(n2306), .Z(n2307) );
  ANDN U1677 ( .B(n2308), .A(n2309), .Z(n2289) );
  NANDN U1678 ( .A(n2310), .B(n2239), .Z(n2308) );
  XOR U1679 ( .A(n2311), .B(n2312), .Z(SUM[611]) );
  NANDN U1680 ( .A(n2313), .B(n2314), .Z(n2312) );
  ANDN U1681 ( .B(n2315), .A(n2316), .Z(n2311) );
  NAND U1682 ( .A(n2317), .B(n2318), .Z(n2315) );
  XNOR U1683 ( .A(n2317), .B(n2319), .Z(SUM[610]) );
  NANDN U1684 ( .A(n2316), .B(n2318), .Z(n2319) );
  NANDN U1685 ( .A(n2320), .B(n2321), .Z(n2317) );
  NAND U1686 ( .A(n2322), .B(n2323), .Z(n2321) );
  XNOR U1687 ( .A(n2267), .B(n2324), .Z(SUM[60]) );
  OR U1688 ( .A(n2266), .B(n2264), .Z(n2324) );
  NANDN U1689 ( .A(n2325), .B(n2326), .Z(n2267) );
  NANDN U1690 ( .A(n2327), .B(n2328), .Z(n2326) );
  XNOR U1691 ( .A(n2322), .B(n2329), .Z(SUM[609]) );
  NANDN U1692 ( .A(n2320), .B(n2323), .Z(n2329) );
  NANDN U1693 ( .A(n2330), .B(n2331), .Z(n2322) );
  NAND U1694 ( .A(n2239), .B(n2332), .Z(n2331) );
  XNOR U1695 ( .A(n2239), .B(n2333), .Z(SUM[608]) );
  NANDN U1696 ( .A(n2330), .B(n2332), .Z(n2333) );
  NANDN U1697 ( .A(n2334), .B(n2335), .Z(n2239) );
  OR U1698 ( .A(n2336), .B(n2337), .Z(n2335) );
  XOR U1699 ( .A(n2338), .B(n2339), .Z(SUM[607]) );
  NANDN U1700 ( .A(n2340), .B(n2341), .Z(n2339) );
  ANDN U1701 ( .B(n2342), .A(n2343), .Z(n2338) );
  NAND U1702 ( .A(n2344), .B(n2345), .Z(n2342) );
  XNOR U1703 ( .A(n2344), .B(n2346), .Z(SUM[606]) );
  NANDN U1704 ( .A(n2343), .B(n2345), .Z(n2346) );
  NANDN U1705 ( .A(n2347), .B(n2348), .Z(n2344) );
  NAND U1706 ( .A(n2349), .B(n2350), .Z(n2348) );
  XNOR U1707 ( .A(n2349), .B(n2351), .Z(SUM[605]) );
  NANDN U1708 ( .A(n2347), .B(n2350), .Z(n2351) );
  NANDN U1709 ( .A(n2352), .B(n2353), .Z(n2349) );
  NAND U1710 ( .A(n2354), .B(n2355), .Z(n2353) );
  XNOR U1711 ( .A(n2354), .B(n2356), .Z(SUM[604]) );
  NANDN U1712 ( .A(n2352), .B(n2355), .Z(n2356) );
  NANDN U1713 ( .A(n2357), .B(n2358), .Z(n2354) );
  NANDN U1714 ( .A(n2359), .B(n2360), .Z(n2358) );
  XOR U1715 ( .A(n2361), .B(n2362), .Z(SUM[603]) );
  NANDN U1716 ( .A(n2363), .B(n2364), .Z(n2362) );
  ANDN U1717 ( .B(n2365), .A(n2366), .Z(n2361) );
  NAND U1718 ( .A(n2367), .B(n2368), .Z(n2365) );
  XNOR U1719 ( .A(n2367), .B(n2369), .Z(SUM[602]) );
  NANDN U1720 ( .A(n2366), .B(n2368), .Z(n2369) );
  NANDN U1721 ( .A(n2370), .B(n2371), .Z(n2367) );
  NAND U1722 ( .A(n2372), .B(n2373), .Z(n2371) );
  XNOR U1723 ( .A(n2372), .B(n2374), .Z(SUM[601]) );
  NANDN U1724 ( .A(n2370), .B(n2373), .Z(n2374) );
  NANDN U1725 ( .A(n2375), .B(n2376), .Z(n2372) );
  NAND U1726 ( .A(n2360), .B(n2377), .Z(n2376) );
  XNOR U1727 ( .A(n2360), .B(n2378), .Z(SUM[600]) );
  NANDN U1728 ( .A(n2375), .B(n2377), .Z(n2378) );
  NANDN U1729 ( .A(n2379), .B(n2380), .Z(n2360) );
  OR U1730 ( .A(n2381), .B(n2382), .Z(n2380) );
  XNOR U1731 ( .A(n2383), .B(n2384), .Z(SUM[5]) );
  OR U1732 ( .A(n2385), .B(n2386), .Z(n2384) );
  XOR U1733 ( .A(n2387), .B(n2388), .Z(SUM[59]) );
  NANDN U1734 ( .A(n2389), .B(n2390), .Z(n2388) );
  ANDN U1735 ( .B(n2391), .A(n2392), .Z(n2387) );
  NAND U1736 ( .A(n2393), .B(n2394), .Z(n2391) );
  XOR U1737 ( .A(n2395), .B(n2396), .Z(SUM[599]) );
  NANDN U1738 ( .A(n2397), .B(n2398), .Z(n2396) );
  ANDN U1739 ( .B(n2399), .A(n2400), .Z(n2395) );
  NAND U1740 ( .A(n2401), .B(n2402), .Z(n2399) );
  XNOR U1741 ( .A(n2401), .B(n2403), .Z(SUM[598]) );
  NANDN U1742 ( .A(n2400), .B(n2402), .Z(n2403) );
  NANDN U1743 ( .A(n2404), .B(n2405), .Z(n2401) );
  NAND U1744 ( .A(n2406), .B(n2407), .Z(n2405) );
  XNOR U1745 ( .A(n2406), .B(n2408), .Z(SUM[597]) );
  NANDN U1746 ( .A(n2404), .B(n2407), .Z(n2408) );
  NANDN U1747 ( .A(n2409), .B(n2410), .Z(n2406) );
  NANDN U1748 ( .A(n2382), .B(n2411), .Z(n2410) );
  XOR U1749 ( .A(n2382), .B(n2412), .Z(SUM[596]) );
  NANDN U1750 ( .A(n2409), .B(n2411), .Z(n2412) );
  ANDN U1751 ( .B(n2413), .A(n2414), .Z(n2382) );
  OR U1752 ( .A(n2415), .B(n2337), .Z(n2413) );
  XOR U1753 ( .A(n2416), .B(n2417), .Z(SUM[595]) );
  NANDN U1754 ( .A(n2418), .B(n2419), .Z(n2417) );
  ANDN U1755 ( .B(n2420), .A(n2421), .Z(n2416) );
  NAND U1756 ( .A(n2422), .B(n2423), .Z(n2420) );
  XNOR U1757 ( .A(n2422), .B(n2424), .Z(SUM[594]) );
  NANDN U1758 ( .A(n2421), .B(n2423), .Z(n2424) );
  NANDN U1759 ( .A(n2425), .B(n2426), .Z(n2422) );
  NAND U1760 ( .A(n2427), .B(n2428), .Z(n2426) );
  XNOR U1761 ( .A(n2427), .B(n2429), .Z(SUM[593]) );
  NANDN U1762 ( .A(n2425), .B(n2428), .Z(n2429) );
  NANDN U1763 ( .A(n2430), .B(n2431), .Z(n2427) );
  NANDN U1764 ( .A(n2337), .B(n2432), .Z(n2431) );
  XOR U1765 ( .A(n2337), .B(n2433), .Z(SUM[592]) );
  NANDN U1766 ( .A(n2430), .B(n2432), .Z(n2433) );
  ANDN U1767 ( .B(n2434), .A(n2435), .Z(n2337) );
  OR U1768 ( .A(n2436), .B(n2137), .Z(n2434) );
  XOR U1769 ( .A(n2437), .B(n2438), .Z(SUM[591]) );
  NANDN U1770 ( .A(n2439), .B(n2440), .Z(n2438) );
  ANDN U1771 ( .B(n2441), .A(n2442), .Z(n2437) );
  NAND U1772 ( .A(n2443), .B(n2444), .Z(n2441) );
  XNOR U1773 ( .A(n2443), .B(n2445), .Z(SUM[590]) );
  NANDN U1774 ( .A(n2442), .B(n2444), .Z(n2445) );
  NANDN U1775 ( .A(n2446), .B(n2447), .Z(n2443) );
  NAND U1776 ( .A(n2448), .B(n2449), .Z(n2447) );
  XNOR U1777 ( .A(n2393), .B(n2450), .Z(SUM[58]) );
  NANDN U1778 ( .A(n2392), .B(n2394), .Z(n2450) );
  NANDN U1779 ( .A(n2451), .B(n2452), .Z(n2393) );
  NAND U1780 ( .A(n2453), .B(n2454), .Z(n2452) );
  XNOR U1781 ( .A(n2448), .B(n2455), .Z(SUM[589]) );
  NANDN U1782 ( .A(n2446), .B(n2449), .Z(n2455) );
  NANDN U1783 ( .A(n2456), .B(n2457), .Z(n2448) );
  NAND U1784 ( .A(n2458), .B(n2459), .Z(n2457) );
  XNOR U1785 ( .A(n2458), .B(n2460), .Z(SUM[588]) );
  NANDN U1786 ( .A(n2456), .B(n2459), .Z(n2460) );
  NANDN U1787 ( .A(n2461), .B(n2462), .Z(n2458) );
  NANDN U1788 ( .A(n2463), .B(n2464), .Z(n2462) );
  XOR U1789 ( .A(n2465), .B(n2466), .Z(SUM[587]) );
  NANDN U1790 ( .A(n2467), .B(n2468), .Z(n2466) );
  ANDN U1791 ( .B(n2469), .A(n2470), .Z(n2465) );
  NAND U1792 ( .A(n2471), .B(n2472), .Z(n2469) );
  XNOR U1793 ( .A(n2471), .B(n2473), .Z(SUM[586]) );
  NANDN U1794 ( .A(n2470), .B(n2472), .Z(n2473) );
  NANDN U1795 ( .A(n2474), .B(n2475), .Z(n2471) );
  NAND U1796 ( .A(n2476), .B(n2477), .Z(n2475) );
  XNOR U1797 ( .A(n2476), .B(n2478), .Z(SUM[585]) );
  NANDN U1798 ( .A(n2474), .B(n2477), .Z(n2478) );
  NANDN U1799 ( .A(n2479), .B(n2480), .Z(n2476) );
  NAND U1800 ( .A(n2464), .B(n2481), .Z(n2480) );
  XNOR U1801 ( .A(n2464), .B(n2482), .Z(SUM[584]) );
  NANDN U1802 ( .A(n2479), .B(n2481), .Z(n2482) );
  NANDN U1803 ( .A(n2483), .B(n2484), .Z(n2464) );
  OR U1804 ( .A(n2485), .B(n2486), .Z(n2484) );
  XOR U1805 ( .A(n2487), .B(n2488), .Z(SUM[583]) );
  NANDN U1806 ( .A(n2489), .B(n2490), .Z(n2488) );
  ANDN U1807 ( .B(n2491), .A(n2492), .Z(n2487) );
  NAND U1808 ( .A(n2493), .B(n2494), .Z(n2491) );
  XNOR U1809 ( .A(n2493), .B(n2495), .Z(SUM[582]) );
  NANDN U1810 ( .A(n2492), .B(n2494), .Z(n2495) );
  NANDN U1811 ( .A(n2496), .B(n2497), .Z(n2493) );
  NAND U1812 ( .A(n2498), .B(n2499), .Z(n2497) );
  XNOR U1813 ( .A(n2498), .B(n2500), .Z(SUM[581]) );
  NANDN U1814 ( .A(n2496), .B(n2499), .Z(n2500) );
  NANDN U1815 ( .A(n2501), .B(n2502), .Z(n2498) );
  NANDN U1816 ( .A(n2486), .B(n2503), .Z(n2502) );
  XOR U1817 ( .A(n2486), .B(n2504), .Z(SUM[580]) );
  NANDN U1818 ( .A(n2501), .B(n2503), .Z(n2504) );
  ANDN U1819 ( .B(n2505), .A(n2506), .Z(n2486) );
  OR U1820 ( .A(n2507), .B(n2137), .Z(n2505) );
  XNOR U1821 ( .A(n2453), .B(n2508), .Z(SUM[57]) );
  NANDN U1822 ( .A(n2451), .B(n2454), .Z(n2508) );
  NANDN U1823 ( .A(n2509), .B(n2510), .Z(n2453) );
  NAND U1824 ( .A(n2328), .B(n2511), .Z(n2510) );
  XOR U1825 ( .A(n2512), .B(n2513), .Z(SUM[579]) );
  NANDN U1826 ( .A(n2514), .B(n2515), .Z(n2513) );
  ANDN U1827 ( .B(n2516), .A(n2517), .Z(n2512) );
  NAND U1828 ( .A(n2518), .B(n2519), .Z(n2516) );
  XNOR U1829 ( .A(n2518), .B(n2520), .Z(SUM[578]) );
  NANDN U1830 ( .A(n2517), .B(n2519), .Z(n2520) );
  NANDN U1831 ( .A(n2521), .B(n2522), .Z(n2518) );
  NAND U1832 ( .A(n2523), .B(n2524), .Z(n2522) );
  XNOR U1833 ( .A(n2523), .B(n2525), .Z(SUM[577]) );
  NANDN U1834 ( .A(n2521), .B(n2524), .Z(n2525) );
  NANDN U1835 ( .A(n2526), .B(n2527), .Z(n2523) );
  NANDN U1836 ( .A(n2137), .B(n2528), .Z(n2527) );
  XOR U1837 ( .A(n2137), .B(n2529), .Z(SUM[576]) );
  NANDN U1838 ( .A(n2526), .B(n2528), .Z(n2529) );
  NOR U1839 ( .A(n2530), .B(n2531), .Z(n2137) );
  XOR U1840 ( .A(n2532), .B(n2533), .Z(SUM[575]) );
  NANDN U1841 ( .A(n2534), .B(n2535), .Z(n2533) );
  ANDN U1842 ( .B(n2536), .A(n2537), .Z(n2532) );
  NAND U1843 ( .A(n2538), .B(n2539), .Z(n2536) );
  XNOR U1844 ( .A(n2538), .B(n2540), .Z(SUM[574]) );
  NANDN U1845 ( .A(n2537), .B(n2539), .Z(n2540) );
  NANDN U1846 ( .A(n2541), .B(n2542), .Z(n2538) );
  NAND U1847 ( .A(n2543), .B(n2544), .Z(n2542) );
  XNOR U1848 ( .A(n2543), .B(n2545), .Z(SUM[573]) );
  NANDN U1849 ( .A(n2541), .B(n2544), .Z(n2545) );
  NANDN U1850 ( .A(n2546), .B(n2547), .Z(n2543) );
  NAND U1851 ( .A(n2548), .B(n2549), .Z(n2547) );
  XNOR U1852 ( .A(n2548), .B(n2550), .Z(SUM[572]) );
  NANDN U1853 ( .A(n2546), .B(n2549), .Z(n2550) );
  NANDN U1854 ( .A(n2551), .B(n2552), .Z(n2548) );
  NANDN U1855 ( .A(n2553), .B(n2554), .Z(n2552) );
  XOR U1856 ( .A(n2555), .B(n2556), .Z(SUM[571]) );
  NANDN U1857 ( .A(n2557), .B(n2558), .Z(n2556) );
  ANDN U1858 ( .B(n2559), .A(n2560), .Z(n2555) );
  NAND U1859 ( .A(n2561), .B(n2562), .Z(n2559) );
  XNOR U1860 ( .A(n2561), .B(n2563), .Z(SUM[570]) );
  NANDN U1861 ( .A(n2560), .B(n2562), .Z(n2563) );
  NANDN U1862 ( .A(n2564), .B(n2565), .Z(n2561) );
  NAND U1863 ( .A(n2566), .B(n2567), .Z(n2565) );
  XNOR U1864 ( .A(n2328), .B(n2568), .Z(SUM[56]) );
  NANDN U1865 ( .A(n2509), .B(n2511), .Z(n2568) );
  NANDN U1866 ( .A(n2569), .B(n2570), .Z(n2328) );
  OR U1867 ( .A(n2571), .B(n2572), .Z(n2570) );
  XNOR U1868 ( .A(n2566), .B(n2573), .Z(SUM[569]) );
  NANDN U1869 ( .A(n2564), .B(n2567), .Z(n2573) );
  NANDN U1870 ( .A(n2574), .B(n2575), .Z(n2566) );
  NAND U1871 ( .A(n2554), .B(n2576), .Z(n2575) );
  XNOR U1872 ( .A(n2554), .B(n2577), .Z(SUM[568]) );
  NANDN U1873 ( .A(n2574), .B(n2576), .Z(n2577) );
  NANDN U1874 ( .A(n2578), .B(n2579), .Z(n2554) );
  OR U1875 ( .A(n2580), .B(n2581), .Z(n2579) );
  XOR U1876 ( .A(n2582), .B(n2583), .Z(SUM[567]) );
  NANDN U1877 ( .A(n2584), .B(n2585), .Z(n2583) );
  ANDN U1878 ( .B(n2586), .A(n2587), .Z(n2582) );
  NAND U1879 ( .A(n2588), .B(n2589), .Z(n2586) );
  XNOR U1880 ( .A(n2588), .B(n2590), .Z(SUM[566]) );
  NANDN U1881 ( .A(n2587), .B(n2589), .Z(n2590) );
  NANDN U1882 ( .A(n2591), .B(n2592), .Z(n2588) );
  NAND U1883 ( .A(n2593), .B(n2594), .Z(n2592) );
  XNOR U1884 ( .A(n2593), .B(n2595), .Z(SUM[565]) );
  NANDN U1885 ( .A(n2591), .B(n2594), .Z(n2595) );
  NANDN U1886 ( .A(n2596), .B(n2597), .Z(n2593) );
  NANDN U1887 ( .A(n2581), .B(n2598), .Z(n2597) );
  XOR U1888 ( .A(n2581), .B(n2599), .Z(SUM[564]) );
  NANDN U1889 ( .A(n2596), .B(n2598), .Z(n2599) );
  ANDN U1890 ( .B(n2600), .A(n2601), .Z(n2581) );
  NANDN U1891 ( .A(n2602), .B(n2603), .Z(n2600) );
  XOR U1892 ( .A(n2604), .B(n2605), .Z(SUM[563]) );
  NANDN U1893 ( .A(n2606), .B(n2607), .Z(n2605) );
  ANDN U1894 ( .B(n2608), .A(n2609), .Z(n2604) );
  NAND U1895 ( .A(n2610), .B(n2611), .Z(n2608) );
  XNOR U1896 ( .A(n2610), .B(n2612), .Z(SUM[562]) );
  NANDN U1897 ( .A(n2609), .B(n2611), .Z(n2612) );
  NANDN U1898 ( .A(n2613), .B(n2614), .Z(n2610) );
  NAND U1899 ( .A(n2615), .B(n2616), .Z(n2614) );
  XNOR U1900 ( .A(n2615), .B(n2617), .Z(SUM[561]) );
  NANDN U1901 ( .A(n2613), .B(n2616), .Z(n2617) );
  NANDN U1902 ( .A(n2618), .B(n2619), .Z(n2615) );
  NAND U1903 ( .A(n2603), .B(n2620), .Z(n2619) );
  XNOR U1904 ( .A(n2603), .B(n2621), .Z(SUM[560]) );
  NANDN U1905 ( .A(n2618), .B(n2620), .Z(n2621) );
  NANDN U1906 ( .A(n2622), .B(n2623), .Z(n2603) );
  NANDN U1907 ( .A(n2624), .B(n2625), .Z(n2623) );
  XOR U1908 ( .A(n2626), .B(n2627), .Z(SUM[55]) );
  NANDN U1909 ( .A(n2628), .B(n2629), .Z(n2627) );
  ANDN U1910 ( .B(n2630), .A(n2631), .Z(n2626) );
  NAND U1911 ( .A(n2632), .B(n2633), .Z(n2630) );
  XOR U1912 ( .A(n2634), .B(n2635), .Z(SUM[559]) );
  NANDN U1913 ( .A(n2636), .B(n2637), .Z(n2635) );
  ANDN U1914 ( .B(n2638), .A(n2639), .Z(n2634) );
  NAND U1915 ( .A(n2640), .B(n2641), .Z(n2638) );
  XNOR U1916 ( .A(n2640), .B(n2642), .Z(SUM[558]) );
  NANDN U1917 ( .A(n2639), .B(n2641), .Z(n2642) );
  NANDN U1918 ( .A(n2643), .B(n2644), .Z(n2640) );
  NAND U1919 ( .A(n2645), .B(n2646), .Z(n2644) );
  XNOR U1920 ( .A(n2645), .B(n2647), .Z(SUM[557]) );
  NANDN U1921 ( .A(n2643), .B(n2646), .Z(n2647) );
  NANDN U1922 ( .A(n2648), .B(n2649), .Z(n2645) );
  NAND U1923 ( .A(n2650), .B(n2651), .Z(n2649) );
  XNOR U1924 ( .A(n2650), .B(n2652), .Z(SUM[556]) );
  NANDN U1925 ( .A(n2648), .B(n2651), .Z(n2652) );
  NANDN U1926 ( .A(n2653), .B(n2654), .Z(n2650) );
  NANDN U1927 ( .A(n2655), .B(n2656), .Z(n2654) );
  XOR U1928 ( .A(n2657), .B(n2658), .Z(SUM[555]) );
  NANDN U1929 ( .A(n2659), .B(n2660), .Z(n2658) );
  ANDN U1930 ( .B(n2661), .A(n2662), .Z(n2657) );
  NAND U1931 ( .A(n2663), .B(n2664), .Z(n2661) );
  XNOR U1932 ( .A(n2663), .B(n2665), .Z(SUM[554]) );
  NANDN U1933 ( .A(n2662), .B(n2664), .Z(n2665) );
  NANDN U1934 ( .A(n2666), .B(n2667), .Z(n2663) );
  NAND U1935 ( .A(n2668), .B(n2669), .Z(n2667) );
  XNOR U1936 ( .A(n2668), .B(n2670), .Z(SUM[553]) );
  NANDN U1937 ( .A(n2666), .B(n2669), .Z(n2670) );
  NANDN U1938 ( .A(n2671), .B(n2672), .Z(n2668) );
  NAND U1939 ( .A(n2656), .B(n2673), .Z(n2672) );
  XNOR U1940 ( .A(n2656), .B(n2674), .Z(SUM[552]) );
  NANDN U1941 ( .A(n2671), .B(n2673), .Z(n2674) );
  NANDN U1942 ( .A(n2675), .B(n2676), .Z(n2656) );
  OR U1943 ( .A(n2677), .B(n2678), .Z(n2676) );
  XOR U1944 ( .A(n2679), .B(n2680), .Z(SUM[551]) );
  NANDN U1945 ( .A(n2681), .B(n2682), .Z(n2680) );
  ANDN U1946 ( .B(n2683), .A(n2684), .Z(n2679) );
  NAND U1947 ( .A(n2685), .B(n2686), .Z(n2683) );
  XNOR U1948 ( .A(n2685), .B(n2687), .Z(SUM[550]) );
  NANDN U1949 ( .A(n2684), .B(n2686), .Z(n2687) );
  NANDN U1950 ( .A(n2688), .B(n2689), .Z(n2685) );
  NAND U1951 ( .A(n2690), .B(n2691), .Z(n2689) );
  XNOR U1952 ( .A(n2632), .B(n2692), .Z(SUM[54]) );
  NANDN U1953 ( .A(n2631), .B(n2633), .Z(n2692) );
  NANDN U1954 ( .A(n2693), .B(n2694), .Z(n2632) );
  NAND U1955 ( .A(n2695), .B(n2696), .Z(n2694) );
  XNOR U1956 ( .A(n2690), .B(n2697), .Z(SUM[549]) );
  NANDN U1957 ( .A(n2688), .B(n2691), .Z(n2697) );
  NANDN U1958 ( .A(n2698), .B(n2699), .Z(n2690) );
  NANDN U1959 ( .A(n2678), .B(n2700), .Z(n2699) );
  XOR U1960 ( .A(n2678), .B(n2701), .Z(SUM[548]) );
  NANDN U1961 ( .A(n2698), .B(n2700), .Z(n2701) );
  ANDN U1962 ( .B(n2702), .A(n2703), .Z(n2678) );
  NANDN U1963 ( .A(n2704), .B(n2625), .Z(n2702) );
  XOR U1964 ( .A(n2705), .B(n2706), .Z(SUM[547]) );
  NANDN U1965 ( .A(n2707), .B(n2708), .Z(n2706) );
  ANDN U1966 ( .B(n2709), .A(n2710), .Z(n2705) );
  NAND U1967 ( .A(n2711), .B(n2712), .Z(n2709) );
  XNOR U1968 ( .A(n2711), .B(n2713), .Z(SUM[546]) );
  NANDN U1969 ( .A(n2710), .B(n2712), .Z(n2713) );
  NANDN U1970 ( .A(n2714), .B(n2715), .Z(n2711) );
  NAND U1971 ( .A(n2716), .B(n2717), .Z(n2715) );
  XNOR U1972 ( .A(n2716), .B(n2718), .Z(SUM[545]) );
  NANDN U1973 ( .A(n2714), .B(n2717), .Z(n2718) );
  NANDN U1974 ( .A(n2719), .B(n2720), .Z(n2716) );
  NAND U1975 ( .A(n2625), .B(n2721), .Z(n2720) );
  XNOR U1976 ( .A(n2625), .B(n2722), .Z(SUM[544]) );
  NANDN U1977 ( .A(n2719), .B(n2721), .Z(n2722) );
  NANDN U1978 ( .A(n2723), .B(n2724), .Z(n2625) );
  OR U1979 ( .A(n2725), .B(n2726), .Z(n2724) );
  XOR U1980 ( .A(n2727), .B(n2728), .Z(SUM[543]) );
  NANDN U1981 ( .A(n2729), .B(n2730), .Z(n2728) );
  ANDN U1982 ( .B(n2731), .A(n2732), .Z(n2727) );
  NAND U1983 ( .A(n2733), .B(n2734), .Z(n2731) );
  XNOR U1984 ( .A(n2733), .B(n2735), .Z(SUM[542]) );
  NANDN U1985 ( .A(n2732), .B(n2734), .Z(n2735) );
  NANDN U1986 ( .A(n2736), .B(n2737), .Z(n2733) );
  NAND U1987 ( .A(n2738), .B(n2739), .Z(n2737) );
  XNOR U1988 ( .A(n2738), .B(n2740), .Z(SUM[541]) );
  NANDN U1989 ( .A(n2736), .B(n2739), .Z(n2740) );
  NANDN U1990 ( .A(n2741), .B(n2742), .Z(n2738) );
  NAND U1991 ( .A(n2743), .B(n2744), .Z(n2742) );
  XNOR U1992 ( .A(n2743), .B(n2745), .Z(SUM[540]) );
  NANDN U1993 ( .A(n2741), .B(n2744), .Z(n2745) );
  NANDN U1994 ( .A(n2746), .B(n2747), .Z(n2743) );
  NANDN U1995 ( .A(n2748), .B(n2749), .Z(n2747) );
  XNOR U1996 ( .A(n2695), .B(n2750), .Z(SUM[53]) );
  NANDN U1997 ( .A(n2693), .B(n2696), .Z(n2750) );
  NANDN U1998 ( .A(n2751), .B(n2752), .Z(n2695) );
  NANDN U1999 ( .A(n2572), .B(n2753), .Z(n2752) );
  XOR U2000 ( .A(n2754), .B(n2755), .Z(SUM[539]) );
  NANDN U2001 ( .A(n2756), .B(n2757), .Z(n2755) );
  ANDN U2002 ( .B(n2758), .A(n2759), .Z(n2754) );
  NAND U2003 ( .A(n2760), .B(n2761), .Z(n2758) );
  XNOR U2004 ( .A(n2760), .B(n2762), .Z(SUM[538]) );
  NANDN U2005 ( .A(n2759), .B(n2761), .Z(n2762) );
  NANDN U2006 ( .A(n2763), .B(n2764), .Z(n2760) );
  NAND U2007 ( .A(n2765), .B(n2766), .Z(n2764) );
  XNOR U2008 ( .A(n2765), .B(n2767), .Z(SUM[537]) );
  NANDN U2009 ( .A(n2763), .B(n2766), .Z(n2767) );
  NANDN U2010 ( .A(n2768), .B(n2769), .Z(n2765) );
  NAND U2011 ( .A(n2749), .B(n2770), .Z(n2769) );
  XNOR U2012 ( .A(n2749), .B(n2771), .Z(SUM[536]) );
  NANDN U2013 ( .A(n2768), .B(n2770), .Z(n2771) );
  NANDN U2014 ( .A(n2772), .B(n2773), .Z(n2749) );
  OR U2015 ( .A(n2774), .B(n2775), .Z(n2773) );
  XOR U2016 ( .A(n2776), .B(n2777), .Z(SUM[535]) );
  NANDN U2017 ( .A(n2778), .B(n2779), .Z(n2777) );
  ANDN U2018 ( .B(n2780), .A(n2781), .Z(n2776) );
  NAND U2019 ( .A(n2782), .B(n2783), .Z(n2780) );
  XNOR U2020 ( .A(n2782), .B(n2784), .Z(SUM[534]) );
  NANDN U2021 ( .A(n2781), .B(n2783), .Z(n2784) );
  NANDN U2022 ( .A(n2785), .B(n2786), .Z(n2782) );
  NAND U2023 ( .A(n2787), .B(n2788), .Z(n2786) );
  XNOR U2024 ( .A(n2787), .B(n2789), .Z(SUM[533]) );
  NANDN U2025 ( .A(n2785), .B(n2788), .Z(n2789) );
  NANDN U2026 ( .A(n2790), .B(n2791), .Z(n2787) );
  NANDN U2027 ( .A(n2775), .B(n2792), .Z(n2791) );
  XOR U2028 ( .A(n2775), .B(n2793), .Z(SUM[532]) );
  NANDN U2029 ( .A(n2790), .B(n2792), .Z(n2793) );
  ANDN U2030 ( .B(n2794), .A(n2795), .Z(n2775) );
  OR U2031 ( .A(n2796), .B(n2726), .Z(n2794) );
  XOR U2032 ( .A(n2797), .B(n2798), .Z(SUM[531]) );
  NANDN U2033 ( .A(n2799), .B(n2800), .Z(n2798) );
  ANDN U2034 ( .B(n2801), .A(n2802), .Z(n2797) );
  NAND U2035 ( .A(n2803), .B(n2804), .Z(n2801) );
  XNOR U2036 ( .A(n2803), .B(n2805), .Z(SUM[530]) );
  NANDN U2037 ( .A(n2802), .B(n2804), .Z(n2805) );
  NANDN U2038 ( .A(n2806), .B(n2807), .Z(n2803) );
  NAND U2039 ( .A(n2808), .B(n2809), .Z(n2807) );
  XOR U2040 ( .A(n2572), .B(n2810), .Z(SUM[52]) );
  NANDN U2041 ( .A(n2751), .B(n2753), .Z(n2810) );
  NOR U2042 ( .A(n2811), .B(n2812), .Z(n2572) );
  XNOR U2043 ( .A(n2808), .B(n2813), .Z(SUM[529]) );
  NANDN U2044 ( .A(n2806), .B(n2809), .Z(n2813) );
  NANDN U2045 ( .A(n2814), .B(n2815), .Z(n2808) );
  NANDN U2046 ( .A(n2726), .B(n2816), .Z(n2815) );
  XOR U2047 ( .A(n2726), .B(n2817), .Z(SUM[528]) );
  NANDN U2048 ( .A(n2814), .B(n2816), .Z(n2817) );
  ANDN U2049 ( .B(n2818), .A(n2819), .Z(n2726) );
  OR U2050 ( .A(n2820), .B(n2821), .Z(n2818) );
  XOR U2051 ( .A(n2822), .B(n2823), .Z(SUM[527]) );
  NANDN U2052 ( .A(n2824), .B(n2825), .Z(n2823) );
  ANDN U2053 ( .B(n2826), .A(n2827), .Z(n2822) );
  NAND U2054 ( .A(n2828), .B(n2829), .Z(n2826) );
  XNOR U2055 ( .A(n2828), .B(n2830), .Z(SUM[526]) );
  NANDN U2056 ( .A(n2827), .B(n2829), .Z(n2830) );
  NANDN U2057 ( .A(n2831), .B(n2832), .Z(n2828) );
  NAND U2058 ( .A(n2833), .B(n2834), .Z(n2832) );
  XNOR U2059 ( .A(n2833), .B(n2835), .Z(SUM[525]) );
  NANDN U2060 ( .A(n2831), .B(n2834), .Z(n2835) );
  NANDN U2061 ( .A(n2836), .B(n2837), .Z(n2833) );
  NAND U2062 ( .A(n2838), .B(n2839), .Z(n2837) );
  XNOR U2063 ( .A(n2838), .B(n2840), .Z(SUM[524]) );
  NANDN U2064 ( .A(n2836), .B(n2839), .Z(n2840) );
  NANDN U2065 ( .A(n2841), .B(n2842), .Z(n2838) );
  NANDN U2066 ( .A(n2843), .B(n2844), .Z(n2842) );
  XOR U2067 ( .A(n2845), .B(n2846), .Z(SUM[523]) );
  NANDN U2068 ( .A(n2847), .B(n2848), .Z(n2846) );
  ANDN U2069 ( .B(n2849), .A(n2850), .Z(n2845) );
  NAND U2070 ( .A(n2851), .B(n2852), .Z(n2849) );
  XNOR U2071 ( .A(n2851), .B(n2853), .Z(SUM[522]) );
  NANDN U2072 ( .A(n2850), .B(n2852), .Z(n2853) );
  NANDN U2073 ( .A(n2854), .B(n2855), .Z(n2851) );
  NAND U2074 ( .A(n2856), .B(n2857), .Z(n2855) );
  XNOR U2075 ( .A(n2856), .B(n2858), .Z(SUM[521]) );
  NANDN U2076 ( .A(n2854), .B(n2857), .Z(n2858) );
  NANDN U2077 ( .A(n2859), .B(n2860), .Z(n2856) );
  NAND U2078 ( .A(n2844), .B(n2861), .Z(n2860) );
  XNOR U2079 ( .A(n2844), .B(n2862), .Z(SUM[520]) );
  NANDN U2080 ( .A(n2859), .B(n2861), .Z(n2862) );
  NANDN U2081 ( .A(n2863), .B(n2864), .Z(n2844) );
  OR U2082 ( .A(n2865), .B(n2866), .Z(n2864) );
  XOR U2083 ( .A(n2867), .B(n2868), .Z(SUM[51]) );
  NANDN U2084 ( .A(n2869), .B(n2870), .Z(n2868) );
  ANDN U2085 ( .B(n2871), .A(n2872), .Z(n2867) );
  NAND U2086 ( .A(n2873), .B(n2874), .Z(n2871) );
  XOR U2087 ( .A(n2875), .B(n2876), .Z(SUM[519]) );
  NANDN U2088 ( .A(n2877), .B(n2878), .Z(n2876) );
  ANDN U2089 ( .B(n2879), .A(n2880), .Z(n2875) );
  NAND U2090 ( .A(n2881), .B(n2882), .Z(n2879) );
  XNOR U2091 ( .A(n2881), .B(n2883), .Z(SUM[518]) );
  NANDN U2092 ( .A(n2880), .B(n2882), .Z(n2883) );
  NANDN U2093 ( .A(n2884), .B(n2885), .Z(n2881) );
  NAND U2094 ( .A(n2886), .B(n2887), .Z(n2885) );
  XNOR U2095 ( .A(n2886), .B(n2888), .Z(SUM[517]) );
  NANDN U2096 ( .A(n2884), .B(n2887), .Z(n2888) );
  NANDN U2097 ( .A(n2889), .B(n2890), .Z(n2886) );
  NANDN U2098 ( .A(n2866), .B(n2891), .Z(n2890) );
  XOR U2099 ( .A(n2866), .B(n2892), .Z(SUM[516]) );
  NANDN U2100 ( .A(n2889), .B(n2891), .Z(n2892) );
  ANDN U2101 ( .B(n2893), .A(n2894), .Z(n2866) );
  OR U2102 ( .A(n2895), .B(n2821), .Z(n2893) );
  XOR U2103 ( .A(n2896), .B(n2897), .Z(SUM[515]) );
  NANDN U2104 ( .A(n2898), .B(n2899), .Z(n2897) );
  ANDN U2105 ( .B(n2900), .A(n2901), .Z(n2896) );
  NAND U2106 ( .A(n2902), .B(n2903), .Z(n2900) );
  XNOR U2107 ( .A(n2902), .B(n2904), .Z(SUM[514]) );
  NANDN U2108 ( .A(n2901), .B(n2903), .Z(n2904) );
  NANDN U2109 ( .A(n2905), .B(n2906), .Z(n2902) );
  NAND U2110 ( .A(n2907), .B(n2908), .Z(n2906) );
  XNOR U2111 ( .A(n2907), .B(n2909), .Z(SUM[513]) );
  NANDN U2112 ( .A(n2905), .B(n2908), .Z(n2909) );
  NANDN U2113 ( .A(n2910), .B(n2911), .Z(n2907) );
  NANDN U2114 ( .A(n2821), .B(n2912), .Z(n2911) );
  XOR U2115 ( .A(n2821), .B(n2913), .Z(SUM[512]) );
  NANDN U2116 ( .A(n2910), .B(n2912), .Z(n2913) );
  XOR U2117 ( .A(n2914), .B(n2915), .Z(SUM[511]) );
  OR U2118 ( .A(n2916), .B(n2917), .Z(n2915) );
  ANDN U2119 ( .B(n2918), .A(n2919), .Z(n2914) );
  NAND U2120 ( .A(n2920), .B(n2921), .Z(n2918) );
  XNOR U2121 ( .A(n2920), .B(n2922), .Z(SUM[510]) );
  NANDN U2122 ( .A(n2919), .B(n2921), .Z(n2922) );
  NANDN U2123 ( .A(n2923), .B(n2924), .Z(n2920) );
  NAND U2124 ( .A(n2925), .B(n2926), .Z(n2924) );
  XNOR U2125 ( .A(n2873), .B(n2927), .Z(SUM[50]) );
  NANDN U2126 ( .A(n2872), .B(n2874), .Z(n2927) );
  NANDN U2127 ( .A(n2928), .B(n2929), .Z(n2873) );
  NAND U2128 ( .A(n2930), .B(n2931), .Z(n2929) );
  XNOR U2129 ( .A(n2925), .B(n2932), .Z(SUM[509]) );
  NANDN U2130 ( .A(n2923), .B(n2926), .Z(n2932) );
  NANDN U2131 ( .A(n2933), .B(n2934), .Z(n2925) );
  NANDN U2132 ( .A(n2935), .B(n2936), .Z(n2934) );
  XNOR U2133 ( .A(n2936), .B(n2937), .Z(SUM[508]) );
  OR U2134 ( .A(n2935), .B(n2933), .Z(n2937) );
  NANDN U2135 ( .A(n2938), .B(n2939), .Z(n2936) );
  NANDN U2136 ( .A(n2940), .B(n2941), .Z(n2939) );
  XOR U2137 ( .A(n2942), .B(n2943), .Z(SUM[507]) );
  NANDN U2138 ( .A(n2944), .B(n2945), .Z(n2943) );
  ANDN U2139 ( .B(n2946), .A(n2947), .Z(n2942) );
  NAND U2140 ( .A(n2948), .B(n2949), .Z(n2946) );
  XNOR U2141 ( .A(n2948), .B(n2950), .Z(SUM[506]) );
  NANDN U2142 ( .A(n2947), .B(n2949), .Z(n2950) );
  NANDN U2143 ( .A(n2951), .B(n2952), .Z(n2948) );
  NAND U2144 ( .A(n2953), .B(n2954), .Z(n2952) );
  XNOR U2145 ( .A(n2953), .B(n2955), .Z(SUM[505]) );
  NANDN U2146 ( .A(n2951), .B(n2954), .Z(n2955) );
  NANDN U2147 ( .A(n2956), .B(n2957), .Z(n2953) );
  NAND U2148 ( .A(n2941), .B(n2958), .Z(n2957) );
  XNOR U2149 ( .A(n2941), .B(n2959), .Z(SUM[504]) );
  NANDN U2150 ( .A(n2956), .B(n2958), .Z(n2959) );
  NANDN U2151 ( .A(n2960), .B(n2961), .Z(n2941) );
  NANDN U2152 ( .A(n2962), .B(n2963), .Z(n2961) );
  XOR U2153 ( .A(n2964), .B(n2965), .Z(SUM[503]) );
  NANDN U2154 ( .A(n2966), .B(n2967), .Z(n2965) );
  ANDN U2155 ( .B(n2968), .A(n2969), .Z(n2964) );
  NAND U2156 ( .A(n2970), .B(n2971), .Z(n2968) );
  XNOR U2157 ( .A(n2970), .B(n2972), .Z(SUM[502]) );
  NANDN U2158 ( .A(n2969), .B(n2971), .Z(n2972) );
  NANDN U2159 ( .A(n2973), .B(n2974), .Z(n2970) );
  NAND U2160 ( .A(n2975), .B(n2976), .Z(n2974) );
  XNOR U2161 ( .A(n2975), .B(n2977), .Z(SUM[501]) );
  NANDN U2162 ( .A(n2973), .B(n2976), .Z(n2977) );
  NANDN U2163 ( .A(n2978), .B(n2979), .Z(n2975) );
  NANDN U2164 ( .A(n2962), .B(n2980), .Z(n2979) );
  XOR U2165 ( .A(n2962), .B(n2981), .Z(SUM[500]) );
  NANDN U2166 ( .A(n2978), .B(n2980), .Z(n2981) );
  ANDN U2167 ( .B(n2982), .A(n2983), .Z(n2962) );
  NANDN U2168 ( .A(n2984), .B(n2985), .Z(n2982) );
  XOR U2169 ( .A(n2986), .B(n2987), .Z(SUM[4]) );
  OR U2170 ( .A(n2988), .B(n2989), .Z(n2987) );
  XNOR U2171 ( .A(n2930), .B(n2990), .Z(SUM[49]) );
  NANDN U2172 ( .A(n2928), .B(n2931), .Z(n2990) );
  NANDN U2173 ( .A(n2991), .B(n2992), .Z(n2930) );
  NANDN U2174 ( .A(n2993), .B(n2994), .Z(n2992) );
  XOR U2175 ( .A(n2995), .B(n2996), .Z(SUM[499]) );
  NANDN U2176 ( .A(n2997), .B(n2998), .Z(n2996) );
  ANDN U2177 ( .B(n2999), .A(n3000), .Z(n2995) );
  NANDN U2178 ( .A(n3001), .B(n3002), .Z(n2999) );
  XNOR U2179 ( .A(n3002), .B(n3003), .Z(SUM[498]) );
  OR U2180 ( .A(n3001), .B(n3000), .Z(n3003) );
  NANDN U2181 ( .A(n3004), .B(n3005), .Z(n3002) );
  NAND U2182 ( .A(n3006), .B(n3007), .Z(n3005) );
  XNOR U2183 ( .A(n3006), .B(n3008), .Z(SUM[497]) );
  NANDN U2184 ( .A(n3004), .B(n3007), .Z(n3008) );
  NANDN U2185 ( .A(n3009), .B(n3010), .Z(n3006) );
  NAND U2186 ( .A(n2985), .B(n3011), .Z(n3010) );
  XNOR U2187 ( .A(n2985), .B(n3012), .Z(SUM[496]) );
  NANDN U2188 ( .A(n3009), .B(n3011), .Z(n3012) );
  NANDN U2189 ( .A(n3013), .B(n3014), .Z(n2985) );
  NANDN U2190 ( .A(n3015), .B(n3016), .Z(n3014) );
  XOR U2191 ( .A(n3017), .B(n3018), .Z(SUM[495]) );
  NANDN U2192 ( .A(n3019), .B(n3020), .Z(n3018) );
  ANDN U2193 ( .B(n3021), .A(n3022), .Z(n3017) );
  NAND U2194 ( .A(n3023), .B(n3024), .Z(n3021) );
  XNOR U2195 ( .A(n3023), .B(n3025), .Z(SUM[494]) );
  NANDN U2196 ( .A(n3022), .B(n3024), .Z(n3025) );
  NANDN U2197 ( .A(n3026), .B(n3027), .Z(n3023) );
  NAND U2198 ( .A(n3028), .B(n3029), .Z(n3027) );
  XNOR U2199 ( .A(n3028), .B(n3030), .Z(SUM[493]) );
  NANDN U2200 ( .A(n3026), .B(n3029), .Z(n3030) );
  NANDN U2201 ( .A(n3031), .B(n3032), .Z(n3028) );
  NAND U2202 ( .A(n3033), .B(n3034), .Z(n3032) );
  XNOR U2203 ( .A(n3033), .B(n3035), .Z(SUM[492]) );
  NANDN U2204 ( .A(n3031), .B(n3034), .Z(n3035) );
  NANDN U2205 ( .A(n3036), .B(n3037), .Z(n3033) );
  NAND U2206 ( .A(n3038), .B(n3039), .Z(n3037) );
  XOR U2207 ( .A(n3040), .B(n3041), .Z(SUM[491]) );
  NANDN U2208 ( .A(n3042), .B(n3043), .Z(n3041) );
  ANDN U2209 ( .B(n3044), .A(n3045), .Z(n3040) );
  NAND U2210 ( .A(n3046), .B(n3047), .Z(n3044) );
  XNOR U2211 ( .A(n3046), .B(n3048), .Z(SUM[490]) );
  NANDN U2212 ( .A(n3045), .B(n3047), .Z(n3048) );
  NANDN U2213 ( .A(n3049), .B(n3050), .Z(n3046) );
  NAND U2214 ( .A(n3051), .B(n3052), .Z(n3050) );
  XOR U2215 ( .A(n2993), .B(n3053), .Z(SUM[48]) );
  NANDN U2216 ( .A(n2991), .B(n2994), .Z(n3053) );
  XNOR U2217 ( .A(n3051), .B(n3054), .Z(SUM[489]) );
  NANDN U2218 ( .A(n3049), .B(n3052), .Z(n3054) );
  NANDN U2219 ( .A(n3055), .B(n3056), .Z(n3051) );
  NAND U2220 ( .A(n3039), .B(n3057), .Z(n3056) );
  XNOR U2221 ( .A(n3039), .B(n3058), .Z(SUM[488]) );
  NANDN U2222 ( .A(n3055), .B(n3057), .Z(n3058) );
  NANDN U2223 ( .A(n3059), .B(n3060), .Z(n3039) );
  OR U2224 ( .A(n3061), .B(n3062), .Z(n3060) );
  XOR U2225 ( .A(n3063), .B(n3064), .Z(SUM[487]) );
  NANDN U2226 ( .A(n3065), .B(n3066), .Z(n3064) );
  ANDN U2227 ( .B(n3067), .A(n3068), .Z(n3063) );
  NAND U2228 ( .A(n3069), .B(n3070), .Z(n3067) );
  XNOR U2229 ( .A(n3069), .B(n3071), .Z(SUM[486]) );
  NANDN U2230 ( .A(n3068), .B(n3070), .Z(n3071) );
  NANDN U2231 ( .A(n3072), .B(n3073), .Z(n3069) );
  NAND U2232 ( .A(n3074), .B(n3075), .Z(n3073) );
  XNOR U2233 ( .A(n3074), .B(n3076), .Z(SUM[485]) );
  NANDN U2234 ( .A(n3072), .B(n3075), .Z(n3076) );
  NANDN U2235 ( .A(n3077), .B(n3078), .Z(n3074) );
  NANDN U2236 ( .A(n3062), .B(n3079), .Z(n3078) );
  XOR U2237 ( .A(n3062), .B(n3080), .Z(SUM[484]) );
  NANDN U2238 ( .A(n3077), .B(n3079), .Z(n3080) );
  ANDN U2239 ( .B(n3081), .A(n3082), .Z(n3062) );
  NANDN U2240 ( .A(n3083), .B(n3016), .Z(n3081) );
  XOR U2241 ( .A(n3084), .B(n3085), .Z(SUM[483]) );
  NANDN U2242 ( .A(n3086), .B(n3087), .Z(n3085) );
  ANDN U2243 ( .B(n3088), .A(n3089), .Z(n3084) );
  NAND U2244 ( .A(n3090), .B(n3091), .Z(n3088) );
  XNOR U2245 ( .A(n3090), .B(n3092), .Z(SUM[482]) );
  NANDN U2246 ( .A(n3089), .B(n3091), .Z(n3092) );
  NANDN U2247 ( .A(n3093), .B(n3094), .Z(n3090) );
  NAND U2248 ( .A(n3095), .B(n3096), .Z(n3094) );
  XNOR U2249 ( .A(n3095), .B(n3097), .Z(SUM[481]) );
  NANDN U2250 ( .A(n3093), .B(n3096), .Z(n3097) );
  NANDN U2251 ( .A(n3098), .B(n3099), .Z(n3095) );
  NAND U2252 ( .A(n3016), .B(n3100), .Z(n3099) );
  XNOR U2253 ( .A(n3016), .B(n3101), .Z(SUM[480]) );
  NANDN U2254 ( .A(n3098), .B(n3100), .Z(n3101) );
  NANDN U2255 ( .A(n3102), .B(n3103), .Z(n3016) );
  NANDN U2256 ( .A(n3104), .B(n3105), .Z(n3103) );
  XOR U2257 ( .A(n3106), .B(n3107), .Z(SUM[47]) );
  OR U2258 ( .A(n3108), .B(n3109), .Z(n3107) );
  ANDN U2259 ( .B(n3110), .A(n3111), .Z(n3106) );
  NANDN U2260 ( .A(n3112), .B(n3113), .Z(n3110) );
  XOR U2261 ( .A(n3114), .B(n3115), .Z(SUM[479]) );
  NANDN U2262 ( .A(n3116), .B(n3117), .Z(n3115) );
  ANDN U2263 ( .B(n3118), .A(n3119), .Z(n3114) );
  NAND U2264 ( .A(n3120), .B(n3121), .Z(n3118) );
  XNOR U2265 ( .A(n3120), .B(n3122), .Z(SUM[478]) );
  NANDN U2266 ( .A(n3119), .B(n3121), .Z(n3122) );
  NANDN U2267 ( .A(n3123), .B(n3124), .Z(n3120) );
  NAND U2268 ( .A(n3125), .B(n3126), .Z(n3124) );
  XNOR U2269 ( .A(n3125), .B(n3127), .Z(SUM[477]) );
  NANDN U2270 ( .A(n3123), .B(n3126), .Z(n3127) );
  NANDN U2271 ( .A(n3128), .B(n3129), .Z(n3125) );
  NAND U2272 ( .A(n3130), .B(n3131), .Z(n3129) );
  XNOR U2273 ( .A(n3130), .B(n3132), .Z(SUM[476]) );
  NANDN U2274 ( .A(n3128), .B(n3131), .Z(n3132) );
  NANDN U2275 ( .A(n3133), .B(n3134), .Z(n3130) );
  NAND U2276 ( .A(n3135), .B(n3136), .Z(n3134) );
  XOR U2277 ( .A(n3137), .B(n3138), .Z(SUM[475]) );
  NANDN U2278 ( .A(n3139), .B(n3140), .Z(n3138) );
  ANDN U2279 ( .B(n3141), .A(n3142), .Z(n3137) );
  NAND U2280 ( .A(n3143), .B(n3144), .Z(n3141) );
  XNOR U2281 ( .A(n3143), .B(n3145), .Z(SUM[474]) );
  NANDN U2282 ( .A(n3142), .B(n3144), .Z(n3145) );
  NANDN U2283 ( .A(n3146), .B(n3147), .Z(n3143) );
  NAND U2284 ( .A(n3148), .B(n3149), .Z(n3147) );
  XNOR U2285 ( .A(n3148), .B(n3150), .Z(SUM[473]) );
  NANDN U2286 ( .A(n3146), .B(n3149), .Z(n3150) );
  NANDN U2287 ( .A(n3151), .B(n3152), .Z(n3148) );
  NAND U2288 ( .A(n3136), .B(n3153), .Z(n3152) );
  XNOR U2289 ( .A(n3136), .B(n3154), .Z(SUM[472]) );
  NANDN U2290 ( .A(n3151), .B(n3153), .Z(n3154) );
  NANDN U2291 ( .A(n3155), .B(n3156), .Z(n3136) );
  OR U2292 ( .A(n3157), .B(n3158), .Z(n3156) );
  XOR U2293 ( .A(n3159), .B(n3160), .Z(SUM[471]) );
  NANDN U2294 ( .A(n3161), .B(n3162), .Z(n3160) );
  ANDN U2295 ( .B(n3163), .A(n3164), .Z(n3159) );
  NAND U2296 ( .A(n3165), .B(n3166), .Z(n3163) );
  XNOR U2297 ( .A(n3165), .B(n3167), .Z(SUM[470]) );
  NANDN U2298 ( .A(n3164), .B(n3166), .Z(n3167) );
  NANDN U2299 ( .A(n3168), .B(n3169), .Z(n3165) );
  NAND U2300 ( .A(n3170), .B(n3171), .Z(n3169) );
  XNOR U2301 ( .A(n3113), .B(n3172), .Z(SUM[46]) );
  OR U2302 ( .A(n3112), .B(n3111), .Z(n3172) );
  NANDN U2303 ( .A(n3173), .B(n3174), .Z(n3113) );
  NANDN U2304 ( .A(n3175), .B(n3176), .Z(n3174) );
  XNOR U2305 ( .A(n3170), .B(n3177), .Z(SUM[469]) );
  NANDN U2306 ( .A(n3168), .B(n3171), .Z(n3177) );
  NANDN U2307 ( .A(n3178), .B(n3179), .Z(n3170) );
  NANDN U2308 ( .A(n3158), .B(n3180), .Z(n3179) );
  XOR U2309 ( .A(n3158), .B(n3181), .Z(SUM[468]) );
  NANDN U2310 ( .A(n3178), .B(n3180), .Z(n3181) );
  ANDN U2311 ( .B(n3182), .A(n3183), .Z(n3158) );
  NANDN U2312 ( .A(n3184), .B(n3105), .Z(n3182) );
  XOR U2313 ( .A(n3185), .B(n3186), .Z(SUM[467]) );
  NANDN U2314 ( .A(n3187), .B(n3188), .Z(n3186) );
  ANDN U2315 ( .B(n3189), .A(n3190), .Z(n3185) );
  NAND U2316 ( .A(n3191), .B(n3192), .Z(n3189) );
  XNOR U2317 ( .A(n3191), .B(n3193), .Z(SUM[466]) );
  NANDN U2318 ( .A(n3190), .B(n3192), .Z(n3193) );
  NANDN U2319 ( .A(n3194), .B(n3195), .Z(n3191) );
  NAND U2320 ( .A(n3196), .B(n3197), .Z(n3195) );
  XNOR U2321 ( .A(n3196), .B(n3198), .Z(SUM[465]) );
  NANDN U2322 ( .A(n3194), .B(n3197), .Z(n3198) );
  NANDN U2323 ( .A(n3199), .B(n3200), .Z(n3196) );
  NAND U2324 ( .A(n3105), .B(n3201), .Z(n3200) );
  XNOR U2325 ( .A(n3105), .B(n3202), .Z(SUM[464]) );
  NANDN U2326 ( .A(n3199), .B(n3201), .Z(n3202) );
  NANDN U2327 ( .A(n3203), .B(n3204), .Z(n3105) );
  NANDN U2328 ( .A(n3205), .B(n3206), .Z(n3204) );
  XOR U2329 ( .A(n3207), .B(n3208), .Z(SUM[463]) );
  NANDN U2330 ( .A(n3209), .B(n3210), .Z(n3208) );
  ANDN U2331 ( .B(n3211), .A(n3212), .Z(n3207) );
  NAND U2332 ( .A(n3213), .B(n3214), .Z(n3211) );
  XNOR U2333 ( .A(n3213), .B(n3215), .Z(SUM[462]) );
  NANDN U2334 ( .A(n3212), .B(n3214), .Z(n3215) );
  NANDN U2335 ( .A(n3216), .B(n3217), .Z(n3213) );
  NAND U2336 ( .A(n3218), .B(n3219), .Z(n3217) );
  XNOR U2337 ( .A(n3218), .B(n3220), .Z(SUM[461]) );
  NANDN U2338 ( .A(n3216), .B(n3219), .Z(n3220) );
  NANDN U2339 ( .A(n3221), .B(n3222), .Z(n3218) );
  NAND U2340 ( .A(n3223), .B(n3224), .Z(n3222) );
  XNOR U2341 ( .A(n3223), .B(n3225), .Z(SUM[460]) );
  NANDN U2342 ( .A(n3221), .B(n3224), .Z(n3225) );
  NANDN U2343 ( .A(n3226), .B(n3227), .Z(n3223) );
  NAND U2344 ( .A(n3228), .B(n3229), .Z(n3227) );
  XNOR U2345 ( .A(n3176), .B(n3230), .Z(SUM[45]) );
  OR U2346 ( .A(n3175), .B(n3173), .Z(n3230) );
  NANDN U2347 ( .A(n3231), .B(n3232), .Z(n3176) );
  NAND U2348 ( .A(n3233), .B(n3234), .Z(n3232) );
  XOR U2349 ( .A(n3235), .B(n3236), .Z(SUM[459]) );
  NANDN U2350 ( .A(n3237), .B(n3238), .Z(n3236) );
  ANDN U2351 ( .B(n3239), .A(n3240), .Z(n3235) );
  NAND U2352 ( .A(n3241), .B(n3242), .Z(n3239) );
  XNOR U2353 ( .A(n3241), .B(n3243), .Z(SUM[458]) );
  NANDN U2354 ( .A(n3240), .B(n3242), .Z(n3243) );
  NANDN U2355 ( .A(n3244), .B(n3245), .Z(n3241) );
  NAND U2356 ( .A(n3246), .B(n3247), .Z(n3245) );
  XNOR U2357 ( .A(n3246), .B(n3248), .Z(SUM[457]) );
  NANDN U2358 ( .A(n3244), .B(n3247), .Z(n3248) );
  NANDN U2359 ( .A(n3249), .B(n3250), .Z(n3246) );
  NAND U2360 ( .A(n3229), .B(n3251), .Z(n3250) );
  XNOR U2361 ( .A(n3229), .B(n3252), .Z(SUM[456]) );
  NANDN U2362 ( .A(n3249), .B(n3251), .Z(n3252) );
  NANDN U2363 ( .A(n3253), .B(n3254), .Z(n3229) );
  OR U2364 ( .A(n3255), .B(n3256), .Z(n3254) );
  XOR U2365 ( .A(n3257), .B(n3258), .Z(SUM[455]) );
  NANDN U2366 ( .A(n3259), .B(n3260), .Z(n3258) );
  ANDN U2367 ( .B(n3261), .A(n3262), .Z(n3257) );
  NAND U2368 ( .A(n3263), .B(n3264), .Z(n3261) );
  XNOR U2369 ( .A(n3263), .B(n3265), .Z(SUM[454]) );
  NANDN U2370 ( .A(n3262), .B(n3264), .Z(n3265) );
  NANDN U2371 ( .A(n3266), .B(n3267), .Z(n3263) );
  NAND U2372 ( .A(n3268), .B(n3269), .Z(n3267) );
  XNOR U2373 ( .A(n3268), .B(n3270), .Z(SUM[453]) );
  NANDN U2374 ( .A(n3266), .B(n3269), .Z(n3270) );
  NANDN U2375 ( .A(n3271), .B(n3272), .Z(n3268) );
  NANDN U2376 ( .A(n3256), .B(n3273), .Z(n3272) );
  XOR U2377 ( .A(n3256), .B(n3274), .Z(SUM[452]) );
  NANDN U2378 ( .A(n3271), .B(n3273), .Z(n3274) );
  ANDN U2379 ( .B(n3275), .A(n3276), .Z(n3256) );
  NANDN U2380 ( .A(n3277), .B(n3206), .Z(n3275) );
  XOR U2381 ( .A(n3278), .B(n3279), .Z(SUM[451]) );
  NANDN U2382 ( .A(n3280), .B(n3281), .Z(n3279) );
  ANDN U2383 ( .B(n3282), .A(n3283), .Z(n3278) );
  NAND U2384 ( .A(n3284), .B(n3285), .Z(n3282) );
  XNOR U2385 ( .A(n3284), .B(n3286), .Z(SUM[450]) );
  NANDN U2386 ( .A(n3283), .B(n3285), .Z(n3286) );
  NANDN U2387 ( .A(n3287), .B(n3288), .Z(n3284) );
  NAND U2388 ( .A(n3289), .B(n3290), .Z(n3288) );
  XNOR U2389 ( .A(n3233), .B(n3291), .Z(SUM[44]) );
  NANDN U2390 ( .A(n3231), .B(n3234), .Z(n3291) );
  NANDN U2391 ( .A(n3292), .B(n3293), .Z(n3233) );
  NANDN U2392 ( .A(n3294), .B(n3295), .Z(n3293) );
  XNOR U2393 ( .A(n3289), .B(n3296), .Z(SUM[449]) );
  NANDN U2394 ( .A(n3287), .B(n3290), .Z(n3296) );
  NANDN U2395 ( .A(n3297), .B(n3298), .Z(n3289) );
  NAND U2396 ( .A(n3206), .B(n3299), .Z(n3298) );
  XNOR U2397 ( .A(n3206), .B(n3300), .Z(SUM[448]) );
  NANDN U2398 ( .A(n3297), .B(n3299), .Z(n3300) );
  NANDN U2399 ( .A(n3301), .B(n3302), .Z(n3206) );
  NANDN U2400 ( .A(n3303), .B(n3304), .Z(n3302) );
  XOR U2401 ( .A(n3305), .B(n3306), .Z(SUM[447]) );
  NANDN U2402 ( .A(n3307), .B(n3308), .Z(n3306) );
  ANDN U2403 ( .B(n3309), .A(n3310), .Z(n3305) );
  NAND U2404 ( .A(n3311), .B(n3312), .Z(n3309) );
  XNOR U2405 ( .A(n3311), .B(n3313), .Z(SUM[446]) );
  NANDN U2406 ( .A(n3310), .B(n3312), .Z(n3313) );
  NANDN U2407 ( .A(n3314), .B(n3315), .Z(n3311) );
  NAND U2408 ( .A(n3316), .B(n3317), .Z(n3315) );
  XNOR U2409 ( .A(n3316), .B(n3318), .Z(SUM[445]) );
  NANDN U2410 ( .A(n3314), .B(n3317), .Z(n3318) );
  NANDN U2411 ( .A(n3319), .B(n3320), .Z(n3316) );
  NAND U2412 ( .A(n3321), .B(n3322), .Z(n3320) );
  XNOR U2413 ( .A(n3321), .B(n3323), .Z(SUM[444]) );
  NANDN U2414 ( .A(n3319), .B(n3322), .Z(n3323) );
  NANDN U2415 ( .A(n3324), .B(n3325), .Z(n3321) );
  NANDN U2416 ( .A(n3326), .B(n3327), .Z(n3325) );
  XOR U2417 ( .A(n3328), .B(n3329), .Z(SUM[443]) );
  NANDN U2418 ( .A(n3330), .B(n3331), .Z(n3329) );
  ANDN U2419 ( .B(n3332), .A(n3333), .Z(n3328) );
  NAND U2420 ( .A(n3334), .B(n3335), .Z(n3332) );
  XNOR U2421 ( .A(n3334), .B(n3336), .Z(SUM[442]) );
  NANDN U2422 ( .A(n3333), .B(n3335), .Z(n3336) );
  NANDN U2423 ( .A(n3337), .B(n3338), .Z(n3334) );
  NAND U2424 ( .A(n3339), .B(n3340), .Z(n3338) );
  XNOR U2425 ( .A(n3339), .B(n3341), .Z(SUM[441]) );
  NANDN U2426 ( .A(n3337), .B(n3340), .Z(n3341) );
  NANDN U2427 ( .A(n3342), .B(n3343), .Z(n3339) );
  NAND U2428 ( .A(n3327), .B(n3344), .Z(n3343) );
  XNOR U2429 ( .A(n3327), .B(n3345), .Z(SUM[440]) );
  NANDN U2430 ( .A(n3342), .B(n3344), .Z(n3345) );
  NANDN U2431 ( .A(n3346), .B(n3347), .Z(n3327) );
  OR U2432 ( .A(n3348), .B(n3349), .Z(n3347) );
  XOR U2433 ( .A(n3350), .B(n3351), .Z(SUM[43]) );
  NANDN U2434 ( .A(n3352), .B(n3353), .Z(n3351) );
  ANDN U2435 ( .B(n3354), .A(n3355), .Z(n3350) );
  NAND U2436 ( .A(n3356), .B(n3357), .Z(n3354) );
  XOR U2437 ( .A(n3358), .B(n3359), .Z(SUM[439]) );
  NANDN U2438 ( .A(n3360), .B(n3361), .Z(n3359) );
  ANDN U2439 ( .B(n3362), .A(n3363), .Z(n3358) );
  NAND U2440 ( .A(n3364), .B(n3365), .Z(n3362) );
  XNOR U2441 ( .A(n3364), .B(n3366), .Z(SUM[438]) );
  NANDN U2442 ( .A(n3363), .B(n3365), .Z(n3366) );
  NANDN U2443 ( .A(n3367), .B(n3368), .Z(n3364) );
  NAND U2444 ( .A(n3369), .B(n3370), .Z(n3368) );
  XNOR U2445 ( .A(n3369), .B(n3371), .Z(SUM[437]) );
  NANDN U2446 ( .A(n3367), .B(n3370), .Z(n3371) );
  NANDN U2447 ( .A(n3372), .B(n3373), .Z(n3369) );
  NANDN U2448 ( .A(n3349), .B(n3374), .Z(n3373) );
  XOR U2449 ( .A(n3349), .B(n3375), .Z(SUM[436]) );
  NANDN U2450 ( .A(n3372), .B(n3374), .Z(n3375) );
  ANDN U2451 ( .B(n3376), .A(n3377), .Z(n3349) );
  NANDN U2452 ( .A(n3378), .B(n3379), .Z(n3376) );
  XOR U2453 ( .A(n3380), .B(n3381), .Z(SUM[435]) );
  NANDN U2454 ( .A(n3382), .B(n3383), .Z(n3381) );
  ANDN U2455 ( .B(n3384), .A(n3385), .Z(n3380) );
  NAND U2456 ( .A(n3386), .B(n3387), .Z(n3384) );
  XNOR U2457 ( .A(n3386), .B(n3388), .Z(SUM[434]) );
  NANDN U2458 ( .A(n3385), .B(n3387), .Z(n3388) );
  NANDN U2459 ( .A(n3389), .B(n3390), .Z(n3386) );
  NAND U2460 ( .A(n3391), .B(n3392), .Z(n3390) );
  XNOR U2461 ( .A(n3391), .B(n3393), .Z(SUM[433]) );
  NANDN U2462 ( .A(n3389), .B(n3392), .Z(n3393) );
  NANDN U2463 ( .A(n3394), .B(n3395), .Z(n3391) );
  NAND U2464 ( .A(n3379), .B(n3396), .Z(n3395) );
  XNOR U2465 ( .A(n3379), .B(n3397), .Z(SUM[432]) );
  NANDN U2466 ( .A(n3394), .B(n3396), .Z(n3397) );
  NANDN U2467 ( .A(n3398), .B(n3399), .Z(n3379) );
  NAND U2468 ( .A(n3400), .B(n3401), .Z(n3399) );
  XOR U2469 ( .A(n3402), .B(n3403), .Z(SUM[431]) );
  NANDN U2470 ( .A(n3404), .B(n3405), .Z(n3403) );
  ANDN U2471 ( .B(n3406), .A(n3407), .Z(n3402) );
  NAND U2472 ( .A(n3408), .B(n3409), .Z(n3406) );
  XNOR U2473 ( .A(n3408), .B(n3410), .Z(SUM[430]) );
  NANDN U2474 ( .A(n3407), .B(n3409), .Z(n3410) );
  NANDN U2475 ( .A(n3411), .B(n3412), .Z(n3408) );
  NAND U2476 ( .A(n3413), .B(n3414), .Z(n3412) );
  XNOR U2477 ( .A(n3356), .B(n3415), .Z(SUM[42]) );
  NANDN U2478 ( .A(n3355), .B(n3357), .Z(n3415) );
  NANDN U2479 ( .A(n3416), .B(n3417), .Z(n3356) );
  NAND U2480 ( .A(n3418), .B(n3419), .Z(n3417) );
  XNOR U2481 ( .A(n3413), .B(n3420), .Z(SUM[429]) );
  NANDN U2482 ( .A(n3411), .B(n3414), .Z(n3420) );
  NANDN U2483 ( .A(n3421), .B(n3422), .Z(n3413) );
  NAND U2484 ( .A(n3423), .B(n3424), .Z(n3422) );
  XNOR U2485 ( .A(n3423), .B(n3425), .Z(SUM[428]) );
  NANDN U2486 ( .A(n3421), .B(n3424), .Z(n3425) );
  NANDN U2487 ( .A(n3426), .B(n3427), .Z(n3423) );
  NAND U2488 ( .A(n3428), .B(n3429), .Z(n3427) );
  XOR U2489 ( .A(n3430), .B(n3431), .Z(SUM[427]) );
  NANDN U2490 ( .A(n3432), .B(n3433), .Z(n3431) );
  ANDN U2491 ( .B(n3434), .A(n3435), .Z(n3430) );
  NAND U2492 ( .A(n3436), .B(n3437), .Z(n3434) );
  XNOR U2493 ( .A(n3436), .B(n3438), .Z(SUM[426]) );
  NANDN U2494 ( .A(n3435), .B(n3437), .Z(n3438) );
  NANDN U2495 ( .A(n3439), .B(n3440), .Z(n3436) );
  NAND U2496 ( .A(n3441), .B(n3442), .Z(n3440) );
  XNOR U2497 ( .A(n3441), .B(n3443), .Z(SUM[425]) );
  NANDN U2498 ( .A(n3439), .B(n3442), .Z(n3443) );
  NANDN U2499 ( .A(n3444), .B(n3445), .Z(n3441) );
  NAND U2500 ( .A(n3429), .B(n3446), .Z(n3445) );
  XNOR U2501 ( .A(n3429), .B(n3447), .Z(SUM[424]) );
  NANDN U2502 ( .A(n3444), .B(n3446), .Z(n3447) );
  NANDN U2503 ( .A(n3448), .B(n3449), .Z(n3429) );
  OR U2504 ( .A(n3450), .B(n3451), .Z(n3449) );
  XOR U2505 ( .A(n3452), .B(n3453), .Z(SUM[423]) );
  NANDN U2506 ( .A(n3454), .B(n3455), .Z(n3453) );
  ANDN U2507 ( .B(n3456), .A(n3457), .Z(n3452) );
  NAND U2508 ( .A(n3458), .B(n3459), .Z(n3456) );
  XNOR U2509 ( .A(n3458), .B(n3460), .Z(SUM[422]) );
  NANDN U2510 ( .A(n3457), .B(n3459), .Z(n3460) );
  NANDN U2511 ( .A(n3461), .B(n3462), .Z(n3458) );
  NAND U2512 ( .A(n3463), .B(n3464), .Z(n3462) );
  XNOR U2513 ( .A(n3463), .B(n3465), .Z(SUM[421]) );
  NANDN U2514 ( .A(n3461), .B(n3464), .Z(n3465) );
  NANDN U2515 ( .A(n3466), .B(n3467), .Z(n3463) );
  NANDN U2516 ( .A(n3451), .B(n3468), .Z(n3467) );
  XOR U2517 ( .A(n3451), .B(n3469), .Z(SUM[420]) );
  NANDN U2518 ( .A(n3466), .B(n3468), .Z(n3469) );
  ANDN U2519 ( .B(n3470), .A(n3471), .Z(n3451) );
  NANDN U2520 ( .A(n3472), .B(n3401), .Z(n3470) );
  XNOR U2521 ( .A(n3418), .B(n3473), .Z(SUM[41]) );
  NANDN U2522 ( .A(n3416), .B(n3419), .Z(n3473) );
  NANDN U2523 ( .A(n3474), .B(n3475), .Z(n3418) );
  NAND U2524 ( .A(n3295), .B(n3476), .Z(n3475) );
  XOR U2525 ( .A(n3477), .B(n3478), .Z(SUM[419]) );
  NANDN U2526 ( .A(n3479), .B(n3480), .Z(n3478) );
  ANDN U2527 ( .B(n3481), .A(n3482), .Z(n3477) );
  NAND U2528 ( .A(n3483), .B(n3484), .Z(n3481) );
  XNOR U2529 ( .A(n3483), .B(n3485), .Z(SUM[418]) );
  NANDN U2530 ( .A(n3482), .B(n3484), .Z(n3485) );
  NANDN U2531 ( .A(n3486), .B(n3487), .Z(n3483) );
  NAND U2532 ( .A(n3488), .B(n3489), .Z(n3487) );
  XNOR U2533 ( .A(n3488), .B(n3490), .Z(SUM[417]) );
  NANDN U2534 ( .A(n3486), .B(n3489), .Z(n3490) );
  NANDN U2535 ( .A(n3491), .B(n3492), .Z(n3488) );
  NAND U2536 ( .A(n3401), .B(n3493), .Z(n3492) );
  XNOR U2537 ( .A(n3401), .B(n3494), .Z(SUM[416]) );
  NANDN U2538 ( .A(n3491), .B(n3493), .Z(n3494) );
  NANDN U2539 ( .A(n3495), .B(n3496), .Z(n3401) );
  OR U2540 ( .A(n3497), .B(n3498), .Z(n3496) );
  XOR U2541 ( .A(n3499), .B(n3500), .Z(SUM[415]) );
  NANDN U2542 ( .A(n3501), .B(n3502), .Z(n3500) );
  ANDN U2543 ( .B(n3503), .A(n3504), .Z(n3499) );
  NAND U2544 ( .A(n3505), .B(n3506), .Z(n3503) );
  XNOR U2545 ( .A(n3505), .B(n3507), .Z(SUM[414]) );
  NANDN U2546 ( .A(n3504), .B(n3506), .Z(n3507) );
  NANDN U2547 ( .A(n3508), .B(n3509), .Z(n3505) );
  NAND U2548 ( .A(n3510), .B(n3511), .Z(n3509) );
  XNOR U2549 ( .A(n3510), .B(n3512), .Z(SUM[413]) );
  NANDN U2550 ( .A(n3508), .B(n3511), .Z(n3512) );
  NANDN U2551 ( .A(n3513), .B(n3514), .Z(n3510) );
  NAND U2552 ( .A(n3515), .B(n3516), .Z(n3514) );
  XNOR U2553 ( .A(n3515), .B(n3517), .Z(SUM[412]) );
  NANDN U2554 ( .A(n3513), .B(n3516), .Z(n3517) );
  NANDN U2555 ( .A(n3518), .B(n3519), .Z(n3515) );
  NAND U2556 ( .A(n3520), .B(n3521), .Z(n3519) );
  XOR U2557 ( .A(n3522), .B(n3523), .Z(SUM[411]) );
  NANDN U2558 ( .A(n3524), .B(n3525), .Z(n3523) );
  ANDN U2559 ( .B(n3526), .A(n3527), .Z(n3522) );
  NAND U2560 ( .A(n3528), .B(n3529), .Z(n3526) );
  XNOR U2561 ( .A(n3528), .B(n3530), .Z(SUM[410]) );
  NANDN U2562 ( .A(n3527), .B(n3529), .Z(n3530) );
  NANDN U2563 ( .A(n3531), .B(n3532), .Z(n3528) );
  NAND U2564 ( .A(n3533), .B(n3534), .Z(n3532) );
  XNOR U2565 ( .A(n3295), .B(n3535), .Z(SUM[40]) );
  NANDN U2566 ( .A(n3474), .B(n3476), .Z(n3535) );
  NANDN U2567 ( .A(n3536), .B(n3537), .Z(n3295) );
  NANDN U2568 ( .A(n3538), .B(n3539), .Z(n3537) );
  XNOR U2569 ( .A(n3533), .B(n3540), .Z(SUM[409]) );
  NANDN U2570 ( .A(n3531), .B(n3534), .Z(n3540) );
  NANDN U2571 ( .A(n3541), .B(n3542), .Z(n3533) );
  NAND U2572 ( .A(n3521), .B(n3543), .Z(n3542) );
  XNOR U2573 ( .A(n3521), .B(n3544), .Z(SUM[408]) );
  NANDN U2574 ( .A(n3541), .B(n3543), .Z(n3544) );
  NANDN U2575 ( .A(n3545), .B(n3546), .Z(n3521) );
  OR U2576 ( .A(n3547), .B(n3548), .Z(n3546) );
  XOR U2577 ( .A(n3549), .B(n3550), .Z(SUM[407]) );
  NANDN U2578 ( .A(n3551), .B(n3552), .Z(n3550) );
  ANDN U2579 ( .B(n3553), .A(n3554), .Z(n3549) );
  NAND U2580 ( .A(n3555), .B(n3556), .Z(n3553) );
  XNOR U2581 ( .A(n3555), .B(n3557), .Z(SUM[406]) );
  NANDN U2582 ( .A(n3554), .B(n3556), .Z(n3557) );
  NANDN U2583 ( .A(n3558), .B(n3559), .Z(n3555) );
  NAND U2584 ( .A(n3560), .B(n3561), .Z(n3559) );
  XNOR U2585 ( .A(n3560), .B(n3562), .Z(SUM[405]) );
  NANDN U2586 ( .A(n3558), .B(n3561), .Z(n3562) );
  NANDN U2587 ( .A(n3563), .B(n3564), .Z(n3560) );
  NANDN U2588 ( .A(n3548), .B(n3565), .Z(n3564) );
  XOR U2589 ( .A(n3548), .B(n3566), .Z(SUM[404]) );
  NANDN U2590 ( .A(n3563), .B(n3565), .Z(n3566) );
  ANDN U2591 ( .B(n3567), .A(n3568), .Z(n3548) );
  OR U2592 ( .A(n3569), .B(n3498), .Z(n3567) );
  XOR U2593 ( .A(n3570), .B(n3571), .Z(SUM[403]) );
  NANDN U2594 ( .A(n3572), .B(n3573), .Z(n3571) );
  ANDN U2595 ( .B(n3574), .A(n3575), .Z(n3570) );
  NAND U2596 ( .A(n3576), .B(n3577), .Z(n3574) );
  XNOR U2597 ( .A(n3576), .B(n3578), .Z(SUM[402]) );
  NANDN U2598 ( .A(n3575), .B(n3577), .Z(n3578) );
  NANDN U2599 ( .A(n3579), .B(n3580), .Z(n3576) );
  NAND U2600 ( .A(n3581), .B(n3582), .Z(n3580) );
  XNOR U2601 ( .A(n3581), .B(n3583), .Z(SUM[401]) );
  NANDN U2602 ( .A(n3579), .B(n3582), .Z(n3583) );
  NANDN U2603 ( .A(n3584), .B(n3585), .Z(n3581) );
  NANDN U2604 ( .A(n3498), .B(n3586), .Z(n3585) );
  XOR U2605 ( .A(n3498), .B(n3587), .Z(SUM[400]) );
  NANDN U2606 ( .A(n3584), .B(n3586), .Z(n3587) );
  ANDN U2607 ( .B(n3588), .A(n3589), .Z(n3498) );
  NANDN U2608 ( .A(n3590), .B(n3304), .Z(n3588) );
  XOR U2609 ( .A(n3591), .B(n3592), .Z(SUM[3]) );
  XNOR U2610 ( .A(B[3]), .B(A[3]), .Z(n3592) );
  XOR U2611 ( .A(n3593), .B(n3594), .Z(SUM[39]) );
  NANDN U2612 ( .A(n3595), .B(n3596), .Z(n3594) );
  ANDN U2613 ( .B(n3597), .A(n3598), .Z(n3593) );
  NAND U2614 ( .A(n3599), .B(n3600), .Z(n3597) );
  XOR U2615 ( .A(n3601), .B(n3602), .Z(SUM[399]) );
  NANDN U2616 ( .A(n3603), .B(n3604), .Z(n3602) );
  ANDN U2617 ( .B(n3605), .A(n3606), .Z(n3601) );
  NAND U2618 ( .A(n3607), .B(n3608), .Z(n3605) );
  XNOR U2619 ( .A(n3607), .B(n3609), .Z(SUM[398]) );
  NANDN U2620 ( .A(n3606), .B(n3608), .Z(n3609) );
  NANDN U2621 ( .A(n3610), .B(n3611), .Z(n3607) );
  NAND U2622 ( .A(n3612), .B(n3613), .Z(n3611) );
  XNOR U2623 ( .A(n3612), .B(n3614), .Z(SUM[397]) );
  NANDN U2624 ( .A(n3610), .B(n3613), .Z(n3614) );
  NANDN U2625 ( .A(n3615), .B(n3616), .Z(n3612) );
  NAND U2626 ( .A(n3617), .B(n3618), .Z(n3616) );
  XNOR U2627 ( .A(n3617), .B(n3619), .Z(SUM[396]) );
  NANDN U2628 ( .A(n3615), .B(n3618), .Z(n3619) );
  NANDN U2629 ( .A(n3620), .B(n3621), .Z(n3617) );
  NAND U2630 ( .A(n3622), .B(n3623), .Z(n3621) );
  XOR U2631 ( .A(n3624), .B(n3625), .Z(SUM[395]) );
  NANDN U2632 ( .A(n3626), .B(n3627), .Z(n3625) );
  ANDN U2633 ( .B(n3628), .A(n3629), .Z(n3624) );
  NAND U2634 ( .A(n3630), .B(n3631), .Z(n3628) );
  XNOR U2635 ( .A(n3630), .B(n3632), .Z(SUM[394]) );
  NANDN U2636 ( .A(n3629), .B(n3631), .Z(n3632) );
  NANDN U2637 ( .A(n3633), .B(n3634), .Z(n3630) );
  NAND U2638 ( .A(n3635), .B(n3636), .Z(n3634) );
  XNOR U2639 ( .A(n3635), .B(n3637), .Z(SUM[393]) );
  NANDN U2640 ( .A(n3633), .B(n3636), .Z(n3637) );
  NANDN U2641 ( .A(n3638), .B(n3639), .Z(n3635) );
  NAND U2642 ( .A(n3623), .B(n3640), .Z(n3639) );
  XNOR U2643 ( .A(n3623), .B(n3641), .Z(SUM[392]) );
  NANDN U2644 ( .A(n3638), .B(n3640), .Z(n3641) );
  NANDN U2645 ( .A(n3642), .B(n3643), .Z(n3623) );
  OR U2646 ( .A(n3644), .B(n3645), .Z(n3643) );
  XOR U2647 ( .A(n3646), .B(n3647), .Z(SUM[391]) );
  NANDN U2648 ( .A(n3648), .B(n3649), .Z(n3647) );
  ANDN U2649 ( .B(n3650), .A(n3651), .Z(n3646) );
  NAND U2650 ( .A(n3652), .B(n3653), .Z(n3650) );
  XNOR U2651 ( .A(n3652), .B(n3654), .Z(SUM[390]) );
  NANDN U2652 ( .A(n3651), .B(n3653), .Z(n3654) );
  NANDN U2653 ( .A(n3655), .B(n3656), .Z(n3652) );
  NAND U2654 ( .A(n3657), .B(n3658), .Z(n3656) );
  XNOR U2655 ( .A(n3599), .B(n3659), .Z(SUM[38]) );
  NANDN U2656 ( .A(n3598), .B(n3600), .Z(n3659) );
  NANDN U2657 ( .A(n3660), .B(n3661), .Z(n3599) );
  NAND U2658 ( .A(n3662), .B(n3663), .Z(n3661) );
  XNOR U2659 ( .A(n3657), .B(n3664), .Z(SUM[389]) );
  NANDN U2660 ( .A(n3655), .B(n3658), .Z(n3664) );
  NANDN U2661 ( .A(n3665), .B(n3666), .Z(n3657) );
  NANDN U2662 ( .A(n3645), .B(n3667), .Z(n3666) );
  XOR U2663 ( .A(n3645), .B(n3668), .Z(SUM[388]) );
  NANDN U2664 ( .A(n3665), .B(n3667), .Z(n3668) );
  ANDN U2665 ( .B(n3669), .A(n3670), .Z(n3645) );
  NANDN U2666 ( .A(n3671), .B(n3304), .Z(n3669) );
  XOR U2667 ( .A(n3672), .B(n3673), .Z(SUM[387]) );
  NANDN U2668 ( .A(n3674), .B(n3675), .Z(n3673) );
  ANDN U2669 ( .B(n3676), .A(n3677), .Z(n3672) );
  NAND U2670 ( .A(n3678), .B(n3679), .Z(n3676) );
  XNOR U2671 ( .A(n3678), .B(n3680), .Z(SUM[386]) );
  NANDN U2672 ( .A(n3677), .B(n3679), .Z(n3680) );
  NANDN U2673 ( .A(n3681), .B(n3682), .Z(n3678) );
  NAND U2674 ( .A(n3683), .B(n3684), .Z(n3682) );
  XNOR U2675 ( .A(n3683), .B(n3685), .Z(SUM[385]) );
  NANDN U2676 ( .A(n3681), .B(n3684), .Z(n3685) );
  NANDN U2677 ( .A(n3686), .B(n3687), .Z(n3683) );
  NAND U2678 ( .A(n3304), .B(n3688), .Z(n3687) );
  XNOR U2679 ( .A(n3304), .B(n3689), .Z(SUM[384]) );
  NANDN U2680 ( .A(n3686), .B(n3688), .Z(n3689) );
  NANDN U2681 ( .A(n3690), .B(n3691), .Z(n3304) );
  OR U2682 ( .A(n3692), .B(n3693), .Z(n3691) );
  XOR U2683 ( .A(n3694), .B(n3695), .Z(SUM[383]) );
  NANDN U2684 ( .A(n3696), .B(n3697), .Z(n3695) );
  ANDN U2685 ( .B(n3698), .A(n3699), .Z(n3694) );
  NAND U2686 ( .A(n3700), .B(n3701), .Z(n3698) );
  XNOR U2687 ( .A(n3700), .B(n3702), .Z(SUM[382]) );
  NANDN U2688 ( .A(n3699), .B(n3701), .Z(n3702) );
  NANDN U2689 ( .A(n3703), .B(n3704), .Z(n3700) );
  NAND U2690 ( .A(n3705), .B(n3706), .Z(n3704) );
  XNOR U2691 ( .A(n3705), .B(n3707), .Z(SUM[381]) );
  NANDN U2692 ( .A(n3703), .B(n3706), .Z(n3707) );
  NANDN U2693 ( .A(n3708), .B(n3709), .Z(n3705) );
  NAND U2694 ( .A(n3710), .B(n3711), .Z(n3709) );
  XNOR U2695 ( .A(n3710), .B(n3712), .Z(SUM[380]) );
  NANDN U2696 ( .A(n3708), .B(n3711), .Z(n3712) );
  NANDN U2697 ( .A(n3713), .B(n3714), .Z(n3710) );
  NANDN U2698 ( .A(n3715), .B(n3716), .Z(n3714) );
  XNOR U2699 ( .A(n3662), .B(n3717), .Z(SUM[37]) );
  NANDN U2700 ( .A(n3660), .B(n3663), .Z(n3717) );
  NANDN U2701 ( .A(n3718), .B(n3719), .Z(n3662) );
  NANDN U2702 ( .A(n3538), .B(n3720), .Z(n3719) );
  XOR U2703 ( .A(n3721), .B(n3722), .Z(SUM[379]) );
  NANDN U2704 ( .A(n3723), .B(n3724), .Z(n3722) );
  ANDN U2705 ( .B(n3725), .A(n3726), .Z(n3721) );
  NAND U2706 ( .A(n3727), .B(n3728), .Z(n3725) );
  XNOR U2707 ( .A(n3727), .B(n3729), .Z(SUM[378]) );
  NANDN U2708 ( .A(n3726), .B(n3728), .Z(n3729) );
  NANDN U2709 ( .A(n3730), .B(n3731), .Z(n3727) );
  NAND U2710 ( .A(n3732), .B(n3733), .Z(n3731) );
  XNOR U2711 ( .A(n3732), .B(n3734), .Z(SUM[377]) );
  NANDN U2712 ( .A(n3730), .B(n3733), .Z(n3734) );
  NANDN U2713 ( .A(n3735), .B(n3736), .Z(n3732) );
  NAND U2714 ( .A(n3716), .B(n3737), .Z(n3736) );
  XNOR U2715 ( .A(n3716), .B(n3738), .Z(SUM[376]) );
  NANDN U2716 ( .A(n3735), .B(n3737), .Z(n3738) );
  NANDN U2717 ( .A(n3739), .B(n3740), .Z(n3716) );
  OR U2718 ( .A(n3741), .B(n3742), .Z(n3740) );
  XOR U2719 ( .A(n3743), .B(n3744), .Z(SUM[375]) );
  NANDN U2720 ( .A(n3745), .B(n3746), .Z(n3744) );
  ANDN U2721 ( .B(n3747), .A(n3748), .Z(n3743) );
  NAND U2722 ( .A(n3749), .B(n3750), .Z(n3747) );
  XNOR U2723 ( .A(n3749), .B(n3751), .Z(SUM[374]) );
  NANDN U2724 ( .A(n3748), .B(n3750), .Z(n3751) );
  NANDN U2725 ( .A(n3752), .B(n3753), .Z(n3749) );
  NAND U2726 ( .A(n3754), .B(n3755), .Z(n3753) );
  XNOR U2727 ( .A(n3754), .B(n3756), .Z(SUM[373]) );
  NANDN U2728 ( .A(n3752), .B(n3755), .Z(n3756) );
  NANDN U2729 ( .A(n3757), .B(n3758), .Z(n3754) );
  NANDN U2730 ( .A(n3742), .B(n3759), .Z(n3758) );
  XOR U2731 ( .A(n3742), .B(n3760), .Z(SUM[372]) );
  NANDN U2732 ( .A(n3757), .B(n3759), .Z(n3760) );
  ANDN U2733 ( .B(n3761), .A(n3762), .Z(n3742) );
  NANDN U2734 ( .A(n3763), .B(n3764), .Z(n3761) );
  XOR U2735 ( .A(n3765), .B(n3766), .Z(SUM[371]) );
  NANDN U2736 ( .A(n3767), .B(n3768), .Z(n3766) );
  ANDN U2737 ( .B(n3769), .A(n3770), .Z(n3765) );
  NAND U2738 ( .A(n3771), .B(n3772), .Z(n3769) );
  XNOR U2739 ( .A(n3771), .B(n3773), .Z(SUM[370]) );
  NANDN U2740 ( .A(n3770), .B(n3772), .Z(n3773) );
  NANDN U2741 ( .A(n3774), .B(n3775), .Z(n3771) );
  NAND U2742 ( .A(n3776), .B(n3777), .Z(n3775) );
  XOR U2743 ( .A(n3538), .B(n3778), .Z(SUM[36]) );
  NANDN U2744 ( .A(n3718), .B(n3720), .Z(n3778) );
  ANDN U2745 ( .B(n3779), .A(n3780), .Z(n3538) );
  OR U2746 ( .A(n3781), .B(n3782), .Z(n3779) );
  XNOR U2747 ( .A(n3776), .B(n3783), .Z(SUM[369]) );
  NANDN U2748 ( .A(n3774), .B(n3777), .Z(n3783) );
  NANDN U2749 ( .A(n3784), .B(n3785), .Z(n3776) );
  NAND U2750 ( .A(n3764), .B(n3786), .Z(n3785) );
  XNOR U2751 ( .A(n3764), .B(n3787), .Z(SUM[368]) );
  NANDN U2752 ( .A(n3784), .B(n3786), .Z(n3787) );
  NANDN U2753 ( .A(n3788), .B(n3789), .Z(n3764) );
  NANDN U2754 ( .A(n3790), .B(n3791), .Z(n3789) );
  XOR U2755 ( .A(n3792), .B(n3793), .Z(SUM[367]) );
  NANDN U2756 ( .A(n3794), .B(n3795), .Z(n3793) );
  ANDN U2757 ( .B(n3796), .A(n3797), .Z(n3792) );
  NAND U2758 ( .A(n3798), .B(n3799), .Z(n3796) );
  XNOR U2759 ( .A(n3798), .B(n3800), .Z(SUM[366]) );
  NANDN U2760 ( .A(n3797), .B(n3799), .Z(n3800) );
  NANDN U2761 ( .A(n3801), .B(n3802), .Z(n3798) );
  NAND U2762 ( .A(n3803), .B(n3804), .Z(n3802) );
  XNOR U2763 ( .A(n3803), .B(n3805), .Z(SUM[365]) );
  NANDN U2764 ( .A(n3801), .B(n3804), .Z(n3805) );
  NANDN U2765 ( .A(n3806), .B(n3807), .Z(n3803) );
  NAND U2766 ( .A(n3808), .B(n3809), .Z(n3807) );
  XNOR U2767 ( .A(n3808), .B(n3810), .Z(SUM[364]) );
  NANDN U2768 ( .A(n3806), .B(n3809), .Z(n3810) );
  NANDN U2769 ( .A(n3811), .B(n3812), .Z(n3808) );
  NANDN U2770 ( .A(n3813), .B(n3814), .Z(n3812) );
  XOR U2771 ( .A(n3815), .B(n3816), .Z(SUM[363]) );
  NANDN U2772 ( .A(n3817), .B(n3818), .Z(n3816) );
  ANDN U2773 ( .B(n3819), .A(n3820), .Z(n3815) );
  NAND U2774 ( .A(n3821), .B(n3822), .Z(n3819) );
  XNOR U2775 ( .A(n3821), .B(n3823), .Z(SUM[362]) );
  NANDN U2776 ( .A(n3820), .B(n3822), .Z(n3823) );
  NANDN U2777 ( .A(n3824), .B(n3825), .Z(n3821) );
  NAND U2778 ( .A(n3826), .B(n3827), .Z(n3825) );
  XNOR U2779 ( .A(n3826), .B(n3828), .Z(SUM[361]) );
  NANDN U2780 ( .A(n3824), .B(n3827), .Z(n3828) );
  NANDN U2781 ( .A(n3829), .B(n3830), .Z(n3826) );
  NAND U2782 ( .A(n3814), .B(n3831), .Z(n3830) );
  XNOR U2783 ( .A(n3814), .B(n3832), .Z(SUM[360]) );
  NANDN U2784 ( .A(n3829), .B(n3831), .Z(n3832) );
  NANDN U2785 ( .A(n3833), .B(n3834), .Z(n3814) );
  OR U2786 ( .A(n3835), .B(n3836), .Z(n3834) );
  XOR U2787 ( .A(n3837), .B(n3838), .Z(SUM[35]) );
  NANDN U2788 ( .A(n3839), .B(n3840), .Z(n3838) );
  ANDN U2789 ( .B(n3841), .A(n3842), .Z(n3837) );
  NANDN U2790 ( .A(n3843), .B(n3844), .Z(n3841) );
  XOR U2791 ( .A(n3845), .B(n3846), .Z(SUM[359]) );
  NANDN U2792 ( .A(n3847), .B(n3848), .Z(n3846) );
  ANDN U2793 ( .B(n3849), .A(n3850), .Z(n3845) );
  NAND U2794 ( .A(n3851), .B(n3852), .Z(n3849) );
  XNOR U2795 ( .A(n3851), .B(n3853), .Z(SUM[358]) );
  NANDN U2796 ( .A(n3850), .B(n3852), .Z(n3853) );
  NANDN U2797 ( .A(n3854), .B(n3855), .Z(n3851) );
  NAND U2798 ( .A(n3856), .B(n3857), .Z(n3855) );
  XNOR U2799 ( .A(n3856), .B(n3858), .Z(SUM[357]) );
  NANDN U2800 ( .A(n3854), .B(n3857), .Z(n3858) );
  NANDN U2801 ( .A(n3859), .B(n3860), .Z(n3856) );
  NANDN U2802 ( .A(n3836), .B(n3861), .Z(n3860) );
  XOR U2803 ( .A(n3836), .B(n3862), .Z(SUM[356]) );
  NANDN U2804 ( .A(n3859), .B(n3861), .Z(n3862) );
  ANDN U2805 ( .B(n3863), .A(n3864), .Z(n3836) );
  NANDN U2806 ( .A(n3865), .B(n3791), .Z(n3863) );
  XOR U2807 ( .A(n3866), .B(n3867), .Z(SUM[355]) );
  NANDN U2808 ( .A(n3868), .B(n3869), .Z(n3867) );
  ANDN U2809 ( .B(n3870), .A(n3871), .Z(n3866) );
  NAND U2810 ( .A(n3872), .B(n3873), .Z(n3870) );
  XNOR U2811 ( .A(n3872), .B(n3874), .Z(SUM[354]) );
  NANDN U2812 ( .A(n3871), .B(n3873), .Z(n3874) );
  NANDN U2813 ( .A(n3875), .B(n3876), .Z(n3872) );
  NAND U2814 ( .A(n3877), .B(n3878), .Z(n3876) );
  XNOR U2815 ( .A(n3877), .B(n3879), .Z(SUM[353]) );
  NANDN U2816 ( .A(n3875), .B(n3878), .Z(n3879) );
  NANDN U2817 ( .A(n3880), .B(n3881), .Z(n3877) );
  NAND U2818 ( .A(n3791), .B(n3882), .Z(n3881) );
  XNOR U2819 ( .A(n3791), .B(n3883), .Z(SUM[352]) );
  NANDN U2820 ( .A(n3880), .B(n3882), .Z(n3883) );
  NANDN U2821 ( .A(n3884), .B(n3885), .Z(n3791) );
  OR U2822 ( .A(n3886), .B(n3887), .Z(n3885) );
  XOR U2823 ( .A(n3888), .B(n3889), .Z(SUM[351]) );
  NANDN U2824 ( .A(n3890), .B(n3891), .Z(n3889) );
  ANDN U2825 ( .B(n3892), .A(n3893), .Z(n3888) );
  NAND U2826 ( .A(n3894), .B(n3895), .Z(n3892) );
  XNOR U2827 ( .A(n3894), .B(n3896), .Z(SUM[350]) );
  NANDN U2828 ( .A(n3893), .B(n3895), .Z(n3896) );
  NANDN U2829 ( .A(n3897), .B(n3898), .Z(n3894) );
  NAND U2830 ( .A(n3899), .B(n3900), .Z(n3898) );
  XNOR U2831 ( .A(n3844), .B(n3901), .Z(SUM[34]) );
  OR U2832 ( .A(n3843), .B(n3842), .Z(n3901) );
  NANDN U2833 ( .A(n3902), .B(n3903), .Z(n3844) );
  NAND U2834 ( .A(n3904), .B(n3905), .Z(n3903) );
  XNOR U2835 ( .A(n3899), .B(n3906), .Z(SUM[349]) );
  NANDN U2836 ( .A(n3897), .B(n3900), .Z(n3906) );
  NANDN U2837 ( .A(n3907), .B(n3908), .Z(n3899) );
  NAND U2838 ( .A(n3909), .B(n3910), .Z(n3908) );
  XNOR U2839 ( .A(n3909), .B(n3911), .Z(SUM[348]) );
  NANDN U2840 ( .A(n3907), .B(n3910), .Z(n3911) );
  NANDN U2841 ( .A(n3912), .B(n3913), .Z(n3909) );
  NANDN U2842 ( .A(n3914), .B(n3915), .Z(n3913) );
  XOR U2843 ( .A(n3916), .B(n3917), .Z(SUM[347]) );
  NANDN U2844 ( .A(n3918), .B(n3919), .Z(n3917) );
  ANDN U2845 ( .B(n3920), .A(n3921), .Z(n3916) );
  NAND U2846 ( .A(n3922), .B(n3923), .Z(n3920) );
  XNOR U2847 ( .A(n3922), .B(n3924), .Z(SUM[346]) );
  NANDN U2848 ( .A(n3921), .B(n3923), .Z(n3924) );
  NANDN U2849 ( .A(n3925), .B(n3926), .Z(n3922) );
  NAND U2850 ( .A(n3927), .B(n3928), .Z(n3926) );
  XNOR U2851 ( .A(n3927), .B(n3929), .Z(SUM[345]) );
  NANDN U2852 ( .A(n3925), .B(n3928), .Z(n3929) );
  NANDN U2853 ( .A(n3930), .B(n3931), .Z(n3927) );
  NAND U2854 ( .A(n3915), .B(n3932), .Z(n3931) );
  XNOR U2855 ( .A(n3915), .B(n3933), .Z(SUM[344]) );
  NANDN U2856 ( .A(n3930), .B(n3932), .Z(n3933) );
  NANDN U2857 ( .A(n3934), .B(n3935), .Z(n3915) );
  OR U2858 ( .A(n3936), .B(n3937), .Z(n3935) );
  XOR U2859 ( .A(n3938), .B(n3939), .Z(SUM[343]) );
  NANDN U2860 ( .A(n3940), .B(n3941), .Z(n3939) );
  ANDN U2861 ( .B(n3942), .A(n3943), .Z(n3938) );
  NAND U2862 ( .A(n3944), .B(n3945), .Z(n3942) );
  XNOR U2863 ( .A(n3944), .B(n3946), .Z(SUM[342]) );
  NANDN U2864 ( .A(n3943), .B(n3945), .Z(n3946) );
  NANDN U2865 ( .A(n3947), .B(n3948), .Z(n3944) );
  NAND U2866 ( .A(n3949), .B(n3950), .Z(n3948) );
  XNOR U2867 ( .A(n3949), .B(n3951), .Z(SUM[341]) );
  NANDN U2868 ( .A(n3947), .B(n3950), .Z(n3951) );
  NANDN U2869 ( .A(n3952), .B(n3953), .Z(n3949) );
  NANDN U2870 ( .A(n3937), .B(n3954), .Z(n3953) );
  XOR U2871 ( .A(n3937), .B(n3955), .Z(SUM[340]) );
  NANDN U2872 ( .A(n3952), .B(n3954), .Z(n3955) );
  ANDN U2873 ( .B(n3956), .A(n3957), .Z(n3937) );
  OR U2874 ( .A(n3958), .B(n3887), .Z(n3956) );
  XNOR U2875 ( .A(n3904), .B(n3959), .Z(SUM[33]) );
  NANDN U2876 ( .A(n3902), .B(n3905), .Z(n3959) );
  NANDN U2877 ( .A(n3960), .B(n3961), .Z(n3904) );
  NANDN U2878 ( .A(n3782), .B(n3962), .Z(n3961) );
  XOR U2879 ( .A(n3963), .B(n3964), .Z(SUM[339]) );
  NANDN U2880 ( .A(n3965), .B(n3966), .Z(n3964) );
  ANDN U2881 ( .B(n3967), .A(n3968), .Z(n3963) );
  NAND U2882 ( .A(n3969), .B(n3970), .Z(n3967) );
  XNOR U2883 ( .A(n3969), .B(n3971), .Z(SUM[338]) );
  NANDN U2884 ( .A(n3968), .B(n3970), .Z(n3971) );
  NANDN U2885 ( .A(n3972), .B(n3973), .Z(n3969) );
  NAND U2886 ( .A(n3974), .B(n3975), .Z(n3973) );
  XNOR U2887 ( .A(n3974), .B(n3976), .Z(SUM[337]) );
  NANDN U2888 ( .A(n3972), .B(n3975), .Z(n3976) );
  NANDN U2889 ( .A(n3977), .B(n3978), .Z(n3974) );
  NANDN U2890 ( .A(n3887), .B(n3979), .Z(n3978) );
  XOR U2891 ( .A(n3887), .B(n3980), .Z(SUM[336]) );
  NANDN U2892 ( .A(n3977), .B(n3979), .Z(n3980) );
  ANDN U2893 ( .B(n3981), .A(n3982), .Z(n3887) );
  OR U2894 ( .A(n3983), .B(n3693), .Z(n3981) );
  XOR U2895 ( .A(n3984), .B(n3985), .Z(SUM[335]) );
  NANDN U2896 ( .A(n3986), .B(n3987), .Z(n3985) );
  ANDN U2897 ( .B(n3988), .A(n3989), .Z(n3984) );
  NAND U2898 ( .A(n3990), .B(n3991), .Z(n3988) );
  XNOR U2899 ( .A(n3990), .B(n3992), .Z(SUM[334]) );
  NANDN U2900 ( .A(n3989), .B(n3991), .Z(n3992) );
  NANDN U2901 ( .A(n3993), .B(n3994), .Z(n3990) );
  NAND U2902 ( .A(n3995), .B(n3996), .Z(n3994) );
  XNOR U2903 ( .A(n3995), .B(n3997), .Z(SUM[333]) );
  NANDN U2904 ( .A(n3993), .B(n3996), .Z(n3997) );
  NANDN U2905 ( .A(n3998), .B(n3999), .Z(n3995) );
  NAND U2906 ( .A(n4000), .B(n4001), .Z(n3999) );
  XNOR U2907 ( .A(n4000), .B(n4002), .Z(SUM[332]) );
  NANDN U2908 ( .A(n3998), .B(n4001), .Z(n4002) );
  NANDN U2909 ( .A(n4003), .B(n4004), .Z(n4000) );
  NANDN U2910 ( .A(n4005), .B(n4006), .Z(n4004) );
  XOR U2911 ( .A(n4007), .B(n4008), .Z(SUM[331]) );
  NANDN U2912 ( .A(n4009), .B(n4010), .Z(n4008) );
  ANDN U2913 ( .B(n4011), .A(n4012), .Z(n4007) );
  NAND U2914 ( .A(n4013), .B(n4014), .Z(n4011) );
  XNOR U2915 ( .A(n4013), .B(n4015), .Z(SUM[330]) );
  NANDN U2916 ( .A(n4012), .B(n4014), .Z(n4015) );
  NANDN U2917 ( .A(n4016), .B(n4017), .Z(n4013) );
  NAND U2918 ( .A(n4018), .B(n4019), .Z(n4017) );
  XOR U2919 ( .A(n3782), .B(n4020), .Z(SUM[32]) );
  NANDN U2920 ( .A(n3960), .B(n3962), .Z(n4020) );
  XNOR U2921 ( .A(n4018), .B(n4021), .Z(SUM[329]) );
  NANDN U2922 ( .A(n4016), .B(n4019), .Z(n4021) );
  NANDN U2923 ( .A(n4022), .B(n4023), .Z(n4018) );
  NAND U2924 ( .A(n4006), .B(n4024), .Z(n4023) );
  XNOR U2925 ( .A(n4006), .B(n4025), .Z(SUM[328]) );
  NANDN U2926 ( .A(n4022), .B(n4024), .Z(n4025) );
  NANDN U2927 ( .A(n4026), .B(n4027), .Z(n4006) );
  OR U2928 ( .A(n4028), .B(n4029), .Z(n4027) );
  XOR U2929 ( .A(n4030), .B(n4031), .Z(SUM[327]) );
  NANDN U2930 ( .A(n4032), .B(n4033), .Z(n4031) );
  ANDN U2931 ( .B(n4034), .A(n4035), .Z(n4030) );
  NAND U2932 ( .A(n4036), .B(n4037), .Z(n4034) );
  XNOR U2933 ( .A(n4036), .B(n4038), .Z(SUM[326]) );
  NANDN U2934 ( .A(n4035), .B(n4037), .Z(n4038) );
  NANDN U2935 ( .A(n4039), .B(n4040), .Z(n4036) );
  NAND U2936 ( .A(n4041), .B(n4042), .Z(n4040) );
  XNOR U2937 ( .A(n4041), .B(n4043), .Z(SUM[325]) );
  NANDN U2938 ( .A(n4039), .B(n4042), .Z(n4043) );
  NANDN U2939 ( .A(n4044), .B(n4045), .Z(n4041) );
  NANDN U2940 ( .A(n4029), .B(n4046), .Z(n4045) );
  XOR U2941 ( .A(n4029), .B(n4047), .Z(SUM[324]) );
  NANDN U2942 ( .A(n4044), .B(n4046), .Z(n4047) );
  ANDN U2943 ( .B(n4048), .A(n4049), .Z(n4029) );
  OR U2944 ( .A(n4050), .B(n3693), .Z(n4048) );
  XOR U2945 ( .A(n4051), .B(n4052), .Z(SUM[323]) );
  NANDN U2946 ( .A(n4053), .B(n4054), .Z(n4052) );
  ANDN U2947 ( .B(n4055), .A(n4056), .Z(n4051) );
  NAND U2948 ( .A(n4057), .B(n4058), .Z(n4055) );
  XNOR U2949 ( .A(n4057), .B(n4059), .Z(SUM[322]) );
  NANDN U2950 ( .A(n4056), .B(n4058), .Z(n4059) );
  NANDN U2951 ( .A(n4060), .B(n4061), .Z(n4057) );
  NAND U2952 ( .A(n4062), .B(n4063), .Z(n4061) );
  XNOR U2953 ( .A(n4062), .B(n4064), .Z(SUM[321]) );
  NANDN U2954 ( .A(n4060), .B(n4063), .Z(n4064) );
  NANDN U2955 ( .A(n4065), .B(n4066), .Z(n4062) );
  NANDN U2956 ( .A(n3693), .B(n4067), .Z(n4066) );
  XOR U2957 ( .A(n3693), .B(n4068), .Z(SUM[320]) );
  NANDN U2958 ( .A(n4065), .B(n4067), .Z(n4068) );
  NOR U2959 ( .A(n4069), .B(n4070), .Z(n3693) );
  XOR U2960 ( .A(n4071), .B(n4072), .Z(SUM[31]) );
  OR U2961 ( .A(n4073), .B(n4074), .Z(n4072) );
  ANDN U2962 ( .B(n4075), .A(n4076), .Z(n4071) );
  NANDN U2963 ( .A(n4077), .B(n4078), .Z(n4075) );
  XOR U2964 ( .A(n4079), .B(n4080), .Z(SUM[319]) );
  NANDN U2965 ( .A(n4081), .B(n4082), .Z(n4080) );
  ANDN U2966 ( .B(n4083), .A(n4084), .Z(n4079) );
  NAND U2967 ( .A(n4085), .B(n4086), .Z(n4083) );
  XNOR U2968 ( .A(n4085), .B(n4087), .Z(SUM[318]) );
  NANDN U2969 ( .A(n4084), .B(n4086), .Z(n4087) );
  NANDN U2970 ( .A(n4088), .B(n4089), .Z(n4085) );
  NAND U2971 ( .A(n4090), .B(n4091), .Z(n4089) );
  XNOR U2972 ( .A(n4090), .B(n4092), .Z(SUM[317]) );
  NANDN U2973 ( .A(n4088), .B(n4091), .Z(n4092) );
  NANDN U2974 ( .A(n4093), .B(n4094), .Z(n4090) );
  NAND U2975 ( .A(n4095), .B(n4096), .Z(n4094) );
  XNOR U2976 ( .A(n4095), .B(n4097), .Z(SUM[316]) );
  NANDN U2977 ( .A(n4093), .B(n4096), .Z(n4097) );
  NANDN U2978 ( .A(n4098), .B(n4099), .Z(n4095) );
  NANDN U2979 ( .A(n4100), .B(n4101), .Z(n4099) );
  XOR U2980 ( .A(n4102), .B(n4103), .Z(SUM[315]) );
  NANDN U2981 ( .A(n4104), .B(n4105), .Z(n4103) );
  ANDN U2982 ( .B(n4106), .A(n4107), .Z(n4102) );
  NAND U2983 ( .A(n4108), .B(n4109), .Z(n4106) );
  XNOR U2984 ( .A(n4108), .B(n4110), .Z(SUM[314]) );
  NANDN U2985 ( .A(n4107), .B(n4109), .Z(n4110) );
  NANDN U2986 ( .A(n4111), .B(n4112), .Z(n4108) );
  NAND U2987 ( .A(n4113), .B(n4114), .Z(n4112) );
  XNOR U2988 ( .A(n4113), .B(n4115), .Z(SUM[313]) );
  NANDN U2989 ( .A(n4111), .B(n4114), .Z(n4115) );
  NANDN U2990 ( .A(n4116), .B(n4117), .Z(n4113) );
  NAND U2991 ( .A(n4101), .B(n4118), .Z(n4117) );
  XNOR U2992 ( .A(n4101), .B(n4119), .Z(SUM[312]) );
  NANDN U2993 ( .A(n4116), .B(n4118), .Z(n4119) );
  NANDN U2994 ( .A(n4120), .B(n4121), .Z(n4101) );
  OR U2995 ( .A(n4122), .B(n4123), .Z(n4121) );
  XOR U2996 ( .A(n4124), .B(n4125), .Z(SUM[311]) );
  NANDN U2997 ( .A(n4126), .B(n4127), .Z(n4125) );
  ANDN U2998 ( .B(n4128), .A(n4129), .Z(n4124) );
  NAND U2999 ( .A(n4130), .B(n4131), .Z(n4128) );
  XNOR U3000 ( .A(n4130), .B(n4132), .Z(SUM[310]) );
  NANDN U3001 ( .A(n4129), .B(n4131), .Z(n4132) );
  NANDN U3002 ( .A(n4133), .B(n4134), .Z(n4130) );
  NAND U3003 ( .A(n4135), .B(n4136), .Z(n4134) );
  XNOR U3004 ( .A(n4078), .B(n4137), .Z(SUM[30]) );
  OR U3005 ( .A(n4077), .B(n4076), .Z(n4137) );
  NANDN U3006 ( .A(n4138), .B(n4139), .Z(n4078) );
  NANDN U3007 ( .A(n4140), .B(n4141), .Z(n4139) );
  XNOR U3008 ( .A(n4135), .B(n4142), .Z(SUM[309]) );
  NANDN U3009 ( .A(n4133), .B(n4136), .Z(n4142) );
  NANDN U3010 ( .A(n4143), .B(n4144), .Z(n4135) );
  NANDN U3011 ( .A(n4123), .B(n4145), .Z(n4144) );
  XOR U3012 ( .A(n4123), .B(n4146), .Z(SUM[308]) );
  NANDN U3013 ( .A(n4143), .B(n4145), .Z(n4146) );
  ANDN U3014 ( .B(n4147), .A(n4148), .Z(n4123) );
  NANDN U3015 ( .A(n4149), .B(n4150), .Z(n4147) );
  XOR U3016 ( .A(n4151), .B(n4152), .Z(SUM[307]) );
  NANDN U3017 ( .A(n4153), .B(n4154), .Z(n4152) );
  ANDN U3018 ( .B(n4155), .A(n4156), .Z(n4151) );
  NAND U3019 ( .A(n4157), .B(n4158), .Z(n4155) );
  XNOR U3020 ( .A(n4157), .B(n4159), .Z(SUM[306]) );
  NANDN U3021 ( .A(n4156), .B(n4158), .Z(n4159) );
  NANDN U3022 ( .A(n4160), .B(n4161), .Z(n4157) );
  NAND U3023 ( .A(n4162), .B(n4163), .Z(n4161) );
  XNOR U3024 ( .A(n4162), .B(n4164), .Z(SUM[305]) );
  NANDN U3025 ( .A(n4160), .B(n4163), .Z(n4164) );
  NANDN U3026 ( .A(n4165), .B(n4166), .Z(n4162) );
  NAND U3027 ( .A(n4150), .B(n4167), .Z(n4166) );
  XNOR U3028 ( .A(n4150), .B(n4168), .Z(SUM[304]) );
  NANDN U3029 ( .A(n4165), .B(n4167), .Z(n4168) );
  NANDN U3030 ( .A(n4169), .B(n4170), .Z(n4150) );
  NANDN U3031 ( .A(n4171), .B(n4172), .Z(n4170) );
  XOR U3032 ( .A(n4173), .B(n4174), .Z(SUM[303]) );
  NANDN U3033 ( .A(n4175), .B(n4176), .Z(n4174) );
  ANDN U3034 ( .B(n4177), .A(n4178), .Z(n4173) );
  NAND U3035 ( .A(n4179), .B(n4180), .Z(n4177) );
  XNOR U3036 ( .A(n4179), .B(n4181), .Z(SUM[302]) );
  NANDN U3037 ( .A(n4178), .B(n4180), .Z(n4181) );
  NANDN U3038 ( .A(n4182), .B(n4183), .Z(n4179) );
  NAND U3039 ( .A(n4184), .B(n4185), .Z(n4183) );
  XNOR U3040 ( .A(n4184), .B(n4186), .Z(SUM[301]) );
  NANDN U3041 ( .A(n4182), .B(n4185), .Z(n4186) );
  NANDN U3042 ( .A(n4187), .B(n4188), .Z(n4184) );
  NAND U3043 ( .A(n4189), .B(n4190), .Z(n4188) );
  XNOR U3044 ( .A(n4189), .B(n4191), .Z(SUM[300]) );
  NANDN U3045 ( .A(n4187), .B(n4190), .Z(n4191) );
  NANDN U3046 ( .A(n4192), .B(n4193), .Z(n4189) );
  NANDN U3047 ( .A(n4194), .B(n4195), .Z(n4193) );
  XNOR U3048 ( .A(n4196), .B(n4197), .Z(SUM[2]) );
  NANDN U3049 ( .A(n4198), .B(n4199), .Z(n4197) );
  XNOR U3050 ( .A(n4141), .B(n4200), .Z(SUM[29]) );
  OR U3051 ( .A(n4140), .B(n4138), .Z(n4200) );
  NANDN U3052 ( .A(n4201), .B(n4202), .Z(n4141) );
  NAND U3053 ( .A(n4203), .B(n4204), .Z(n4202) );
  XOR U3054 ( .A(n4205), .B(n4206), .Z(SUM[299]) );
  NANDN U3055 ( .A(n4207), .B(n4208), .Z(n4206) );
  ANDN U3056 ( .B(n4209), .A(n4210), .Z(n4205) );
  NAND U3057 ( .A(n4211), .B(n4212), .Z(n4209) );
  XNOR U3058 ( .A(n4211), .B(n4213), .Z(SUM[298]) );
  NANDN U3059 ( .A(n4210), .B(n4212), .Z(n4213) );
  NANDN U3060 ( .A(n4214), .B(n4215), .Z(n4211) );
  NAND U3061 ( .A(n4216), .B(n4217), .Z(n4215) );
  XNOR U3062 ( .A(n4216), .B(n4218), .Z(SUM[297]) );
  NANDN U3063 ( .A(n4214), .B(n4217), .Z(n4218) );
  NANDN U3064 ( .A(n4219), .B(n4220), .Z(n4216) );
  NAND U3065 ( .A(n4195), .B(n4221), .Z(n4220) );
  XNOR U3066 ( .A(n4195), .B(n4222), .Z(SUM[296]) );
  NANDN U3067 ( .A(n4219), .B(n4221), .Z(n4222) );
  NANDN U3068 ( .A(n4223), .B(n4224), .Z(n4195) );
  OR U3069 ( .A(n4225), .B(n4226), .Z(n4224) );
  XOR U3070 ( .A(n4227), .B(n4228), .Z(SUM[295]) );
  NANDN U3071 ( .A(n4229), .B(n4230), .Z(n4228) );
  ANDN U3072 ( .B(n4231), .A(n4232), .Z(n4227) );
  NAND U3073 ( .A(n4233), .B(n4234), .Z(n4231) );
  XNOR U3074 ( .A(n4233), .B(n4235), .Z(SUM[294]) );
  NANDN U3075 ( .A(n4232), .B(n4234), .Z(n4235) );
  NANDN U3076 ( .A(n4236), .B(n4237), .Z(n4233) );
  NAND U3077 ( .A(n4238), .B(n4239), .Z(n4237) );
  XNOR U3078 ( .A(n4238), .B(n4240), .Z(SUM[293]) );
  NANDN U3079 ( .A(n4236), .B(n4239), .Z(n4240) );
  NANDN U3080 ( .A(n4241), .B(n4242), .Z(n4238) );
  NANDN U3081 ( .A(n4226), .B(n4243), .Z(n4242) );
  XOR U3082 ( .A(n4226), .B(n4244), .Z(SUM[292]) );
  NANDN U3083 ( .A(n4241), .B(n4243), .Z(n4244) );
  ANDN U3084 ( .B(n4245), .A(n4246), .Z(n4226) );
  NANDN U3085 ( .A(n4247), .B(n4172), .Z(n4245) );
  XOR U3086 ( .A(n4248), .B(n4249), .Z(SUM[291]) );
  NANDN U3087 ( .A(n4250), .B(n4251), .Z(n4249) );
  ANDN U3088 ( .B(n4252), .A(n4253), .Z(n4248) );
  NAND U3089 ( .A(n4254), .B(n4255), .Z(n4252) );
  XNOR U3090 ( .A(n4254), .B(n4256), .Z(SUM[290]) );
  NANDN U3091 ( .A(n4253), .B(n4255), .Z(n4256) );
  NANDN U3092 ( .A(n4257), .B(n4258), .Z(n4254) );
  NAND U3093 ( .A(n4259), .B(n4260), .Z(n4258) );
  XNOR U3094 ( .A(n4203), .B(n4261), .Z(SUM[28]) );
  NANDN U3095 ( .A(n4201), .B(n4204), .Z(n4261) );
  NANDN U3096 ( .A(n4262), .B(n4263), .Z(n4203) );
  NANDN U3097 ( .A(n4264), .B(n4265), .Z(n4263) );
  XNOR U3098 ( .A(n4259), .B(n4266), .Z(SUM[289]) );
  NANDN U3099 ( .A(n4257), .B(n4260), .Z(n4266) );
  NANDN U3100 ( .A(n4267), .B(n4268), .Z(n4259) );
  NAND U3101 ( .A(n4172), .B(n4269), .Z(n4268) );
  XNOR U3102 ( .A(n4172), .B(n4270), .Z(SUM[288]) );
  NANDN U3103 ( .A(n4267), .B(n4269), .Z(n4270) );
  NANDN U3104 ( .A(n4271), .B(n4272), .Z(n4172) );
  OR U3105 ( .A(n4273), .B(n4274), .Z(n4272) );
  XOR U3106 ( .A(n4275), .B(n4276), .Z(SUM[287]) );
  NANDN U3107 ( .A(n4277), .B(n4278), .Z(n4276) );
  ANDN U3108 ( .B(n4279), .A(n4280), .Z(n4275) );
  NAND U3109 ( .A(n4281), .B(n4282), .Z(n4279) );
  XNOR U3110 ( .A(n4281), .B(n4283), .Z(SUM[286]) );
  NANDN U3111 ( .A(n4280), .B(n4282), .Z(n4283) );
  NANDN U3112 ( .A(n4284), .B(n4285), .Z(n4281) );
  NAND U3113 ( .A(n4286), .B(n4287), .Z(n4285) );
  XNOR U3114 ( .A(n4286), .B(n4288), .Z(SUM[285]) );
  NANDN U3115 ( .A(n4284), .B(n4287), .Z(n4288) );
  NANDN U3116 ( .A(n4289), .B(n4290), .Z(n4286) );
  NAND U3117 ( .A(n4291), .B(n4292), .Z(n4290) );
  XNOR U3118 ( .A(n4291), .B(n4293), .Z(SUM[284]) );
  NANDN U3119 ( .A(n4289), .B(n4292), .Z(n4293) );
  NANDN U3120 ( .A(n4294), .B(n4295), .Z(n4291) );
  NANDN U3121 ( .A(n4296), .B(n4297), .Z(n4295) );
  XOR U3122 ( .A(n4298), .B(n4299), .Z(SUM[283]) );
  NANDN U3123 ( .A(n4300), .B(n4301), .Z(n4299) );
  ANDN U3124 ( .B(n4302), .A(n4303), .Z(n4298) );
  NAND U3125 ( .A(n4304), .B(n4305), .Z(n4302) );
  XNOR U3126 ( .A(n4304), .B(n4306), .Z(SUM[282]) );
  NANDN U3127 ( .A(n4303), .B(n4305), .Z(n4306) );
  NANDN U3128 ( .A(n4307), .B(n4308), .Z(n4304) );
  NAND U3129 ( .A(n4309), .B(n4310), .Z(n4308) );
  XNOR U3130 ( .A(n4309), .B(n4311), .Z(SUM[281]) );
  NANDN U3131 ( .A(n4307), .B(n4310), .Z(n4311) );
  NANDN U3132 ( .A(n4312), .B(n4313), .Z(n4309) );
  NAND U3133 ( .A(n4297), .B(n4314), .Z(n4313) );
  XNOR U3134 ( .A(n4297), .B(n4315), .Z(SUM[280]) );
  NANDN U3135 ( .A(n4312), .B(n4314), .Z(n4315) );
  NANDN U3136 ( .A(n4316), .B(n4317), .Z(n4297) );
  OR U3137 ( .A(n4318), .B(n4319), .Z(n4317) );
  XOR U3138 ( .A(n4320), .B(n4321), .Z(SUM[27]) );
  NANDN U3139 ( .A(n4322), .B(n4323), .Z(n4321) );
  ANDN U3140 ( .B(n4324), .A(n4325), .Z(n4320) );
  NAND U3141 ( .A(n4326), .B(n4327), .Z(n4324) );
  XOR U3142 ( .A(n4328), .B(n4329), .Z(SUM[279]) );
  NANDN U3143 ( .A(n4330), .B(n4331), .Z(n4329) );
  ANDN U3144 ( .B(n4332), .A(n4333), .Z(n4328) );
  NAND U3145 ( .A(n4334), .B(n4335), .Z(n4332) );
  XNOR U3146 ( .A(n4334), .B(n4336), .Z(SUM[278]) );
  NANDN U3147 ( .A(n4333), .B(n4335), .Z(n4336) );
  NANDN U3148 ( .A(n4337), .B(n4338), .Z(n4334) );
  NAND U3149 ( .A(n4339), .B(n4340), .Z(n4338) );
  XNOR U3150 ( .A(n4339), .B(n4341), .Z(SUM[277]) );
  NANDN U3151 ( .A(n4337), .B(n4340), .Z(n4341) );
  NANDN U3152 ( .A(n4342), .B(n4343), .Z(n4339) );
  NANDN U3153 ( .A(n4319), .B(n4344), .Z(n4343) );
  XOR U3154 ( .A(n4319), .B(n4345), .Z(SUM[276]) );
  NANDN U3155 ( .A(n4342), .B(n4344), .Z(n4345) );
  ANDN U3156 ( .B(n4346), .A(n4347), .Z(n4319) );
  OR U3157 ( .A(n4348), .B(n4274), .Z(n4346) );
  XOR U3158 ( .A(n4349), .B(n4350), .Z(SUM[275]) );
  NANDN U3159 ( .A(n4351), .B(n4352), .Z(n4350) );
  ANDN U3160 ( .B(n4353), .A(n4354), .Z(n4349) );
  NAND U3161 ( .A(n4355), .B(n4356), .Z(n4353) );
  XNOR U3162 ( .A(n4355), .B(n4357), .Z(SUM[274]) );
  NANDN U3163 ( .A(n4354), .B(n4356), .Z(n4357) );
  NANDN U3164 ( .A(n4358), .B(n4359), .Z(n4355) );
  NAND U3165 ( .A(n4360), .B(n4361), .Z(n4359) );
  XNOR U3166 ( .A(n4360), .B(n4362), .Z(SUM[273]) );
  NANDN U3167 ( .A(n4358), .B(n4361), .Z(n4362) );
  NANDN U3168 ( .A(n4363), .B(n4364), .Z(n4360) );
  NANDN U3169 ( .A(n4274), .B(n4365), .Z(n4364) );
  XOR U3170 ( .A(n4274), .B(n4366), .Z(SUM[272]) );
  NANDN U3171 ( .A(n4363), .B(n4365), .Z(n4366) );
  ANDN U3172 ( .B(n4367), .A(n4368), .Z(n4274) );
  OR U3173 ( .A(n4369), .B(n4370), .Z(n4367) );
  XOR U3174 ( .A(n4371), .B(n4372), .Z(SUM[271]) );
  NANDN U3175 ( .A(n4373), .B(n4374), .Z(n4372) );
  ANDN U3176 ( .B(n4375), .A(n4376), .Z(n4371) );
  NAND U3177 ( .A(n4377), .B(n4378), .Z(n4375) );
  XNOR U3178 ( .A(n4377), .B(n4379), .Z(SUM[270]) );
  NANDN U3179 ( .A(n4376), .B(n4378), .Z(n4379) );
  NANDN U3180 ( .A(n4380), .B(n4381), .Z(n4377) );
  NAND U3181 ( .A(n4382), .B(n4383), .Z(n4381) );
  XNOR U3182 ( .A(n4326), .B(n4384), .Z(SUM[26]) );
  NANDN U3183 ( .A(n4325), .B(n4327), .Z(n4384) );
  NANDN U3184 ( .A(n4385), .B(n4386), .Z(n4326) );
  NAND U3185 ( .A(n4387), .B(n4388), .Z(n4386) );
  XNOR U3186 ( .A(n4382), .B(n4389), .Z(SUM[269]) );
  NANDN U3187 ( .A(n4380), .B(n4383), .Z(n4389) );
  NANDN U3188 ( .A(n4390), .B(n4391), .Z(n4382) );
  NAND U3189 ( .A(n4392), .B(n4393), .Z(n4391) );
  XNOR U3190 ( .A(n4392), .B(n4394), .Z(SUM[268]) );
  NANDN U3191 ( .A(n4390), .B(n4393), .Z(n4394) );
  NANDN U3192 ( .A(n4395), .B(n4396), .Z(n4392) );
  NANDN U3193 ( .A(n4397), .B(n4398), .Z(n4396) );
  XOR U3194 ( .A(n4399), .B(n4400), .Z(SUM[267]) );
  NANDN U3195 ( .A(n4401), .B(n4402), .Z(n4400) );
  ANDN U3196 ( .B(n4403), .A(n4404), .Z(n4399) );
  NAND U3197 ( .A(n4405), .B(n4406), .Z(n4403) );
  XNOR U3198 ( .A(n4405), .B(n4407), .Z(SUM[266]) );
  NANDN U3199 ( .A(n4404), .B(n4406), .Z(n4407) );
  NANDN U3200 ( .A(n4408), .B(n4409), .Z(n4405) );
  NAND U3201 ( .A(n4410), .B(n4411), .Z(n4409) );
  XNOR U3202 ( .A(n4410), .B(n4412), .Z(SUM[265]) );
  NANDN U3203 ( .A(n4408), .B(n4411), .Z(n4412) );
  NANDN U3204 ( .A(n4413), .B(n4414), .Z(n4410) );
  NAND U3205 ( .A(n4398), .B(n4415), .Z(n4414) );
  XNOR U3206 ( .A(n4398), .B(n4416), .Z(SUM[264]) );
  NANDN U3207 ( .A(n4413), .B(n4415), .Z(n4416) );
  NANDN U3208 ( .A(n4417), .B(n4418), .Z(n4398) );
  OR U3209 ( .A(n4419), .B(n4420), .Z(n4418) );
  XOR U3210 ( .A(n4421), .B(n4422), .Z(SUM[263]) );
  NANDN U3211 ( .A(n4423), .B(n4424), .Z(n4422) );
  ANDN U3212 ( .B(n4425), .A(n4426), .Z(n4421) );
  NAND U3213 ( .A(n4427), .B(n4428), .Z(n4425) );
  XNOR U3214 ( .A(n4427), .B(n4429), .Z(SUM[262]) );
  NANDN U3215 ( .A(n4426), .B(n4428), .Z(n4429) );
  NANDN U3216 ( .A(n4430), .B(n4431), .Z(n4427) );
  NAND U3217 ( .A(n4432), .B(n4433), .Z(n4431) );
  XNOR U3218 ( .A(n4432), .B(n4434), .Z(SUM[261]) );
  NANDN U3219 ( .A(n4430), .B(n4433), .Z(n4434) );
  NANDN U3220 ( .A(n4435), .B(n4436), .Z(n4432) );
  NANDN U3221 ( .A(n4420), .B(n4437), .Z(n4436) );
  XOR U3222 ( .A(n4420), .B(n4438), .Z(SUM[260]) );
  NANDN U3223 ( .A(n4435), .B(n4437), .Z(n4438) );
  ANDN U3224 ( .B(n4439), .A(n4440), .Z(n4420) );
  OR U3225 ( .A(n4441), .B(n4370), .Z(n4439) );
  XNOR U3226 ( .A(n4387), .B(n4442), .Z(SUM[25]) );
  NANDN U3227 ( .A(n4385), .B(n4388), .Z(n4442) );
  NANDN U3228 ( .A(n4443), .B(n4444), .Z(n4387) );
  NAND U3229 ( .A(n4265), .B(n4445), .Z(n4444) );
  XOR U3230 ( .A(n4446), .B(n4447), .Z(SUM[259]) );
  NANDN U3231 ( .A(n4448), .B(n4449), .Z(n4447) );
  ANDN U3232 ( .B(n4450), .A(n4451), .Z(n4446) );
  NAND U3233 ( .A(n4452), .B(n4453), .Z(n4450) );
  XNOR U3234 ( .A(n4452), .B(n4454), .Z(SUM[258]) );
  NANDN U3235 ( .A(n4451), .B(n4453), .Z(n4454) );
  NANDN U3236 ( .A(n4455), .B(n4456), .Z(n4452) );
  NAND U3237 ( .A(n4457), .B(n4458), .Z(n4456) );
  XNOR U3238 ( .A(n4457), .B(n4459), .Z(SUM[257]) );
  NANDN U3239 ( .A(n4455), .B(n4458), .Z(n4459) );
  NANDN U3240 ( .A(n4460), .B(n4461), .Z(n4457) );
  NANDN U3241 ( .A(n4370), .B(n4462), .Z(n4461) );
  XOR U3242 ( .A(n4370), .B(n4463), .Z(SUM[256]) );
  NANDN U3243 ( .A(n4460), .B(n4462), .Z(n4463) );
  XOR U3244 ( .A(n4464), .B(n4465), .Z(SUM[255]) );
  OR U3245 ( .A(n4466), .B(n4467), .Z(n4465) );
  ANDN U3246 ( .B(n4468), .A(n4469), .Z(n4464) );
  NANDN U3247 ( .A(n4470), .B(n4471), .Z(n4468) );
  XNOR U3248 ( .A(n4471), .B(n4472), .Z(SUM[254]) );
  OR U3249 ( .A(n4470), .B(n4469), .Z(n4472) );
  NANDN U3250 ( .A(n4473), .B(n4474), .Z(n4471) );
  NANDN U3251 ( .A(n4475), .B(n4476), .Z(n4474) );
  XNOR U3252 ( .A(n4476), .B(n4477), .Z(SUM[253]) );
  OR U3253 ( .A(n4475), .B(n4473), .Z(n4477) );
  NANDN U3254 ( .A(n4478), .B(n4479), .Z(n4476) );
  NAND U3255 ( .A(n4480), .B(n4481), .Z(n4479) );
  XNOR U3256 ( .A(n4480), .B(n4482), .Z(SUM[252]) );
  NANDN U3257 ( .A(n4478), .B(n4481), .Z(n4482) );
  NANDN U3258 ( .A(n4483), .B(n4484), .Z(n4480) );
  NANDN U3259 ( .A(n4485), .B(n4486), .Z(n4484) );
  XOR U3260 ( .A(n4487), .B(n4488), .Z(SUM[251]) );
  NANDN U3261 ( .A(n4489), .B(n4490), .Z(n4488) );
  ANDN U3262 ( .B(n4491), .A(n4492), .Z(n4487) );
  NAND U3263 ( .A(n4493), .B(n4494), .Z(n4491) );
  XNOR U3264 ( .A(n4493), .B(n4495), .Z(SUM[250]) );
  NANDN U3265 ( .A(n4492), .B(n4494), .Z(n4495) );
  NANDN U3266 ( .A(n4496), .B(n4497), .Z(n4493) );
  NAND U3267 ( .A(n4498), .B(n4499), .Z(n4497) );
  XNOR U3268 ( .A(n4265), .B(n4500), .Z(SUM[24]) );
  NANDN U3269 ( .A(n4443), .B(n4445), .Z(n4500) );
  NANDN U3270 ( .A(n4501), .B(n4502), .Z(n4265) );
  NANDN U3271 ( .A(n4503), .B(n4504), .Z(n4502) );
  XNOR U3272 ( .A(n4498), .B(n4505), .Z(SUM[249]) );
  NANDN U3273 ( .A(n4496), .B(n4499), .Z(n4505) );
  NANDN U3274 ( .A(n4506), .B(n4507), .Z(n4498) );
  NAND U3275 ( .A(n4486), .B(n4508), .Z(n4507) );
  XNOR U3276 ( .A(n4486), .B(n4509), .Z(SUM[248]) );
  NANDN U3277 ( .A(n4506), .B(n4508), .Z(n4509) );
  NANDN U3278 ( .A(n4510), .B(n4511), .Z(n4486) );
  NANDN U3279 ( .A(n4512), .B(n4513), .Z(n4511) );
  XOR U3280 ( .A(n4514), .B(n4515), .Z(SUM[247]) );
  NANDN U3281 ( .A(n4516), .B(n4517), .Z(n4515) );
  ANDN U3282 ( .B(n4518), .A(n4519), .Z(n4514) );
  NAND U3283 ( .A(n4520), .B(n4521), .Z(n4518) );
  XNOR U3284 ( .A(n4520), .B(n4522), .Z(SUM[246]) );
  NANDN U3285 ( .A(n4519), .B(n4521), .Z(n4522) );
  NANDN U3286 ( .A(n4523), .B(n4524), .Z(n4520) );
  NAND U3287 ( .A(n4525), .B(n4526), .Z(n4524) );
  XNOR U3288 ( .A(n4525), .B(n4527), .Z(SUM[245]) );
  NANDN U3289 ( .A(n4523), .B(n4526), .Z(n4527) );
  NANDN U3290 ( .A(n4528), .B(n4529), .Z(n4525) );
  NANDN U3291 ( .A(n4512), .B(n4530), .Z(n4529) );
  XOR U3292 ( .A(n4512), .B(n4531), .Z(SUM[244]) );
  NANDN U3293 ( .A(n4528), .B(n4530), .Z(n4531) );
  ANDN U3294 ( .B(n4532), .A(n4533), .Z(n4512) );
  OR U3295 ( .A(n4534), .B(n4535), .Z(n4532) );
  XOR U3296 ( .A(n4536), .B(n4537), .Z(SUM[243]) );
  NANDN U3297 ( .A(n4538), .B(n4539), .Z(n4537) );
  ANDN U3298 ( .B(n4540), .A(n4541), .Z(n4536) );
  NANDN U3299 ( .A(n4542), .B(n4543), .Z(n4540) );
  XNOR U3300 ( .A(n4543), .B(n4544), .Z(SUM[242]) );
  OR U3301 ( .A(n4542), .B(n4541), .Z(n4544) );
  NANDN U3302 ( .A(n4545), .B(n4546), .Z(n4543) );
  NAND U3303 ( .A(n4547), .B(n4548), .Z(n4546) );
  XNOR U3304 ( .A(n4547), .B(n4549), .Z(SUM[241]) );
  NANDN U3305 ( .A(n4545), .B(n4548), .Z(n4549) );
  NANDN U3306 ( .A(n4550), .B(n4551), .Z(n4547) );
  NANDN U3307 ( .A(n4535), .B(n4552), .Z(n4551) );
  XOR U3308 ( .A(n4535), .B(n4553), .Z(SUM[240]) );
  NANDN U3309 ( .A(n4550), .B(n4552), .Z(n4553) );
  XOR U3310 ( .A(n4554), .B(n4555), .Z(SUM[23]) );
  NANDN U3311 ( .A(n4556), .B(n4557), .Z(n4555) );
  ANDN U3312 ( .B(n4558), .A(n4559), .Z(n4554) );
  NAND U3313 ( .A(n4560), .B(n4561), .Z(n4558) );
  XOR U3314 ( .A(n4562), .B(n4563), .Z(SUM[239]) );
  OR U3315 ( .A(n4564), .B(n4565), .Z(n4563) );
  ANDN U3316 ( .B(n4566), .A(n4567), .Z(n4562) );
  NANDN U3317 ( .A(n4568), .B(n4569), .Z(n4566) );
  XNOR U3318 ( .A(n4569), .B(n4570), .Z(SUM[238]) );
  OR U3319 ( .A(n4568), .B(n4567), .Z(n4570) );
  NANDN U3320 ( .A(n4571), .B(n4572), .Z(n4569) );
  NANDN U3321 ( .A(n4573), .B(n4574), .Z(n4572) );
  XNOR U3322 ( .A(n4574), .B(n4575), .Z(SUM[237]) );
  OR U3323 ( .A(n4573), .B(n4571), .Z(n4575) );
  NANDN U3324 ( .A(n4576), .B(n4577), .Z(n4574) );
  NAND U3325 ( .A(n4578), .B(n4579), .Z(n4577) );
  XNOR U3326 ( .A(n4578), .B(n4580), .Z(SUM[236]) );
  NANDN U3327 ( .A(n4576), .B(n4579), .Z(n4580) );
  NANDN U3328 ( .A(n4581), .B(n4582), .Z(n4578) );
  NANDN U3329 ( .A(n4583), .B(n4584), .Z(n4582) );
  XOR U3330 ( .A(n4585), .B(n4586), .Z(SUM[235]) );
  NANDN U3331 ( .A(n4587), .B(n4588), .Z(n4586) );
  ANDN U3332 ( .B(n4589), .A(n4590), .Z(n4585) );
  NAND U3333 ( .A(n4591), .B(n4592), .Z(n4589) );
  XNOR U3334 ( .A(n4591), .B(n4593), .Z(SUM[234]) );
  NANDN U3335 ( .A(n4590), .B(n4592), .Z(n4593) );
  NANDN U3336 ( .A(n4594), .B(n4595), .Z(n4591) );
  NAND U3337 ( .A(n4596), .B(n4597), .Z(n4595) );
  XNOR U3338 ( .A(n4596), .B(n4598), .Z(SUM[233]) );
  NANDN U3339 ( .A(n4594), .B(n4597), .Z(n4598) );
  NANDN U3340 ( .A(n4599), .B(n4600), .Z(n4596) );
  NAND U3341 ( .A(n4584), .B(n4601), .Z(n4600) );
  XNOR U3342 ( .A(n4584), .B(n4602), .Z(SUM[232]) );
  NANDN U3343 ( .A(n4599), .B(n4601), .Z(n4602) );
  NANDN U3344 ( .A(n4603), .B(n4604), .Z(n4584) );
  NANDN U3345 ( .A(n4605), .B(n4606), .Z(n4604) );
  XOR U3346 ( .A(n4607), .B(n4608), .Z(SUM[231]) );
  NANDN U3347 ( .A(n4609), .B(n4610), .Z(n4608) );
  ANDN U3348 ( .B(n4611), .A(n4612), .Z(n4607) );
  NAND U3349 ( .A(n4613), .B(n4614), .Z(n4611) );
  XNOR U3350 ( .A(n4613), .B(n4615), .Z(SUM[230]) );
  NANDN U3351 ( .A(n4612), .B(n4614), .Z(n4615) );
  NANDN U3352 ( .A(n4616), .B(n4617), .Z(n4613) );
  NAND U3353 ( .A(n4618), .B(n4619), .Z(n4617) );
  XNOR U3354 ( .A(n4560), .B(n4620), .Z(SUM[22]) );
  NANDN U3355 ( .A(n4559), .B(n4561), .Z(n4620) );
  NANDN U3356 ( .A(n4621), .B(n4622), .Z(n4560) );
  NAND U3357 ( .A(n4623), .B(n4624), .Z(n4622) );
  XNOR U3358 ( .A(n4618), .B(n4625), .Z(SUM[229]) );
  NANDN U3359 ( .A(n4616), .B(n4619), .Z(n4625) );
  NANDN U3360 ( .A(n4626), .B(n4627), .Z(n4618) );
  NANDN U3361 ( .A(n4605), .B(n4628), .Z(n4627) );
  XOR U3362 ( .A(n4605), .B(n4629), .Z(SUM[228]) );
  NANDN U3363 ( .A(n4626), .B(n4628), .Z(n4629) );
  ANDN U3364 ( .B(n4630), .A(n4631), .Z(n4605) );
  OR U3365 ( .A(n4632), .B(n4633), .Z(n4630) );
  XOR U3366 ( .A(n4634), .B(n4635), .Z(SUM[227]) );
  NANDN U3367 ( .A(n4636), .B(n4637), .Z(n4635) );
  ANDN U3368 ( .B(n4638), .A(n4639), .Z(n4634) );
  NANDN U3369 ( .A(n4640), .B(n4641), .Z(n4638) );
  XNOR U3370 ( .A(n4641), .B(n4642), .Z(SUM[226]) );
  OR U3371 ( .A(n4640), .B(n4639), .Z(n4642) );
  NANDN U3372 ( .A(n4643), .B(n4644), .Z(n4641) );
  NAND U3373 ( .A(n4645), .B(n4646), .Z(n4644) );
  XNOR U3374 ( .A(n4645), .B(n4647), .Z(SUM[225]) );
  NANDN U3375 ( .A(n4643), .B(n4646), .Z(n4647) );
  NANDN U3376 ( .A(n4648), .B(n4649), .Z(n4645) );
  NANDN U3377 ( .A(n4633), .B(n4650), .Z(n4649) );
  XOR U3378 ( .A(n4633), .B(n4651), .Z(SUM[224]) );
  NANDN U3379 ( .A(n4648), .B(n4650), .Z(n4651) );
  XOR U3380 ( .A(n4652), .B(n4653), .Z(SUM[223]) );
  OR U3381 ( .A(n4654), .B(n4655), .Z(n4653) );
  ANDN U3382 ( .B(n4656), .A(n4657), .Z(n4652) );
  NANDN U3383 ( .A(n4658), .B(n4659), .Z(n4656) );
  XNOR U3384 ( .A(n4659), .B(n4660), .Z(SUM[222]) );
  OR U3385 ( .A(n4658), .B(n4657), .Z(n4660) );
  NANDN U3386 ( .A(n4661), .B(n4662), .Z(n4659) );
  NANDN U3387 ( .A(n4663), .B(n4664), .Z(n4662) );
  XNOR U3388 ( .A(n4664), .B(n4665), .Z(SUM[221]) );
  OR U3389 ( .A(n4663), .B(n4661), .Z(n4665) );
  NANDN U3390 ( .A(n4666), .B(n4667), .Z(n4664) );
  NAND U3391 ( .A(n4668), .B(n4669), .Z(n4667) );
  XNOR U3392 ( .A(n4668), .B(n4670), .Z(SUM[220]) );
  NANDN U3393 ( .A(n4666), .B(n4669), .Z(n4670) );
  NANDN U3394 ( .A(n4671), .B(n4672), .Z(n4668) );
  NANDN U3395 ( .A(n4673), .B(n4674), .Z(n4672) );
  XNOR U3396 ( .A(n4623), .B(n4675), .Z(SUM[21]) );
  NANDN U3397 ( .A(n4621), .B(n4624), .Z(n4675) );
  NANDN U3398 ( .A(n4676), .B(n4677), .Z(n4623) );
  NANDN U3399 ( .A(n4503), .B(n4678), .Z(n4677) );
  XOR U3400 ( .A(n4679), .B(n4680), .Z(SUM[219]) );
  NANDN U3401 ( .A(n4681), .B(n4682), .Z(n4680) );
  ANDN U3402 ( .B(n4683), .A(n4684), .Z(n4679) );
  NAND U3403 ( .A(n4685), .B(n4686), .Z(n4683) );
  XNOR U3404 ( .A(n4685), .B(n4687), .Z(SUM[218]) );
  NANDN U3405 ( .A(n4684), .B(n4686), .Z(n4687) );
  NANDN U3406 ( .A(n4688), .B(n4689), .Z(n4685) );
  NAND U3407 ( .A(n4690), .B(n4691), .Z(n4689) );
  XNOR U3408 ( .A(n4690), .B(n4692), .Z(SUM[217]) );
  NANDN U3409 ( .A(n4688), .B(n4691), .Z(n4692) );
  NANDN U3410 ( .A(n4693), .B(n4694), .Z(n4690) );
  NAND U3411 ( .A(n4674), .B(n4695), .Z(n4694) );
  XNOR U3412 ( .A(n4674), .B(n4696), .Z(SUM[216]) );
  NANDN U3413 ( .A(n4693), .B(n4695), .Z(n4696) );
  NANDN U3414 ( .A(n4697), .B(n4698), .Z(n4674) );
  NANDN U3415 ( .A(n4699), .B(n4700), .Z(n4698) );
  XOR U3416 ( .A(n4701), .B(n4702), .Z(SUM[215]) );
  NANDN U3417 ( .A(n4703), .B(n4704), .Z(n4702) );
  ANDN U3418 ( .B(n4705), .A(n4706), .Z(n4701) );
  NAND U3419 ( .A(n4707), .B(n4708), .Z(n4705) );
  XNOR U3420 ( .A(n4707), .B(n4709), .Z(SUM[214]) );
  NANDN U3421 ( .A(n4706), .B(n4708), .Z(n4709) );
  NANDN U3422 ( .A(n4710), .B(n4711), .Z(n4707) );
  NAND U3423 ( .A(n4712), .B(n4713), .Z(n4711) );
  XNOR U3424 ( .A(n4712), .B(n4714), .Z(SUM[213]) );
  NANDN U3425 ( .A(n4710), .B(n4713), .Z(n4714) );
  NANDN U3426 ( .A(n4715), .B(n4716), .Z(n4712) );
  NANDN U3427 ( .A(n4699), .B(n4717), .Z(n4716) );
  XOR U3428 ( .A(n4699), .B(n4718), .Z(SUM[212]) );
  NANDN U3429 ( .A(n4715), .B(n4717), .Z(n4718) );
  ANDN U3430 ( .B(n4719), .A(n4720), .Z(n4699) );
  OR U3431 ( .A(n4721), .B(n4722), .Z(n4719) );
  XOR U3432 ( .A(n4723), .B(n4724), .Z(SUM[211]) );
  NANDN U3433 ( .A(n4725), .B(n4726), .Z(n4724) );
  ANDN U3434 ( .B(n4727), .A(n4728), .Z(n4723) );
  NANDN U3435 ( .A(n4729), .B(n4730), .Z(n4727) );
  XNOR U3436 ( .A(n4730), .B(n4731), .Z(SUM[210]) );
  OR U3437 ( .A(n4729), .B(n4728), .Z(n4731) );
  NANDN U3438 ( .A(n4732), .B(n4733), .Z(n4730) );
  NAND U3439 ( .A(n4734), .B(n4735), .Z(n4733) );
  XOR U3440 ( .A(n4503), .B(n4736), .Z(SUM[20]) );
  NANDN U3441 ( .A(n4676), .B(n4678), .Z(n4736) );
  ANDN U3442 ( .B(n4737), .A(n4738), .Z(n4503) );
  OR U3443 ( .A(n4739), .B(n4740), .Z(n4737) );
  XNOR U3444 ( .A(n4734), .B(n4741), .Z(SUM[209]) );
  NANDN U3445 ( .A(n4732), .B(n4735), .Z(n4741) );
  NANDN U3446 ( .A(n4742), .B(n4743), .Z(n4734) );
  NANDN U3447 ( .A(n4722), .B(n4744), .Z(n4743) );
  XOR U3448 ( .A(n4722), .B(n4745), .Z(SUM[208]) );
  NANDN U3449 ( .A(n4742), .B(n4744), .Z(n4745) );
  XOR U3450 ( .A(n4746), .B(n4747), .Z(SUM[207]) );
  OR U3451 ( .A(n4748), .B(n4749), .Z(n4747) );
  ANDN U3452 ( .B(n4750), .A(n4751), .Z(n4746) );
  NANDN U3453 ( .A(n4752), .B(n4753), .Z(n4750) );
  XNOR U3454 ( .A(n4753), .B(n4754), .Z(SUM[206]) );
  OR U3455 ( .A(n4752), .B(n4751), .Z(n4754) );
  NANDN U3456 ( .A(n4755), .B(n4756), .Z(n4753) );
  NANDN U3457 ( .A(n4757), .B(n4758), .Z(n4756) );
  XNOR U3458 ( .A(n4758), .B(n4759), .Z(SUM[205]) );
  OR U3459 ( .A(n4757), .B(n4755), .Z(n4759) );
  NANDN U3460 ( .A(n4760), .B(n4761), .Z(n4758) );
  NAND U3461 ( .A(n4762), .B(n4763), .Z(n4761) );
  XNOR U3462 ( .A(n4762), .B(n4764), .Z(SUM[204]) );
  NANDN U3463 ( .A(n4760), .B(n4763), .Z(n4764) );
  NANDN U3464 ( .A(n4765), .B(n4766), .Z(n4762) );
  NANDN U3465 ( .A(n4767), .B(n4768), .Z(n4766) );
  XOR U3466 ( .A(n4769), .B(n4770), .Z(SUM[203]) );
  NANDN U3467 ( .A(n4771), .B(n4772), .Z(n4770) );
  ANDN U3468 ( .B(n4773), .A(n4774), .Z(n4769) );
  NAND U3469 ( .A(n4775), .B(n4776), .Z(n4773) );
  XNOR U3470 ( .A(n4775), .B(n4777), .Z(SUM[202]) );
  NANDN U3471 ( .A(n4774), .B(n4776), .Z(n4777) );
  NANDN U3472 ( .A(n4778), .B(n4779), .Z(n4775) );
  NAND U3473 ( .A(n4780), .B(n4781), .Z(n4779) );
  XNOR U3474 ( .A(n4780), .B(n4782), .Z(SUM[201]) );
  NANDN U3475 ( .A(n4778), .B(n4781), .Z(n4782) );
  NANDN U3476 ( .A(n4783), .B(n4784), .Z(n4780) );
  NAND U3477 ( .A(n4768), .B(n4785), .Z(n4784) );
  XNOR U3478 ( .A(n4768), .B(n4786), .Z(SUM[200]) );
  NANDN U3479 ( .A(n4783), .B(n4785), .Z(n4786) );
  NANDN U3480 ( .A(n4787), .B(n4788), .Z(n4768) );
  NANDN U3481 ( .A(n4789), .B(n4790), .Z(n4788) );
  XOR U3482 ( .A(n4791), .B(n4792), .Z(SUM[1]) );
  NOR U3483 ( .A(n4793), .B(n4794), .Z(n4792) );
  XOR U3484 ( .A(n4795), .B(n4796), .Z(SUM[19]) );
  NANDN U3485 ( .A(n4797), .B(n4798), .Z(n4796) );
  ANDN U3486 ( .B(n4799), .A(n4800), .Z(n4795) );
  NANDN U3487 ( .A(n4801), .B(n4802), .Z(n4799) );
  XOR U3488 ( .A(n4803), .B(n4804), .Z(SUM[199]) );
  NANDN U3489 ( .A(n4805), .B(n4806), .Z(n4804) );
  ANDN U3490 ( .B(n4807), .A(n4808), .Z(n4803) );
  NAND U3491 ( .A(n4809), .B(n4810), .Z(n4807) );
  XNOR U3492 ( .A(n4809), .B(n4811), .Z(SUM[198]) );
  NANDN U3493 ( .A(n4808), .B(n4810), .Z(n4811) );
  NANDN U3494 ( .A(n4812), .B(n4813), .Z(n4809) );
  NAND U3495 ( .A(n4814), .B(n4815), .Z(n4813) );
  XNOR U3496 ( .A(n4814), .B(n4816), .Z(SUM[197]) );
  NANDN U3497 ( .A(n4812), .B(n4815), .Z(n4816) );
  NANDN U3498 ( .A(n4817), .B(n4818), .Z(n4814) );
  NANDN U3499 ( .A(n4789), .B(n4819), .Z(n4818) );
  XOR U3500 ( .A(n4789), .B(n4820), .Z(SUM[196]) );
  NANDN U3501 ( .A(n4817), .B(n4819), .Z(n4820) );
  ANDN U3502 ( .B(n4821), .A(n4822), .Z(n4789) );
  OR U3503 ( .A(n4823), .B(n4824), .Z(n4821) );
  XOR U3504 ( .A(n4825), .B(n4826), .Z(SUM[195]) );
  NANDN U3505 ( .A(n4827), .B(n4828), .Z(n4826) );
  ANDN U3506 ( .B(n4829), .A(n4830), .Z(n4825) );
  NANDN U3507 ( .A(n4831), .B(n4832), .Z(n4829) );
  XNOR U3508 ( .A(n4832), .B(n4833), .Z(SUM[194]) );
  OR U3509 ( .A(n4831), .B(n4830), .Z(n4833) );
  NANDN U3510 ( .A(n4834), .B(n4835), .Z(n4832) );
  NAND U3511 ( .A(n4836), .B(n4837), .Z(n4835) );
  XNOR U3512 ( .A(n4836), .B(n4838), .Z(SUM[193]) );
  NANDN U3513 ( .A(n4834), .B(n4837), .Z(n4838) );
  NANDN U3514 ( .A(n4839), .B(n4840), .Z(n4836) );
  NANDN U3515 ( .A(n4824), .B(n4841), .Z(n4840) );
  XOR U3516 ( .A(n4824), .B(n4842), .Z(SUM[192]) );
  NANDN U3517 ( .A(n4839), .B(n4841), .Z(n4842) );
  XOR U3518 ( .A(n4843), .B(n4844), .Z(SUM[191]) );
  OR U3519 ( .A(n4845), .B(n4846), .Z(n4844) );
  ANDN U3520 ( .B(n4847), .A(n4848), .Z(n4843) );
  NAND U3521 ( .A(n4849), .B(n4850), .Z(n4847) );
  XNOR U3522 ( .A(n4849), .B(n4851), .Z(SUM[190]) );
  NANDN U3523 ( .A(n4848), .B(n4850), .Z(n4851) );
  NANDN U3524 ( .A(n4852), .B(n4853), .Z(n4849) );
  NAND U3525 ( .A(n4854), .B(n4855), .Z(n4853) );
  XNOR U3526 ( .A(n4802), .B(n4856), .Z(SUM[18]) );
  OR U3527 ( .A(n4801), .B(n4800), .Z(n4856) );
  NANDN U3528 ( .A(n4857), .B(n4858), .Z(n4802) );
  NAND U3529 ( .A(n4859), .B(n4860), .Z(n4858) );
  XNOR U3530 ( .A(n4854), .B(n4861), .Z(SUM[189]) );
  NANDN U3531 ( .A(n4852), .B(n4855), .Z(n4861) );
  NANDN U3532 ( .A(n4862), .B(n4863), .Z(n4854) );
  NANDN U3533 ( .A(n4864), .B(n4865), .Z(n4863) );
  XNOR U3534 ( .A(n4865), .B(n4866), .Z(SUM[188]) );
  OR U3535 ( .A(n4864), .B(n4862), .Z(n4866) );
  NANDN U3536 ( .A(n4867), .B(n4868), .Z(n4865) );
  NANDN U3537 ( .A(n4869), .B(n4870), .Z(n4868) );
  XOR U3538 ( .A(n4871), .B(n4872), .Z(SUM[187]) );
  NANDN U3539 ( .A(n4873), .B(n4874), .Z(n4872) );
  ANDN U3540 ( .B(n4875), .A(n4876), .Z(n4871) );
  NAND U3541 ( .A(n4877), .B(n4878), .Z(n4875) );
  XNOR U3542 ( .A(n4877), .B(n4879), .Z(SUM[186]) );
  NANDN U3543 ( .A(n4876), .B(n4878), .Z(n4879) );
  NANDN U3544 ( .A(n4880), .B(n4881), .Z(n4877) );
  NAND U3545 ( .A(n4882), .B(n4883), .Z(n4881) );
  XNOR U3546 ( .A(n4882), .B(n4884), .Z(SUM[185]) );
  NANDN U3547 ( .A(n4880), .B(n4883), .Z(n4884) );
  NANDN U3548 ( .A(n4885), .B(n4886), .Z(n4882) );
  NAND U3549 ( .A(n4870), .B(n4887), .Z(n4886) );
  XNOR U3550 ( .A(n4870), .B(n4888), .Z(SUM[184]) );
  NANDN U3551 ( .A(n4885), .B(n4887), .Z(n4888) );
  NANDN U3552 ( .A(n4889), .B(n4890), .Z(n4870) );
  NANDN U3553 ( .A(n4891), .B(n4892), .Z(n4890) );
  XOR U3554 ( .A(n4893), .B(n4894), .Z(SUM[183]) );
  NANDN U3555 ( .A(n4895), .B(n4896), .Z(n4894) );
  ANDN U3556 ( .B(n4897), .A(n4898), .Z(n4893) );
  NAND U3557 ( .A(n4899), .B(n4900), .Z(n4897) );
  XNOR U3558 ( .A(n4899), .B(n4901), .Z(SUM[182]) );
  NANDN U3559 ( .A(n4898), .B(n4900), .Z(n4901) );
  NANDN U3560 ( .A(n4902), .B(n4903), .Z(n4899) );
  NAND U3561 ( .A(n4904), .B(n4905), .Z(n4903) );
  XNOR U3562 ( .A(n4904), .B(n4906), .Z(SUM[181]) );
  NANDN U3563 ( .A(n4902), .B(n4905), .Z(n4906) );
  NANDN U3564 ( .A(n4907), .B(n4908), .Z(n4904) );
  NANDN U3565 ( .A(n4891), .B(n4909), .Z(n4908) );
  XOR U3566 ( .A(n4891), .B(n4910), .Z(SUM[180]) );
  NANDN U3567 ( .A(n4907), .B(n4909), .Z(n4910) );
  ANDN U3568 ( .B(n4911), .A(n4912), .Z(n4891) );
  NANDN U3569 ( .A(n4913), .B(n4914), .Z(n4911) );
  XNOR U3570 ( .A(n4859), .B(n4915), .Z(SUM[17]) );
  NANDN U3571 ( .A(n4857), .B(n4860), .Z(n4915) );
  NANDN U3572 ( .A(n4916), .B(n4917), .Z(n4859) );
  NANDN U3573 ( .A(n4740), .B(n4918), .Z(n4917) );
  XOR U3574 ( .A(n4919), .B(n4920), .Z(SUM[179]) );
  NANDN U3575 ( .A(n4921), .B(n4922), .Z(n4920) );
  ANDN U3576 ( .B(n4923), .A(n4924), .Z(n4919) );
  NANDN U3577 ( .A(n4925), .B(n4926), .Z(n4923) );
  XNOR U3578 ( .A(n4926), .B(n4927), .Z(SUM[178]) );
  OR U3579 ( .A(n4925), .B(n4924), .Z(n4927) );
  NANDN U3580 ( .A(n4928), .B(n4929), .Z(n4926) );
  NAND U3581 ( .A(n4930), .B(n4931), .Z(n4929) );
  XNOR U3582 ( .A(n4930), .B(n4932), .Z(SUM[177]) );
  NANDN U3583 ( .A(n4928), .B(n4931), .Z(n4932) );
  NANDN U3584 ( .A(n4933), .B(n4934), .Z(n4930) );
  NAND U3585 ( .A(n4914), .B(n4935), .Z(n4934) );
  XNOR U3586 ( .A(n4914), .B(n4936), .Z(SUM[176]) );
  NANDN U3587 ( .A(n4933), .B(n4935), .Z(n4936) );
  XOR U3588 ( .A(n4937), .B(n4938), .Z(SUM[175]) );
  NANDN U3589 ( .A(n4939), .B(n4940), .Z(n4938) );
  ANDN U3590 ( .B(n4941), .A(n4942), .Z(n4937) );
  NAND U3591 ( .A(n4943), .B(n4944), .Z(n4941) );
  XNOR U3592 ( .A(n4943), .B(n4945), .Z(SUM[174]) );
  NANDN U3593 ( .A(n4942), .B(n4944), .Z(n4945) );
  NANDN U3594 ( .A(n4946), .B(n4947), .Z(n4943) );
  NAND U3595 ( .A(n4948), .B(n4949), .Z(n4947) );
  XNOR U3596 ( .A(n4948), .B(n4950), .Z(SUM[173]) );
  NANDN U3597 ( .A(n4946), .B(n4949), .Z(n4950) );
  NANDN U3598 ( .A(n4951), .B(n4952), .Z(n4948) );
  NAND U3599 ( .A(n4953), .B(n4954), .Z(n4952) );
  XNOR U3600 ( .A(n4953), .B(n4955), .Z(SUM[172]) );
  NANDN U3601 ( .A(n4951), .B(n4954), .Z(n4955) );
  NANDN U3602 ( .A(n4956), .B(n4957), .Z(n4953) );
  NAND U3603 ( .A(n4958), .B(n4959), .Z(n4957) );
  XOR U3604 ( .A(n4960), .B(n4961), .Z(SUM[171]) );
  NANDN U3605 ( .A(n4962), .B(n4963), .Z(n4961) );
  ANDN U3606 ( .B(n4964), .A(n4965), .Z(n4960) );
  NAND U3607 ( .A(n4966), .B(n4967), .Z(n4964) );
  XNOR U3608 ( .A(n4966), .B(n4968), .Z(SUM[170]) );
  NANDN U3609 ( .A(n4965), .B(n4967), .Z(n4968) );
  NANDN U3610 ( .A(n4969), .B(n4970), .Z(n4966) );
  NAND U3611 ( .A(n4971), .B(n4972), .Z(n4970) );
  XOR U3612 ( .A(n4740), .B(n4973), .Z(SUM[16]) );
  NANDN U3613 ( .A(n4916), .B(n4918), .Z(n4973) );
  XNOR U3614 ( .A(n4971), .B(n4974), .Z(SUM[169]) );
  NANDN U3615 ( .A(n4969), .B(n4972), .Z(n4974) );
  NANDN U3616 ( .A(n4975), .B(n4976), .Z(n4971) );
  NAND U3617 ( .A(n4959), .B(n4977), .Z(n4976) );
  XNOR U3618 ( .A(n4959), .B(n4978), .Z(SUM[168]) );
  NANDN U3619 ( .A(n4975), .B(n4977), .Z(n4978) );
  NANDN U3620 ( .A(n4979), .B(n4980), .Z(n4959) );
  OR U3621 ( .A(n4981), .B(n4982), .Z(n4980) );
  XOR U3622 ( .A(n4983), .B(n4984), .Z(SUM[167]) );
  NANDN U3623 ( .A(n4985), .B(n4986), .Z(n4984) );
  ANDN U3624 ( .B(n4987), .A(n4988), .Z(n4983) );
  NAND U3625 ( .A(n4989), .B(n4990), .Z(n4987) );
  XNOR U3626 ( .A(n4989), .B(n4991), .Z(SUM[166]) );
  NANDN U3627 ( .A(n4988), .B(n4990), .Z(n4991) );
  NANDN U3628 ( .A(n4992), .B(n4993), .Z(n4989) );
  NAND U3629 ( .A(n4994), .B(n4995), .Z(n4993) );
  XNOR U3630 ( .A(n4994), .B(n4996), .Z(SUM[165]) );
  NANDN U3631 ( .A(n4992), .B(n4995), .Z(n4996) );
  NANDN U3632 ( .A(n4997), .B(n4998), .Z(n4994) );
  NANDN U3633 ( .A(n4982), .B(n4999), .Z(n4998) );
  XOR U3634 ( .A(n4982), .B(n5000), .Z(SUM[164]) );
  NANDN U3635 ( .A(n4997), .B(n4999), .Z(n5000) );
  ANDN U3636 ( .B(n5001), .A(n5002), .Z(n4982) );
  NANDN U3637 ( .A(n5003), .B(n5004), .Z(n5001) );
  XOR U3638 ( .A(n5005), .B(n5006), .Z(SUM[163]) );
  NANDN U3639 ( .A(n5007), .B(n5008), .Z(n5006) );
  ANDN U3640 ( .B(n5009), .A(n5010), .Z(n5005) );
  NAND U3641 ( .A(n5011), .B(n5012), .Z(n5009) );
  XNOR U3642 ( .A(n5011), .B(n5013), .Z(SUM[162]) );
  NANDN U3643 ( .A(n5010), .B(n5012), .Z(n5013) );
  NANDN U3644 ( .A(n5014), .B(n5015), .Z(n5011) );
  NAND U3645 ( .A(n5016), .B(n5017), .Z(n5015) );
  XNOR U3646 ( .A(n5016), .B(n5018), .Z(SUM[161]) );
  NANDN U3647 ( .A(n5014), .B(n5017), .Z(n5018) );
  NANDN U3648 ( .A(n5019), .B(n5020), .Z(n5016) );
  NAND U3649 ( .A(n5004), .B(n5021), .Z(n5020) );
  XNOR U3650 ( .A(n5004), .B(n5022), .Z(SUM[160]) );
  NANDN U3651 ( .A(n5019), .B(n5021), .Z(n5022) );
  XNOR U3652 ( .A(n5023), .B(n5024), .Z(SUM[15]) );
  NANDN U3653 ( .A(n5025), .B(n5026), .Z(n5024) );
  XOR U3654 ( .A(n5027), .B(n5028), .Z(SUM[159]) );
  NANDN U3655 ( .A(n5029), .B(n5030), .Z(n5028) );
  ANDN U3656 ( .B(n5031), .A(n5032), .Z(n5027) );
  NAND U3657 ( .A(n5033), .B(n5034), .Z(n5031) );
  XNOR U3658 ( .A(n5033), .B(n5035), .Z(SUM[158]) );
  NANDN U3659 ( .A(n5032), .B(n5034), .Z(n5035) );
  NANDN U3660 ( .A(n5036), .B(n5037), .Z(n5033) );
  NAND U3661 ( .A(n5038), .B(n5039), .Z(n5037) );
  XNOR U3662 ( .A(n5038), .B(n5040), .Z(SUM[157]) );
  NANDN U3663 ( .A(n5036), .B(n5039), .Z(n5040) );
  NANDN U3664 ( .A(n5041), .B(n5042), .Z(n5038) );
  NAND U3665 ( .A(n5043), .B(n5044), .Z(n5042) );
  XNOR U3666 ( .A(n5043), .B(n5045), .Z(SUM[156]) );
  NANDN U3667 ( .A(n5041), .B(n5044), .Z(n5045) );
  NANDN U3668 ( .A(n5046), .B(n5047), .Z(n5043) );
  NAND U3669 ( .A(n5048), .B(n5049), .Z(n5047) );
  XOR U3670 ( .A(n5050), .B(n5051), .Z(SUM[155]) );
  NANDN U3671 ( .A(n5052), .B(n5053), .Z(n5051) );
  ANDN U3672 ( .B(n5054), .A(n5055), .Z(n5050) );
  NAND U3673 ( .A(n5056), .B(n5057), .Z(n5054) );
  XNOR U3674 ( .A(n5056), .B(n5058), .Z(SUM[154]) );
  NANDN U3675 ( .A(n5055), .B(n5057), .Z(n5058) );
  NANDN U3676 ( .A(n5059), .B(n5060), .Z(n5056) );
  NAND U3677 ( .A(n5061), .B(n5062), .Z(n5060) );
  XNOR U3678 ( .A(n5061), .B(n5063), .Z(SUM[153]) );
  NANDN U3679 ( .A(n5059), .B(n5062), .Z(n5063) );
  NANDN U3680 ( .A(n5064), .B(n5065), .Z(n5061) );
  NAND U3681 ( .A(n5049), .B(n5066), .Z(n5065) );
  XNOR U3682 ( .A(n5049), .B(n5067), .Z(SUM[152]) );
  NANDN U3683 ( .A(n5064), .B(n5066), .Z(n5067) );
  NANDN U3684 ( .A(n5068), .B(n5069), .Z(n5049) );
  OR U3685 ( .A(n5070), .B(n5071), .Z(n5069) );
  XOR U3686 ( .A(n5072), .B(n5073), .Z(SUM[151]) );
  NANDN U3687 ( .A(n5074), .B(n5075), .Z(n5073) );
  ANDN U3688 ( .B(n5076), .A(n5077), .Z(n5072) );
  NAND U3689 ( .A(n5078), .B(n5079), .Z(n5076) );
  XNOR U3690 ( .A(n5078), .B(n5080), .Z(SUM[150]) );
  NANDN U3691 ( .A(n5077), .B(n5079), .Z(n5080) );
  NANDN U3692 ( .A(n5081), .B(n5082), .Z(n5078) );
  NAND U3693 ( .A(n5083), .B(n5084), .Z(n5082) );
  XNOR U3694 ( .A(n5085), .B(n5086), .Z(SUM[14]) );
  NANDN U3695 ( .A(n5087), .B(n5088), .Z(n5086) );
  XNOR U3696 ( .A(n5083), .B(n5089), .Z(SUM[149]) );
  NANDN U3697 ( .A(n5081), .B(n5084), .Z(n5089) );
  NANDN U3698 ( .A(n5090), .B(n5091), .Z(n5083) );
  NANDN U3699 ( .A(n5071), .B(n5092), .Z(n5091) );
  XOR U3700 ( .A(n5071), .B(n5093), .Z(SUM[148]) );
  NANDN U3701 ( .A(n5090), .B(n5092), .Z(n5093) );
  ANDN U3702 ( .B(n5094), .A(n5095), .Z(n5071) );
  NANDN U3703 ( .A(n5096), .B(n5097), .Z(n5094) );
  XOR U3704 ( .A(n5098), .B(n5099), .Z(SUM[147]) );
  NANDN U3705 ( .A(n5100), .B(n5101), .Z(n5099) );
  ANDN U3706 ( .B(n5102), .A(n5103), .Z(n5098) );
  NAND U3707 ( .A(n5104), .B(n5105), .Z(n5102) );
  XNOR U3708 ( .A(n5104), .B(n5106), .Z(SUM[146]) );
  NANDN U3709 ( .A(n5103), .B(n5105), .Z(n5106) );
  NANDN U3710 ( .A(n5107), .B(n5108), .Z(n5104) );
  NAND U3711 ( .A(n5109), .B(n5110), .Z(n5108) );
  XNOR U3712 ( .A(n5109), .B(n5111), .Z(SUM[145]) );
  NANDN U3713 ( .A(n5107), .B(n5110), .Z(n5111) );
  NANDN U3714 ( .A(n5112), .B(n5113), .Z(n5109) );
  NAND U3715 ( .A(n5097), .B(n5114), .Z(n5113) );
  XNOR U3716 ( .A(n5097), .B(n5115), .Z(SUM[144]) );
  NANDN U3717 ( .A(n5112), .B(n5114), .Z(n5115) );
  XOR U3718 ( .A(n5116), .B(n5117), .Z(SUM[143]) );
  NANDN U3719 ( .A(n5118), .B(n5119), .Z(n5117) );
  ANDN U3720 ( .B(n5120), .A(n5121), .Z(n5116) );
  NAND U3721 ( .A(n5122), .B(n5123), .Z(n5120) );
  XNOR U3722 ( .A(n5122), .B(n5124), .Z(SUM[142]) );
  NANDN U3723 ( .A(n5121), .B(n5123), .Z(n5124) );
  NANDN U3724 ( .A(n5125), .B(n5126), .Z(n5122) );
  NAND U3725 ( .A(n5127), .B(n5128), .Z(n5126) );
  XNOR U3726 ( .A(n5127), .B(n5129), .Z(SUM[141]) );
  NANDN U3727 ( .A(n5125), .B(n5128), .Z(n5129) );
  NANDN U3728 ( .A(n5130), .B(n5131), .Z(n5127) );
  NAND U3729 ( .A(n5132), .B(n5133), .Z(n5131) );
  XNOR U3730 ( .A(n5132), .B(n5134), .Z(SUM[140]) );
  NANDN U3731 ( .A(n5130), .B(n5133), .Z(n5134) );
  NANDN U3732 ( .A(n5135), .B(n5136), .Z(n5132) );
  NAND U3733 ( .A(n5137), .B(n5138), .Z(n5136) );
  XNOR U3734 ( .A(n5139), .B(n5140), .Z(SUM[13]) );
  NANDN U3735 ( .A(n5141), .B(n5142), .Z(n5140) );
  XOR U3736 ( .A(n5143), .B(n5144), .Z(SUM[139]) );
  NANDN U3737 ( .A(n5145), .B(n5146), .Z(n5144) );
  ANDN U3738 ( .B(n5147), .A(n5148), .Z(n5143) );
  NAND U3739 ( .A(n5149), .B(n5150), .Z(n5147) );
  XNOR U3740 ( .A(n5149), .B(n5151), .Z(SUM[138]) );
  NANDN U3741 ( .A(n5148), .B(n5150), .Z(n5151) );
  NANDN U3742 ( .A(n5152), .B(n5153), .Z(n5149) );
  NAND U3743 ( .A(n5154), .B(n5155), .Z(n5153) );
  XNOR U3744 ( .A(n5154), .B(n5156), .Z(SUM[137]) );
  NANDN U3745 ( .A(n5152), .B(n5155), .Z(n5156) );
  NANDN U3746 ( .A(n5157), .B(n5158), .Z(n5154) );
  NAND U3747 ( .A(n5138), .B(n5159), .Z(n5158) );
  XNOR U3748 ( .A(n5138), .B(n5160), .Z(SUM[136]) );
  NANDN U3749 ( .A(n5157), .B(n5159), .Z(n5160) );
  NANDN U3750 ( .A(n5161), .B(n5162), .Z(n5138) );
  OR U3751 ( .A(n5163), .B(n5164), .Z(n5162) );
  XOR U3752 ( .A(n5165), .B(n5166), .Z(SUM[135]) );
  NANDN U3753 ( .A(n5167), .B(n5168), .Z(n5166) );
  ANDN U3754 ( .B(n5169), .A(n5170), .Z(n5165) );
  NAND U3755 ( .A(n5171), .B(n5172), .Z(n5169) );
  XNOR U3756 ( .A(n5171), .B(n5173), .Z(SUM[134]) );
  NANDN U3757 ( .A(n5170), .B(n5172), .Z(n5173) );
  NANDN U3758 ( .A(n5174), .B(n5175), .Z(n5171) );
  NAND U3759 ( .A(n5176), .B(n5177), .Z(n5175) );
  XNOR U3760 ( .A(n5176), .B(n5178), .Z(SUM[133]) );
  NANDN U3761 ( .A(n5174), .B(n5177), .Z(n5178) );
  NANDN U3762 ( .A(n5179), .B(n5180), .Z(n5176) );
  NANDN U3763 ( .A(n5164), .B(n5181), .Z(n5180) );
  XOR U3764 ( .A(n5164), .B(n5182), .Z(SUM[132]) );
  NANDN U3765 ( .A(n5179), .B(n5181), .Z(n5182) );
  ANDN U3766 ( .B(n5183), .A(n5184), .Z(n5164) );
  OR U3767 ( .A(n5185), .B(n5186), .Z(n5183) );
  XOR U3768 ( .A(n5187), .B(n5188), .Z(SUM[131]) );
  NANDN U3769 ( .A(n5189), .B(n5190), .Z(n5188) );
  ANDN U3770 ( .B(n5191), .A(n5192), .Z(n5187) );
  NAND U3771 ( .A(n5193), .B(n5194), .Z(n5191) );
  XNOR U3772 ( .A(n5193), .B(n5195), .Z(SUM[130]) );
  NANDN U3773 ( .A(n5192), .B(n5194), .Z(n5195) );
  NANDN U3774 ( .A(n5196), .B(n5197), .Z(n5193) );
  NAND U3775 ( .A(n5198), .B(n5199), .Z(n5197) );
  XNOR U3776 ( .A(n5200), .B(n5201), .Z(SUM[12]) );
  NANDN U3777 ( .A(n5202), .B(n5203), .Z(n5201) );
  XNOR U3778 ( .A(n5198), .B(n5204), .Z(SUM[129]) );
  NANDN U3779 ( .A(n5196), .B(n5199), .Z(n5204) );
  NANDN U3780 ( .A(n5205), .B(n5206), .Z(n5198) );
  NANDN U3781 ( .A(n5186), .B(n5207), .Z(n5206) );
  XOR U3782 ( .A(n5186), .B(n5208), .Z(SUM[128]) );
  NANDN U3783 ( .A(n5205), .B(n5207), .Z(n5208) );
  XOR U3784 ( .A(n5209), .B(n5210), .Z(SUM[127]) );
  OR U3785 ( .A(n5211), .B(n5212), .Z(n5210) );
  ANDN U3786 ( .B(n5213), .A(n5214), .Z(n5209) );
  NAND U3787 ( .A(n5215), .B(n5216), .Z(n5213) );
  XNOR U3788 ( .A(n5215), .B(n5217), .Z(SUM[126]) );
  NANDN U3789 ( .A(n5214), .B(n5216), .Z(n5217) );
  NANDN U3790 ( .A(n5218), .B(n5219), .Z(n5215) );
  NAND U3791 ( .A(n5220), .B(n5221), .Z(n5219) );
  XNOR U3792 ( .A(n5220), .B(n5222), .Z(SUM[125]) );
  NANDN U3793 ( .A(n5218), .B(n5221), .Z(n5222) );
  NANDN U3794 ( .A(n5223), .B(n5224), .Z(n5220) );
  NANDN U3795 ( .A(n5225), .B(n5226), .Z(n5224) );
  XNOR U3796 ( .A(n5226), .B(n5227), .Z(SUM[124]) );
  OR U3797 ( .A(n5225), .B(n5223), .Z(n5227) );
  NANDN U3798 ( .A(n5228), .B(n5229), .Z(n5226) );
  NANDN U3799 ( .A(n5230), .B(n5231), .Z(n5229) );
  XOR U3800 ( .A(n5232), .B(n5233), .Z(SUM[123]) );
  NANDN U3801 ( .A(n5234), .B(n5235), .Z(n5233) );
  ANDN U3802 ( .B(n5236), .A(n5237), .Z(n5232) );
  NAND U3803 ( .A(n5238), .B(n5239), .Z(n5236) );
  XNOR U3804 ( .A(n5238), .B(n5240), .Z(SUM[122]) );
  NANDN U3805 ( .A(n5237), .B(n5239), .Z(n5240) );
  NANDN U3806 ( .A(n5241), .B(n5242), .Z(n5238) );
  NAND U3807 ( .A(n5243), .B(n5244), .Z(n5242) );
  XNOR U3808 ( .A(n5243), .B(n5245), .Z(SUM[121]) );
  NANDN U3809 ( .A(n5241), .B(n5244), .Z(n5245) );
  NANDN U3810 ( .A(n5246), .B(n5247), .Z(n5243) );
  NAND U3811 ( .A(n5231), .B(n5248), .Z(n5247) );
  XNOR U3812 ( .A(n5231), .B(n5249), .Z(SUM[120]) );
  NANDN U3813 ( .A(n5246), .B(n5248), .Z(n5249) );
  NANDN U3814 ( .A(n5250), .B(n5251), .Z(n5231) );
  NANDN U3815 ( .A(n5252), .B(n5253), .Z(n5251) );
  XOR U3816 ( .A(n5254), .B(n5255), .Z(SUM[11]) );
  OR U3817 ( .A(n5256), .B(n5257), .Z(n5255) );
  ANDN U3818 ( .B(n5258), .A(n5259), .Z(n5254) );
  NANDN U3819 ( .A(n5260), .B(n5261), .Z(n5258) );
  XOR U3820 ( .A(n5262), .B(n5263), .Z(SUM[119]) );
  NANDN U3821 ( .A(n5264), .B(n5265), .Z(n5263) );
  ANDN U3822 ( .B(n5266), .A(n5267), .Z(n5262) );
  NAND U3823 ( .A(n5268), .B(n5269), .Z(n5266) );
  XNOR U3824 ( .A(n5268), .B(n5270), .Z(SUM[118]) );
  NANDN U3825 ( .A(n5267), .B(n5269), .Z(n5270) );
  NANDN U3826 ( .A(n5271), .B(n5272), .Z(n5268) );
  NAND U3827 ( .A(n5273), .B(n5274), .Z(n5272) );
  XNOR U3828 ( .A(n5273), .B(n5275), .Z(SUM[117]) );
  NANDN U3829 ( .A(n5271), .B(n5274), .Z(n5275) );
  NANDN U3830 ( .A(n5276), .B(n5277), .Z(n5273) );
  NANDN U3831 ( .A(n5252), .B(n5278), .Z(n5277) );
  XOR U3832 ( .A(n5252), .B(n5279), .Z(SUM[116]) );
  NANDN U3833 ( .A(n5276), .B(n5278), .Z(n5279) );
  ANDN U3834 ( .B(n5280), .A(n5281), .Z(n5252) );
  NANDN U3835 ( .A(n5282), .B(n5283), .Z(n5280) );
  XOR U3836 ( .A(n5284), .B(n5285), .Z(SUM[115]) );
  NANDN U3837 ( .A(n5286), .B(n5287), .Z(n5285) );
  ANDN U3838 ( .B(n5288), .A(n5289), .Z(n5284) );
  NANDN U3839 ( .A(n5290), .B(n5291), .Z(n5288) );
  XNOR U3840 ( .A(n5291), .B(n5292), .Z(SUM[114]) );
  OR U3841 ( .A(n5290), .B(n5289), .Z(n5292) );
  NANDN U3842 ( .A(n5293), .B(n5294), .Z(n5291) );
  NAND U3843 ( .A(n5295), .B(n5296), .Z(n5294) );
  XNOR U3844 ( .A(n5295), .B(n5297), .Z(SUM[113]) );
  NANDN U3845 ( .A(n5293), .B(n5296), .Z(n5297) );
  NANDN U3846 ( .A(n5298), .B(n5299), .Z(n5295) );
  NAND U3847 ( .A(n5283), .B(n5300), .Z(n5299) );
  XNOR U3848 ( .A(n5283), .B(n5301), .Z(SUM[112]) );
  NANDN U3849 ( .A(n5298), .B(n5300), .Z(n5301) );
  NANDN U3850 ( .A(n5302), .B(n5303), .Z(n5283) );
  OR U3851 ( .A(n5304), .B(n125), .Z(n5303) );
  XOR U3852 ( .A(n5305), .B(n5306), .Z(SUM[111]) );
  NANDN U3853 ( .A(n5307), .B(n5308), .Z(n5306) );
  ANDN U3854 ( .B(n5309), .A(n5310), .Z(n5305) );
  NAND U3855 ( .A(n5311), .B(n5312), .Z(n5309) );
  XNOR U3856 ( .A(n5311), .B(n5313), .Z(SUM[110]) );
  NANDN U3857 ( .A(n5310), .B(n5312), .Z(n5313) );
  NANDN U3858 ( .A(n5314), .B(n5315), .Z(n5311) );
  NAND U3859 ( .A(n5316), .B(n5317), .Z(n5315) );
  XNOR U3860 ( .A(n5261), .B(n5318), .Z(SUM[10]) );
  OR U3861 ( .A(n5260), .B(n5259), .Z(n5318) );
  NANDN U3862 ( .A(n3), .B(n5319), .Z(n5261) );
  NANDN U3863 ( .A(n1), .B(n4), .Z(n5319) );
  ANDN U3864 ( .B(n5320), .A(n591), .Z(n1) );
  XNOR U3865 ( .A(n5316), .B(n5321), .Z(SUM[109]) );
  NANDN U3866 ( .A(n5314), .B(n5317), .Z(n5321) );
  NANDN U3867 ( .A(n5322), .B(n5323), .Z(n5316) );
  NAND U3868 ( .A(n5324), .B(n5325), .Z(n5323) );
  XNOR U3869 ( .A(n5324), .B(n5326), .Z(SUM[108]) );
  NANDN U3870 ( .A(n5322), .B(n5325), .Z(n5326) );
  NANDN U3871 ( .A(n5327), .B(n5328), .Z(n5324) );
  NAND U3872 ( .A(n5329), .B(n5330), .Z(n5328) );
  XOR U3873 ( .A(n5331), .B(n5332), .Z(SUM[107]) );
  NANDN U3874 ( .A(n5333), .B(n5334), .Z(n5332) );
  ANDN U3875 ( .B(n5335), .A(n5336), .Z(n5331) );
  NAND U3876 ( .A(n5337), .B(n5338), .Z(n5335) );
  XNOR U3877 ( .A(n5337), .B(n5339), .Z(SUM[106]) );
  NANDN U3878 ( .A(n5336), .B(n5338), .Z(n5339) );
  NANDN U3879 ( .A(n5340), .B(n5341), .Z(n5337) );
  NAND U3880 ( .A(n5342), .B(n5343), .Z(n5341) );
  XNOR U3881 ( .A(n5342), .B(n5344), .Z(SUM[105]) );
  NANDN U3882 ( .A(n5340), .B(n5343), .Z(n5344) );
  NANDN U3883 ( .A(n5345), .B(n5346), .Z(n5342) );
  NAND U3884 ( .A(n5330), .B(n5347), .Z(n5346) );
  XNOR U3885 ( .A(n5330), .B(n5348), .Z(SUM[104]) );
  NANDN U3886 ( .A(n5345), .B(n5347), .Z(n5348) );
  NANDN U3887 ( .A(n5349), .B(n5350), .Z(n5330) );
  OR U3888 ( .A(n5351), .B(n5352), .Z(n5350) );
  XOR U3889 ( .A(n5353), .B(n5354), .Z(SUM[103]) );
  NANDN U3890 ( .A(n5355), .B(n5356), .Z(n5354) );
  ANDN U3891 ( .B(n5357), .A(n5358), .Z(n5353) );
  NAND U3892 ( .A(n5359), .B(n5360), .Z(n5357) );
  XNOR U3893 ( .A(n5359), .B(n5361), .Z(SUM[102]) );
  NANDN U3894 ( .A(n5358), .B(n5360), .Z(n5361) );
  NANDN U3895 ( .A(n5362), .B(n5363), .Z(n5359) );
  NAND U3896 ( .A(n5364), .B(n5365), .Z(n5363) );
  XOR U3897 ( .A(n5366), .B(n5367), .Z(SUM[1022]) );
  XNOR U3898 ( .A(B[1022]), .B(A[1022]), .Z(n5367) );
  ANDN U3899 ( .B(n5368), .A(n5369), .Z(n5366) );
  NAND U3900 ( .A(n5370), .B(n5371), .Z(n5368) );
  XNOR U3901 ( .A(n5370), .B(n5372), .Z(SUM[1021]) );
  NANDN U3902 ( .A(n5369), .B(n5371), .Z(n5372) );
  OR U3903 ( .A(B[1021]), .B(A[1021]), .Z(n5371) );
  AND U3904 ( .A(B[1021]), .B(A[1021]), .Z(n5369) );
  NANDN U3905 ( .A(n5373), .B(n5374), .Z(n5370) );
  NAND U3906 ( .A(n5375), .B(n5376), .Z(n5374) );
  XNOR U3907 ( .A(n5375), .B(n5377), .Z(SUM[1020]) );
  NANDN U3908 ( .A(n5373), .B(n5376), .Z(n5377) );
  OR U3909 ( .A(B[1020]), .B(A[1020]), .Z(n5376) );
  AND U3910 ( .A(B[1020]), .B(A[1020]), .Z(n5373) );
  NANDN U3911 ( .A(n5378), .B(n5379), .Z(n5375) );
  NAND U3912 ( .A(n5380), .B(n5381), .Z(n5379) );
  XNOR U3913 ( .A(n5364), .B(n5382), .Z(SUM[101]) );
  NANDN U3914 ( .A(n5362), .B(n5365), .Z(n5382) );
  NANDN U3915 ( .A(n5383), .B(n5384), .Z(n5364) );
  NANDN U3916 ( .A(n5352), .B(n5385), .Z(n5384) );
  XNOR U3917 ( .A(n5380), .B(n5386), .Z(SUM[1019]) );
  NANDN U3918 ( .A(n5378), .B(n5381), .Z(n5386) );
  OR U3919 ( .A(B[1019]), .B(A[1019]), .Z(n5381) );
  AND U3920 ( .A(B[1019]), .B(A[1019]), .Z(n5378) );
  NANDN U3921 ( .A(n5387), .B(n5388), .Z(n5380) );
  NAND U3922 ( .A(n5389), .B(n5390), .Z(n5388) );
  XNOR U3923 ( .A(n5389), .B(n5391), .Z(SUM[1018]) );
  NANDN U3924 ( .A(n5387), .B(n5390), .Z(n5391) );
  OR U3925 ( .A(B[1018]), .B(A[1018]), .Z(n5390) );
  AND U3926 ( .A(B[1018]), .B(A[1018]), .Z(n5387) );
  NANDN U3927 ( .A(n5392), .B(n5393), .Z(n5389) );
  NAND U3928 ( .A(n5394), .B(n5395), .Z(n5393) );
  XNOR U3929 ( .A(n5394), .B(n5396), .Z(SUM[1017]) );
  NANDN U3930 ( .A(n5392), .B(n5395), .Z(n5396) );
  OR U3931 ( .A(B[1017]), .B(A[1017]), .Z(n5395) );
  AND U3932 ( .A(B[1017]), .B(A[1017]), .Z(n5392) );
  NANDN U3933 ( .A(n5397), .B(n5398), .Z(n5394) );
  NAND U3934 ( .A(n5399), .B(n5400), .Z(n5398) );
  XNOR U3935 ( .A(n5399), .B(n5401), .Z(SUM[1016]) );
  NANDN U3936 ( .A(n5397), .B(n5400), .Z(n5401) );
  OR U3937 ( .A(B[1016]), .B(A[1016]), .Z(n5400) );
  AND U3938 ( .A(B[1016]), .B(A[1016]), .Z(n5397) );
  NANDN U3939 ( .A(n5402), .B(n5403), .Z(n5399) );
  NAND U3940 ( .A(n5404), .B(n5405), .Z(n5403) );
  XNOR U3941 ( .A(n5404), .B(n5406), .Z(SUM[1015]) );
  NANDN U3942 ( .A(n5402), .B(n5405), .Z(n5406) );
  OR U3943 ( .A(B[1015]), .B(A[1015]), .Z(n5405) );
  AND U3944 ( .A(B[1015]), .B(A[1015]), .Z(n5402) );
  NANDN U3945 ( .A(n5407), .B(n5408), .Z(n5404) );
  NAND U3946 ( .A(n5409), .B(n5410), .Z(n5408) );
  XNOR U3947 ( .A(n5409), .B(n5411), .Z(SUM[1014]) );
  NANDN U3948 ( .A(n5407), .B(n5410), .Z(n5411) );
  OR U3949 ( .A(B[1014]), .B(A[1014]), .Z(n5410) );
  AND U3950 ( .A(B[1014]), .B(A[1014]), .Z(n5407) );
  NANDN U3951 ( .A(n5412), .B(n5413), .Z(n5409) );
  NAND U3952 ( .A(n5414), .B(n5415), .Z(n5413) );
  XNOR U3953 ( .A(n5414), .B(n5416), .Z(SUM[1013]) );
  NANDN U3954 ( .A(n5412), .B(n5415), .Z(n5416) );
  OR U3955 ( .A(B[1013]), .B(A[1013]), .Z(n5415) );
  AND U3956 ( .A(B[1013]), .B(A[1013]), .Z(n5412) );
  NANDN U3957 ( .A(n5417), .B(n5418), .Z(n5414) );
  NAND U3958 ( .A(n5419), .B(n5420), .Z(n5418) );
  XNOR U3959 ( .A(n5419), .B(n5421), .Z(SUM[1012]) );
  NANDN U3960 ( .A(n5417), .B(n5420), .Z(n5421) );
  OR U3961 ( .A(B[1012]), .B(A[1012]), .Z(n5420) );
  AND U3962 ( .A(B[1012]), .B(A[1012]), .Z(n5417) );
  NANDN U3963 ( .A(n5422), .B(n5423), .Z(n5419) );
  NAND U3964 ( .A(n5424), .B(n5425), .Z(n5423) );
  XNOR U3965 ( .A(n5424), .B(n5426), .Z(SUM[1011]) );
  NANDN U3966 ( .A(n5422), .B(n5425), .Z(n5426) );
  OR U3967 ( .A(B[1011]), .B(A[1011]), .Z(n5425) );
  AND U3968 ( .A(B[1011]), .B(A[1011]), .Z(n5422) );
  NANDN U3969 ( .A(n5427), .B(n5428), .Z(n5424) );
  NAND U3970 ( .A(n5429), .B(n5430), .Z(n5428) );
  XNOR U3971 ( .A(n5429), .B(n5431), .Z(SUM[1010]) );
  NANDN U3972 ( .A(n5427), .B(n5430), .Z(n5431) );
  OR U3973 ( .A(B[1010]), .B(A[1010]), .Z(n5430) );
  AND U3974 ( .A(B[1010]), .B(A[1010]), .Z(n5427) );
  NANDN U3975 ( .A(n5432), .B(n5433), .Z(n5429) );
  NAND U3976 ( .A(n5434), .B(n5435), .Z(n5433) );
  XOR U3977 ( .A(n5352), .B(n5436), .Z(SUM[100]) );
  NANDN U3978 ( .A(n5383), .B(n5385), .Z(n5436) );
  ANDN U3979 ( .B(n5437), .A(n5438), .Z(n5352) );
  OR U3980 ( .A(n5439), .B(n125), .Z(n5437) );
  ANDN U3981 ( .B(n5440), .A(n5441), .Z(n125) );
  OR U3982 ( .A(n890), .B(n5442), .Z(n5440) );
  ANDN U3983 ( .B(n5443), .A(n5444), .Z(n890) );
  XNOR U3984 ( .A(n5434), .B(n5445), .Z(SUM[1009]) );
  NANDN U3985 ( .A(n5432), .B(n5435), .Z(n5445) );
  OR U3986 ( .A(B[1009]), .B(A[1009]), .Z(n5435) );
  AND U3987 ( .A(B[1009]), .B(A[1009]), .Z(n5432) );
  NANDN U3988 ( .A(n5446), .B(n5447), .Z(n5434) );
  NAND U3989 ( .A(n5448), .B(n5449), .Z(n5447) );
  XNOR U3990 ( .A(n5448), .B(n5450), .Z(SUM[1008]) );
  NANDN U3991 ( .A(n5446), .B(n5449), .Z(n5450) );
  OR U3992 ( .A(B[1008]), .B(A[1008]), .Z(n5449) );
  AND U3993 ( .A(B[1008]), .B(A[1008]), .Z(n5446) );
  NANDN U3994 ( .A(n5451), .B(n5452), .Z(n5448) );
  NANDN U3995 ( .A(n5453), .B(n5454), .Z(n5452) );
  NANDN U3996 ( .A(n5455), .B(n5456), .Z(n5454) );
  NANDN U3997 ( .A(n5457), .B(n5458), .Z(n5456) );
  NANDN U3998 ( .A(n5459), .B(n5460), .Z(n5458) );
  NANDN U3999 ( .A(n5461), .B(n5462), .Z(n5460) );
  NANDN U4000 ( .A(n5463), .B(n5464), .Z(n5462) );
  NANDN U4001 ( .A(n5465), .B(n5466), .Z(n5464) );
  NANDN U4002 ( .A(n5467), .B(n5468), .Z(n5466) );
  NANDN U4003 ( .A(n5469), .B(n5470), .Z(n5468) );
  NANDN U4004 ( .A(n5471), .B(n5472), .Z(n5470) );
  AND U4005 ( .A(n5473), .B(n5474), .Z(n5472) );
  OR U4006 ( .A(n5475), .B(n5476), .Z(n5474) );
  OR U4007 ( .A(n5475), .B(n5477), .Z(n5473) );
  XOR U4008 ( .A(n5478), .B(n5479), .Z(SUM[1007]) );
  OR U4009 ( .A(n5453), .B(n5451), .Z(n5479) );
  AND U4010 ( .A(B[1007]), .B(A[1007]), .Z(n5451) );
  NOR U4011 ( .A(B[1007]), .B(A[1007]), .Z(n5453) );
  ANDN U4012 ( .B(n5480), .A(n5455), .Z(n5478) );
  NANDN U4013 ( .A(n5457), .B(n5481), .Z(n5480) );
  XNOR U4014 ( .A(n5481), .B(n5482), .Z(SUM[1006]) );
  OR U4015 ( .A(n5457), .B(n5455), .Z(n5482) );
  AND U4016 ( .A(B[1006]), .B(A[1006]), .Z(n5455) );
  NOR U4017 ( .A(B[1006]), .B(A[1006]), .Z(n5457) );
  NANDN U4018 ( .A(n5459), .B(n5483), .Z(n5481) );
  NANDN U4019 ( .A(n5461), .B(n5484), .Z(n5483) );
  XNOR U4020 ( .A(n5484), .B(n5485), .Z(SUM[1005]) );
  OR U4021 ( .A(n5461), .B(n5459), .Z(n5485) );
  AND U4022 ( .A(B[1005]), .B(A[1005]), .Z(n5459) );
  NOR U4023 ( .A(B[1005]), .B(A[1005]), .Z(n5461) );
  NANDN U4024 ( .A(n5463), .B(n5486), .Z(n5484) );
  NANDN U4025 ( .A(n5465), .B(n5487), .Z(n5486) );
  XNOR U4026 ( .A(n5487), .B(n5488), .Z(SUM[1004]) );
  OR U4027 ( .A(n5465), .B(n5463), .Z(n5488) );
  AND U4028 ( .A(B[1004]), .B(A[1004]), .Z(n5463) );
  NOR U4029 ( .A(B[1004]), .B(A[1004]), .Z(n5465) );
  NANDN U4030 ( .A(n5467), .B(n5489), .Z(n5487) );
  NANDN U4031 ( .A(n5469), .B(n5490), .Z(n5489) );
  NAND U4032 ( .A(n5491), .B(n5492), .Z(n5469) );
  AND U4033 ( .A(n5493), .B(n5494), .Z(n5492) );
  AND U4034 ( .A(n5495), .B(n5496), .Z(n5491) );
  NANDN U4035 ( .A(n5497), .B(n5498), .Z(n5467) );
  NAND U4036 ( .A(n5499), .B(n5496), .Z(n5498) );
  NANDN U4037 ( .A(n5500), .B(n5501), .Z(n5499) );
  NAND U4038 ( .A(n5502), .B(n5495), .Z(n5501) );
  NANDN U4039 ( .A(n5503), .B(n5504), .Z(n5502) );
  NAND U4040 ( .A(n5494), .B(n5505), .Z(n5504) );
  XOR U4041 ( .A(n5506), .B(n5507), .Z(SUM[1003]) );
  NANDN U4042 ( .A(n5497), .B(n5496), .Z(n5507) );
  OR U4043 ( .A(B[1003]), .B(A[1003]), .Z(n5496) );
  AND U4044 ( .A(B[1003]), .B(A[1003]), .Z(n5497) );
  ANDN U4045 ( .B(n5508), .A(n5500), .Z(n5506) );
  NAND U4046 ( .A(n5509), .B(n5495), .Z(n5508) );
  XNOR U4047 ( .A(n5509), .B(n5510), .Z(SUM[1002]) );
  NANDN U4048 ( .A(n5500), .B(n5495), .Z(n5510) );
  OR U4049 ( .A(B[1002]), .B(A[1002]), .Z(n5495) );
  AND U4050 ( .A(B[1002]), .B(A[1002]), .Z(n5500) );
  NANDN U4051 ( .A(n5503), .B(n5511), .Z(n5509) );
  NAND U4052 ( .A(n5512), .B(n5494), .Z(n5511) );
  XNOR U4053 ( .A(n5512), .B(n5513), .Z(SUM[1001]) );
  NANDN U4054 ( .A(n5503), .B(n5494), .Z(n5513) );
  OR U4055 ( .A(B[1001]), .B(A[1001]), .Z(n5494) );
  AND U4056 ( .A(B[1001]), .B(A[1001]), .Z(n5503) );
  NANDN U4057 ( .A(n5505), .B(n5514), .Z(n5512) );
  NAND U4058 ( .A(n5490), .B(n5493), .Z(n5514) );
  XNOR U4059 ( .A(n5490), .B(n5515), .Z(SUM[1000]) );
  NANDN U4060 ( .A(n5505), .B(n5493), .Z(n5515) );
  OR U4061 ( .A(B[1000]), .B(A[1000]), .Z(n5493) );
  AND U4062 ( .A(B[1000]), .B(A[1000]), .Z(n5505) );
  NANDN U4063 ( .A(n5471), .B(n5516), .Z(n5490) );
  OR U4064 ( .A(n5475), .B(n29), .Z(n5516) );
  AND U4065 ( .A(n5477), .B(n5476), .Z(n29) );
  ANDN U4066 ( .B(n5517), .A(n34), .Z(n5476) );
  AND U4067 ( .A(B[995]), .B(A[995]), .Z(n34) );
  NAND U4068 ( .A(n5518), .B(n35), .Z(n5517) );
  NANDN U4069 ( .A(n37), .B(n5519), .Z(n5518) );
  NAND U4070 ( .A(n5520), .B(n39), .Z(n5519) );
  NANDN U4071 ( .A(n41), .B(n5521), .Z(n5520) );
  NAND U4072 ( .A(n44), .B(n46), .Z(n5521) );
  AND U4073 ( .A(B[992]), .B(A[992]), .Z(n46) );
  AND U4074 ( .A(B[993]), .B(A[993]), .Z(n41) );
  AND U4075 ( .A(B[994]), .B(A[994]), .Z(n37) );
  NAND U4076 ( .A(n5522), .B(n5523), .Z(n5477) );
  AND U4077 ( .A(n44), .B(n5524), .Z(n5523) );
  AND U4078 ( .A(n35), .B(n39), .Z(n5524) );
  OR U4079 ( .A(B[994]), .B(A[994]), .Z(n39) );
  OR U4080 ( .A(B[995]), .B(A[995]), .Z(n35) );
  OR U4081 ( .A(B[993]), .B(A[993]), .Z(n44) );
  NOR U4082 ( .A(n48), .B(n49), .Z(n5522) );
  NOR U4083 ( .A(B[992]), .B(A[992]), .Z(n49) );
  ANDN U4084 ( .B(n5525), .A(n54), .Z(n48) );
  AND U4085 ( .A(B[991]), .B(A[991]), .Z(n54) );
  NANDN U4086 ( .A(n53), .B(n5526), .Z(n5525) );
  NANDN U4087 ( .A(n56), .B(n5527), .Z(n5526) );
  NANDN U4088 ( .A(n57), .B(n5528), .Z(n5527) );
  NANDN U4089 ( .A(n60), .B(n5529), .Z(n5528) );
  NANDN U4090 ( .A(n62), .B(n5530), .Z(n5529) );
  NANDN U4091 ( .A(n70), .B(n5531), .Z(n5530) );
  NANDN U4092 ( .A(n72), .B(n5532), .Z(n5531) );
  NANDN U4093 ( .A(n75), .B(n5533), .Z(n5532) );
  NANDN U4094 ( .A(n77), .B(n5534), .Z(n5533) );
  NANDN U4095 ( .A(n97), .B(n5535), .Z(n5534) );
  AND U4096 ( .A(n5536), .B(n5537), .Z(n5535) );
  NANDN U4097 ( .A(n99), .B(n119), .Z(n5537) );
  NANDN U4098 ( .A(n128), .B(n5538), .Z(n119) );
  NAND U4099 ( .A(n5539), .B(n129), .Z(n5538) );
  NANDN U4100 ( .A(n131), .B(n5540), .Z(n5539) );
  NAND U4101 ( .A(n5541), .B(n133), .Z(n5540) );
  NANDN U4102 ( .A(n135), .B(n5542), .Z(n5541) );
  NAND U4103 ( .A(n138), .B(n140), .Z(n5542) );
  AND U4104 ( .A(A[976]), .B(B[976]), .Z(n140) );
  AND U4105 ( .A(A[977]), .B(B[977]), .Z(n135) );
  AND U4106 ( .A(A[978]), .B(B[978]), .Z(n131) );
  AND U4107 ( .A(B[979]), .B(A[979]), .Z(n128) );
  NANDN U4108 ( .A(n99), .B(n120), .Z(n5536) );
  AND U4109 ( .A(n5543), .B(n5544), .Z(n120) );
  AND U4110 ( .A(n138), .B(n5545), .Z(n5544) );
  NOR U4111 ( .A(n142), .B(n143), .Z(n5545) );
  NOR U4112 ( .A(B[976]), .B(A[976]), .Z(n143) );
  ANDN U4113 ( .B(n5546), .A(n148), .Z(n142) );
  AND U4114 ( .A(B[975]), .B(A[975]), .Z(n148) );
  NANDN U4115 ( .A(n147), .B(n5547), .Z(n5546) );
  NANDN U4116 ( .A(n150), .B(n5548), .Z(n5547) );
  NANDN U4117 ( .A(n151), .B(n5549), .Z(n5548) );
  NANDN U4118 ( .A(n154), .B(n5550), .Z(n5549) );
  NANDN U4119 ( .A(n156), .B(n5551), .Z(n5550) );
  NANDN U4120 ( .A(n159), .B(n5552), .Z(n5551) );
  NANDN U4121 ( .A(n161), .B(n5553), .Z(n5552) );
  NANDN U4122 ( .A(n164), .B(n5554), .Z(n5553) );
  NANDN U4123 ( .A(n166), .B(n5555), .Z(n5554) );
  NANDN U4124 ( .A(n187), .B(n5556), .Z(n5555) );
  AND U4125 ( .A(n5557), .B(n5558), .Z(n5556) );
  NANDN U4126 ( .A(n189), .B(n209), .Z(n5558) );
  NANDN U4127 ( .A(n213), .B(n5559), .Z(n209) );
  NAND U4128 ( .A(n5560), .B(n214), .Z(n5559) );
  NANDN U4129 ( .A(n216), .B(n5561), .Z(n5560) );
  NAND U4130 ( .A(n5562), .B(n218), .Z(n5561) );
  NANDN U4131 ( .A(n220), .B(n5563), .Z(n5562) );
  NAND U4132 ( .A(n223), .B(n225), .Z(n5563) );
  AND U4133 ( .A(A[960]), .B(B[960]), .Z(n225) );
  AND U4134 ( .A(A[961]), .B(B[961]), .Z(n220) );
  AND U4135 ( .A(A[962]), .B(B[962]), .Z(n216) );
  AND U4136 ( .A(B[963]), .B(A[963]), .Z(n213) );
  NANDN U4137 ( .A(n189), .B(n210), .Z(n5557) );
  AND U4138 ( .A(n5564), .B(n5565), .Z(n210) );
  AND U4139 ( .A(n223), .B(n5566), .Z(n5565) );
  NOR U4140 ( .A(n227), .B(n228), .Z(n5566) );
  NOR U4141 ( .A(B[960]), .B(A[960]), .Z(n228) );
  ANDN U4142 ( .B(n5567), .A(n241), .Z(n227) );
  AND U4143 ( .A(B[959]), .B(A[959]), .Z(n241) );
  NANDN U4144 ( .A(n240), .B(n5568), .Z(n5567) );
  NANDN U4145 ( .A(n243), .B(n5569), .Z(n5568) );
  NANDN U4146 ( .A(n244), .B(n5570), .Z(n5569) );
  NANDN U4147 ( .A(n247), .B(n5571), .Z(n5570) );
  NANDN U4148 ( .A(n249), .B(n5572), .Z(n5571) );
  NAND U4149 ( .A(n5573), .B(n5574), .Z(n5572) );
  NAND U4150 ( .A(n5575), .B(n5576), .Z(n5574) );
  AND U4151 ( .A(n282), .B(n5577), .Z(n5576) );
  ANDN U4152 ( .B(n255), .A(n309), .Z(n5577) );
  ANDN U4153 ( .B(n5578), .A(n331), .Z(n309) );
  AND U4154 ( .A(B[943]), .B(A[943]), .Z(n331) );
  NANDN U4155 ( .A(n330), .B(n5579), .Z(n5578) );
  NANDN U4156 ( .A(n333), .B(n5580), .Z(n5579) );
  NANDN U4157 ( .A(n334), .B(n5581), .Z(n5580) );
  NANDN U4158 ( .A(n337), .B(n5582), .Z(n5581) );
  NANDN U4159 ( .A(n339), .B(n5583), .Z(n5582) );
  NAND U4160 ( .A(n5584), .B(n5585), .Z(n5583) );
  NAND U4161 ( .A(n5586), .B(n5587), .Z(n5585) );
  AND U4162 ( .A(n377), .B(n5588), .Z(n5587) );
  ANDN U4163 ( .B(n345), .A(n399), .Z(n5588) );
  ANDN U4164 ( .B(n5589), .A(n426), .Z(n399) );
  AND U4165 ( .A(B[927]), .B(A[927]), .Z(n426) );
  NANDN U4166 ( .A(n425), .B(n5590), .Z(n5589) );
  NANDN U4167 ( .A(n428), .B(n5591), .Z(n5590) );
  NANDN U4168 ( .A(n429), .B(n5592), .Z(n5591) );
  NANDN U4169 ( .A(n432), .B(n5593), .Z(n5592) );
  NANDN U4170 ( .A(n434), .B(n5594), .Z(n5593) );
  NAND U4171 ( .A(n5595), .B(n5596), .Z(n5594) );
  NAND U4172 ( .A(n5597), .B(n5598), .Z(n5596) );
  AND U4173 ( .A(n467), .B(n5599), .Z(n5598) );
  ANDN U4174 ( .B(n440), .A(n497), .Z(n5599) );
  ANDN U4175 ( .B(n5600), .A(n519), .Z(n497) );
  AND U4176 ( .A(B[911]), .B(A[911]), .Z(n519) );
  NANDN U4177 ( .A(n518), .B(n5601), .Z(n5600) );
  NANDN U4178 ( .A(n521), .B(n5602), .Z(n5601) );
  NANDN U4179 ( .A(n522), .B(n5603), .Z(n5602) );
  NANDN U4180 ( .A(n525), .B(n5604), .Z(n5603) );
  NANDN U4181 ( .A(n527), .B(n5605), .Z(n5604) );
  NAND U4182 ( .A(n5606), .B(n5607), .Z(n5605) );
  NAND U4183 ( .A(n5608), .B(n5609), .Z(n5607) );
  AND U4184 ( .A(n565), .B(n5610), .Z(n5609) );
  ANDN U4185 ( .B(n538), .A(n587), .Z(n5610) );
  ANDN U4186 ( .B(n5611), .A(n617), .Z(n587) );
  AND U4187 ( .A(B[895]), .B(A[895]), .Z(n617) );
  NANDN U4188 ( .A(n616), .B(n5612), .Z(n5611) );
  NANDN U4189 ( .A(n619), .B(n5613), .Z(n5612) );
  NANDN U4190 ( .A(n620), .B(n5614), .Z(n5613) );
  NANDN U4191 ( .A(n623), .B(n5615), .Z(n5614) );
  NANDN U4192 ( .A(n625), .B(n5616), .Z(n5615) );
  NAND U4193 ( .A(n5617), .B(n5618), .Z(n5616) );
  NAND U4194 ( .A(n5619), .B(n5620), .Z(n5618) );
  AND U4195 ( .A(n663), .B(n5621), .Z(n5620) );
  ANDN U4196 ( .B(n631), .A(n685), .Z(n5621) );
  ANDN U4197 ( .B(n5622), .A(n715), .Z(n685) );
  AND U4198 ( .A(B[879]), .B(A[879]), .Z(n715) );
  NANDN U4199 ( .A(n714), .B(n5623), .Z(n5622) );
  NANDN U4200 ( .A(n717), .B(n5624), .Z(n5623) );
  NANDN U4201 ( .A(n718), .B(n5625), .Z(n5624) );
  NANDN U4202 ( .A(n721), .B(n5626), .Z(n5625) );
  NANDN U4203 ( .A(n723), .B(n5627), .Z(n5626) );
  NAND U4204 ( .A(n5628), .B(n5629), .Z(n5627) );
  NAND U4205 ( .A(n5630), .B(n5631), .Z(n5629) );
  AND U4206 ( .A(n756), .B(n5632), .Z(n5631) );
  ANDN U4207 ( .B(n729), .A(n783), .Z(n5632) );
  ANDN U4208 ( .B(n5633), .A(n805), .Z(n783) );
  AND U4209 ( .A(B[863]), .B(A[863]), .Z(n805) );
  NANDN U4210 ( .A(n804), .B(n5634), .Z(n5633) );
  NANDN U4211 ( .A(n807), .B(n5635), .Z(n5634) );
  NANDN U4212 ( .A(n808), .B(n5636), .Z(n5635) );
  NANDN U4213 ( .A(n811), .B(n5637), .Z(n5636) );
  NANDN U4214 ( .A(n813), .B(n5638), .Z(n5637) );
  NAND U4215 ( .A(n5639), .B(n5640), .Z(n5638) );
  NAND U4216 ( .A(n5641), .B(n5642), .Z(n5640) );
  AND U4217 ( .A(n850), .B(n5643), .Z(n5642) );
  ANDN U4218 ( .B(n819), .A(n872), .Z(n5643) );
  ANDN U4219 ( .B(n5644), .A(n899), .Z(n872) );
  AND U4220 ( .A(B[847]), .B(A[847]), .Z(n899) );
  NANDN U4221 ( .A(n898), .B(n5645), .Z(n5644) );
  NANDN U4222 ( .A(n901), .B(n5646), .Z(n5645) );
  NANDN U4223 ( .A(n902), .B(n5647), .Z(n5646) );
  NANDN U4224 ( .A(n905), .B(n5648), .Z(n5647) );
  NANDN U4225 ( .A(n907), .B(n5649), .Z(n5648) );
  NAND U4226 ( .A(n5650), .B(n5651), .Z(n5649) );
  NAND U4227 ( .A(n5652), .B(n5653), .Z(n5651) );
  AND U4228 ( .A(n940), .B(n5654), .Z(n5653) );
  ANDN U4229 ( .B(n913), .A(n970), .Z(n5654) );
  ANDN U4230 ( .B(n5655), .A(n992), .Z(n970) );
  AND U4231 ( .A(B[831]), .B(A[831]), .Z(n992) );
  NANDN U4232 ( .A(n991), .B(n5656), .Z(n5655) );
  NANDN U4233 ( .A(n994), .B(n5657), .Z(n5656) );
  NANDN U4234 ( .A(n995), .B(n5658), .Z(n5657) );
  NANDN U4235 ( .A(n998), .B(n5659), .Z(n5658) );
  NANDN U4236 ( .A(n1000), .B(n5660), .Z(n5659) );
  NAND U4237 ( .A(n5661), .B(n5662), .Z(n5660) );
  NAND U4238 ( .A(n5663), .B(n5664), .Z(n5662) );
  AND U4239 ( .A(n1038), .B(n5665), .Z(n5664) );
  ANDN U4240 ( .B(n1011), .A(n1060), .Z(n5665) );
  ANDN U4241 ( .B(n5666), .A(n1086), .Z(n1060) );
  AND U4242 ( .A(B[815]), .B(A[815]), .Z(n1086) );
  NANDN U4243 ( .A(n1085), .B(n5667), .Z(n5666) );
  NANDN U4244 ( .A(n1088), .B(n5668), .Z(n5667) );
  NANDN U4245 ( .A(n1089), .B(n5669), .Z(n5668) );
  NANDN U4246 ( .A(n1092), .B(n5670), .Z(n5669) );
  NANDN U4247 ( .A(n1094), .B(n5671), .Z(n5670) );
  NAND U4248 ( .A(n5672), .B(n5673), .Z(n5671) );
  NAND U4249 ( .A(n5674), .B(n5675), .Z(n5673) );
  AND U4250 ( .A(n1128), .B(n5676), .Z(n5675) );
  ANDN U4251 ( .B(n1100), .A(n1150), .Z(n5676) );
  ANDN U4252 ( .B(n5677), .A(n1186), .Z(n1150) );
  AND U4253 ( .A(B[799]), .B(A[799]), .Z(n1186) );
  NANDN U4254 ( .A(n1185), .B(n5678), .Z(n5677) );
  NANDN U4255 ( .A(n1188), .B(n5679), .Z(n5678) );
  NANDN U4256 ( .A(n1189), .B(n5680), .Z(n5679) );
  NANDN U4257 ( .A(n1192), .B(n5681), .Z(n5680) );
  NANDN U4258 ( .A(n1194), .B(n5682), .Z(n5681) );
  NAND U4259 ( .A(n5683), .B(n5684), .Z(n5682) );
  NAND U4260 ( .A(n5685), .B(n5686), .Z(n5684) );
  AND U4261 ( .A(n1227), .B(n5687), .Z(n5686) );
  ANDN U4262 ( .B(n1200), .A(n1254), .Z(n5687) );
  ANDN U4263 ( .B(n5688), .A(n1276), .Z(n1254) );
  AND U4264 ( .A(B[783]), .B(A[783]), .Z(n1276) );
  NANDN U4265 ( .A(n1275), .B(n5689), .Z(n5688) );
  NANDN U4266 ( .A(n1278), .B(n5690), .Z(n5689) );
  NANDN U4267 ( .A(n1279), .B(n5691), .Z(n5690) );
  NANDN U4268 ( .A(n1282), .B(n5692), .Z(n5691) );
  NANDN U4269 ( .A(n1284), .B(n5693), .Z(n5692) );
  NAND U4270 ( .A(n5694), .B(n5695), .Z(n5693) );
  NAND U4271 ( .A(n5696), .B(n5697), .Z(n5695) );
  AND U4272 ( .A(n1322), .B(n5698), .Z(n5697) );
  ANDN U4273 ( .B(n1290), .A(n1344), .Z(n5698) );
  ANDN U4274 ( .B(n5699), .A(n1371), .Z(n1344) );
  AND U4275 ( .A(B[767]), .B(A[767]), .Z(n1371) );
  NANDN U4276 ( .A(n1370), .B(n5700), .Z(n5699) );
  NAND U4277 ( .A(n5701), .B(n5702), .Z(n5700) );
  NAND U4278 ( .A(n5703), .B(n5704), .Z(n5702) );
  AND U4279 ( .A(n5705), .B(n5706), .Z(n5704) );
  ANDN U4280 ( .B(n1380), .A(n1384), .Z(n5706) );
  AND U4281 ( .A(n1375), .B(n5707), .Z(n5705) );
  NANDN U4282 ( .A(n1461), .B(n5708), .Z(n5707) );
  NANDN U4283 ( .A(n1463), .B(n5709), .Z(n5708) );
  NANDN U4284 ( .A(n1558), .B(n5710), .Z(n5709) );
  NANDN U4285 ( .A(n1560), .B(n5711), .Z(n5710) );
  NANDN U4286 ( .A(n1651), .B(n5712), .Z(n5711) );
  NANDN U4287 ( .A(n1653), .B(n5713), .Z(n5712) );
  NANDN U4288 ( .A(n1752), .B(n5714), .Z(n5713) );
  NANDN U4289 ( .A(n1754), .B(n5715), .Z(n5714) );
  NANDN U4290 ( .A(n2134), .B(n5716), .Z(n5715) );
  AND U4291 ( .A(n5717), .B(n5718), .Z(n5716) );
  NANDN U4292 ( .A(n2136), .B(n2530), .Z(n5718) );
  NAND U4293 ( .A(n5719), .B(n5720), .Z(n2530) );
  NAND U4294 ( .A(n5721), .B(n2535), .Z(n5720) );
  NANDN U4295 ( .A(n2537), .B(n5722), .Z(n5721) );
  NAND U4296 ( .A(n5723), .B(n2539), .Z(n5722) );
  NANDN U4297 ( .A(n2541), .B(n5724), .Z(n5723) );
  NAND U4298 ( .A(n5725), .B(n2544), .Z(n5724) );
  NANDN U4299 ( .A(n2546), .B(n5726), .Z(n5725) );
  NAND U4300 ( .A(n5727), .B(n2549), .Z(n5726) );
  NANDN U4301 ( .A(n2551), .B(n5728), .Z(n5727) );
  NANDN U4302 ( .A(n2553), .B(n5729), .Z(n5728) );
  NANDN U4303 ( .A(n2578), .B(n5730), .Z(n5729) );
  NANDN U4304 ( .A(n2580), .B(n2601), .Z(n5730) );
  NANDN U4305 ( .A(n2606), .B(n5731), .Z(n2601) );
  NAND U4306 ( .A(n5732), .B(n2607), .Z(n5731) );
  NANDN U4307 ( .A(n2609), .B(n5733), .Z(n5732) );
  NAND U4308 ( .A(n5734), .B(n2611), .Z(n5733) );
  NANDN U4309 ( .A(n2613), .B(n5735), .Z(n5734) );
  NAND U4310 ( .A(n2616), .B(n2618), .Z(n5735) );
  AND U4311 ( .A(A[560]), .B(B[560]), .Z(n2618) );
  AND U4312 ( .A(A[561]), .B(B[561]), .Z(n2613) );
  AND U4313 ( .A(A[562]), .B(B[562]), .Z(n2609) );
  AND U4314 ( .A(B[563]), .B(A[563]), .Z(n2606) );
  NANDN U4315 ( .A(n2584), .B(n5736), .Z(n2578) );
  NAND U4316 ( .A(n5737), .B(n2585), .Z(n5736) );
  NANDN U4317 ( .A(n2587), .B(n5738), .Z(n5737) );
  NAND U4318 ( .A(n5739), .B(n2589), .Z(n5738) );
  NANDN U4319 ( .A(n2591), .B(n5740), .Z(n5739) );
  NAND U4320 ( .A(n2594), .B(n2596), .Z(n5740) );
  AND U4321 ( .A(A[564]), .B(B[564]), .Z(n2596) );
  AND U4322 ( .A(A[565]), .B(B[565]), .Z(n2591) );
  AND U4323 ( .A(A[566]), .B(B[566]), .Z(n2587) );
  AND U4324 ( .A(B[567]), .B(A[567]), .Z(n2584) );
  NANDN U4325 ( .A(n2557), .B(n5741), .Z(n2551) );
  NAND U4326 ( .A(n5742), .B(n2558), .Z(n5741) );
  NANDN U4327 ( .A(n2560), .B(n5743), .Z(n5742) );
  NAND U4328 ( .A(n5744), .B(n2562), .Z(n5743) );
  NANDN U4329 ( .A(n2564), .B(n5745), .Z(n5744) );
  NAND U4330 ( .A(n2567), .B(n2574), .Z(n5745) );
  AND U4331 ( .A(A[568]), .B(B[568]), .Z(n2574) );
  AND U4332 ( .A(A[569]), .B(B[569]), .Z(n2564) );
  AND U4333 ( .A(A[570]), .B(B[570]), .Z(n2560) );
  AND U4334 ( .A(B[571]), .B(A[571]), .Z(n2557) );
  AND U4335 ( .A(A[572]), .B(B[572]), .Z(n2546) );
  AND U4336 ( .A(A[573]), .B(B[573]), .Z(n2541) );
  AND U4337 ( .A(A[574]), .B(B[574]), .Z(n2537) );
  ANDN U4338 ( .B(n5746), .A(n2534), .Z(n5719) );
  AND U4339 ( .A(B[575]), .B(A[575]), .Z(n2534) );
  NANDN U4340 ( .A(n5747), .B(n5748), .Z(n5746) );
  NANDN U4341 ( .A(n2622), .B(n5749), .Z(n5748) );
  NANDN U4342 ( .A(n2624), .B(n5750), .Z(n5749) );
  NANDN U4343 ( .A(n2723), .B(n5751), .Z(n5750) );
  NANDN U4344 ( .A(n2725), .B(n2819), .Z(n5751) );
  NANDN U4345 ( .A(n2824), .B(n5752), .Z(n2819) );
  NAND U4346 ( .A(n5753), .B(n2825), .Z(n5752) );
  NANDN U4347 ( .A(n2827), .B(n5754), .Z(n5753) );
  NAND U4348 ( .A(n5755), .B(n2829), .Z(n5754) );
  NANDN U4349 ( .A(n2831), .B(n5756), .Z(n5755) );
  NAND U4350 ( .A(n5757), .B(n2834), .Z(n5756) );
  NANDN U4351 ( .A(n2836), .B(n5758), .Z(n5757) );
  NAND U4352 ( .A(n5759), .B(n2839), .Z(n5758) );
  NANDN U4353 ( .A(n2841), .B(n5760), .Z(n5759) );
  NANDN U4354 ( .A(n2843), .B(n5761), .Z(n5760) );
  NANDN U4355 ( .A(n2863), .B(n5762), .Z(n5761) );
  NANDN U4356 ( .A(n2865), .B(n2894), .Z(n5762) );
  NANDN U4357 ( .A(n2898), .B(n5763), .Z(n2894) );
  NAND U4358 ( .A(n5764), .B(n2899), .Z(n5763) );
  NANDN U4359 ( .A(n2901), .B(n5765), .Z(n5764) );
  NAND U4360 ( .A(n5766), .B(n2903), .Z(n5765) );
  NANDN U4361 ( .A(n2905), .B(n5767), .Z(n5766) );
  NAND U4362 ( .A(n2908), .B(n2910), .Z(n5767) );
  AND U4363 ( .A(A[512]), .B(B[512]), .Z(n2910) );
  AND U4364 ( .A(A[513]), .B(B[513]), .Z(n2905) );
  AND U4365 ( .A(A[514]), .B(B[514]), .Z(n2901) );
  AND U4366 ( .A(B[515]), .B(A[515]), .Z(n2898) );
  NANDN U4367 ( .A(n2877), .B(n5768), .Z(n2863) );
  NAND U4368 ( .A(n5769), .B(n2878), .Z(n5768) );
  NANDN U4369 ( .A(n2880), .B(n5770), .Z(n5769) );
  NAND U4370 ( .A(n5771), .B(n2882), .Z(n5770) );
  NANDN U4371 ( .A(n2884), .B(n5772), .Z(n5771) );
  NAND U4372 ( .A(n2887), .B(n2889), .Z(n5772) );
  AND U4373 ( .A(A[516]), .B(B[516]), .Z(n2889) );
  AND U4374 ( .A(A[517]), .B(B[517]), .Z(n2884) );
  AND U4375 ( .A(A[518]), .B(B[518]), .Z(n2880) );
  AND U4376 ( .A(B[519]), .B(A[519]), .Z(n2877) );
  NANDN U4377 ( .A(n2847), .B(n5773), .Z(n2841) );
  NAND U4378 ( .A(n5774), .B(n2848), .Z(n5773) );
  NANDN U4379 ( .A(n2850), .B(n5775), .Z(n5774) );
  NAND U4380 ( .A(n5776), .B(n2852), .Z(n5775) );
  NANDN U4381 ( .A(n2854), .B(n5777), .Z(n5776) );
  NAND U4382 ( .A(n2857), .B(n2859), .Z(n5777) );
  AND U4383 ( .A(A[520]), .B(B[520]), .Z(n2859) );
  AND U4384 ( .A(A[521]), .B(B[521]), .Z(n2854) );
  AND U4385 ( .A(A[522]), .B(B[522]), .Z(n2850) );
  AND U4386 ( .A(B[523]), .B(A[523]), .Z(n2847) );
  AND U4387 ( .A(A[524]), .B(B[524]), .Z(n2836) );
  AND U4388 ( .A(A[525]), .B(B[525]), .Z(n2831) );
  AND U4389 ( .A(A[526]), .B(B[526]), .Z(n2827) );
  AND U4390 ( .A(B[527]), .B(A[527]), .Z(n2824) );
  NANDN U4391 ( .A(n2729), .B(n5778), .Z(n2723) );
  NAND U4392 ( .A(n5779), .B(n2730), .Z(n5778) );
  NANDN U4393 ( .A(n2732), .B(n5780), .Z(n5779) );
  NAND U4394 ( .A(n5781), .B(n2734), .Z(n5780) );
  NANDN U4395 ( .A(n2736), .B(n5782), .Z(n5781) );
  NAND U4396 ( .A(n5783), .B(n2739), .Z(n5782) );
  NANDN U4397 ( .A(n2741), .B(n5784), .Z(n5783) );
  NAND U4398 ( .A(n5785), .B(n2744), .Z(n5784) );
  NANDN U4399 ( .A(n2746), .B(n5786), .Z(n5785) );
  NANDN U4400 ( .A(n2748), .B(n5787), .Z(n5786) );
  NANDN U4401 ( .A(n2772), .B(n5788), .Z(n5787) );
  NANDN U4402 ( .A(n2774), .B(n2795), .Z(n5788) );
  NANDN U4403 ( .A(n2799), .B(n5789), .Z(n2795) );
  NAND U4404 ( .A(n5790), .B(n2800), .Z(n5789) );
  NANDN U4405 ( .A(n2802), .B(n5791), .Z(n5790) );
  NAND U4406 ( .A(n5792), .B(n2804), .Z(n5791) );
  NANDN U4407 ( .A(n2806), .B(n5793), .Z(n5792) );
  NAND U4408 ( .A(n2809), .B(n2814), .Z(n5793) );
  AND U4409 ( .A(A[528]), .B(B[528]), .Z(n2814) );
  AND U4410 ( .A(A[529]), .B(B[529]), .Z(n2806) );
  AND U4411 ( .A(A[530]), .B(B[530]), .Z(n2802) );
  AND U4412 ( .A(B[531]), .B(A[531]), .Z(n2799) );
  NANDN U4413 ( .A(n2778), .B(n5794), .Z(n2772) );
  NAND U4414 ( .A(n5795), .B(n2779), .Z(n5794) );
  NANDN U4415 ( .A(n2781), .B(n5796), .Z(n5795) );
  NAND U4416 ( .A(n5797), .B(n2783), .Z(n5796) );
  NANDN U4417 ( .A(n2785), .B(n5798), .Z(n5797) );
  NAND U4418 ( .A(n2788), .B(n2790), .Z(n5798) );
  AND U4419 ( .A(A[532]), .B(B[532]), .Z(n2790) );
  AND U4420 ( .A(A[533]), .B(B[533]), .Z(n2785) );
  AND U4421 ( .A(A[534]), .B(B[534]), .Z(n2781) );
  AND U4422 ( .A(B[535]), .B(A[535]), .Z(n2778) );
  NANDN U4423 ( .A(n2756), .B(n5799), .Z(n2746) );
  NAND U4424 ( .A(n5800), .B(n2757), .Z(n5799) );
  NANDN U4425 ( .A(n2759), .B(n5801), .Z(n5800) );
  NAND U4426 ( .A(n5802), .B(n2761), .Z(n5801) );
  NANDN U4427 ( .A(n2763), .B(n5803), .Z(n5802) );
  NAND U4428 ( .A(n2766), .B(n2768), .Z(n5803) );
  AND U4429 ( .A(A[536]), .B(B[536]), .Z(n2768) );
  AND U4430 ( .A(A[537]), .B(B[537]), .Z(n2763) );
  AND U4431 ( .A(A[538]), .B(B[538]), .Z(n2759) );
  AND U4432 ( .A(B[539]), .B(A[539]), .Z(n2756) );
  AND U4433 ( .A(A[540]), .B(B[540]), .Z(n2741) );
  AND U4434 ( .A(A[541]), .B(B[541]), .Z(n2736) );
  AND U4435 ( .A(A[542]), .B(B[542]), .Z(n2732) );
  AND U4436 ( .A(B[543]), .B(A[543]), .Z(n2729) );
  NANDN U4437 ( .A(n2636), .B(n5804), .Z(n2622) );
  NAND U4438 ( .A(n5805), .B(n2637), .Z(n5804) );
  NANDN U4439 ( .A(n2639), .B(n5806), .Z(n5805) );
  NAND U4440 ( .A(n5807), .B(n2641), .Z(n5806) );
  NANDN U4441 ( .A(n2643), .B(n5808), .Z(n5807) );
  NAND U4442 ( .A(n5809), .B(n2646), .Z(n5808) );
  NANDN U4443 ( .A(n2648), .B(n5810), .Z(n5809) );
  NAND U4444 ( .A(n5811), .B(n2651), .Z(n5810) );
  NANDN U4445 ( .A(n2653), .B(n5812), .Z(n5811) );
  NANDN U4446 ( .A(n2655), .B(n5813), .Z(n5812) );
  NANDN U4447 ( .A(n2675), .B(n5814), .Z(n5813) );
  NANDN U4448 ( .A(n2677), .B(n2703), .Z(n5814) );
  NANDN U4449 ( .A(n2707), .B(n5815), .Z(n2703) );
  NAND U4450 ( .A(n5816), .B(n2708), .Z(n5815) );
  NANDN U4451 ( .A(n2710), .B(n5817), .Z(n5816) );
  NAND U4452 ( .A(n5818), .B(n2712), .Z(n5817) );
  NANDN U4453 ( .A(n2714), .B(n5819), .Z(n5818) );
  NAND U4454 ( .A(n2717), .B(n2719), .Z(n5819) );
  AND U4455 ( .A(A[544]), .B(B[544]), .Z(n2719) );
  AND U4456 ( .A(A[545]), .B(B[545]), .Z(n2714) );
  AND U4457 ( .A(A[546]), .B(B[546]), .Z(n2710) );
  AND U4458 ( .A(B[547]), .B(A[547]), .Z(n2707) );
  NANDN U4459 ( .A(n2681), .B(n5820), .Z(n2675) );
  NAND U4460 ( .A(n5821), .B(n2682), .Z(n5820) );
  NANDN U4461 ( .A(n2684), .B(n5822), .Z(n5821) );
  NAND U4462 ( .A(n5823), .B(n2686), .Z(n5822) );
  NANDN U4463 ( .A(n2688), .B(n5824), .Z(n5823) );
  NAND U4464 ( .A(n2691), .B(n2698), .Z(n5824) );
  AND U4465 ( .A(A[548]), .B(B[548]), .Z(n2698) );
  AND U4466 ( .A(A[549]), .B(B[549]), .Z(n2688) );
  AND U4467 ( .A(A[550]), .B(B[550]), .Z(n2684) );
  AND U4468 ( .A(B[551]), .B(A[551]), .Z(n2681) );
  NANDN U4469 ( .A(n2659), .B(n5825), .Z(n2653) );
  NAND U4470 ( .A(n5826), .B(n2660), .Z(n5825) );
  NANDN U4471 ( .A(n2662), .B(n5827), .Z(n5826) );
  NAND U4472 ( .A(n5828), .B(n2664), .Z(n5827) );
  NANDN U4473 ( .A(n2666), .B(n5829), .Z(n5828) );
  NAND U4474 ( .A(n2669), .B(n2671), .Z(n5829) );
  AND U4475 ( .A(A[552]), .B(B[552]), .Z(n2671) );
  AND U4476 ( .A(A[553]), .B(B[553]), .Z(n2666) );
  AND U4477 ( .A(A[554]), .B(B[554]), .Z(n2662) );
  AND U4478 ( .A(B[555]), .B(A[555]), .Z(n2659) );
  AND U4479 ( .A(A[556]), .B(B[556]), .Z(n2648) );
  AND U4480 ( .A(A[557]), .B(B[557]), .Z(n2643) );
  AND U4481 ( .A(A[558]), .B(B[558]), .Z(n2639) );
  AND U4482 ( .A(B[559]), .B(A[559]), .Z(n2636) );
  NANDN U4483 ( .A(n2136), .B(n2531), .Z(n5717) );
  AND U4484 ( .A(n5830), .B(n5831), .Z(n2531) );
  ANDN U4485 ( .B(n5832), .A(n2624), .Z(n5831) );
  NAND U4486 ( .A(n5833), .B(n5834), .Z(n2624) );
  AND U4487 ( .A(n5835), .B(n5836), .Z(n5834) );
  AND U4488 ( .A(n2651), .B(n2646), .Z(n5836) );
  OR U4489 ( .A(A[557]), .B(B[557]), .Z(n2646) );
  OR U4490 ( .A(A[556]), .B(B[556]), .Z(n2651) );
  AND U4491 ( .A(n2641), .B(n2637), .Z(n5835) );
  OR U4492 ( .A(B[559]), .B(A[559]), .Z(n2637) );
  OR U4493 ( .A(A[558]), .B(B[558]), .Z(n2641) );
  ANDN U4494 ( .B(n5837), .A(n2704), .Z(n5833) );
  NAND U4495 ( .A(n5838), .B(n5839), .Z(n2704) );
  AND U4496 ( .A(n2721), .B(n2717), .Z(n5839) );
  OR U4497 ( .A(A[545]), .B(B[545]), .Z(n2717) );
  OR U4498 ( .A(A[544]), .B(B[544]), .Z(n2721) );
  AND U4499 ( .A(n2712), .B(n2708), .Z(n5838) );
  OR U4500 ( .A(B[547]), .B(A[547]), .Z(n2708) );
  OR U4501 ( .A(A[546]), .B(B[546]), .Z(n2712) );
  NOR U4502 ( .A(n2677), .B(n2655), .Z(n5837) );
  NAND U4503 ( .A(n5840), .B(n5841), .Z(n2655) );
  AND U4504 ( .A(n2673), .B(n2669), .Z(n5841) );
  OR U4505 ( .A(A[553]), .B(B[553]), .Z(n2669) );
  OR U4506 ( .A(A[552]), .B(B[552]), .Z(n2673) );
  AND U4507 ( .A(n2664), .B(n2660), .Z(n5840) );
  OR U4508 ( .A(B[555]), .B(A[555]), .Z(n2660) );
  OR U4509 ( .A(A[554]), .B(B[554]), .Z(n2664) );
  NAND U4510 ( .A(n5842), .B(n5843), .Z(n2677) );
  AND U4511 ( .A(n2700), .B(n2691), .Z(n5843) );
  OR U4512 ( .A(A[549]), .B(B[549]), .Z(n2691) );
  OR U4513 ( .A(A[548]), .B(B[548]), .Z(n2700) );
  AND U4514 ( .A(n2686), .B(n2682), .Z(n5842) );
  OR U4515 ( .A(B[551]), .B(A[551]), .Z(n2682) );
  OR U4516 ( .A(A[550]), .B(B[550]), .Z(n2686) );
  NOR U4517 ( .A(n2821), .B(n2725), .Z(n5832) );
  NAND U4518 ( .A(n5844), .B(n5845), .Z(n2725) );
  AND U4519 ( .A(n5846), .B(n5847), .Z(n5845) );
  AND U4520 ( .A(n2744), .B(n2739), .Z(n5847) );
  OR U4521 ( .A(A[541]), .B(B[541]), .Z(n2739) );
  OR U4522 ( .A(A[540]), .B(B[540]), .Z(n2744) );
  AND U4523 ( .A(n2734), .B(n2730), .Z(n5846) );
  OR U4524 ( .A(B[543]), .B(A[543]), .Z(n2730) );
  OR U4525 ( .A(A[542]), .B(B[542]), .Z(n2734) );
  ANDN U4526 ( .B(n5848), .A(n2796), .Z(n5844) );
  NAND U4527 ( .A(n5849), .B(n5850), .Z(n2796) );
  AND U4528 ( .A(n2816), .B(n2809), .Z(n5850) );
  OR U4529 ( .A(A[529]), .B(B[529]), .Z(n2809) );
  OR U4530 ( .A(A[528]), .B(B[528]), .Z(n2816) );
  AND U4531 ( .A(n2804), .B(n2800), .Z(n5849) );
  OR U4532 ( .A(B[531]), .B(A[531]), .Z(n2800) );
  OR U4533 ( .A(A[530]), .B(B[530]), .Z(n2804) );
  NOR U4534 ( .A(n2774), .B(n2748), .Z(n5848) );
  NAND U4535 ( .A(n5851), .B(n5852), .Z(n2748) );
  AND U4536 ( .A(n2770), .B(n2766), .Z(n5852) );
  OR U4537 ( .A(A[537]), .B(B[537]), .Z(n2766) );
  OR U4538 ( .A(A[536]), .B(B[536]), .Z(n2770) );
  AND U4539 ( .A(n2761), .B(n2757), .Z(n5851) );
  OR U4540 ( .A(B[539]), .B(A[539]), .Z(n2757) );
  OR U4541 ( .A(A[538]), .B(B[538]), .Z(n2761) );
  NAND U4542 ( .A(n5853), .B(n5854), .Z(n2774) );
  AND U4543 ( .A(n2792), .B(n2788), .Z(n5854) );
  OR U4544 ( .A(A[533]), .B(B[533]), .Z(n2788) );
  OR U4545 ( .A(A[532]), .B(B[532]), .Z(n2792) );
  AND U4546 ( .A(n2783), .B(n2779), .Z(n5853) );
  OR U4547 ( .A(B[535]), .B(A[535]), .Z(n2779) );
  OR U4548 ( .A(A[534]), .B(B[534]), .Z(n2783) );
  ANDN U4549 ( .B(n5855), .A(n2917), .Z(n2821) );
  AND U4550 ( .A(B[511]), .B(A[511]), .Z(n2917) );
  NANDN U4551 ( .A(n2916), .B(n5856), .Z(n5855) );
  NAND U4552 ( .A(n5857), .B(n5858), .Z(n5856) );
  NAND U4553 ( .A(n5859), .B(n5860), .Z(n5858) );
  AND U4554 ( .A(n5861), .B(n5862), .Z(n5860) );
  ANDN U4555 ( .B(n2926), .A(n2935), .Z(n5862) );
  AND U4556 ( .A(n2921), .B(n5863), .Z(n5861) );
  NANDN U4557 ( .A(n3013), .B(n5864), .Z(n5863) );
  NANDN U4558 ( .A(n3015), .B(n5865), .Z(n5864) );
  NANDN U4559 ( .A(n3102), .B(n5866), .Z(n5865) );
  NANDN U4560 ( .A(n3104), .B(n5867), .Z(n5866) );
  NANDN U4561 ( .A(n3203), .B(n5868), .Z(n5867) );
  NANDN U4562 ( .A(n3205), .B(n5869), .Z(n5868) );
  NANDN U4563 ( .A(n3301), .B(n5870), .Z(n5869) );
  NANDN U4564 ( .A(n3303), .B(n5871), .Z(n5870) );
  NANDN U4565 ( .A(n3690), .B(n5872), .Z(n5871) );
  AND U4566 ( .A(n5873), .B(n5874), .Z(n5872) );
  NANDN U4567 ( .A(n3692), .B(n4069), .Z(n5874) );
  NAND U4568 ( .A(n5875), .B(n5876), .Z(n4069) );
  NAND U4569 ( .A(n5877), .B(n4082), .Z(n5876) );
  NANDN U4570 ( .A(n4084), .B(n5878), .Z(n5877) );
  NAND U4571 ( .A(n5879), .B(n4086), .Z(n5878) );
  NANDN U4572 ( .A(n4088), .B(n5880), .Z(n5879) );
  NAND U4573 ( .A(n5881), .B(n4091), .Z(n5880) );
  NANDN U4574 ( .A(n4093), .B(n5882), .Z(n5881) );
  NAND U4575 ( .A(n5883), .B(n4096), .Z(n5882) );
  NANDN U4576 ( .A(n4098), .B(n5884), .Z(n5883) );
  NANDN U4577 ( .A(n4100), .B(n5885), .Z(n5884) );
  NANDN U4578 ( .A(n4120), .B(n5886), .Z(n5885) );
  NANDN U4579 ( .A(n4122), .B(n4148), .Z(n5886) );
  NANDN U4580 ( .A(n4153), .B(n5887), .Z(n4148) );
  NAND U4581 ( .A(n5888), .B(n4154), .Z(n5887) );
  NANDN U4582 ( .A(n4156), .B(n5889), .Z(n5888) );
  NAND U4583 ( .A(n5890), .B(n4158), .Z(n5889) );
  NANDN U4584 ( .A(n4160), .B(n5891), .Z(n5890) );
  NAND U4585 ( .A(n4163), .B(n4165), .Z(n5891) );
  AND U4586 ( .A(A[304]), .B(B[304]), .Z(n4165) );
  AND U4587 ( .A(A[305]), .B(B[305]), .Z(n4160) );
  AND U4588 ( .A(A[306]), .B(B[306]), .Z(n4156) );
  AND U4589 ( .A(B[307]), .B(A[307]), .Z(n4153) );
  NANDN U4590 ( .A(n4126), .B(n5892), .Z(n4120) );
  NAND U4591 ( .A(n5893), .B(n4127), .Z(n5892) );
  NANDN U4592 ( .A(n4129), .B(n5894), .Z(n5893) );
  NAND U4593 ( .A(n5895), .B(n4131), .Z(n5894) );
  NANDN U4594 ( .A(n4133), .B(n5896), .Z(n5895) );
  NAND U4595 ( .A(n4136), .B(n4143), .Z(n5896) );
  AND U4596 ( .A(A[308]), .B(B[308]), .Z(n4143) );
  AND U4597 ( .A(A[309]), .B(B[309]), .Z(n4133) );
  AND U4598 ( .A(A[310]), .B(B[310]), .Z(n4129) );
  AND U4599 ( .A(B[311]), .B(A[311]), .Z(n4126) );
  NANDN U4600 ( .A(n4104), .B(n5897), .Z(n4098) );
  NAND U4601 ( .A(n5898), .B(n4105), .Z(n5897) );
  NANDN U4602 ( .A(n4107), .B(n5899), .Z(n5898) );
  NAND U4603 ( .A(n5900), .B(n4109), .Z(n5899) );
  NANDN U4604 ( .A(n4111), .B(n5901), .Z(n5900) );
  NAND U4605 ( .A(n4114), .B(n4116), .Z(n5901) );
  AND U4606 ( .A(A[312]), .B(B[312]), .Z(n4116) );
  AND U4607 ( .A(A[313]), .B(B[313]), .Z(n4111) );
  AND U4608 ( .A(A[314]), .B(B[314]), .Z(n4107) );
  AND U4609 ( .A(B[315]), .B(A[315]), .Z(n4104) );
  AND U4610 ( .A(A[316]), .B(B[316]), .Z(n4093) );
  AND U4611 ( .A(A[317]), .B(B[317]), .Z(n4088) );
  AND U4612 ( .A(A[318]), .B(B[318]), .Z(n4084) );
  ANDN U4613 ( .B(n5902), .A(n4081), .Z(n5875) );
  AND U4614 ( .A(B[319]), .B(A[319]), .Z(n4081) );
  NANDN U4615 ( .A(n5903), .B(n5904), .Z(n5902) );
  NANDN U4616 ( .A(n4169), .B(n5905), .Z(n5904) );
  NANDN U4617 ( .A(n4171), .B(n5906), .Z(n5905) );
  NANDN U4618 ( .A(n4271), .B(n5907), .Z(n5906) );
  NANDN U4619 ( .A(n4273), .B(n4368), .Z(n5907) );
  NANDN U4620 ( .A(n4373), .B(n5908), .Z(n4368) );
  NAND U4621 ( .A(n5909), .B(n4374), .Z(n5908) );
  NANDN U4622 ( .A(n4376), .B(n5910), .Z(n5909) );
  NAND U4623 ( .A(n5911), .B(n4378), .Z(n5910) );
  NANDN U4624 ( .A(n4380), .B(n5912), .Z(n5911) );
  NAND U4625 ( .A(n5913), .B(n4383), .Z(n5912) );
  NANDN U4626 ( .A(n4390), .B(n5914), .Z(n5913) );
  NAND U4627 ( .A(n5915), .B(n4393), .Z(n5914) );
  NANDN U4628 ( .A(n4395), .B(n5916), .Z(n5915) );
  NANDN U4629 ( .A(n4397), .B(n5917), .Z(n5916) );
  NANDN U4630 ( .A(n4417), .B(n5918), .Z(n5917) );
  NANDN U4631 ( .A(n4419), .B(n4440), .Z(n5918) );
  NANDN U4632 ( .A(n4448), .B(n5919), .Z(n4440) );
  NAND U4633 ( .A(n5920), .B(n4449), .Z(n5919) );
  NANDN U4634 ( .A(n4451), .B(n5921), .Z(n5920) );
  NAND U4635 ( .A(n5922), .B(n4453), .Z(n5921) );
  NANDN U4636 ( .A(n4455), .B(n5923), .Z(n5922) );
  NAND U4637 ( .A(n4458), .B(n4460), .Z(n5923) );
  AND U4638 ( .A(A[256]), .B(B[256]), .Z(n4460) );
  AND U4639 ( .A(A[257]), .B(B[257]), .Z(n4455) );
  AND U4640 ( .A(A[258]), .B(B[258]), .Z(n4451) );
  AND U4641 ( .A(B[259]), .B(A[259]), .Z(n4448) );
  NANDN U4642 ( .A(n4423), .B(n5924), .Z(n4417) );
  NAND U4643 ( .A(n5925), .B(n4424), .Z(n5924) );
  NANDN U4644 ( .A(n4426), .B(n5926), .Z(n5925) );
  NAND U4645 ( .A(n5927), .B(n4428), .Z(n5926) );
  NANDN U4646 ( .A(n4430), .B(n5928), .Z(n5927) );
  NAND U4647 ( .A(n4433), .B(n4435), .Z(n5928) );
  AND U4648 ( .A(A[260]), .B(B[260]), .Z(n4435) );
  AND U4649 ( .A(A[261]), .B(B[261]), .Z(n4430) );
  AND U4650 ( .A(A[262]), .B(B[262]), .Z(n4426) );
  AND U4651 ( .A(B[263]), .B(A[263]), .Z(n4423) );
  NANDN U4652 ( .A(n4401), .B(n5929), .Z(n4395) );
  NAND U4653 ( .A(n5930), .B(n4402), .Z(n5929) );
  NANDN U4654 ( .A(n4404), .B(n5931), .Z(n5930) );
  NAND U4655 ( .A(n5932), .B(n4406), .Z(n5931) );
  NANDN U4656 ( .A(n4408), .B(n5933), .Z(n5932) );
  NAND U4657 ( .A(n4411), .B(n4413), .Z(n5933) );
  AND U4658 ( .A(A[264]), .B(B[264]), .Z(n4413) );
  AND U4659 ( .A(A[265]), .B(B[265]), .Z(n4408) );
  AND U4660 ( .A(A[266]), .B(B[266]), .Z(n4404) );
  AND U4661 ( .A(B[267]), .B(A[267]), .Z(n4401) );
  AND U4662 ( .A(A[268]), .B(B[268]), .Z(n4390) );
  AND U4663 ( .A(A[269]), .B(B[269]), .Z(n4380) );
  AND U4664 ( .A(A[270]), .B(B[270]), .Z(n4376) );
  AND U4665 ( .A(B[271]), .B(A[271]), .Z(n4373) );
  NANDN U4666 ( .A(n4277), .B(n5934), .Z(n4271) );
  NAND U4667 ( .A(n5935), .B(n4278), .Z(n5934) );
  NANDN U4668 ( .A(n4280), .B(n5936), .Z(n5935) );
  NAND U4669 ( .A(n5937), .B(n4282), .Z(n5936) );
  NANDN U4670 ( .A(n4284), .B(n5938), .Z(n5937) );
  NAND U4671 ( .A(n5939), .B(n4287), .Z(n5938) );
  NANDN U4672 ( .A(n4289), .B(n5940), .Z(n5939) );
  NAND U4673 ( .A(n5941), .B(n4292), .Z(n5940) );
  NANDN U4674 ( .A(n4294), .B(n5942), .Z(n5941) );
  NANDN U4675 ( .A(n4296), .B(n5943), .Z(n5942) );
  NANDN U4676 ( .A(n4316), .B(n5944), .Z(n5943) );
  NANDN U4677 ( .A(n4318), .B(n4347), .Z(n5944) );
  NANDN U4678 ( .A(n4351), .B(n5945), .Z(n4347) );
  NAND U4679 ( .A(n5946), .B(n4352), .Z(n5945) );
  NANDN U4680 ( .A(n4354), .B(n5947), .Z(n5946) );
  NAND U4681 ( .A(n5948), .B(n4356), .Z(n5947) );
  NANDN U4682 ( .A(n4358), .B(n5949), .Z(n5948) );
  NAND U4683 ( .A(n4361), .B(n4363), .Z(n5949) );
  AND U4684 ( .A(A[272]), .B(B[272]), .Z(n4363) );
  AND U4685 ( .A(A[273]), .B(B[273]), .Z(n4358) );
  AND U4686 ( .A(A[274]), .B(B[274]), .Z(n4354) );
  AND U4687 ( .A(B[275]), .B(A[275]), .Z(n4351) );
  NANDN U4688 ( .A(n4330), .B(n5950), .Z(n4316) );
  NAND U4689 ( .A(n5951), .B(n4331), .Z(n5950) );
  NANDN U4690 ( .A(n4333), .B(n5952), .Z(n5951) );
  NAND U4691 ( .A(n5953), .B(n4335), .Z(n5952) );
  NANDN U4692 ( .A(n4337), .B(n5954), .Z(n5953) );
  NAND U4693 ( .A(n4340), .B(n4342), .Z(n5954) );
  AND U4694 ( .A(A[276]), .B(B[276]), .Z(n4342) );
  AND U4695 ( .A(A[277]), .B(B[277]), .Z(n4337) );
  AND U4696 ( .A(A[278]), .B(B[278]), .Z(n4333) );
  AND U4697 ( .A(B[279]), .B(A[279]), .Z(n4330) );
  NANDN U4698 ( .A(n4300), .B(n5955), .Z(n4294) );
  NAND U4699 ( .A(n5956), .B(n4301), .Z(n5955) );
  NANDN U4700 ( .A(n4303), .B(n5957), .Z(n5956) );
  NAND U4701 ( .A(n5958), .B(n4305), .Z(n5957) );
  NANDN U4702 ( .A(n4307), .B(n5959), .Z(n5958) );
  NAND U4703 ( .A(n4310), .B(n4312), .Z(n5959) );
  AND U4704 ( .A(A[280]), .B(B[280]), .Z(n4312) );
  AND U4705 ( .A(A[281]), .B(B[281]), .Z(n4307) );
  AND U4706 ( .A(A[282]), .B(B[282]), .Z(n4303) );
  AND U4707 ( .A(B[283]), .B(A[283]), .Z(n4300) );
  AND U4708 ( .A(A[284]), .B(B[284]), .Z(n4289) );
  AND U4709 ( .A(A[285]), .B(B[285]), .Z(n4284) );
  AND U4710 ( .A(A[286]), .B(B[286]), .Z(n4280) );
  AND U4711 ( .A(B[287]), .B(A[287]), .Z(n4277) );
  NANDN U4712 ( .A(n4175), .B(n5960), .Z(n4169) );
  NAND U4713 ( .A(n5961), .B(n4176), .Z(n5960) );
  NANDN U4714 ( .A(n4178), .B(n5962), .Z(n5961) );
  NAND U4715 ( .A(n5963), .B(n4180), .Z(n5962) );
  NANDN U4716 ( .A(n4182), .B(n5964), .Z(n5963) );
  NAND U4717 ( .A(n5965), .B(n4185), .Z(n5964) );
  NANDN U4718 ( .A(n4187), .B(n5966), .Z(n5965) );
  NAND U4719 ( .A(n5967), .B(n4190), .Z(n5966) );
  NANDN U4720 ( .A(n4192), .B(n5968), .Z(n5967) );
  NANDN U4721 ( .A(n4194), .B(n5969), .Z(n5968) );
  NANDN U4722 ( .A(n4223), .B(n5970), .Z(n5969) );
  NANDN U4723 ( .A(n4225), .B(n4246), .Z(n5970) );
  NANDN U4724 ( .A(n4250), .B(n5971), .Z(n4246) );
  NAND U4725 ( .A(n5972), .B(n4251), .Z(n5971) );
  NANDN U4726 ( .A(n4253), .B(n5973), .Z(n5972) );
  NAND U4727 ( .A(n5974), .B(n4255), .Z(n5973) );
  NANDN U4728 ( .A(n4257), .B(n5975), .Z(n5974) );
  NAND U4729 ( .A(n4260), .B(n4267), .Z(n5975) );
  AND U4730 ( .A(A[288]), .B(B[288]), .Z(n4267) );
  AND U4731 ( .A(A[289]), .B(B[289]), .Z(n4257) );
  AND U4732 ( .A(A[290]), .B(B[290]), .Z(n4253) );
  AND U4733 ( .A(B[291]), .B(A[291]), .Z(n4250) );
  NANDN U4734 ( .A(n4229), .B(n5976), .Z(n4223) );
  NAND U4735 ( .A(n5977), .B(n4230), .Z(n5976) );
  NANDN U4736 ( .A(n4232), .B(n5978), .Z(n5977) );
  NAND U4737 ( .A(n5979), .B(n4234), .Z(n5978) );
  NANDN U4738 ( .A(n4236), .B(n5980), .Z(n5979) );
  NAND U4739 ( .A(n4239), .B(n4241), .Z(n5980) );
  AND U4740 ( .A(A[292]), .B(B[292]), .Z(n4241) );
  AND U4741 ( .A(A[293]), .B(B[293]), .Z(n4236) );
  AND U4742 ( .A(A[294]), .B(B[294]), .Z(n4232) );
  AND U4743 ( .A(B[295]), .B(A[295]), .Z(n4229) );
  NANDN U4744 ( .A(n4207), .B(n5981), .Z(n4192) );
  NAND U4745 ( .A(n5982), .B(n4208), .Z(n5981) );
  NANDN U4746 ( .A(n4210), .B(n5983), .Z(n5982) );
  NAND U4747 ( .A(n5984), .B(n4212), .Z(n5983) );
  NANDN U4748 ( .A(n4214), .B(n5985), .Z(n5984) );
  NAND U4749 ( .A(n4217), .B(n4219), .Z(n5985) );
  AND U4750 ( .A(A[296]), .B(B[296]), .Z(n4219) );
  AND U4751 ( .A(A[297]), .B(B[297]), .Z(n4214) );
  AND U4752 ( .A(A[298]), .B(B[298]), .Z(n4210) );
  AND U4753 ( .A(B[299]), .B(A[299]), .Z(n4207) );
  AND U4754 ( .A(A[300]), .B(B[300]), .Z(n4187) );
  AND U4755 ( .A(A[301]), .B(B[301]), .Z(n4182) );
  AND U4756 ( .A(A[302]), .B(B[302]), .Z(n4178) );
  AND U4757 ( .A(B[303]), .B(A[303]), .Z(n4175) );
  NANDN U4758 ( .A(n3692), .B(n4070), .Z(n5873) );
  AND U4759 ( .A(n5986), .B(n5987), .Z(n4070) );
  ANDN U4760 ( .B(n5988), .A(n4171), .Z(n5987) );
  NAND U4761 ( .A(n5989), .B(n5990), .Z(n4171) );
  AND U4762 ( .A(n5991), .B(n5992), .Z(n5990) );
  AND U4763 ( .A(n4190), .B(n4185), .Z(n5992) );
  OR U4764 ( .A(A[301]), .B(B[301]), .Z(n4185) );
  OR U4765 ( .A(A[300]), .B(B[300]), .Z(n4190) );
  AND U4766 ( .A(n4180), .B(n4176), .Z(n5991) );
  OR U4767 ( .A(B[303]), .B(A[303]), .Z(n4176) );
  OR U4768 ( .A(A[302]), .B(B[302]), .Z(n4180) );
  ANDN U4769 ( .B(n5993), .A(n4247), .Z(n5989) );
  NAND U4770 ( .A(n5994), .B(n5995), .Z(n4247) );
  AND U4771 ( .A(n4269), .B(n4260), .Z(n5995) );
  OR U4772 ( .A(A[289]), .B(B[289]), .Z(n4260) );
  OR U4773 ( .A(A[288]), .B(B[288]), .Z(n4269) );
  AND U4774 ( .A(n4255), .B(n4251), .Z(n5994) );
  OR U4775 ( .A(B[291]), .B(A[291]), .Z(n4251) );
  OR U4776 ( .A(A[290]), .B(B[290]), .Z(n4255) );
  NOR U4777 ( .A(n4225), .B(n4194), .Z(n5993) );
  NAND U4778 ( .A(n5996), .B(n5997), .Z(n4194) );
  AND U4779 ( .A(n4221), .B(n4217), .Z(n5997) );
  OR U4780 ( .A(A[297]), .B(B[297]), .Z(n4217) );
  OR U4781 ( .A(A[296]), .B(B[296]), .Z(n4221) );
  AND U4782 ( .A(n4212), .B(n4208), .Z(n5996) );
  OR U4783 ( .A(B[299]), .B(A[299]), .Z(n4208) );
  OR U4784 ( .A(A[298]), .B(B[298]), .Z(n4212) );
  NAND U4785 ( .A(n5998), .B(n5999), .Z(n4225) );
  AND U4786 ( .A(n4243), .B(n4239), .Z(n5999) );
  OR U4787 ( .A(A[293]), .B(B[293]), .Z(n4239) );
  OR U4788 ( .A(A[292]), .B(B[292]), .Z(n4243) );
  AND U4789 ( .A(n4234), .B(n4230), .Z(n5998) );
  OR U4790 ( .A(B[295]), .B(A[295]), .Z(n4230) );
  OR U4791 ( .A(A[294]), .B(B[294]), .Z(n4234) );
  NOR U4792 ( .A(n4370), .B(n4273), .Z(n5988) );
  NAND U4793 ( .A(n6000), .B(n6001), .Z(n4273) );
  AND U4794 ( .A(n6002), .B(n6003), .Z(n6001) );
  AND U4795 ( .A(n4292), .B(n4287), .Z(n6003) );
  OR U4796 ( .A(A[285]), .B(B[285]), .Z(n4287) );
  OR U4797 ( .A(A[284]), .B(B[284]), .Z(n4292) );
  AND U4798 ( .A(n4282), .B(n4278), .Z(n6002) );
  OR U4799 ( .A(B[287]), .B(A[287]), .Z(n4278) );
  OR U4800 ( .A(A[286]), .B(B[286]), .Z(n4282) );
  ANDN U4801 ( .B(n6004), .A(n4348), .Z(n6000) );
  NAND U4802 ( .A(n6005), .B(n6006), .Z(n4348) );
  AND U4803 ( .A(n4365), .B(n4361), .Z(n6006) );
  OR U4804 ( .A(A[273]), .B(B[273]), .Z(n4361) );
  OR U4805 ( .A(A[272]), .B(B[272]), .Z(n4365) );
  AND U4806 ( .A(n4356), .B(n4352), .Z(n6005) );
  OR U4807 ( .A(B[275]), .B(A[275]), .Z(n4352) );
  OR U4808 ( .A(A[274]), .B(B[274]), .Z(n4356) );
  NOR U4809 ( .A(n4318), .B(n4296), .Z(n6004) );
  NAND U4810 ( .A(n6007), .B(n6008), .Z(n4296) );
  AND U4811 ( .A(n4314), .B(n4310), .Z(n6008) );
  OR U4812 ( .A(A[281]), .B(B[281]), .Z(n4310) );
  OR U4813 ( .A(A[280]), .B(B[280]), .Z(n4314) );
  AND U4814 ( .A(n4305), .B(n4301), .Z(n6007) );
  OR U4815 ( .A(B[283]), .B(A[283]), .Z(n4301) );
  OR U4816 ( .A(A[282]), .B(B[282]), .Z(n4305) );
  NAND U4817 ( .A(n6009), .B(n6010), .Z(n4318) );
  AND U4818 ( .A(n4344), .B(n4340), .Z(n6010) );
  OR U4819 ( .A(A[277]), .B(B[277]), .Z(n4340) );
  OR U4820 ( .A(A[276]), .B(B[276]), .Z(n4344) );
  AND U4821 ( .A(n4335), .B(n4331), .Z(n6009) );
  OR U4822 ( .A(B[279]), .B(A[279]), .Z(n4331) );
  OR U4823 ( .A(A[278]), .B(B[278]), .Z(n4335) );
  ANDN U4824 ( .B(n6011), .A(n4467), .Z(n4370) );
  AND U4825 ( .A(B[255]), .B(A[255]), .Z(n4467) );
  NANDN U4826 ( .A(n4466), .B(n6012), .Z(n6011) );
  NANDN U4827 ( .A(n4469), .B(n6013), .Z(n6012) );
  NANDN U4828 ( .A(n4470), .B(n6014), .Z(n6013) );
  NANDN U4829 ( .A(n4473), .B(n6015), .Z(n6014) );
  NANDN U4830 ( .A(n4475), .B(n6016), .Z(n6015) );
  NAND U4831 ( .A(n6017), .B(n6018), .Z(n6016) );
  NAND U4832 ( .A(n6019), .B(n6020), .Z(n6018) );
  AND U4833 ( .A(n4513), .B(n6021), .Z(n6020) );
  ANDN U4834 ( .B(n4481), .A(n4535), .Z(n6021) );
  ANDN U4835 ( .B(n6022), .A(n4565), .Z(n4535) );
  AND U4836 ( .A(B[239]), .B(A[239]), .Z(n4565) );
  NANDN U4837 ( .A(n4564), .B(n6023), .Z(n6022) );
  NANDN U4838 ( .A(n4567), .B(n6024), .Z(n6023) );
  NANDN U4839 ( .A(n4568), .B(n6025), .Z(n6024) );
  NANDN U4840 ( .A(n4571), .B(n6026), .Z(n6025) );
  NANDN U4841 ( .A(n4573), .B(n6027), .Z(n6026) );
  NAND U4842 ( .A(n6028), .B(n6029), .Z(n6027) );
  NAND U4843 ( .A(n6030), .B(n6031), .Z(n6029) );
  AND U4844 ( .A(n4606), .B(n6032), .Z(n6031) );
  ANDN U4845 ( .B(n4579), .A(n4633), .Z(n6032) );
  ANDN U4846 ( .B(n6033), .A(n4655), .Z(n4633) );
  AND U4847 ( .A(B[223]), .B(A[223]), .Z(n4655) );
  NANDN U4848 ( .A(n4654), .B(n6034), .Z(n6033) );
  NANDN U4849 ( .A(n4657), .B(n6035), .Z(n6034) );
  NANDN U4850 ( .A(n4658), .B(n6036), .Z(n6035) );
  NANDN U4851 ( .A(n4661), .B(n6037), .Z(n6036) );
  NANDN U4852 ( .A(n4663), .B(n6038), .Z(n6037) );
  NAND U4853 ( .A(n6039), .B(n6040), .Z(n6038) );
  NAND U4854 ( .A(n6041), .B(n6042), .Z(n6040) );
  AND U4855 ( .A(n4700), .B(n6043), .Z(n6042) );
  ANDN U4856 ( .B(n4669), .A(n4722), .Z(n6043) );
  ANDN U4857 ( .B(n6044), .A(n4749), .Z(n4722) );
  AND U4858 ( .A(B[207]), .B(A[207]), .Z(n4749) );
  NANDN U4859 ( .A(n4748), .B(n6045), .Z(n6044) );
  NANDN U4860 ( .A(n4751), .B(n6046), .Z(n6045) );
  NANDN U4861 ( .A(n4752), .B(n6047), .Z(n6046) );
  NANDN U4862 ( .A(n4755), .B(n6048), .Z(n6047) );
  NANDN U4863 ( .A(n4757), .B(n6049), .Z(n6048) );
  NAND U4864 ( .A(n6050), .B(n6051), .Z(n6049) );
  NAND U4865 ( .A(n6052), .B(n6053), .Z(n6051) );
  AND U4866 ( .A(n4790), .B(n6054), .Z(n6053) );
  ANDN U4867 ( .B(n4763), .A(n4824), .Z(n6054) );
  ANDN U4868 ( .B(n6055), .A(n4846), .Z(n4824) );
  AND U4869 ( .A(B[191]), .B(A[191]), .Z(n4846) );
  NANDN U4870 ( .A(n4845), .B(n6056), .Z(n6055) );
  NAND U4871 ( .A(n6057), .B(n6058), .Z(n6056) );
  NAND U4872 ( .A(n6059), .B(n6060), .Z(n6058) );
  AND U4873 ( .A(n6061), .B(n6062), .Z(n6060) );
  ANDN U4874 ( .B(n4855), .A(n4864), .Z(n6062) );
  AND U4875 ( .A(n4850), .B(n4914), .Z(n6061) );
  NANDN U4876 ( .A(n6063), .B(n6064), .Z(n4914) );
  NANDN U4877 ( .A(n6065), .B(n5004), .Z(n6064) );
  NANDN U4878 ( .A(n6066), .B(n6067), .Z(n5004) );
  NANDN U4879 ( .A(n6068), .B(n5097), .Z(n6067) );
  NANDN U4880 ( .A(n6069), .B(n6070), .Z(n5097) );
  OR U4881 ( .A(n6071), .B(n5186), .Z(n6070) );
  ANDN U4882 ( .B(n6072), .A(n5212), .Z(n5186) );
  AND U4883 ( .A(B[127]), .B(A[127]), .Z(n5212) );
  NANDN U4884 ( .A(n5211), .B(n6073), .Z(n6072) );
  NAND U4885 ( .A(n6074), .B(n6075), .Z(n6073) );
  NAND U4886 ( .A(n6076), .B(n6077), .Z(n6075) );
  AND U4887 ( .A(n6078), .B(n6079), .Z(n6077) );
  ANDN U4888 ( .B(n5221), .A(n5225), .Z(n6079) );
  AND U4889 ( .A(n5216), .B(n6080), .Z(n6078) );
  NANDN U4890 ( .A(n5302), .B(n6081), .Z(n6080) );
  NANDN U4891 ( .A(n5304), .B(n6082), .Z(n6081) );
  NANDN U4892 ( .A(n5441), .B(n6083), .Z(n6082) );
  NANDN U4893 ( .A(n5442), .B(n6084), .Z(n6083) );
  NANDN U4894 ( .A(n5444), .B(n5443), .Z(n6084) );
  OR U4895 ( .A(n6085), .B(n1847), .Z(n5443) );
  ANDN U4896 ( .B(n6086), .A(n2141), .Z(n1847) );
  AND U4897 ( .A(B[63]), .B(A[63]), .Z(n2141) );
  NANDN U4898 ( .A(n2140), .B(n6087), .Z(n6086) );
  NANDN U4899 ( .A(n2143), .B(n6088), .Z(n6087) );
  NANDN U4900 ( .A(n2144), .B(n6089), .Z(n6088) );
  NANDN U4901 ( .A(n2205), .B(n6090), .Z(n6089) );
  NANDN U4902 ( .A(n2207), .B(n6091), .Z(n6090) );
  NANDN U4903 ( .A(n2264), .B(n6092), .Z(n6091) );
  NANDN U4904 ( .A(n2266), .B(n6093), .Z(n6092) );
  NANDN U4905 ( .A(n2325), .B(n6094), .Z(n6093) );
  NANDN U4906 ( .A(n2327), .B(n6095), .Z(n6094) );
  NANDN U4907 ( .A(n2569), .B(n6096), .Z(n6095) );
  AND U4908 ( .A(n6097), .B(n6098), .Z(n6096) );
  NANDN U4909 ( .A(n2571), .B(n2811), .Z(n6098) );
  NANDN U4910 ( .A(n2869), .B(n6099), .Z(n2811) );
  NAND U4911 ( .A(n6100), .B(n2870), .Z(n6099) );
  NANDN U4912 ( .A(n2872), .B(n6101), .Z(n6100) );
  NAND U4913 ( .A(n6102), .B(n2874), .Z(n6101) );
  NANDN U4914 ( .A(n2928), .B(n6103), .Z(n6102) );
  NAND U4915 ( .A(n2931), .B(n2991), .Z(n6103) );
  AND U4916 ( .A(A[48]), .B(B[48]), .Z(n2991) );
  AND U4917 ( .A(A[49]), .B(B[49]), .Z(n2928) );
  AND U4918 ( .A(A[50]), .B(B[50]), .Z(n2872) );
  AND U4919 ( .A(B[51]), .B(A[51]), .Z(n2869) );
  NANDN U4920 ( .A(n2571), .B(n2812), .Z(n6097) );
  AND U4921 ( .A(n6104), .B(n6105), .Z(n2812) );
  AND U4922 ( .A(n2874), .B(n6106), .Z(n6105) );
  AND U4923 ( .A(n2994), .B(n2931), .Z(n6106) );
  OR U4924 ( .A(A[49]), .B(B[49]), .Z(n2931) );
  OR U4925 ( .A(A[48]), .B(B[48]), .Z(n2994) );
  OR U4926 ( .A(A[50]), .B(B[50]), .Z(n2874) );
  ANDN U4927 ( .B(n2870), .A(n2993), .Z(n6104) );
  ANDN U4928 ( .B(n6107), .A(n3109), .Z(n2993) );
  AND U4929 ( .A(B[47]), .B(A[47]), .Z(n3109) );
  NANDN U4930 ( .A(n3108), .B(n6108), .Z(n6107) );
  NANDN U4931 ( .A(n3111), .B(n6109), .Z(n6108) );
  NANDN U4932 ( .A(n3112), .B(n6110), .Z(n6109) );
  NANDN U4933 ( .A(n3173), .B(n6111), .Z(n6110) );
  NANDN U4934 ( .A(n3175), .B(n6112), .Z(n6111) );
  NAND U4935 ( .A(n6113), .B(n6114), .Z(n6112) );
  NAND U4936 ( .A(n6115), .B(n6116), .Z(n6114) );
  AND U4937 ( .A(n3539), .B(n6117), .Z(n6116) );
  ANDN U4938 ( .B(n3234), .A(n3782), .Z(n6117) );
  ANDN U4939 ( .B(n6118), .A(n4074), .Z(n3782) );
  AND U4940 ( .A(B[31]), .B(A[31]), .Z(n4074) );
  NANDN U4941 ( .A(n4073), .B(n6119), .Z(n6118) );
  NANDN U4942 ( .A(n4076), .B(n6120), .Z(n6119) );
  NANDN U4943 ( .A(n4077), .B(n6121), .Z(n6120) );
  NANDN U4944 ( .A(n4138), .B(n6122), .Z(n6121) );
  NANDN U4945 ( .A(n4140), .B(n6123), .Z(n6122) );
  NAND U4946 ( .A(n6124), .B(n6125), .Z(n6123) );
  NAND U4947 ( .A(n6126), .B(n6127), .Z(n6125) );
  AND U4948 ( .A(n4504), .B(n6128), .Z(n6127) );
  ANDN U4949 ( .B(n4204), .A(n4740), .Z(n6128) );
  ANDN U4950 ( .B(n6129), .A(n5025), .Z(n4740) );
  AND U4951 ( .A(B[15]), .B(A[15]), .Z(n5025) );
  NAND U4952 ( .A(n5023), .B(n5026), .Z(n6129) );
  OR U4953 ( .A(B[15]), .B(A[15]), .Z(n5026) );
  NANDN U4954 ( .A(n5087), .B(n6130), .Z(n5023) );
  NAND U4955 ( .A(n5085), .B(n5088), .Z(n6130) );
  OR U4956 ( .A(B[14]), .B(A[14]), .Z(n5088) );
  NANDN U4957 ( .A(n5141), .B(n6131), .Z(n5085) );
  NAND U4958 ( .A(n5139), .B(n5142), .Z(n6131) );
  OR U4959 ( .A(B[13]), .B(A[13]), .Z(n5142) );
  NANDN U4960 ( .A(n5202), .B(n6132), .Z(n5139) );
  NAND U4961 ( .A(n5200), .B(n5203), .Z(n6132) );
  OR U4962 ( .A(B[12]), .B(A[12]), .Z(n5203) );
  NANDN U4963 ( .A(n5257), .B(n6133), .Z(n5200) );
  NANDN U4964 ( .A(n5256), .B(n6134), .Z(n6133) );
  NANDN U4965 ( .A(n5259), .B(n6135), .Z(n6134) );
  NANDN U4966 ( .A(n5260), .B(n6136), .Z(n6135) );
  NANDN U4967 ( .A(n3), .B(n6137), .Z(n6136) );
  NAND U4968 ( .A(n6138), .B(n4), .Z(n6137) );
  OR U4969 ( .A(A[9]), .B(B[9]), .Z(n4) );
  NANDN U4970 ( .A(n591), .B(n5320), .Z(n6138) );
  OR U4971 ( .A(n588), .B(n590), .Z(n5320) );
  NOR U4972 ( .A(B[8]), .B(A[8]), .Z(n590) );
  ANDN U4973 ( .B(n6139), .A(n1172), .Z(n588) );
  AND U4974 ( .A(B[7]), .B(A[7]), .Z(n1172) );
  NANDN U4975 ( .A(n1171), .B(n6140), .Z(n6139) );
  NANDN U4976 ( .A(n1174), .B(n1173), .Z(n6140) );
  NANDN U4977 ( .A(n1781), .B(n1779), .Z(n1173) );
  NANDN U4978 ( .A(n2386), .B(n6141), .Z(n1779) );
  NANDN U4979 ( .A(n2385), .B(n2383), .Z(n6141) );
  NANDN U4980 ( .A(n2989), .B(n6142), .Z(n2383) );
  OR U4981 ( .A(n2986), .B(n2988), .Z(n6142) );
  NOR U4982 ( .A(B[4]), .B(A[4]), .Z(n2988) );
  AND U4983 ( .A(n6143), .B(n6144), .Z(n2986) );
  NAND U4984 ( .A(n6145), .B(B[3]), .Z(n6144) );
  NANDN U4985 ( .A(A[3]), .B(n3591), .Z(n6145) );
  NANDN U4986 ( .A(n3591), .B(A[3]), .Z(n6143) );
  ANDN U4987 ( .B(n6146), .A(n4198), .Z(n3591) );
  AND U4988 ( .A(B[2]), .B(A[2]), .Z(n4198) );
  NAND U4989 ( .A(n4196), .B(n4199), .Z(n6146) );
  OR U4990 ( .A(B[2]), .B(A[2]), .Z(n4199) );
  NANDN U4991 ( .A(n4794), .B(n6147), .Z(n4196) );
  NANDN U4992 ( .A(n4793), .B(n4791), .Z(n6147) );
  NOR U4993 ( .A(B[1]), .B(A[1]), .Z(n4793) );
  AND U4994 ( .A(B[1]), .B(A[1]), .Z(n4794) );
  AND U4995 ( .A(B[4]), .B(A[4]), .Z(n2989) );
  NOR U4996 ( .A(B[5]), .B(A[5]), .Z(n2385) );
  AND U4997 ( .A(B[5]), .B(A[5]), .Z(n2386) );
  NOR U4998 ( .A(B[6]), .B(A[6]), .Z(n1781) );
  AND U4999 ( .A(B[6]), .B(A[6]), .Z(n1174) );
  NOR U5000 ( .A(B[7]), .B(A[7]), .Z(n1171) );
  AND U5001 ( .A(B[8]), .B(A[8]), .Z(n591) );
  AND U5002 ( .A(B[9]), .B(A[9]), .Z(n3) );
  NOR U5003 ( .A(B[10]), .B(A[10]), .Z(n5260) );
  AND U5004 ( .A(B[10]), .B(A[10]), .Z(n5259) );
  NOR U5005 ( .A(B[11]), .B(A[11]), .Z(n5256) );
  AND U5006 ( .A(B[11]), .B(A[11]), .Z(n5257) );
  AND U5007 ( .A(B[12]), .B(A[12]), .Z(n5202) );
  AND U5008 ( .A(B[13]), .B(A[13]), .Z(n5141) );
  AND U5009 ( .A(B[14]), .B(A[14]), .Z(n5087) );
  NOR U5010 ( .A(n4739), .B(n4264), .Z(n6126) );
  NAND U5011 ( .A(n6148), .B(n6149), .Z(n4739) );
  AND U5012 ( .A(n4918), .B(n4860), .Z(n6149) );
  OR U5013 ( .A(B[16]), .B(A[16]), .Z(n4918) );
  ANDN U5014 ( .B(n4798), .A(n4801), .Z(n6148) );
  ANDN U5015 ( .B(n6150), .A(n4201), .Z(n6124) );
  AND U5016 ( .A(B[28]), .B(A[28]), .Z(n4201) );
  NAND U5017 ( .A(n6151), .B(n4204), .Z(n6150) );
  OR U5018 ( .A(A[28]), .B(B[28]), .Z(n4204) );
  NANDN U5019 ( .A(n4262), .B(n6152), .Z(n6151) );
  NANDN U5020 ( .A(n4264), .B(n6153), .Z(n6152) );
  NANDN U5021 ( .A(n4501), .B(n6154), .Z(n6153) );
  NAND U5022 ( .A(n4738), .B(n4504), .Z(n6154) );
  AND U5023 ( .A(n6155), .B(n6156), .Z(n4504) );
  AND U5024 ( .A(n4678), .B(n4624), .Z(n6156) );
  OR U5025 ( .A(B[20]), .B(A[20]), .Z(n4678) );
  AND U5026 ( .A(n4561), .B(n4557), .Z(n6155) );
  NANDN U5027 ( .A(n4797), .B(n6157), .Z(n4738) );
  NAND U5028 ( .A(n6158), .B(n4798), .Z(n6157) );
  OR U5029 ( .A(B[19]), .B(A[19]), .Z(n4798) );
  NANDN U5030 ( .A(n4800), .B(n6159), .Z(n6158) );
  NANDN U5031 ( .A(n4801), .B(n6160), .Z(n6159) );
  NANDN U5032 ( .A(n4857), .B(n6161), .Z(n6160) );
  NAND U5033 ( .A(n4860), .B(n4916), .Z(n6161) );
  AND U5034 ( .A(A[16]), .B(B[16]), .Z(n4916) );
  OR U5035 ( .A(B[17]), .B(A[17]), .Z(n4860) );
  AND U5036 ( .A(B[17]), .B(A[17]), .Z(n4857) );
  NOR U5037 ( .A(B[18]), .B(A[18]), .Z(n4801) );
  AND U5038 ( .A(B[18]), .B(A[18]), .Z(n4800) );
  AND U5039 ( .A(B[19]), .B(A[19]), .Z(n4797) );
  NANDN U5040 ( .A(n4556), .B(n6162), .Z(n4501) );
  NAND U5041 ( .A(n6163), .B(n4557), .Z(n6162) );
  OR U5042 ( .A(B[23]), .B(A[23]), .Z(n4557) );
  NANDN U5043 ( .A(n4559), .B(n6164), .Z(n6163) );
  NAND U5044 ( .A(n6165), .B(n4561), .Z(n6164) );
  OR U5045 ( .A(B[22]), .B(A[22]), .Z(n4561) );
  NANDN U5046 ( .A(n4621), .B(n6166), .Z(n6165) );
  NAND U5047 ( .A(n4624), .B(n4676), .Z(n6166) );
  AND U5048 ( .A(B[20]), .B(A[20]), .Z(n4676) );
  OR U5049 ( .A(B[21]), .B(A[21]), .Z(n4624) );
  AND U5050 ( .A(B[21]), .B(A[21]), .Z(n4621) );
  AND U5051 ( .A(B[22]), .B(A[22]), .Z(n4559) );
  AND U5052 ( .A(B[23]), .B(A[23]), .Z(n4556) );
  NAND U5053 ( .A(n6167), .B(n6168), .Z(n4264) );
  AND U5054 ( .A(n4445), .B(n4388), .Z(n6168) );
  OR U5055 ( .A(B[24]), .B(A[24]), .Z(n4445) );
  AND U5056 ( .A(n4327), .B(n4323), .Z(n6167) );
  NANDN U5057 ( .A(n4322), .B(n6169), .Z(n4262) );
  NAND U5058 ( .A(n6170), .B(n4323), .Z(n6169) );
  OR U5059 ( .A(B[27]), .B(A[27]), .Z(n4323) );
  NANDN U5060 ( .A(n4325), .B(n6171), .Z(n6170) );
  NAND U5061 ( .A(n6172), .B(n4327), .Z(n6171) );
  OR U5062 ( .A(B[26]), .B(A[26]), .Z(n4327) );
  NANDN U5063 ( .A(n4385), .B(n6173), .Z(n6172) );
  NAND U5064 ( .A(n4388), .B(n4443), .Z(n6173) );
  AND U5065 ( .A(B[24]), .B(A[24]), .Z(n4443) );
  OR U5066 ( .A(B[25]), .B(A[25]), .Z(n4388) );
  AND U5067 ( .A(B[25]), .B(A[25]), .Z(n4385) );
  AND U5068 ( .A(B[26]), .B(A[26]), .Z(n4325) );
  AND U5069 ( .A(B[27]), .B(A[27]), .Z(n4322) );
  NOR U5070 ( .A(B[29]), .B(A[29]), .Z(n4140) );
  AND U5071 ( .A(B[29]), .B(A[29]), .Z(n4138) );
  NOR U5072 ( .A(B[30]), .B(A[30]), .Z(n4077) );
  AND U5073 ( .A(B[30]), .B(A[30]), .Z(n4076) );
  NOR U5074 ( .A(B[31]), .B(A[31]), .Z(n4073) );
  NOR U5075 ( .A(n3781), .B(n3294), .Z(n6115) );
  NAND U5076 ( .A(n6174), .B(n6175), .Z(n3781) );
  AND U5077 ( .A(n3962), .B(n3905), .Z(n6175) );
  OR U5078 ( .A(B[32]), .B(A[32]), .Z(n3962) );
  ANDN U5079 ( .B(n3840), .A(n3843), .Z(n6174) );
  ANDN U5080 ( .B(n6176), .A(n3231), .Z(n6113) );
  AND U5081 ( .A(B[44]), .B(A[44]), .Z(n3231) );
  NAND U5082 ( .A(n6177), .B(n3234), .Z(n6176) );
  OR U5083 ( .A(A[44]), .B(B[44]), .Z(n3234) );
  NANDN U5084 ( .A(n3292), .B(n6178), .Z(n6177) );
  NANDN U5085 ( .A(n3294), .B(n6179), .Z(n6178) );
  NANDN U5086 ( .A(n3536), .B(n6180), .Z(n6179) );
  NAND U5087 ( .A(n3780), .B(n3539), .Z(n6180) );
  AND U5088 ( .A(n6181), .B(n6182), .Z(n3539) );
  AND U5089 ( .A(n3720), .B(n3663), .Z(n6182) );
  OR U5090 ( .A(B[36]), .B(A[36]), .Z(n3720) );
  AND U5091 ( .A(n3600), .B(n3596), .Z(n6181) );
  NANDN U5092 ( .A(n3839), .B(n6183), .Z(n3780) );
  NAND U5093 ( .A(n6184), .B(n3840), .Z(n6183) );
  OR U5094 ( .A(B[35]), .B(A[35]), .Z(n3840) );
  NANDN U5095 ( .A(n3842), .B(n6185), .Z(n6184) );
  NANDN U5096 ( .A(n3843), .B(n6186), .Z(n6185) );
  NANDN U5097 ( .A(n3902), .B(n6187), .Z(n6186) );
  NAND U5098 ( .A(n3905), .B(n3960), .Z(n6187) );
  AND U5099 ( .A(A[32]), .B(B[32]), .Z(n3960) );
  OR U5100 ( .A(B[33]), .B(A[33]), .Z(n3905) );
  AND U5101 ( .A(B[33]), .B(A[33]), .Z(n3902) );
  NOR U5102 ( .A(B[34]), .B(A[34]), .Z(n3843) );
  AND U5103 ( .A(B[34]), .B(A[34]), .Z(n3842) );
  AND U5104 ( .A(B[35]), .B(A[35]), .Z(n3839) );
  NANDN U5105 ( .A(n3595), .B(n6188), .Z(n3536) );
  NAND U5106 ( .A(n6189), .B(n3596), .Z(n6188) );
  OR U5107 ( .A(B[39]), .B(A[39]), .Z(n3596) );
  NANDN U5108 ( .A(n3598), .B(n6190), .Z(n6189) );
  NAND U5109 ( .A(n6191), .B(n3600), .Z(n6190) );
  OR U5110 ( .A(B[38]), .B(A[38]), .Z(n3600) );
  NANDN U5111 ( .A(n3660), .B(n6192), .Z(n6191) );
  NAND U5112 ( .A(n3663), .B(n3718), .Z(n6192) );
  AND U5113 ( .A(B[36]), .B(A[36]), .Z(n3718) );
  OR U5114 ( .A(B[37]), .B(A[37]), .Z(n3663) );
  AND U5115 ( .A(B[37]), .B(A[37]), .Z(n3660) );
  AND U5116 ( .A(B[38]), .B(A[38]), .Z(n3598) );
  AND U5117 ( .A(B[39]), .B(A[39]), .Z(n3595) );
  NAND U5118 ( .A(n6193), .B(n6194), .Z(n3294) );
  AND U5119 ( .A(n3476), .B(n3419), .Z(n6194) );
  OR U5120 ( .A(B[40]), .B(A[40]), .Z(n3476) );
  AND U5121 ( .A(n3357), .B(n3353), .Z(n6193) );
  NANDN U5122 ( .A(n3352), .B(n6195), .Z(n3292) );
  NAND U5123 ( .A(n6196), .B(n3353), .Z(n6195) );
  OR U5124 ( .A(B[43]), .B(A[43]), .Z(n3353) );
  NANDN U5125 ( .A(n3355), .B(n6197), .Z(n6196) );
  NAND U5126 ( .A(n6198), .B(n3357), .Z(n6197) );
  OR U5127 ( .A(B[42]), .B(A[42]), .Z(n3357) );
  NANDN U5128 ( .A(n3416), .B(n6199), .Z(n6198) );
  NAND U5129 ( .A(n3419), .B(n3474), .Z(n6199) );
  AND U5130 ( .A(B[40]), .B(A[40]), .Z(n3474) );
  OR U5131 ( .A(B[41]), .B(A[41]), .Z(n3419) );
  AND U5132 ( .A(B[41]), .B(A[41]), .Z(n3416) );
  AND U5133 ( .A(B[42]), .B(A[42]), .Z(n3355) );
  AND U5134 ( .A(B[43]), .B(A[43]), .Z(n3352) );
  NOR U5135 ( .A(B[45]), .B(A[45]), .Z(n3175) );
  AND U5136 ( .A(B[45]), .B(A[45]), .Z(n3173) );
  NOR U5137 ( .A(B[46]), .B(A[46]), .Z(n3112) );
  AND U5138 ( .A(B[46]), .B(A[46]), .Z(n3111) );
  NOR U5139 ( .A(B[47]), .B(A[47]), .Z(n3108) );
  OR U5140 ( .A(B[51]), .B(A[51]), .Z(n2870) );
  NAND U5141 ( .A(n6200), .B(n6201), .Z(n2571) );
  AND U5142 ( .A(n2753), .B(n2696), .Z(n6201) );
  OR U5143 ( .A(A[52]), .B(B[52]), .Z(n2753) );
  AND U5144 ( .A(n2633), .B(n2629), .Z(n6200) );
  NANDN U5145 ( .A(n2628), .B(n6202), .Z(n2569) );
  NAND U5146 ( .A(n6203), .B(n2629), .Z(n6202) );
  OR U5147 ( .A(B[55]), .B(A[55]), .Z(n2629) );
  NANDN U5148 ( .A(n2631), .B(n6204), .Z(n6203) );
  NAND U5149 ( .A(n6205), .B(n2633), .Z(n6204) );
  OR U5150 ( .A(A[54]), .B(B[54]), .Z(n2633) );
  NANDN U5151 ( .A(n2693), .B(n6206), .Z(n6205) );
  NAND U5152 ( .A(n2696), .B(n2751), .Z(n6206) );
  AND U5153 ( .A(A[52]), .B(B[52]), .Z(n2751) );
  OR U5154 ( .A(A[53]), .B(B[53]), .Z(n2696) );
  AND U5155 ( .A(A[53]), .B(B[53]), .Z(n2693) );
  AND U5156 ( .A(A[54]), .B(B[54]), .Z(n2631) );
  AND U5157 ( .A(B[55]), .B(A[55]), .Z(n2628) );
  NAND U5158 ( .A(n6207), .B(n6208), .Z(n2327) );
  AND U5159 ( .A(n2511), .B(n2454), .Z(n6208) );
  OR U5160 ( .A(B[56]), .B(A[56]), .Z(n2511) );
  AND U5161 ( .A(n2394), .B(n2390), .Z(n6207) );
  NANDN U5162 ( .A(n2389), .B(n6209), .Z(n2325) );
  NAND U5163 ( .A(n6210), .B(n2390), .Z(n6209) );
  OR U5164 ( .A(B[59]), .B(A[59]), .Z(n2390) );
  NANDN U5165 ( .A(n2392), .B(n6211), .Z(n6210) );
  NAND U5166 ( .A(n6212), .B(n2394), .Z(n6211) );
  OR U5167 ( .A(B[58]), .B(A[58]), .Z(n2394) );
  NANDN U5168 ( .A(n2451), .B(n6213), .Z(n6212) );
  NAND U5169 ( .A(n2454), .B(n2509), .Z(n6213) );
  AND U5170 ( .A(B[56]), .B(A[56]), .Z(n2509) );
  OR U5171 ( .A(B[57]), .B(A[57]), .Z(n2454) );
  AND U5172 ( .A(B[57]), .B(A[57]), .Z(n2451) );
  AND U5173 ( .A(B[58]), .B(A[58]), .Z(n2392) );
  AND U5174 ( .A(B[59]), .B(A[59]), .Z(n2389) );
  NOR U5175 ( .A(B[60]), .B(A[60]), .Z(n2266) );
  AND U5176 ( .A(B[60]), .B(A[60]), .Z(n2264) );
  NOR U5177 ( .A(B[61]), .B(A[61]), .Z(n2207) );
  AND U5178 ( .A(B[61]), .B(A[61]), .Z(n2205) );
  NOR U5179 ( .A(B[62]), .B(A[62]), .Z(n2144) );
  AND U5180 ( .A(B[62]), .B(A[62]), .Z(n2143) );
  NOR U5181 ( .A(B[63]), .B(A[63]), .Z(n2140) );
  NAND U5182 ( .A(n6214), .B(n6215), .Z(n6085) );
  AND U5183 ( .A(n6216), .B(n6217), .Z(n6215) );
  ANDN U5184 ( .B(n1245), .A(n1299), .Z(n6217) );
  ANDN U5185 ( .B(n1178), .A(n1181), .Z(n6216) );
  ANDN U5186 ( .B(n6218), .A(n1846), .Z(n6214) );
  NAND U5187 ( .A(n6219), .B(n6220), .Z(n1846) );
  AND U5188 ( .A(n2027), .B(n1970), .Z(n6220) );
  OR U5189 ( .A(B[64]), .B(A[64]), .Z(n2027) );
  ANDN U5190 ( .B(n1905), .A(n1908), .Z(n6219) );
  ANDN U5191 ( .B(n1602), .A(n1361), .Z(n6218) );
  NANDN U5192 ( .A(n1177), .B(n6221), .Z(n5444) );
  NAND U5193 ( .A(n6222), .B(n1178), .Z(n6221) );
  OR U5194 ( .A(B[79]), .B(A[79]), .Z(n1178) );
  NANDN U5195 ( .A(n1180), .B(n6223), .Z(n6222) );
  NANDN U5196 ( .A(n1181), .B(n6224), .Z(n6223) );
  NANDN U5197 ( .A(n1242), .B(n6225), .Z(n6224) );
  NAND U5198 ( .A(n6226), .B(n1245), .Z(n6225) );
  OR U5199 ( .A(B[77]), .B(A[77]), .Z(n1245) );
  NANDN U5200 ( .A(n1297), .B(n6227), .Z(n6226) );
  NANDN U5201 ( .A(n1299), .B(n6228), .Z(n6227) );
  NANDN U5202 ( .A(n1359), .B(n6229), .Z(n6228) );
  NANDN U5203 ( .A(n1361), .B(n6230), .Z(n6229) );
  NANDN U5204 ( .A(n1599), .B(n6231), .Z(n6230) );
  NAND U5205 ( .A(n1845), .B(n1602), .Z(n6231) );
  AND U5206 ( .A(n6232), .B(n6233), .Z(n1602) );
  AND U5207 ( .A(n1785), .B(n1725), .Z(n6233) );
  OR U5208 ( .A(B[68]), .B(A[68]), .Z(n1785) );
  AND U5209 ( .A(n1662), .B(n1658), .Z(n6232) );
  NANDN U5210 ( .A(n1904), .B(n6234), .Z(n1845) );
  NAND U5211 ( .A(n6235), .B(n1905), .Z(n6234) );
  OR U5212 ( .A(B[67]), .B(A[67]), .Z(n1905) );
  NANDN U5213 ( .A(n1907), .B(n6236), .Z(n6235) );
  NANDN U5214 ( .A(n1908), .B(n6237), .Z(n6236) );
  NANDN U5215 ( .A(n1967), .B(n6238), .Z(n6237) );
  NAND U5216 ( .A(n1970), .B(n2025), .Z(n6238) );
  AND U5217 ( .A(A[64]), .B(B[64]), .Z(n2025) );
  OR U5218 ( .A(B[65]), .B(A[65]), .Z(n1970) );
  AND U5219 ( .A(B[65]), .B(A[65]), .Z(n1967) );
  NOR U5220 ( .A(B[66]), .B(A[66]), .Z(n1908) );
  AND U5221 ( .A(B[66]), .B(A[66]), .Z(n1907) );
  AND U5222 ( .A(B[67]), .B(A[67]), .Z(n1904) );
  NANDN U5223 ( .A(n1657), .B(n6239), .Z(n1599) );
  NAND U5224 ( .A(n6240), .B(n1658), .Z(n6239) );
  OR U5225 ( .A(B[71]), .B(A[71]), .Z(n1658) );
  NANDN U5226 ( .A(n1660), .B(n6241), .Z(n6240) );
  NAND U5227 ( .A(n6242), .B(n1662), .Z(n6241) );
  OR U5228 ( .A(B[70]), .B(A[70]), .Z(n1662) );
  NANDN U5229 ( .A(n1722), .B(n6243), .Z(n6242) );
  NAND U5230 ( .A(n1725), .B(n1783), .Z(n6243) );
  AND U5231 ( .A(B[68]), .B(A[68]), .Z(n1783) );
  OR U5232 ( .A(B[69]), .B(A[69]), .Z(n1725) );
  AND U5233 ( .A(B[69]), .B(A[69]), .Z(n1722) );
  AND U5234 ( .A(B[70]), .B(A[70]), .Z(n1660) );
  AND U5235 ( .A(B[71]), .B(A[71]), .Z(n1657) );
  NAND U5236 ( .A(n6244), .B(n6245), .Z(n1361) );
  AND U5237 ( .A(n1539), .B(n1482), .Z(n6245) );
  OR U5238 ( .A(B[72]), .B(A[72]), .Z(n1539) );
  AND U5239 ( .A(n1420), .B(n1416), .Z(n6244) );
  NANDN U5240 ( .A(n1415), .B(n6246), .Z(n1359) );
  NAND U5241 ( .A(n6247), .B(n1416), .Z(n6246) );
  OR U5242 ( .A(B[75]), .B(A[75]), .Z(n1416) );
  NANDN U5243 ( .A(n1418), .B(n6248), .Z(n6247) );
  NAND U5244 ( .A(n6249), .B(n1420), .Z(n6248) );
  OR U5245 ( .A(B[74]), .B(A[74]), .Z(n1420) );
  NANDN U5246 ( .A(n1479), .B(n6250), .Z(n6249) );
  NAND U5247 ( .A(n1482), .B(n1537), .Z(n6250) );
  AND U5248 ( .A(B[72]), .B(A[72]), .Z(n1537) );
  OR U5249 ( .A(B[73]), .B(A[73]), .Z(n1482) );
  AND U5250 ( .A(B[73]), .B(A[73]), .Z(n1479) );
  AND U5251 ( .A(B[74]), .B(A[74]), .Z(n1418) );
  AND U5252 ( .A(B[75]), .B(A[75]), .Z(n1415) );
  NOR U5253 ( .A(B[76]), .B(A[76]), .Z(n1299) );
  AND U5254 ( .A(B[76]), .B(A[76]), .Z(n1297) );
  AND U5255 ( .A(B[77]), .B(A[77]), .Z(n1242) );
  NOR U5256 ( .A(B[78]), .B(A[78]), .Z(n1181) );
  AND U5257 ( .A(B[78]), .B(A[78]), .Z(n1180) );
  AND U5258 ( .A(B[79]), .B(A[79]), .Z(n1177) );
  NAND U5259 ( .A(n6251), .B(n6252), .Z(n5442) );
  AND U5260 ( .A(n6253), .B(n6254), .Z(n6252) );
  ANDN U5261 ( .B(n300), .A(n354), .Z(n6254) );
  ANDN U5262 ( .B(n233), .A(n236), .Z(n6253) );
  ANDN U5263 ( .B(n6255), .A(n889), .Z(n6251) );
  NAND U5264 ( .A(n6256), .B(n6257), .Z(n889) );
  AND U5265 ( .A(n1064), .B(n1006), .Z(n6257) );
  OR U5266 ( .A(B[80]), .B(A[80]), .Z(n1064) );
  ANDN U5267 ( .B(n944), .A(n947), .Z(n6256) );
  ANDN U5268 ( .B(n654), .A(n416), .Z(n6255) );
  NANDN U5269 ( .A(n232), .B(n6258), .Z(n5441) );
  NAND U5270 ( .A(n6259), .B(n233), .Z(n6258) );
  OR U5271 ( .A(B[95]), .B(A[95]), .Z(n233) );
  NANDN U5272 ( .A(n235), .B(n6260), .Z(n6259) );
  NANDN U5273 ( .A(n236), .B(n6261), .Z(n6260) );
  NANDN U5274 ( .A(n297), .B(n6262), .Z(n6261) );
  NAND U5275 ( .A(n6263), .B(n300), .Z(n6262) );
  OR U5276 ( .A(B[93]), .B(A[93]), .Z(n300) );
  NANDN U5277 ( .A(n352), .B(n6264), .Z(n6263) );
  NANDN U5278 ( .A(n354), .B(n6265), .Z(n6264) );
  NANDN U5279 ( .A(n414), .B(n6266), .Z(n6265) );
  NANDN U5280 ( .A(n416), .B(n6267), .Z(n6266) );
  NANDN U5281 ( .A(n651), .B(n6268), .Z(n6267) );
  NAND U5282 ( .A(n888), .B(n654), .Z(n6268) );
  AND U5283 ( .A(n6269), .B(n6270), .Z(n654) );
  AND U5284 ( .A(n828), .B(n774), .Z(n6270) );
  OR U5285 ( .A(B[84]), .B(A[84]), .Z(n828) );
  AND U5286 ( .A(n711), .B(n707), .Z(n6269) );
  NANDN U5287 ( .A(n943), .B(n6271), .Z(n888) );
  NAND U5288 ( .A(n6272), .B(n944), .Z(n6271) );
  OR U5289 ( .A(B[83]), .B(A[83]), .Z(n944) );
  NANDN U5290 ( .A(n946), .B(n6273), .Z(n6272) );
  NANDN U5291 ( .A(n947), .B(n6274), .Z(n6273) );
  NANDN U5292 ( .A(n1003), .B(n6275), .Z(n6274) );
  NAND U5293 ( .A(n1006), .B(n1062), .Z(n6275) );
  AND U5294 ( .A(A[80]), .B(B[80]), .Z(n1062) );
  OR U5295 ( .A(B[81]), .B(A[81]), .Z(n1006) );
  AND U5296 ( .A(B[81]), .B(A[81]), .Z(n1003) );
  NOR U5297 ( .A(B[82]), .B(A[82]), .Z(n947) );
  AND U5298 ( .A(B[82]), .B(A[82]), .Z(n946) );
  AND U5299 ( .A(B[83]), .B(A[83]), .Z(n943) );
  NANDN U5300 ( .A(n706), .B(n6276), .Z(n651) );
  NAND U5301 ( .A(n6277), .B(n707), .Z(n6276) );
  OR U5302 ( .A(B[87]), .B(A[87]), .Z(n707) );
  NANDN U5303 ( .A(n709), .B(n6278), .Z(n6277) );
  NAND U5304 ( .A(n6279), .B(n711), .Z(n6278) );
  OR U5305 ( .A(B[86]), .B(A[86]), .Z(n711) );
  NANDN U5306 ( .A(n771), .B(n6280), .Z(n6279) );
  NAND U5307 ( .A(n774), .B(n826), .Z(n6280) );
  AND U5308 ( .A(B[84]), .B(A[84]), .Z(n826) );
  OR U5309 ( .A(B[85]), .B(A[85]), .Z(n774) );
  AND U5310 ( .A(B[85]), .B(A[85]), .Z(n771) );
  AND U5311 ( .A(B[86]), .B(A[86]), .Z(n709) );
  AND U5312 ( .A(B[87]), .B(A[87]), .Z(n706) );
  NAND U5313 ( .A(n6281), .B(n6282), .Z(n416) );
  AND U5314 ( .A(n595), .B(n533), .Z(n6282) );
  OR U5315 ( .A(B[88]), .B(A[88]), .Z(n595) );
  AND U5316 ( .A(n475), .B(n471), .Z(n6281) );
  NANDN U5317 ( .A(n470), .B(n6283), .Z(n414) );
  NAND U5318 ( .A(n6284), .B(n471), .Z(n6283) );
  OR U5319 ( .A(B[91]), .B(A[91]), .Z(n471) );
  NANDN U5320 ( .A(n473), .B(n6285), .Z(n6284) );
  NAND U5321 ( .A(n6286), .B(n475), .Z(n6285) );
  OR U5322 ( .A(B[90]), .B(A[90]), .Z(n475) );
  NANDN U5323 ( .A(n530), .B(n6287), .Z(n6286) );
  NAND U5324 ( .A(n533), .B(n593), .Z(n6287) );
  AND U5325 ( .A(B[88]), .B(A[88]), .Z(n593) );
  OR U5326 ( .A(B[89]), .B(A[89]), .Z(n533) );
  AND U5327 ( .A(B[89]), .B(A[89]), .Z(n530) );
  AND U5328 ( .A(B[90]), .B(A[90]), .Z(n473) );
  AND U5329 ( .A(B[91]), .B(A[91]), .Z(n470) );
  NOR U5330 ( .A(B[92]), .B(A[92]), .Z(n354) );
  AND U5331 ( .A(B[92]), .B(A[92]), .Z(n352) );
  AND U5332 ( .A(B[93]), .B(A[93]), .Z(n297) );
  NOR U5333 ( .A(B[94]), .B(A[94]), .Z(n236) );
  AND U5334 ( .A(B[94]), .B(A[94]), .Z(n235) );
  AND U5335 ( .A(B[95]), .B(A[95]), .Z(n232) );
  NAND U5336 ( .A(n6288), .B(n6289), .Z(n5304) );
  AND U5337 ( .A(n6290), .B(n6291), .Z(n6289) );
  AND U5338 ( .A(n5325), .B(n5317), .Z(n6291) );
  AND U5339 ( .A(n5312), .B(n5308), .Z(n6290) );
  ANDN U5340 ( .B(n6292), .A(n5439), .Z(n6288) );
  NAND U5341 ( .A(n6293), .B(n6294), .Z(n5439) );
  AND U5342 ( .A(n12), .B(n68), .Z(n6294) );
  ANDN U5343 ( .B(n8), .A(n124), .Z(n6293) );
  NOR U5344 ( .A(B[96]), .B(A[96]), .Z(n124) );
  ANDN U5345 ( .B(n5329), .A(n5351), .Z(n6292) );
  NANDN U5346 ( .A(n5307), .B(n6295), .Z(n5302) );
  NAND U5347 ( .A(n6296), .B(n5308), .Z(n6295) );
  OR U5348 ( .A(B[111]), .B(A[111]), .Z(n5308) );
  NANDN U5349 ( .A(n5310), .B(n6297), .Z(n6296) );
  NAND U5350 ( .A(n6298), .B(n5312), .Z(n6297) );
  OR U5351 ( .A(B[110]), .B(A[110]), .Z(n5312) );
  NANDN U5352 ( .A(n5314), .B(n6299), .Z(n6298) );
  NAND U5353 ( .A(n6300), .B(n5317), .Z(n6299) );
  OR U5354 ( .A(B[109]), .B(A[109]), .Z(n5317) );
  NANDN U5355 ( .A(n5322), .B(n6301), .Z(n6300) );
  NAND U5356 ( .A(n6302), .B(n5325), .Z(n6301) );
  OR U5357 ( .A(B[108]), .B(A[108]), .Z(n5325) );
  NANDN U5358 ( .A(n5327), .B(n6303), .Z(n6302) );
  NAND U5359 ( .A(n6304), .B(n5329), .Z(n6303) );
  AND U5360 ( .A(n6305), .B(n6306), .Z(n5329) );
  AND U5361 ( .A(n5347), .B(n5343), .Z(n6306) );
  OR U5362 ( .A(B[104]), .B(A[104]), .Z(n5347) );
  AND U5363 ( .A(n5338), .B(n5334), .Z(n6305) );
  NANDN U5364 ( .A(n5349), .B(n6307), .Z(n6304) );
  NANDN U5365 ( .A(n5351), .B(n5438), .Z(n6307) );
  NANDN U5366 ( .A(n7), .B(n6308), .Z(n5438) );
  NAND U5367 ( .A(n6309), .B(n8), .Z(n6308) );
  OR U5368 ( .A(B[99]), .B(A[99]), .Z(n8) );
  NANDN U5369 ( .A(n10), .B(n6310), .Z(n6309) );
  NAND U5370 ( .A(n6311), .B(n12), .Z(n6310) );
  OR U5371 ( .A(B[98]), .B(A[98]), .Z(n12) );
  NANDN U5372 ( .A(n65), .B(n6312), .Z(n6311) );
  NAND U5373 ( .A(n68), .B(n122), .Z(n6312) );
  AND U5374 ( .A(B[96]), .B(A[96]), .Z(n122) );
  OR U5375 ( .A(B[97]), .B(A[97]), .Z(n68) );
  AND U5376 ( .A(B[97]), .B(A[97]), .Z(n65) );
  AND U5377 ( .A(A[98]), .B(B[98]), .Z(n10) );
  AND U5378 ( .A(B[99]), .B(A[99]), .Z(n7) );
  NAND U5379 ( .A(n6313), .B(n6314), .Z(n5351) );
  AND U5380 ( .A(n5385), .B(n5365), .Z(n6314) );
  OR U5381 ( .A(B[100]), .B(A[100]), .Z(n5385) );
  AND U5382 ( .A(n5360), .B(n5356), .Z(n6313) );
  NANDN U5383 ( .A(n5355), .B(n6315), .Z(n5349) );
  NAND U5384 ( .A(n6316), .B(n5356), .Z(n6315) );
  OR U5385 ( .A(B[103]), .B(A[103]), .Z(n5356) );
  NANDN U5386 ( .A(n5358), .B(n6317), .Z(n6316) );
  NAND U5387 ( .A(n6318), .B(n5360), .Z(n6317) );
  OR U5388 ( .A(B[102]), .B(A[102]), .Z(n5360) );
  NANDN U5389 ( .A(n5362), .B(n6319), .Z(n6318) );
  NAND U5390 ( .A(n5365), .B(n5383), .Z(n6319) );
  AND U5391 ( .A(B[100]), .B(A[100]), .Z(n5383) );
  OR U5392 ( .A(B[101]), .B(A[101]), .Z(n5365) );
  AND U5393 ( .A(B[101]), .B(A[101]), .Z(n5362) );
  AND U5394 ( .A(B[102]), .B(A[102]), .Z(n5358) );
  AND U5395 ( .A(B[103]), .B(A[103]), .Z(n5355) );
  NANDN U5396 ( .A(n5333), .B(n6320), .Z(n5327) );
  NAND U5397 ( .A(n6321), .B(n5334), .Z(n6320) );
  OR U5398 ( .A(B[107]), .B(A[107]), .Z(n5334) );
  NANDN U5399 ( .A(n5336), .B(n6322), .Z(n6321) );
  NAND U5400 ( .A(n6323), .B(n5338), .Z(n6322) );
  OR U5401 ( .A(B[106]), .B(A[106]), .Z(n5338) );
  NANDN U5402 ( .A(n5340), .B(n6324), .Z(n6323) );
  NAND U5403 ( .A(n5343), .B(n5345), .Z(n6324) );
  AND U5404 ( .A(B[104]), .B(A[104]), .Z(n5345) );
  OR U5405 ( .A(B[105]), .B(A[105]), .Z(n5343) );
  AND U5406 ( .A(B[105]), .B(A[105]), .Z(n5340) );
  AND U5407 ( .A(B[106]), .B(A[106]), .Z(n5336) );
  AND U5408 ( .A(B[107]), .B(A[107]), .Z(n5333) );
  AND U5409 ( .A(B[108]), .B(A[108]), .Z(n5322) );
  AND U5410 ( .A(B[109]), .B(A[109]), .Z(n5314) );
  AND U5411 ( .A(B[110]), .B(A[110]), .Z(n5310) );
  AND U5412 ( .A(B[111]), .B(A[111]), .Z(n5307) );
  ANDN U5413 ( .B(n6325), .A(n5282), .Z(n6076) );
  NAND U5414 ( .A(n6326), .B(n6327), .Z(n5282) );
  AND U5415 ( .A(n5300), .B(n5296), .Z(n6327) );
  OR U5416 ( .A(B[112]), .B(A[112]), .Z(n5300) );
  ANDN U5417 ( .B(n5287), .A(n5290), .Z(n6326) );
  ANDN U5418 ( .B(n5253), .A(n5230), .Z(n6325) );
  ANDN U5419 ( .B(n6328), .A(n5214), .Z(n6074) );
  AND U5420 ( .A(B[126]), .B(A[126]), .Z(n5214) );
  NAND U5421 ( .A(n6329), .B(n5216), .Z(n6328) );
  OR U5422 ( .A(A[126]), .B(B[126]), .Z(n5216) );
  NANDN U5423 ( .A(n5218), .B(n6330), .Z(n6329) );
  NAND U5424 ( .A(n6331), .B(n5221), .Z(n6330) );
  OR U5425 ( .A(B[125]), .B(A[125]), .Z(n5221) );
  NANDN U5426 ( .A(n5223), .B(n6332), .Z(n6331) );
  NANDN U5427 ( .A(n5225), .B(n6333), .Z(n6332) );
  NANDN U5428 ( .A(n5228), .B(n6334), .Z(n6333) );
  NANDN U5429 ( .A(n5230), .B(n6335), .Z(n6334) );
  NANDN U5430 ( .A(n5250), .B(n6336), .Z(n6335) );
  NAND U5431 ( .A(n5281), .B(n5253), .Z(n6336) );
  AND U5432 ( .A(n6337), .B(n6338), .Z(n5253) );
  AND U5433 ( .A(n5278), .B(n5274), .Z(n6338) );
  OR U5434 ( .A(B[116]), .B(A[116]), .Z(n5278) );
  AND U5435 ( .A(n5269), .B(n5265), .Z(n6337) );
  NANDN U5436 ( .A(n5286), .B(n6339), .Z(n5281) );
  NAND U5437 ( .A(n6340), .B(n5287), .Z(n6339) );
  OR U5438 ( .A(B[115]), .B(A[115]), .Z(n5287) );
  NANDN U5439 ( .A(n5289), .B(n6341), .Z(n6340) );
  NANDN U5440 ( .A(n5290), .B(n6342), .Z(n6341) );
  NANDN U5441 ( .A(n5293), .B(n6343), .Z(n6342) );
  NAND U5442 ( .A(n5296), .B(n5298), .Z(n6343) );
  AND U5443 ( .A(A[112]), .B(B[112]), .Z(n5298) );
  OR U5444 ( .A(B[113]), .B(A[113]), .Z(n5296) );
  AND U5445 ( .A(B[113]), .B(A[113]), .Z(n5293) );
  NOR U5446 ( .A(B[114]), .B(A[114]), .Z(n5290) );
  AND U5447 ( .A(B[114]), .B(A[114]), .Z(n5289) );
  AND U5448 ( .A(B[115]), .B(A[115]), .Z(n5286) );
  NANDN U5449 ( .A(n5264), .B(n6344), .Z(n5250) );
  NAND U5450 ( .A(n6345), .B(n5265), .Z(n6344) );
  OR U5451 ( .A(B[119]), .B(A[119]), .Z(n5265) );
  NANDN U5452 ( .A(n5267), .B(n6346), .Z(n6345) );
  NAND U5453 ( .A(n6347), .B(n5269), .Z(n6346) );
  OR U5454 ( .A(B[118]), .B(A[118]), .Z(n5269) );
  NANDN U5455 ( .A(n5271), .B(n6348), .Z(n6347) );
  NAND U5456 ( .A(n5274), .B(n5276), .Z(n6348) );
  AND U5457 ( .A(B[116]), .B(A[116]), .Z(n5276) );
  OR U5458 ( .A(B[117]), .B(A[117]), .Z(n5274) );
  AND U5459 ( .A(B[117]), .B(A[117]), .Z(n5271) );
  AND U5460 ( .A(B[118]), .B(A[118]), .Z(n5267) );
  AND U5461 ( .A(B[119]), .B(A[119]), .Z(n5264) );
  NAND U5462 ( .A(n6349), .B(n6350), .Z(n5230) );
  AND U5463 ( .A(n5248), .B(n5244), .Z(n6350) );
  OR U5464 ( .A(B[120]), .B(A[120]), .Z(n5248) );
  AND U5465 ( .A(n5239), .B(n5235), .Z(n6349) );
  NANDN U5466 ( .A(n5234), .B(n6351), .Z(n5228) );
  NAND U5467 ( .A(n6352), .B(n5235), .Z(n6351) );
  OR U5468 ( .A(B[123]), .B(A[123]), .Z(n5235) );
  NANDN U5469 ( .A(n5237), .B(n6353), .Z(n6352) );
  NAND U5470 ( .A(n6354), .B(n5239), .Z(n6353) );
  OR U5471 ( .A(B[122]), .B(A[122]), .Z(n5239) );
  NANDN U5472 ( .A(n5241), .B(n6355), .Z(n6354) );
  NAND U5473 ( .A(n5244), .B(n5246), .Z(n6355) );
  AND U5474 ( .A(B[120]), .B(A[120]), .Z(n5246) );
  OR U5475 ( .A(B[121]), .B(A[121]), .Z(n5244) );
  AND U5476 ( .A(B[121]), .B(A[121]), .Z(n5241) );
  AND U5477 ( .A(B[122]), .B(A[122]), .Z(n5237) );
  AND U5478 ( .A(B[123]), .B(A[123]), .Z(n5234) );
  NOR U5479 ( .A(B[124]), .B(A[124]), .Z(n5225) );
  AND U5480 ( .A(B[124]), .B(A[124]), .Z(n5223) );
  AND U5481 ( .A(B[125]), .B(A[125]), .Z(n5218) );
  NOR U5482 ( .A(B[127]), .B(A[127]), .Z(n5211) );
  NAND U5483 ( .A(n6356), .B(n6357), .Z(n6071) );
  AND U5484 ( .A(n6358), .B(n6359), .Z(n6357) );
  AND U5485 ( .A(n5133), .B(n5128), .Z(n6359) );
  AND U5486 ( .A(n5123), .B(n5119), .Z(n6358) );
  ANDN U5487 ( .B(n6360), .A(n5185), .Z(n6356) );
  NAND U5488 ( .A(n6361), .B(n6362), .Z(n5185) );
  AND U5489 ( .A(n5207), .B(n5199), .Z(n6362) );
  OR U5490 ( .A(B[128]), .B(A[128]), .Z(n5207) );
  AND U5491 ( .A(n5194), .B(n5190), .Z(n6361) );
  ANDN U5492 ( .B(n5137), .A(n5163), .Z(n6360) );
  NANDN U5493 ( .A(n5118), .B(n6363), .Z(n6069) );
  NAND U5494 ( .A(n6364), .B(n5119), .Z(n6363) );
  OR U5495 ( .A(B[143]), .B(A[143]), .Z(n5119) );
  NANDN U5496 ( .A(n5121), .B(n6365), .Z(n6364) );
  NAND U5497 ( .A(n6366), .B(n5123), .Z(n6365) );
  OR U5498 ( .A(B[142]), .B(A[142]), .Z(n5123) );
  NANDN U5499 ( .A(n5125), .B(n6367), .Z(n6366) );
  NAND U5500 ( .A(n6368), .B(n5128), .Z(n6367) );
  OR U5501 ( .A(B[141]), .B(A[141]), .Z(n5128) );
  NANDN U5502 ( .A(n5130), .B(n6369), .Z(n6368) );
  NAND U5503 ( .A(n6370), .B(n5133), .Z(n6369) );
  OR U5504 ( .A(B[140]), .B(A[140]), .Z(n5133) );
  NANDN U5505 ( .A(n5135), .B(n6371), .Z(n6370) );
  NAND U5506 ( .A(n6372), .B(n5137), .Z(n6371) );
  AND U5507 ( .A(n6373), .B(n6374), .Z(n5137) );
  AND U5508 ( .A(n5159), .B(n5155), .Z(n6374) );
  OR U5509 ( .A(B[136]), .B(A[136]), .Z(n5159) );
  AND U5510 ( .A(n5150), .B(n5146), .Z(n6373) );
  NANDN U5511 ( .A(n5161), .B(n6375), .Z(n6372) );
  NANDN U5512 ( .A(n5163), .B(n5184), .Z(n6375) );
  NANDN U5513 ( .A(n5189), .B(n6376), .Z(n5184) );
  NAND U5514 ( .A(n6377), .B(n5190), .Z(n6376) );
  OR U5515 ( .A(B[131]), .B(A[131]), .Z(n5190) );
  NANDN U5516 ( .A(n5192), .B(n6378), .Z(n6377) );
  NAND U5517 ( .A(n6379), .B(n5194), .Z(n6378) );
  OR U5518 ( .A(B[130]), .B(A[130]), .Z(n5194) );
  NANDN U5519 ( .A(n5196), .B(n6380), .Z(n6379) );
  NAND U5520 ( .A(n5199), .B(n5205), .Z(n6380) );
  AND U5521 ( .A(B[128]), .B(A[128]), .Z(n5205) );
  OR U5522 ( .A(B[129]), .B(A[129]), .Z(n5199) );
  AND U5523 ( .A(B[129]), .B(A[129]), .Z(n5196) );
  AND U5524 ( .A(B[130]), .B(A[130]), .Z(n5192) );
  AND U5525 ( .A(B[131]), .B(A[131]), .Z(n5189) );
  NAND U5526 ( .A(n6381), .B(n6382), .Z(n5163) );
  AND U5527 ( .A(n5181), .B(n5177), .Z(n6382) );
  OR U5528 ( .A(B[132]), .B(A[132]), .Z(n5181) );
  AND U5529 ( .A(n5172), .B(n5168), .Z(n6381) );
  NANDN U5530 ( .A(n5167), .B(n6383), .Z(n5161) );
  NAND U5531 ( .A(n6384), .B(n5168), .Z(n6383) );
  OR U5532 ( .A(B[135]), .B(A[135]), .Z(n5168) );
  NANDN U5533 ( .A(n5170), .B(n6385), .Z(n6384) );
  NAND U5534 ( .A(n6386), .B(n5172), .Z(n6385) );
  OR U5535 ( .A(B[134]), .B(A[134]), .Z(n5172) );
  NANDN U5536 ( .A(n5174), .B(n6387), .Z(n6386) );
  NAND U5537 ( .A(n5177), .B(n5179), .Z(n6387) );
  AND U5538 ( .A(B[132]), .B(A[132]), .Z(n5179) );
  OR U5539 ( .A(B[133]), .B(A[133]), .Z(n5177) );
  AND U5540 ( .A(B[133]), .B(A[133]), .Z(n5174) );
  AND U5541 ( .A(B[134]), .B(A[134]), .Z(n5170) );
  AND U5542 ( .A(B[135]), .B(A[135]), .Z(n5167) );
  NANDN U5543 ( .A(n5145), .B(n6388), .Z(n5135) );
  NAND U5544 ( .A(n6389), .B(n5146), .Z(n6388) );
  OR U5545 ( .A(B[139]), .B(A[139]), .Z(n5146) );
  NANDN U5546 ( .A(n5148), .B(n6390), .Z(n6389) );
  NAND U5547 ( .A(n6391), .B(n5150), .Z(n6390) );
  OR U5548 ( .A(B[138]), .B(A[138]), .Z(n5150) );
  NANDN U5549 ( .A(n5152), .B(n6392), .Z(n6391) );
  NAND U5550 ( .A(n5155), .B(n5157), .Z(n6392) );
  AND U5551 ( .A(B[136]), .B(A[136]), .Z(n5157) );
  OR U5552 ( .A(B[137]), .B(A[137]), .Z(n5155) );
  AND U5553 ( .A(B[137]), .B(A[137]), .Z(n5152) );
  AND U5554 ( .A(B[138]), .B(A[138]), .Z(n5148) );
  AND U5555 ( .A(B[139]), .B(A[139]), .Z(n5145) );
  AND U5556 ( .A(B[140]), .B(A[140]), .Z(n5130) );
  AND U5557 ( .A(B[141]), .B(A[141]), .Z(n5125) );
  AND U5558 ( .A(B[142]), .B(A[142]), .Z(n5121) );
  AND U5559 ( .A(B[143]), .B(A[143]), .Z(n5118) );
  NAND U5560 ( .A(n6393), .B(n6394), .Z(n6068) );
  AND U5561 ( .A(n6395), .B(n6396), .Z(n6394) );
  AND U5562 ( .A(n5044), .B(n5039), .Z(n6396) );
  AND U5563 ( .A(n5034), .B(n5030), .Z(n6395) );
  ANDN U5564 ( .B(n6397), .A(n5096), .Z(n6393) );
  NAND U5565 ( .A(n6398), .B(n6399), .Z(n5096) );
  AND U5566 ( .A(n5114), .B(n5110), .Z(n6399) );
  OR U5567 ( .A(B[144]), .B(A[144]), .Z(n5114) );
  AND U5568 ( .A(n5105), .B(n5101), .Z(n6398) );
  ANDN U5569 ( .B(n5048), .A(n5070), .Z(n6397) );
  NANDN U5570 ( .A(n5029), .B(n6400), .Z(n6066) );
  NAND U5571 ( .A(n6401), .B(n5030), .Z(n6400) );
  OR U5572 ( .A(B[159]), .B(A[159]), .Z(n5030) );
  NANDN U5573 ( .A(n5032), .B(n6402), .Z(n6401) );
  NAND U5574 ( .A(n6403), .B(n5034), .Z(n6402) );
  OR U5575 ( .A(B[158]), .B(A[158]), .Z(n5034) );
  NANDN U5576 ( .A(n5036), .B(n6404), .Z(n6403) );
  NAND U5577 ( .A(n6405), .B(n5039), .Z(n6404) );
  OR U5578 ( .A(B[157]), .B(A[157]), .Z(n5039) );
  NANDN U5579 ( .A(n5041), .B(n6406), .Z(n6405) );
  NAND U5580 ( .A(n6407), .B(n5044), .Z(n6406) );
  OR U5581 ( .A(B[156]), .B(A[156]), .Z(n5044) );
  NANDN U5582 ( .A(n5046), .B(n6408), .Z(n6407) );
  NAND U5583 ( .A(n6409), .B(n5048), .Z(n6408) );
  AND U5584 ( .A(n6410), .B(n6411), .Z(n5048) );
  AND U5585 ( .A(n5066), .B(n5062), .Z(n6411) );
  OR U5586 ( .A(B[152]), .B(A[152]), .Z(n5066) );
  AND U5587 ( .A(n5057), .B(n5053), .Z(n6410) );
  NANDN U5588 ( .A(n5068), .B(n6412), .Z(n6409) );
  NANDN U5589 ( .A(n5070), .B(n5095), .Z(n6412) );
  NANDN U5590 ( .A(n5100), .B(n6413), .Z(n5095) );
  NAND U5591 ( .A(n6414), .B(n5101), .Z(n6413) );
  OR U5592 ( .A(B[147]), .B(A[147]), .Z(n5101) );
  NANDN U5593 ( .A(n5103), .B(n6415), .Z(n6414) );
  NAND U5594 ( .A(n6416), .B(n5105), .Z(n6415) );
  OR U5595 ( .A(B[146]), .B(A[146]), .Z(n5105) );
  NANDN U5596 ( .A(n5107), .B(n6417), .Z(n6416) );
  NAND U5597 ( .A(n5110), .B(n5112), .Z(n6417) );
  AND U5598 ( .A(B[144]), .B(A[144]), .Z(n5112) );
  OR U5599 ( .A(B[145]), .B(A[145]), .Z(n5110) );
  AND U5600 ( .A(B[145]), .B(A[145]), .Z(n5107) );
  AND U5601 ( .A(B[146]), .B(A[146]), .Z(n5103) );
  AND U5602 ( .A(B[147]), .B(A[147]), .Z(n5100) );
  NAND U5603 ( .A(n6418), .B(n6419), .Z(n5070) );
  AND U5604 ( .A(n5092), .B(n5084), .Z(n6419) );
  OR U5605 ( .A(B[148]), .B(A[148]), .Z(n5092) );
  AND U5606 ( .A(n5079), .B(n5075), .Z(n6418) );
  NANDN U5607 ( .A(n5074), .B(n6420), .Z(n5068) );
  NAND U5608 ( .A(n6421), .B(n5075), .Z(n6420) );
  OR U5609 ( .A(B[151]), .B(A[151]), .Z(n5075) );
  NANDN U5610 ( .A(n5077), .B(n6422), .Z(n6421) );
  NAND U5611 ( .A(n6423), .B(n5079), .Z(n6422) );
  OR U5612 ( .A(B[150]), .B(A[150]), .Z(n5079) );
  NANDN U5613 ( .A(n5081), .B(n6424), .Z(n6423) );
  NAND U5614 ( .A(n5084), .B(n5090), .Z(n6424) );
  AND U5615 ( .A(B[148]), .B(A[148]), .Z(n5090) );
  OR U5616 ( .A(B[149]), .B(A[149]), .Z(n5084) );
  AND U5617 ( .A(B[149]), .B(A[149]), .Z(n5081) );
  AND U5618 ( .A(B[150]), .B(A[150]), .Z(n5077) );
  AND U5619 ( .A(B[151]), .B(A[151]), .Z(n5074) );
  NANDN U5620 ( .A(n5052), .B(n6425), .Z(n5046) );
  NAND U5621 ( .A(n6426), .B(n5053), .Z(n6425) );
  OR U5622 ( .A(B[155]), .B(A[155]), .Z(n5053) );
  NANDN U5623 ( .A(n5055), .B(n6427), .Z(n6426) );
  NAND U5624 ( .A(n6428), .B(n5057), .Z(n6427) );
  OR U5625 ( .A(B[154]), .B(A[154]), .Z(n5057) );
  NANDN U5626 ( .A(n5059), .B(n6429), .Z(n6428) );
  NAND U5627 ( .A(n5062), .B(n5064), .Z(n6429) );
  AND U5628 ( .A(B[152]), .B(A[152]), .Z(n5064) );
  OR U5629 ( .A(B[153]), .B(A[153]), .Z(n5062) );
  AND U5630 ( .A(B[153]), .B(A[153]), .Z(n5059) );
  AND U5631 ( .A(B[154]), .B(A[154]), .Z(n5055) );
  AND U5632 ( .A(B[155]), .B(A[155]), .Z(n5052) );
  AND U5633 ( .A(B[156]), .B(A[156]), .Z(n5041) );
  AND U5634 ( .A(B[157]), .B(A[157]), .Z(n5036) );
  AND U5635 ( .A(B[158]), .B(A[158]), .Z(n5032) );
  AND U5636 ( .A(B[159]), .B(A[159]), .Z(n5029) );
  NAND U5637 ( .A(n6430), .B(n6431), .Z(n6065) );
  AND U5638 ( .A(n6432), .B(n6433), .Z(n6431) );
  AND U5639 ( .A(n4954), .B(n4949), .Z(n6433) );
  AND U5640 ( .A(n4944), .B(n4940), .Z(n6432) );
  ANDN U5641 ( .B(n6434), .A(n5003), .Z(n6430) );
  NAND U5642 ( .A(n6435), .B(n6436), .Z(n5003) );
  AND U5643 ( .A(n5021), .B(n5017), .Z(n6436) );
  OR U5644 ( .A(B[160]), .B(A[160]), .Z(n5021) );
  AND U5645 ( .A(n5012), .B(n5008), .Z(n6435) );
  ANDN U5646 ( .B(n4958), .A(n4981), .Z(n6434) );
  NANDN U5647 ( .A(n4939), .B(n6437), .Z(n6063) );
  NAND U5648 ( .A(n6438), .B(n4940), .Z(n6437) );
  OR U5649 ( .A(B[175]), .B(A[175]), .Z(n4940) );
  NANDN U5650 ( .A(n4942), .B(n6439), .Z(n6438) );
  NAND U5651 ( .A(n6440), .B(n4944), .Z(n6439) );
  OR U5652 ( .A(B[174]), .B(A[174]), .Z(n4944) );
  NANDN U5653 ( .A(n4946), .B(n6441), .Z(n6440) );
  NAND U5654 ( .A(n6442), .B(n4949), .Z(n6441) );
  OR U5655 ( .A(B[173]), .B(A[173]), .Z(n4949) );
  NANDN U5656 ( .A(n4951), .B(n6443), .Z(n6442) );
  NAND U5657 ( .A(n6444), .B(n4954), .Z(n6443) );
  OR U5658 ( .A(B[172]), .B(A[172]), .Z(n4954) );
  NANDN U5659 ( .A(n4956), .B(n6445), .Z(n6444) );
  NAND U5660 ( .A(n6446), .B(n4958), .Z(n6445) );
  AND U5661 ( .A(n6447), .B(n6448), .Z(n4958) );
  AND U5662 ( .A(n4977), .B(n4972), .Z(n6448) );
  OR U5663 ( .A(B[168]), .B(A[168]), .Z(n4977) );
  AND U5664 ( .A(n4967), .B(n4963), .Z(n6447) );
  NANDN U5665 ( .A(n4979), .B(n6449), .Z(n6446) );
  NANDN U5666 ( .A(n4981), .B(n5002), .Z(n6449) );
  NANDN U5667 ( .A(n5007), .B(n6450), .Z(n5002) );
  NAND U5668 ( .A(n6451), .B(n5008), .Z(n6450) );
  OR U5669 ( .A(B[163]), .B(A[163]), .Z(n5008) );
  NANDN U5670 ( .A(n5010), .B(n6452), .Z(n6451) );
  NAND U5671 ( .A(n6453), .B(n5012), .Z(n6452) );
  OR U5672 ( .A(B[162]), .B(A[162]), .Z(n5012) );
  NANDN U5673 ( .A(n5014), .B(n6454), .Z(n6453) );
  NAND U5674 ( .A(n5017), .B(n5019), .Z(n6454) );
  AND U5675 ( .A(B[160]), .B(A[160]), .Z(n5019) );
  OR U5676 ( .A(B[161]), .B(A[161]), .Z(n5017) );
  AND U5677 ( .A(B[161]), .B(A[161]), .Z(n5014) );
  AND U5678 ( .A(B[162]), .B(A[162]), .Z(n5010) );
  AND U5679 ( .A(B[163]), .B(A[163]), .Z(n5007) );
  NAND U5680 ( .A(n6455), .B(n6456), .Z(n4981) );
  AND U5681 ( .A(n4999), .B(n4995), .Z(n6456) );
  OR U5682 ( .A(B[164]), .B(A[164]), .Z(n4999) );
  AND U5683 ( .A(n4990), .B(n4986), .Z(n6455) );
  NANDN U5684 ( .A(n4985), .B(n6457), .Z(n4979) );
  NAND U5685 ( .A(n6458), .B(n4986), .Z(n6457) );
  OR U5686 ( .A(B[167]), .B(A[167]), .Z(n4986) );
  NANDN U5687 ( .A(n4988), .B(n6459), .Z(n6458) );
  NAND U5688 ( .A(n6460), .B(n4990), .Z(n6459) );
  OR U5689 ( .A(B[166]), .B(A[166]), .Z(n4990) );
  NANDN U5690 ( .A(n4992), .B(n6461), .Z(n6460) );
  NAND U5691 ( .A(n4995), .B(n4997), .Z(n6461) );
  AND U5692 ( .A(B[164]), .B(A[164]), .Z(n4997) );
  OR U5693 ( .A(B[165]), .B(A[165]), .Z(n4995) );
  AND U5694 ( .A(B[165]), .B(A[165]), .Z(n4992) );
  AND U5695 ( .A(B[166]), .B(A[166]), .Z(n4988) );
  AND U5696 ( .A(B[167]), .B(A[167]), .Z(n4985) );
  NANDN U5697 ( .A(n4962), .B(n6462), .Z(n4956) );
  NAND U5698 ( .A(n6463), .B(n4963), .Z(n6462) );
  OR U5699 ( .A(B[171]), .B(A[171]), .Z(n4963) );
  NANDN U5700 ( .A(n4965), .B(n6464), .Z(n6463) );
  NAND U5701 ( .A(n6465), .B(n4967), .Z(n6464) );
  OR U5702 ( .A(B[170]), .B(A[170]), .Z(n4967) );
  NANDN U5703 ( .A(n4969), .B(n6466), .Z(n6465) );
  NAND U5704 ( .A(n4972), .B(n4975), .Z(n6466) );
  AND U5705 ( .A(B[168]), .B(A[168]), .Z(n4975) );
  OR U5706 ( .A(B[169]), .B(A[169]), .Z(n4972) );
  AND U5707 ( .A(B[169]), .B(A[169]), .Z(n4969) );
  AND U5708 ( .A(B[170]), .B(A[170]), .Z(n4965) );
  AND U5709 ( .A(B[171]), .B(A[171]), .Z(n4962) );
  AND U5710 ( .A(B[172]), .B(A[172]), .Z(n4951) );
  AND U5711 ( .A(B[173]), .B(A[173]), .Z(n4946) );
  AND U5712 ( .A(B[174]), .B(A[174]), .Z(n4942) );
  AND U5713 ( .A(B[175]), .B(A[175]), .Z(n4939) );
  ANDN U5714 ( .B(n6467), .A(n4913), .Z(n6059) );
  NAND U5715 ( .A(n6468), .B(n6469), .Z(n4913) );
  AND U5716 ( .A(n4935), .B(n4931), .Z(n6469) );
  OR U5717 ( .A(B[176]), .B(A[176]), .Z(n4935) );
  ANDN U5718 ( .B(n4922), .A(n4925), .Z(n6468) );
  ANDN U5719 ( .B(n4892), .A(n4869), .Z(n6467) );
  ANDN U5720 ( .B(n6470), .A(n4848), .Z(n6057) );
  AND U5721 ( .A(B[190]), .B(A[190]), .Z(n4848) );
  NAND U5722 ( .A(n6471), .B(n4850), .Z(n6470) );
  OR U5723 ( .A(A[190]), .B(B[190]), .Z(n4850) );
  NANDN U5724 ( .A(n4852), .B(n6472), .Z(n6471) );
  NAND U5725 ( .A(n6473), .B(n4855), .Z(n6472) );
  OR U5726 ( .A(B[189]), .B(A[189]), .Z(n4855) );
  NANDN U5727 ( .A(n4862), .B(n6474), .Z(n6473) );
  NANDN U5728 ( .A(n4864), .B(n6475), .Z(n6474) );
  NANDN U5729 ( .A(n4867), .B(n6476), .Z(n6475) );
  NANDN U5730 ( .A(n4869), .B(n6477), .Z(n6476) );
  NANDN U5731 ( .A(n4889), .B(n6478), .Z(n6477) );
  NAND U5732 ( .A(n4912), .B(n4892), .Z(n6478) );
  AND U5733 ( .A(n6479), .B(n6480), .Z(n4892) );
  AND U5734 ( .A(n4909), .B(n4905), .Z(n6480) );
  OR U5735 ( .A(B[180]), .B(A[180]), .Z(n4909) );
  AND U5736 ( .A(n4900), .B(n4896), .Z(n6479) );
  NANDN U5737 ( .A(n4921), .B(n6481), .Z(n4912) );
  NAND U5738 ( .A(n6482), .B(n4922), .Z(n6481) );
  OR U5739 ( .A(B[179]), .B(A[179]), .Z(n4922) );
  NANDN U5740 ( .A(n4924), .B(n6483), .Z(n6482) );
  NANDN U5741 ( .A(n4925), .B(n6484), .Z(n6483) );
  NANDN U5742 ( .A(n4928), .B(n6485), .Z(n6484) );
  NAND U5743 ( .A(n4931), .B(n4933), .Z(n6485) );
  AND U5744 ( .A(A[176]), .B(B[176]), .Z(n4933) );
  OR U5745 ( .A(B[177]), .B(A[177]), .Z(n4931) );
  AND U5746 ( .A(B[177]), .B(A[177]), .Z(n4928) );
  NOR U5747 ( .A(B[178]), .B(A[178]), .Z(n4925) );
  AND U5748 ( .A(B[178]), .B(A[178]), .Z(n4924) );
  AND U5749 ( .A(B[179]), .B(A[179]), .Z(n4921) );
  NANDN U5750 ( .A(n4895), .B(n6486), .Z(n4889) );
  NAND U5751 ( .A(n6487), .B(n4896), .Z(n6486) );
  OR U5752 ( .A(B[183]), .B(A[183]), .Z(n4896) );
  NANDN U5753 ( .A(n4898), .B(n6488), .Z(n6487) );
  NAND U5754 ( .A(n6489), .B(n4900), .Z(n6488) );
  OR U5755 ( .A(B[182]), .B(A[182]), .Z(n4900) );
  NANDN U5756 ( .A(n4902), .B(n6490), .Z(n6489) );
  NAND U5757 ( .A(n4905), .B(n4907), .Z(n6490) );
  AND U5758 ( .A(B[180]), .B(A[180]), .Z(n4907) );
  OR U5759 ( .A(B[181]), .B(A[181]), .Z(n4905) );
  AND U5760 ( .A(B[181]), .B(A[181]), .Z(n4902) );
  AND U5761 ( .A(B[182]), .B(A[182]), .Z(n4898) );
  AND U5762 ( .A(B[183]), .B(A[183]), .Z(n4895) );
  NAND U5763 ( .A(n6491), .B(n6492), .Z(n4869) );
  AND U5764 ( .A(n4887), .B(n4883), .Z(n6492) );
  OR U5765 ( .A(B[184]), .B(A[184]), .Z(n4887) );
  AND U5766 ( .A(n4878), .B(n4874), .Z(n6491) );
  NANDN U5767 ( .A(n4873), .B(n6493), .Z(n4867) );
  NAND U5768 ( .A(n6494), .B(n4874), .Z(n6493) );
  OR U5769 ( .A(B[187]), .B(A[187]), .Z(n4874) );
  NANDN U5770 ( .A(n4876), .B(n6495), .Z(n6494) );
  NAND U5771 ( .A(n6496), .B(n4878), .Z(n6495) );
  OR U5772 ( .A(B[186]), .B(A[186]), .Z(n4878) );
  NANDN U5773 ( .A(n4880), .B(n6497), .Z(n6496) );
  NAND U5774 ( .A(n4883), .B(n4885), .Z(n6497) );
  AND U5775 ( .A(B[184]), .B(A[184]), .Z(n4885) );
  OR U5776 ( .A(B[185]), .B(A[185]), .Z(n4883) );
  AND U5777 ( .A(B[185]), .B(A[185]), .Z(n4880) );
  AND U5778 ( .A(B[186]), .B(A[186]), .Z(n4876) );
  AND U5779 ( .A(B[187]), .B(A[187]), .Z(n4873) );
  NOR U5780 ( .A(B[188]), .B(A[188]), .Z(n4864) );
  AND U5781 ( .A(B[188]), .B(A[188]), .Z(n4862) );
  AND U5782 ( .A(B[189]), .B(A[189]), .Z(n4852) );
  NOR U5783 ( .A(B[191]), .B(A[191]), .Z(n4845) );
  NOR U5784 ( .A(n4823), .B(n4767), .Z(n6052) );
  NAND U5785 ( .A(n6498), .B(n6499), .Z(n4823) );
  AND U5786 ( .A(n4841), .B(n4837), .Z(n6499) );
  OR U5787 ( .A(B[192]), .B(A[192]), .Z(n4841) );
  ANDN U5788 ( .B(n4828), .A(n4831), .Z(n6498) );
  ANDN U5789 ( .B(n6500), .A(n4760), .Z(n6050) );
  AND U5790 ( .A(B[204]), .B(A[204]), .Z(n4760) );
  NAND U5791 ( .A(n6501), .B(n4763), .Z(n6500) );
  OR U5792 ( .A(A[204]), .B(B[204]), .Z(n4763) );
  NANDN U5793 ( .A(n4765), .B(n6502), .Z(n6501) );
  NANDN U5794 ( .A(n4767), .B(n6503), .Z(n6502) );
  NANDN U5795 ( .A(n4787), .B(n6504), .Z(n6503) );
  NAND U5796 ( .A(n4822), .B(n4790), .Z(n6504) );
  AND U5797 ( .A(n6505), .B(n6506), .Z(n4790) );
  AND U5798 ( .A(n4819), .B(n4815), .Z(n6506) );
  OR U5799 ( .A(B[196]), .B(A[196]), .Z(n4819) );
  AND U5800 ( .A(n4810), .B(n4806), .Z(n6505) );
  NANDN U5801 ( .A(n4827), .B(n6507), .Z(n4822) );
  NAND U5802 ( .A(n6508), .B(n4828), .Z(n6507) );
  OR U5803 ( .A(B[195]), .B(A[195]), .Z(n4828) );
  NANDN U5804 ( .A(n4830), .B(n6509), .Z(n6508) );
  NANDN U5805 ( .A(n4831), .B(n6510), .Z(n6509) );
  NANDN U5806 ( .A(n4834), .B(n6511), .Z(n6510) );
  NAND U5807 ( .A(n4837), .B(n4839), .Z(n6511) );
  AND U5808 ( .A(A[192]), .B(B[192]), .Z(n4839) );
  OR U5809 ( .A(B[193]), .B(A[193]), .Z(n4837) );
  AND U5810 ( .A(B[193]), .B(A[193]), .Z(n4834) );
  NOR U5811 ( .A(B[194]), .B(A[194]), .Z(n4831) );
  AND U5812 ( .A(B[194]), .B(A[194]), .Z(n4830) );
  AND U5813 ( .A(B[195]), .B(A[195]), .Z(n4827) );
  NANDN U5814 ( .A(n4805), .B(n6512), .Z(n4787) );
  NAND U5815 ( .A(n6513), .B(n4806), .Z(n6512) );
  OR U5816 ( .A(B[199]), .B(A[199]), .Z(n4806) );
  NANDN U5817 ( .A(n4808), .B(n6514), .Z(n6513) );
  NAND U5818 ( .A(n6515), .B(n4810), .Z(n6514) );
  OR U5819 ( .A(B[198]), .B(A[198]), .Z(n4810) );
  NANDN U5820 ( .A(n4812), .B(n6516), .Z(n6515) );
  NAND U5821 ( .A(n4815), .B(n4817), .Z(n6516) );
  AND U5822 ( .A(B[196]), .B(A[196]), .Z(n4817) );
  OR U5823 ( .A(B[197]), .B(A[197]), .Z(n4815) );
  AND U5824 ( .A(B[197]), .B(A[197]), .Z(n4812) );
  AND U5825 ( .A(B[198]), .B(A[198]), .Z(n4808) );
  AND U5826 ( .A(B[199]), .B(A[199]), .Z(n4805) );
  NAND U5827 ( .A(n6517), .B(n6518), .Z(n4767) );
  AND U5828 ( .A(n4785), .B(n4781), .Z(n6518) );
  OR U5829 ( .A(B[200]), .B(A[200]), .Z(n4785) );
  AND U5830 ( .A(n4776), .B(n4772), .Z(n6517) );
  NANDN U5831 ( .A(n4771), .B(n6519), .Z(n4765) );
  NAND U5832 ( .A(n6520), .B(n4772), .Z(n6519) );
  OR U5833 ( .A(B[203]), .B(A[203]), .Z(n4772) );
  NANDN U5834 ( .A(n4774), .B(n6521), .Z(n6520) );
  NAND U5835 ( .A(n6522), .B(n4776), .Z(n6521) );
  OR U5836 ( .A(B[202]), .B(A[202]), .Z(n4776) );
  NANDN U5837 ( .A(n4778), .B(n6523), .Z(n6522) );
  NAND U5838 ( .A(n4781), .B(n4783), .Z(n6523) );
  AND U5839 ( .A(B[200]), .B(A[200]), .Z(n4783) );
  OR U5840 ( .A(B[201]), .B(A[201]), .Z(n4781) );
  AND U5841 ( .A(B[201]), .B(A[201]), .Z(n4778) );
  AND U5842 ( .A(B[202]), .B(A[202]), .Z(n4774) );
  AND U5843 ( .A(B[203]), .B(A[203]), .Z(n4771) );
  NOR U5844 ( .A(B[205]), .B(A[205]), .Z(n4757) );
  AND U5845 ( .A(B[205]), .B(A[205]), .Z(n4755) );
  NOR U5846 ( .A(B[206]), .B(A[206]), .Z(n4752) );
  AND U5847 ( .A(B[206]), .B(A[206]), .Z(n4751) );
  NOR U5848 ( .A(B[207]), .B(A[207]), .Z(n4748) );
  NOR U5849 ( .A(n4721), .B(n4673), .Z(n6041) );
  NAND U5850 ( .A(n6524), .B(n6525), .Z(n4721) );
  AND U5851 ( .A(n4744), .B(n4735), .Z(n6525) );
  OR U5852 ( .A(B[208]), .B(A[208]), .Z(n4744) );
  ANDN U5853 ( .B(n4726), .A(n4729), .Z(n6524) );
  ANDN U5854 ( .B(n6526), .A(n4666), .Z(n6039) );
  AND U5855 ( .A(B[220]), .B(A[220]), .Z(n4666) );
  NAND U5856 ( .A(n6527), .B(n4669), .Z(n6526) );
  OR U5857 ( .A(A[220]), .B(B[220]), .Z(n4669) );
  NANDN U5858 ( .A(n4671), .B(n6528), .Z(n6527) );
  NANDN U5859 ( .A(n4673), .B(n6529), .Z(n6528) );
  NANDN U5860 ( .A(n4697), .B(n6530), .Z(n6529) );
  NAND U5861 ( .A(n4720), .B(n4700), .Z(n6530) );
  AND U5862 ( .A(n6531), .B(n6532), .Z(n4700) );
  AND U5863 ( .A(n4717), .B(n4713), .Z(n6532) );
  OR U5864 ( .A(B[212]), .B(A[212]), .Z(n4717) );
  AND U5865 ( .A(n4708), .B(n4704), .Z(n6531) );
  NANDN U5866 ( .A(n4725), .B(n6533), .Z(n4720) );
  NAND U5867 ( .A(n6534), .B(n4726), .Z(n6533) );
  OR U5868 ( .A(B[211]), .B(A[211]), .Z(n4726) );
  NANDN U5869 ( .A(n4728), .B(n6535), .Z(n6534) );
  NANDN U5870 ( .A(n4729), .B(n6536), .Z(n6535) );
  NANDN U5871 ( .A(n4732), .B(n6537), .Z(n6536) );
  NAND U5872 ( .A(n4735), .B(n4742), .Z(n6537) );
  AND U5873 ( .A(A[208]), .B(B[208]), .Z(n4742) );
  OR U5874 ( .A(B[209]), .B(A[209]), .Z(n4735) );
  AND U5875 ( .A(B[209]), .B(A[209]), .Z(n4732) );
  NOR U5876 ( .A(B[210]), .B(A[210]), .Z(n4729) );
  AND U5877 ( .A(B[210]), .B(A[210]), .Z(n4728) );
  AND U5878 ( .A(B[211]), .B(A[211]), .Z(n4725) );
  NANDN U5879 ( .A(n4703), .B(n6538), .Z(n4697) );
  NAND U5880 ( .A(n6539), .B(n4704), .Z(n6538) );
  OR U5881 ( .A(B[215]), .B(A[215]), .Z(n4704) );
  NANDN U5882 ( .A(n4706), .B(n6540), .Z(n6539) );
  NAND U5883 ( .A(n6541), .B(n4708), .Z(n6540) );
  OR U5884 ( .A(B[214]), .B(A[214]), .Z(n4708) );
  NANDN U5885 ( .A(n4710), .B(n6542), .Z(n6541) );
  NAND U5886 ( .A(n4713), .B(n4715), .Z(n6542) );
  AND U5887 ( .A(B[212]), .B(A[212]), .Z(n4715) );
  OR U5888 ( .A(B[213]), .B(A[213]), .Z(n4713) );
  AND U5889 ( .A(B[213]), .B(A[213]), .Z(n4710) );
  AND U5890 ( .A(B[214]), .B(A[214]), .Z(n4706) );
  AND U5891 ( .A(B[215]), .B(A[215]), .Z(n4703) );
  NAND U5892 ( .A(n6543), .B(n6544), .Z(n4673) );
  AND U5893 ( .A(n4695), .B(n4691), .Z(n6544) );
  OR U5894 ( .A(B[216]), .B(A[216]), .Z(n4695) );
  AND U5895 ( .A(n4686), .B(n4682), .Z(n6543) );
  NANDN U5896 ( .A(n4681), .B(n6545), .Z(n4671) );
  NAND U5897 ( .A(n6546), .B(n4682), .Z(n6545) );
  OR U5898 ( .A(B[219]), .B(A[219]), .Z(n4682) );
  NANDN U5899 ( .A(n4684), .B(n6547), .Z(n6546) );
  NAND U5900 ( .A(n6548), .B(n4686), .Z(n6547) );
  OR U5901 ( .A(B[218]), .B(A[218]), .Z(n4686) );
  NANDN U5902 ( .A(n4688), .B(n6549), .Z(n6548) );
  NAND U5903 ( .A(n4691), .B(n4693), .Z(n6549) );
  AND U5904 ( .A(B[216]), .B(A[216]), .Z(n4693) );
  OR U5905 ( .A(B[217]), .B(A[217]), .Z(n4691) );
  AND U5906 ( .A(B[217]), .B(A[217]), .Z(n4688) );
  AND U5907 ( .A(B[218]), .B(A[218]), .Z(n4684) );
  AND U5908 ( .A(B[219]), .B(A[219]), .Z(n4681) );
  NOR U5909 ( .A(B[221]), .B(A[221]), .Z(n4663) );
  AND U5910 ( .A(B[221]), .B(A[221]), .Z(n4661) );
  NOR U5911 ( .A(B[222]), .B(A[222]), .Z(n4658) );
  AND U5912 ( .A(B[222]), .B(A[222]), .Z(n4657) );
  NOR U5913 ( .A(B[223]), .B(A[223]), .Z(n4654) );
  NOR U5914 ( .A(n4632), .B(n4583), .Z(n6030) );
  NAND U5915 ( .A(n6550), .B(n6551), .Z(n4632) );
  AND U5916 ( .A(n4650), .B(n4646), .Z(n6551) );
  OR U5917 ( .A(B[224]), .B(A[224]), .Z(n4650) );
  ANDN U5918 ( .B(n4637), .A(n4640), .Z(n6550) );
  ANDN U5919 ( .B(n6552), .A(n4576), .Z(n6028) );
  AND U5920 ( .A(B[236]), .B(A[236]), .Z(n4576) );
  NAND U5921 ( .A(n6553), .B(n4579), .Z(n6552) );
  OR U5922 ( .A(A[236]), .B(B[236]), .Z(n4579) );
  NANDN U5923 ( .A(n4581), .B(n6554), .Z(n6553) );
  NANDN U5924 ( .A(n4583), .B(n6555), .Z(n6554) );
  NANDN U5925 ( .A(n4603), .B(n6556), .Z(n6555) );
  NAND U5926 ( .A(n4631), .B(n4606), .Z(n6556) );
  AND U5927 ( .A(n6557), .B(n6558), .Z(n4606) );
  AND U5928 ( .A(n4628), .B(n4619), .Z(n6558) );
  OR U5929 ( .A(B[228]), .B(A[228]), .Z(n4628) );
  AND U5930 ( .A(n4614), .B(n4610), .Z(n6557) );
  NANDN U5931 ( .A(n4636), .B(n6559), .Z(n4631) );
  NAND U5932 ( .A(n6560), .B(n4637), .Z(n6559) );
  OR U5933 ( .A(B[227]), .B(A[227]), .Z(n4637) );
  NANDN U5934 ( .A(n4639), .B(n6561), .Z(n6560) );
  NANDN U5935 ( .A(n4640), .B(n6562), .Z(n6561) );
  NANDN U5936 ( .A(n4643), .B(n6563), .Z(n6562) );
  NAND U5937 ( .A(n4646), .B(n4648), .Z(n6563) );
  AND U5938 ( .A(A[224]), .B(B[224]), .Z(n4648) );
  OR U5939 ( .A(B[225]), .B(A[225]), .Z(n4646) );
  AND U5940 ( .A(B[225]), .B(A[225]), .Z(n4643) );
  NOR U5941 ( .A(B[226]), .B(A[226]), .Z(n4640) );
  AND U5942 ( .A(B[226]), .B(A[226]), .Z(n4639) );
  AND U5943 ( .A(B[227]), .B(A[227]), .Z(n4636) );
  NANDN U5944 ( .A(n4609), .B(n6564), .Z(n4603) );
  NAND U5945 ( .A(n6565), .B(n4610), .Z(n6564) );
  OR U5946 ( .A(B[231]), .B(A[231]), .Z(n4610) );
  NANDN U5947 ( .A(n4612), .B(n6566), .Z(n6565) );
  NAND U5948 ( .A(n6567), .B(n4614), .Z(n6566) );
  OR U5949 ( .A(B[230]), .B(A[230]), .Z(n4614) );
  NANDN U5950 ( .A(n4616), .B(n6568), .Z(n6567) );
  NAND U5951 ( .A(n4619), .B(n4626), .Z(n6568) );
  AND U5952 ( .A(B[228]), .B(A[228]), .Z(n4626) );
  OR U5953 ( .A(B[229]), .B(A[229]), .Z(n4619) );
  AND U5954 ( .A(B[229]), .B(A[229]), .Z(n4616) );
  AND U5955 ( .A(B[230]), .B(A[230]), .Z(n4612) );
  AND U5956 ( .A(B[231]), .B(A[231]), .Z(n4609) );
  NAND U5957 ( .A(n6569), .B(n6570), .Z(n4583) );
  AND U5958 ( .A(n4601), .B(n4597), .Z(n6570) );
  OR U5959 ( .A(B[232]), .B(A[232]), .Z(n4601) );
  AND U5960 ( .A(n4592), .B(n4588), .Z(n6569) );
  NANDN U5961 ( .A(n4587), .B(n6571), .Z(n4581) );
  NAND U5962 ( .A(n6572), .B(n4588), .Z(n6571) );
  OR U5963 ( .A(B[235]), .B(A[235]), .Z(n4588) );
  NANDN U5964 ( .A(n4590), .B(n6573), .Z(n6572) );
  NAND U5965 ( .A(n6574), .B(n4592), .Z(n6573) );
  OR U5966 ( .A(B[234]), .B(A[234]), .Z(n4592) );
  NANDN U5967 ( .A(n4594), .B(n6575), .Z(n6574) );
  NAND U5968 ( .A(n4597), .B(n4599), .Z(n6575) );
  AND U5969 ( .A(B[232]), .B(A[232]), .Z(n4599) );
  OR U5970 ( .A(B[233]), .B(A[233]), .Z(n4597) );
  AND U5971 ( .A(B[233]), .B(A[233]), .Z(n4594) );
  AND U5972 ( .A(B[234]), .B(A[234]), .Z(n4590) );
  AND U5973 ( .A(B[235]), .B(A[235]), .Z(n4587) );
  NOR U5974 ( .A(B[237]), .B(A[237]), .Z(n4573) );
  AND U5975 ( .A(B[237]), .B(A[237]), .Z(n4571) );
  NOR U5976 ( .A(B[238]), .B(A[238]), .Z(n4568) );
  AND U5977 ( .A(B[238]), .B(A[238]), .Z(n4567) );
  NOR U5978 ( .A(B[239]), .B(A[239]), .Z(n4564) );
  NOR U5979 ( .A(n4534), .B(n4485), .Z(n6019) );
  NAND U5980 ( .A(n6576), .B(n6577), .Z(n4534) );
  AND U5981 ( .A(n4552), .B(n4548), .Z(n6577) );
  OR U5982 ( .A(B[240]), .B(A[240]), .Z(n4552) );
  ANDN U5983 ( .B(n4539), .A(n4542), .Z(n6576) );
  ANDN U5984 ( .B(n6578), .A(n4478), .Z(n6017) );
  AND U5985 ( .A(B[252]), .B(A[252]), .Z(n4478) );
  NAND U5986 ( .A(n6579), .B(n4481), .Z(n6578) );
  OR U5987 ( .A(A[252]), .B(B[252]), .Z(n4481) );
  NANDN U5988 ( .A(n4483), .B(n6580), .Z(n6579) );
  NANDN U5989 ( .A(n4485), .B(n6581), .Z(n6580) );
  NANDN U5990 ( .A(n4510), .B(n6582), .Z(n6581) );
  NAND U5991 ( .A(n4533), .B(n4513), .Z(n6582) );
  AND U5992 ( .A(n6583), .B(n6584), .Z(n4513) );
  AND U5993 ( .A(n4530), .B(n4526), .Z(n6584) );
  OR U5994 ( .A(B[244]), .B(A[244]), .Z(n4530) );
  AND U5995 ( .A(n4521), .B(n4517), .Z(n6583) );
  NANDN U5996 ( .A(n4538), .B(n6585), .Z(n4533) );
  NAND U5997 ( .A(n6586), .B(n4539), .Z(n6585) );
  OR U5998 ( .A(B[243]), .B(A[243]), .Z(n4539) );
  NANDN U5999 ( .A(n4541), .B(n6587), .Z(n6586) );
  NANDN U6000 ( .A(n4542), .B(n6588), .Z(n6587) );
  NANDN U6001 ( .A(n4545), .B(n6589), .Z(n6588) );
  NAND U6002 ( .A(n4548), .B(n4550), .Z(n6589) );
  AND U6003 ( .A(A[240]), .B(B[240]), .Z(n4550) );
  OR U6004 ( .A(B[241]), .B(A[241]), .Z(n4548) );
  AND U6005 ( .A(B[241]), .B(A[241]), .Z(n4545) );
  NOR U6006 ( .A(B[242]), .B(A[242]), .Z(n4542) );
  AND U6007 ( .A(B[242]), .B(A[242]), .Z(n4541) );
  AND U6008 ( .A(B[243]), .B(A[243]), .Z(n4538) );
  NANDN U6009 ( .A(n4516), .B(n6590), .Z(n4510) );
  NAND U6010 ( .A(n6591), .B(n4517), .Z(n6590) );
  OR U6011 ( .A(B[247]), .B(A[247]), .Z(n4517) );
  NANDN U6012 ( .A(n4519), .B(n6592), .Z(n6591) );
  NAND U6013 ( .A(n6593), .B(n4521), .Z(n6592) );
  OR U6014 ( .A(B[246]), .B(A[246]), .Z(n4521) );
  NANDN U6015 ( .A(n4523), .B(n6594), .Z(n6593) );
  NAND U6016 ( .A(n4526), .B(n4528), .Z(n6594) );
  AND U6017 ( .A(B[244]), .B(A[244]), .Z(n4528) );
  OR U6018 ( .A(B[245]), .B(A[245]), .Z(n4526) );
  AND U6019 ( .A(B[245]), .B(A[245]), .Z(n4523) );
  AND U6020 ( .A(B[246]), .B(A[246]), .Z(n4519) );
  AND U6021 ( .A(B[247]), .B(A[247]), .Z(n4516) );
  NAND U6022 ( .A(n6595), .B(n6596), .Z(n4485) );
  AND U6023 ( .A(n4508), .B(n4499), .Z(n6596) );
  OR U6024 ( .A(B[248]), .B(A[248]), .Z(n4508) );
  AND U6025 ( .A(n4494), .B(n4490), .Z(n6595) );
  NANDN U6026 ( .A(n4489), .B(n6597), .Z(n4483) );
  NAND U6027 ( .A(n6598), .B(n4490), .Z(n6597) );
  OR U6028 ( .A(B[251]), .B(A[251]), .Z(n4490) );
  NANDN U6029 ( .A(n4492), .B(n6599), .Z(n6598) );
  NAND U6030 ( .A(n6600), .B(n4494), .Z(n6599) );
  OR U6031 ( .A(B[250]), .B(A[250]), .Z(n4494) );
  NANDN U6032 ( .A(n4496), .B(n6601), .Z(n6600) );
  NAND U6033 ( .A(n4499), .B(n4506), .Z(n6601) );
  AND U6034 ( .A(B[248]), .B(A[248]), .Z(n4506) );
  OR U6035 ( .A(B[249]), .B(A[249]), .Z(n4499) );
  AND U6036 ( .A(B[249]), .B(A[249]), .Z(n4496) );
  AND U6037 ( .A(B[250]), .B(A[250]), .Z(n4492) );
  AND U6038 ( .A(B[251]), .B(A[251]), .Z(n4489) );
  NOR U6039 ( .A(B[253]), .B(A[253]), .Z(n4475) );
  AND U6040 ( .A(B[253]), .B(A[253]), .Z(n4473) );
  NOR U6041 ( .A(B[254]), .B(A[254]), .Z(n4470) );
  AND U6042 ( .A(B[254]), .B(A[254]), .Z(n4469) );
  NOR U6043 ( .A(B[255]), .B(A[255]), .Z(n4466) );
  NOR U6044 ( .A(n4369), .B(n5903), .Z(n5986) );
  NAND U6045 ( .A(n6602), .B(n6603), .Z(n5903) );
  AND U6046 ( .A(n6604), .B(n6605), .Z(n6603) );
  AND U6047 ( .A(n4096), .B(n4091), .Z(n6605) );
  OR U6048 ( .A(A[317]), .B(B[317]), .Z(n4091) );
  OR U6049 ( .A(A[316]), .B(B[316]), .Z(n4096) );
  AND U6050 ( .A(n4086), .B(n4082), .Z(n6604) );
  OR U6051 ( .A(B[319]), .B(A[319]), .Z(n4082) );
  OR U6052 ( .A(A[318]), .B(B[318]), .Z(n4086) );
  ANDN U6053 ( .B(n6606), .A(n4122), .Z(n6602) );
  NAND U6054 ( .A(n6607), .B(n6608), .Z(n4122) );
  AND U6055 ( .A(n4145), .B(n4136), .Z(n6608) );
  OR U6056 ( .A(A[309]), .B(B[309]), .Z(n4136) );
  OR U6057 ( .A(A[308]), .B(B[308]), .Z(n4145) );
  AND U6058 ( .A(n4131), .B(n4127), .Z(n6607) );
  OR U6059 ( .A(B[311]), .B(A[311]), .Z(n4127) );
  OR U6060 ( .A(A[310]), .B(B[310]), .Z(n4131) );
  NOR U6061 ( .A(n4149), .B(n4100), .Z(n6606) );
  NAND U6062 ( .A(n6609), .B(n6610), .Z(n4100) );
  AND U6063 ( .A(n4118), .B(n4114), .Z(n6610) );
  OR U6064 ( .A(A[313]), .B(B[313]), .Z(n4114) );
  OR U6065 ( .A(A[312]), .B(B[312]), .Z(n4118) );
  AND U6066 ( .A(n4109), .B(n4105), .Z(n6609) );
  OR U6067 ( .A(B[315]), .B(A[315]), .Z(n4105) );
  OR U6068 ( .A(A[314]), .B(B[314]), .Z(n4109) );
  NAND U6069 ( .A(n6611), .B(n6612), .Z(n4149) );
  AND U6070 ( .A(n4167), .B(n4163), .Z(n6612) );
  OR U6071 ( .A(A[305]), .B(B[305]), .Z(n4163) );
  OR U6072 ( .A(A[304]), .B(B[304]), .Z(n4167) );
  AND U6073 ( .A(n4158), .B(n4154), .Z(n6611) );
  OR U6074 ( .A(B[307]), .B(A[307]), .Z(n4154) );
  OR U6075 ( .A(A[306]), .B(B[306]), .Z(n4158) );
  NAND U6076 ( .A(n6613), .B(n6614), .Z(n4369) );
  AND U6077 ( .A(n6615), .B(n6616), .Z(n6614) );
  AND U6078 ( .A(n4393), .B(n4383), .Z(n6616) );
  OR U6079 ( .A(A[269]), .B(B[269]), .Z(n4383) );
  OR U6080 ( .A(A[268]), .B(B[268]), .Z(n4393) );
  AND U6081 ( .A(n4378), .B(n4374), .Z(n6615) );
  OR U6082 ( .A(B[271]), .B(A[271]), .Z(n4374) );
  OR U6083 ( .A(A[270]), .B(B[270]), .Z(n4378) );
  ANDN U6084 ( .B(n6617), .A(n4441), .Z(n6613) );
  NAND U6085 ( .A(n6618), .B(n6619), .Z(n4441) );
  AND U6086 ( .A(n4462), .B(n4458), .Z(n6619) );
  OR U6087 ( .A(A[257]), .B(B[257]), .Z(n4458) );
  OR U6088 ( .A(A[256]), .B(B[256]), .Z(n4462) );
  AND U6089 ( .A(n4453), .B(n4449), .Z(n6618) );
  OR U6090 ( .A(B[259]), .B(A[259]), .Z(n4449) );
  OR U6091 ( .A(A[258]), .B(B[258]), .Z(n4453) );
  NOR U6092 ( .A(n4419), .B(n4397), .Z(n6617) );
  NAND U6093 ( .A(n6620), .B(n6621), .Z(n4397) );
  AND U6094 ( .A(n4415), .B(n4411), .Z(n6621) );
  OR U6095 ( .A(A[265]), .B(B[265]), .Z(n4411) );
  OR U6096 ( .A(A[264]), .B(B[264]), .Z(n4415) );
  AND U6097 ( .A(n4406), .B(n4402), .Z(n6620) );
  OR U6098 ( .A(B[267]), .B(A[267]), .Z(n4402) );
  OR U6099 ( .A(A[266]), .B(B[266]), .Z(n4406) );
  NAND U6100 ( .A(n6622), .B(n6623), .Z(n4419) );
  AND U6101 ( .A(n4437), .B(n4433), .Z(n6623) );
  OR U6102 ( .A(A[261]), .B(B[261]), .Z(n4433) );
  OR U6103 ( .A(A[260]), .B(B[260]), .Z(n4437) );
  AND U6104 ( .A(n4428), .B(n4424), .Z(n6622) );
  OR U6105 ( .A(B[263]), .B(A[263]), .Z(n4424) );
  OR U6106 ( .A(A[262]), .B(B[262]), .Z(n4428) );
  NAND U6107 ( .A(n6624), .B(n6625), .Z(n3692) );
  NOR U6108 ( .A(n3886), .B(n3790), .Z(n6625) );
  NOR U6109 ( .A(n3983), .B(n6626), .Z(n6624) );
  NAND U6110 ( .A(n6627), .B(n6628), .Z(n3983) );
  AND U6111 ( .A(n6629), .B(n6630), .Z(n6628) );
  AND U6112 ( .A(n4001), .B(n3996), .Z(n6630) );
  AND U6113 ( .A(n3991), .B(n3987), .Z(n6629) );
  ANDN U6114 ( .B(n6631), .A(n4050), .Z(n6627) );
  NAND U6115 ( .A(n6632), .B(n6633), .Z(n4050) );
  AND U6116 ( .A(n4067), .B(n4063), .Z(n6633) );
  OR U6117 ( .A(A[320]), .B(B[320]), .Z(n4067) );
  AND U6118 ( .A(n4058), .B(n4054), .Z(n6632) );
  NOR U6119 ( .A(n4028), .B(n4005), .Z(n6631) );
  NAND U6120 ( .A(n6634), .B(n6635), .Z(n3690) );
  NAND U6121 ( .A(n6636), .B(n3697), .Z(n6635) );
  NANDN U6122 ( .A(n3699), .B(n6637), .Z(n6636) );
  NAND U6123 ( .A(n6638), .B(n3701), .Z(n6637) );
  NANDN U6124 ( .A(n3703), .B(n6639), .Z(n6638) );
  NAND U6125 ( .A(n6640), .B(n3706), .Z(n6639) );
  NANDN U6126 ( .A(n3708), .B(n6641), .Z(n6640) );
  NAND U6127 ( .A(n6642), .B(n3711), .Z(n6641) );
  NANDN U6128 ( .A(n3713), .B(n6643), .Z(n6642) );
  NANDN U6129 ( .A(n3715), .B(n6644), .Z(n6643) );
  NANDN U6130 ( .A(n3739), .B(n6645), .Z(n6644) );
  NANDN U6131 ( .A(n3741), .B(n3762), .Z(n6645) );
  NANDN U6132 ( .A(n3767), .B(n6646), .Z(n3762) );
  NAND U6133 ( .A(n6647), .B(n3768), .Z(n6646) );
  NANDN U6134 ( .A(n3770), .B(n6648), .Z(n6647) );
  NAND U6135 ( .A(n6649), .B(n3772), .Z(n6648) );
  NANDN U6136 ( .A(n3774), .B(n6650), .Z(n6649) );
  NAND U6137 ( .A(n3777), .B(n3784), .Z(n6650) );
  AND U6138 ( .A(A[368]), .B(B[368]), .Z(n3784) );
  AND U6139 ( .A(A[369]), .B(B[369]), .Z(n3774) );
  AND U6140 ( .A(A[370]), .B(B[370]), .Z(n3770) );
  AND U6141 ( .A(B[371]), .B(A[371]), .Z(n3767) );
  NANDN U6142 ( .A(n3745), .B(n6651), .Z(n3739) );
  NAND U6143 ( .A(n6652), .B(n3746), .Z(n6651) );
  NANDN U6144 ( .A(n3748), .B(n6653), .Z(n6652) );
  NAND U6145 ( .A(n6654), .B(n3750), .Z(n6653) );
  NANDN U6146 ( .A(n3752), .B(n6655), .Z(n6654) );
  NAND U6147 ( .A(n3755), .B(n3757), .Z(n6655) );
  AND U6148 ( .A(A[372]), .B(B[372]), .Z(n3757) );
  AND U6149 ( .A(A[373]), .B(B[373]), .Z(n3752) );
  AND U6150 ( .A(A[374]), .B(B[374]), .Z(n3748) );
  AND U6151 ( .A(B[375]), .B(A[375]), .Z(n3745) );
  NANDN U6152 ( .A(n3723), .B(n6656), .Z(n3713) );
  NAND U6153 ( .A(n6657), .B(n3724), .Z(n6656) );
  NANDN U6154 ( .A(n3726), .B(n6658), .Z(n6657) );
  NAND U6155 ( .A(n6659), .B(n3728), .Z(n6658) );
  NANDN U6156 ( .A(n3730), .B(n6660), .Z(n6659) );
  NAND U6157 ( .A(n3733), .B(n3735), .Z(n6660) );
  AND U6158 ( .A(A[376]), .B(B[376]), .Z(n3735) );
  AND U6159 ( .A(A[377]), .B(B[377]), .Z(n3730) );
  AND U6160 ( .A(A[378]), .B(B[378]), .Z(n3726) );
  AND U6161 ( .A(B[379]), .B(A[379]), .Z(n3723) );
  AND U6162 ( .A(A[380]), .B(B[380]), .Z(n3708) );
  AND U6163 ( .A(A[381]), .B(B[381]), .Z(n3703) );
  AND U6164 ( .A(A[382]), .B(B[382]), .Z(n3699) );
  ANDN U6165 ( .B(n6661), .A(n3696), .Z(n6634) );
  AND U6166 ( .A(B[383]), .B(A[383]), .Z(n3696) );
  NANDN U6167 ( .A(n6626), .B(n6662), .Z(n6661) );
  NANDN U6168 ( .A(n3788), .B(n6663), .Z(n6662) );
  NANDN U6169 ( .A(n3790), .B(n6664), .Z(n6663) );
  NANDN U6170 ( .A(n3884), .B(n6665), .Z(n6664) );
  NANDN U6171 ( .A(n3886), .B(n3982), .Z(n6665) );
  NANDN U6172 ( .A(n3986), .B(n6666), .Z(n3982) );
  NAND U6173 ( .A(n6667), .B(n3987), .Z(n6666) );
  OR U6174 ( .A(B[335]), .B(A[335]), .Z(n3987) );
  NANDN U6175 ( .A(n3989), .B(n6668), .Z(n6667) );
  NAND U6176 ( .A(n6669), .B(n3991), .Z(n6668) );
  OR U6177 ( .A(A[334]), .B(B[334]), .Z(n3991) );
  NANDN U6178 ( .A(n3993), .B(n6670), .Z(n6669) );
  NAND U6179 ( .A(n6671), .B(n3996), .Z(n6670) );
  OR U6180 ( .A(A[333]), .B(B[333]), .Z(n3996) );
  NANDN U6181 ( .A(n3998), .B(n6672), .Z(n6671) );
  NAND U6182 ( .A(n6673), .B(n4001), .Z(n6672) );
  OR U6183 ( .A(A[332]), .B(B[332]), .Z(n4001) );
  NANDN U6184 ( .A(n4003), .B(n6674), .Z(n6673) );
  NANDN U6185 ( .A(n4005), .B(n6675), .Z(n6674) );
  NANDN U6186 ( .A(n4026), .B(n6676), .Z(n6675) );
  NANDN U6187 ( .A(n4028), .B(n4049), .Z(n6676) );
  NANDN U6188 ( .A(n4053), .B(n6677), .Z(n4049) );
  NAND U6189 ( .A(n6678), .B(n4054), .Z(n6677) );
  OR U6190 ( .A(B[323]), .B(A[323]), .Z(n4054) );
  NANDN U6191 ( .A(n4056), .B(n6679), .Z(n6678) );
  NAND U6192 ( .A(n6680), .B(n4058), .Z(n6679) );
  OR U6193 ( .A(A[322]), .B(B[322]), .Z(n4058) );
  NANDN U6194 ( .A(n4060), .B(n6681), .Z(n6680) );
  NAND U6195 ( .A(n4063), .B(n4065), .Z(n6681) );
  AND U6196 ( .A(A[320]), .B(B[320]), .Z(n4065) );
  OR U6197 ( .A(A[321]), .B(B[321]), .Z(n4063) );
  AND U6198 ( .A(A[321]), .B(B[321]), .Z(n4060) );
  AND U6199 ( .A(A[322]), .B(B[322]), .Z(n4056) );
  AND U6200 ( .A(B[323]), .B(A[323]), .Z(n4053) );
  NAND U6201 ( .A(n6682), .B(n6683), .Z(n4028) );
  AND U6202 ( .A(n4046), .B(n4042), .Z(n6683) );
  OR U6203 ( .A(A[324]), .B(B[324]), .Z(n4046) );
  AND U6204 ( .A(n4037), .B(n4033), .Z(n6682) );
  NANDN U6205 ( .A(n4032), .B(n6684), .Z(n4026) );
  NAND U6206 ( .A(n6685), .B(n4033), .Z(n6684) );
  OR U6207 ( .A(B[327]), .B(A[327]), .Z(n4033) );
  NANDN U6208 ( .A(n4035), .B(n6686), .Z(n6685) );
  NAND U6209 ( .A(n6687), .B(n4037), .Z(n6686) );
  OR U6210 ( .A(A[326]), .B(B[326]), .Z(n4037) );
  NANDN U6211 ( .A(n4039), .B(n6688), .Z(n6687) );
  NAND U6212 ( .A(n4042), .B(n4044), .Z(n6688) );
  AND U6213 ( .A(A[324]), .B(B[324]), .Z(n4044) );
  OR U6214 ( .A(A[325]), .B(B[325]), .Z(n4042) );
  AND U6215 ( .A(A[325]), .B(B[325]), .Z(n4039) );
  AND U6216 ( .A(A[326]), .B(B[326]), .Z(n4035) );
  AND U6217 ( .A(B[327]), .B(A[327]), .Z(n4032) );
  NAND U6218 ( .A(n6689), .B(n6690), .Z(n4005) );
  AND U6219 ( .A(n4024), .B(n4019), .Z(n6690) );
  OR U6220 ( .A(A[328]), .B(B[328]), .Z(n4024) );
  AND U6221 ( .A(n4014), .B(n4010), .Z(n6689) );
  NANDN U6222 ( .A(n4009), .B(n6691), .Z(n4003) );
  NAND U6223 ( .A(n6692), .B(n4010), .Z(n6691) );
  OR U6224 ( .A(B[331]), .B(A[331]), .Z(n4010) );
  NANDN U6225 ( .A(n4012), .B(n6693), .Z(n6692) );
  NAND U6226 ( .A(n6694), .B(n4014), .Z(n6693) );
  OR U6227 ( .A(A[330]), .B(B[330]), .Z(n4014) );
  NANDN U6228 ( .A(n4016), .B(n6695), .Z(n6694) );
  NAND U6229 ( .A(n4019), .B(n4022), .Z(n6695) );
  AND U6230 ( .A(A[328]), .B(B[328]), .Z(n4022) );
  OR U6231 ( .A(A[329]), .B(B[329]), .Z(n4019) );
  AND U6232 ( .A(A[329]), .B(B[329]), .Z(n4016) );
  AND U6233 ( .A(A[330]), .B(B[330]), .Z(n4012) );
  AND U6234 ( .A(B[331]), .B(A[331]), .Z(n4009) );
  AND U6235 ( .A(A[332]), .B(B[332]), .Z(n3998) );
  AND U6236 ( .A(A[333]), .B(B[333]), .Z(n3993) );
  AND U6237 ( .A(A[334]), .B(B[334]), .Z(n3989) );
  AND U6238 ( .A(B[335]), .B(A[335]), .Z(n3986) );
  NAND U6239 ( .A(n6696), .B(n6697), .Z(n3886) );
  AND U6240 ( .A(n6698), .B(n6699), .Z(n6697) );
  AND U6241 ( .A(n3910), .B(n3900), .Z(n6699) );
  AND U6242 ( .A(n3895), .B(n3891), .Z(n6698) );
  ANDN U6243 ( .B(n6700), .A(n3958), .Z(n6696) );
  NAND U6244 ( .A(n6701), .B(n6702), .Z(n3958) );
  AND U6245 ( .A(n3979), .B(n3975), .Z(n6702) );
  OR U6246 ( .A(A[336]), .B(B[336]), .Z(n3979) );
  AND U6247 ( .A(n3970), .B(n3966), .Z(n6701) );
  NOR U6248 ( .A(n3936), .B(n3914), .Z(n6700) );
  NANDN U6249 ( .A(n3890), .B(n6703), .Z(n3884) );
  NAND U6250 ( .A(n6704), .B(n3891), .Z(n6703) );
  OR U6251 ( .A(B[351]), .B(A[351]), .Z(n3891) );
  NANDN U6252 ( .A(n3893), .B(n6705), .Z(n6704) );
  NAND U6253 ( .A(n6706), .B(n3895), .Z(n6705) );
  OR U6254 ( .A(A[350]), .B(B[350]), .Z(n3895) );
  NANDN U6255 ( .A(n3897), .B(n6707), .Z(n6706) );
  NAND U6256 ( .A(n6708), .B(n3900), .Z(n6707) );
  OR U6257 ( .A(A[349]), .B(B[349]), .Z(n3900) );
  NANDN U6258 ( .A(n3907), .B(n6709), .Z(n6708) );
  NAND U6259 ( .A(n6710), .B(n3910), .Z(n6709) );
  OR U6260 ( .A(A[348]), .B(B[348]), .Z(n3910) );
  NANDN U6261 ( .A(n3912), .B(n6711), .Z(n6710) );
  NANDN U6262 ( .A(n3914), .B(n6712), .Z(n6711) );
  NANDN U6263 ( .A(n3934), .B(n6713), .Z(n6712) );
  NANDN U6264 ( .A(n3936), .B(n3957), .Z(n6713) );
  NANDN U6265 ( .A(n3965), .B(n6714), .Z(n3957) );
  NAND U6266 ( .A(n6715), .B(n3966), .Z(n6714) );
  OR U6267 ( .A(B[339]), .B(A[339]), .Z(n3966) );
  NANDN U6268 ( .A(n3968), .B(n6716), .Z(n6715) );
  NAND U6269 ( .A(n6717), .B(n3970), .Z(n6716) );
  OR U6270 ( .A(A[338]), .B(B[338]), .Z(n3970) );
  NANDN U6271 ( .A(n3972), .B(n6718), .Z(n6717) );
  NAND U6272 ( .A(n3975), .B(n3977), .Z(n6718) );
  AND U6273 ( .A(A[336]), .B(B[336]), .Z(n3977) );
  OR U6274 ( .A(A[337]), .B(B[337]), .Z(n3975) );
  AND U6275 ( .A(A[337]), .B(B[337]), .Z(n3972) );
  AND U6276 ( .A(A[338]), .B(B[338]), .Z(n3968) );
  AND U6277 ( .A(B[339]), .B(A[339]), .Z(n3965) );
  NAND U6278 ( .A(n6719), .B(n6720), .Z(n3936) );
  AND U6279 ( .A(n3954), .B(n3950), .Z(n6720) );
  OR U6280 ( .A(A[340]), .B(B[340]), .Z(n3954) );
  AND U6281 ( .A(n3945), .B(n3941), .Z(n6719) );
  NANDN U6282 ( .A(n3940), .B(n6721), .Z(n3934) );
  NAND U6283 ( .A(n6722), .B(n3941), .Z(n6721) );
  OR U6284 ( .A(B[343]), .B(A[343]), .Z(n3941) );
  NANDN U6285 ( .A(n3943), .B(n6723), .Z(n6722) );
  NAND U6286 ( .A(n6724), .B(n3945), .Z(n6723) );
  OR U6287 ( .A(A[342]), .B(B[342]), .Z(n3945) );
  NANDN U6288 ( .A(n3947), .B(n6725), .Z(n6724) );
  NAND U6289 ( .A(n3950), .B(n3952), .Z(n6725) );
  AND U6290 ( .A(A[340]), .B(B[340]), .Z(n3952) );
  OR U6291 ( .A(A[341]), .B(B[341]), .Z(n3950) );
  AND U6292 ( .A(A[341]), .B(B[341]), .Z(n3947) );
  AND U6293 ( .A(A[342]), .B(B[342]), .Z(n3943) );
  AND U6294 ( .A(B[343]), .B(A[343]), .Z(n3940) );
  NAND U6295 ( .A(n6726), .B(n6727), .Z(n3914) );
  AND U6296 ( .A(n3932), .B(n3928), .Z(n6727) );
  OR U6297 ( .A(A[344]), .B(B[344]), .Z(n3932) );
  AND U6298 ( .A(n3923), .B(n3919), .Z(n6726) );
  NANDN U6299 ( .A(n3918), .B(n6728), .Z(n3912) );
  NAND U6300 ( .A(n6729), .B(n3919), .Z(n6728) );
  OR U6301 ( .A(B[347]), .B(A[347]), .Z(n3919) );
  NANDN U6302 ( .A(n3921), .B(n6730), .Z(n6729) );
  NAND U6303 ( .A(n6731), .B(n3923), .Z(n6730) );
  OR U6304 ( .A(A[346]), .B(B[346]), .Z(n3923) );
  NANDN U6305 ( .A(n3925), .B(n6732), .Z(n6731) );
  NAND U6306 ( .A(n3928), .B(n3930), .Z(n6732) );
  AND U6307 ( .A(A[344]), .B(B[344]), .Z(n3930) );
  OR U6308 ( .A(A[345]), .B(B[345]), .Z(n3928) );
  AND U6309 ( .A(A[345]), .B(B[345]), .Z(n3925) );
  AND U6310 ( .A(A[346]), .B(B[346]), .Z(n3921) );
  AND U6311 ( .A(B[347]), .B(A[347]), .Z(n3918) );
  AND U6312 ( .A(A[348]), .B(B[348]), .Z(n3907) );
  AND U6313 ( .A(A[349]), .B(B[349]), .Z(n3897) );
  AND U6314 ( .A(A[350]), .B(B[350]), .Z(n3893) );
  AND U6315 ( .A(B[351]), .B(A[351]), .Z(n3890) );
  NAND U6316 ( .A(n6733), .B(n6734), .Z(n3790) );
  AND U6317 ( .A(n6735), .B(n6736), .Z(n6734) );
  AND U6318 ( .A(n3809), .B(n3804), .Z(n6736) );
  AND U6319 ( .A(n3799), .B(n3795), .Z(n6735) );
  ANDN U6320 ( .B(n6737), .A(n3865), .Z(n6733) );
  NAND U6321 ( .A(n6738), .B(n6739), .Z(n3865) );
  AND U6322 ( .A(n3882), .B(n3878), .Z(n6739) );
  OR U6323 ( .A(A[352]), .B(B[352]), .Z(n3882) );
  AND U6324 ( .A(n3873), .B(n3869), .Z(n6738) );
  NOR U6325 ( .A(n3835), .B(n3813), .Z(n6737) );
  NANDN U6326 ( .A(n3794), .B(n6740), .Z(n3788) );
  NAND U6327 ( .A(n6741), .B(n3795), .Z(n6740) );
  OR U6328 ( .A(B[367]), .B(A[367]), .Z(n3795) );
  NANDN U6329 ( .A(n3797), .B(n6742), .Z(n6741) );
  NAND U6330 ( .A(n6743), .B(n3799), .Z(n6742) );
  OR U6331 ( .A(A[366]), .B(B[366]), .Z(n3799) );
  NANDN U6332 ( .A(n3801), .B(n6744), .Z(n6743) );
  NAND U6333 ( .A(n6745), .B(n3804), .Z(n6744) );
  OR U6334 ( .A(A[365]), .B(B[365]), .Z(n3804) );
  NANDN U6335 ( .A(n3806), .B(n6746), .Z(n6745) );
  NAND U6336 ( .A(n6747), .B(n3809), .Z(n6746) );
  OR U6337 ( .A(A[364]), .B(B[364]), .Z(n3809) );
  NANDN U6338 ( .A(n3811), .B(n6748), .Z(n6747) );
  NANDN U6339 ( .A(n3813), .B(n6749), .Z(n6748) );
  NANDN U6340 ( .A(n3833), .B(n6750), .Z(n6749) );
  NANDN U6341 ( .A(n3835), .B(n3864), .Z(n6750) );
  NANDN U6342 ( .A(n3868), .B(n6751), .Z(n3864) );
  NAND U6343 ( .A(n6752), .B(n3869), .Z(n6751) );
  OR U6344 ( .A(B[355]), .B(A[355]), .Z(n3869) );
  NANDN U6345 ( .A(n3871), .B(n6753), .Z(n6752) );
  NAND U6346 ( .A(n6754), .B(n3873), .Z(n6753) );
  OR U6347 ( .A(A[354]), .B(B[354]), .Z(n3873) );
  NANDN U6348 ( .A(n3875), .B(n6755), .Z(n6754) );
  NAND U6349 ( .A(n3878), .B(n3880), .Z(n6755) );
  AND U6350 ( .A(A[352]), .B(B[352]), .Z(n3880) );
  OR U6351 ( .A(A[353]), .B(B[353]), .Z(n3878) );
  AND U6352 ( .A(A[353]), .B(B[353]), .Z(n3875) );
  AND U6353 ( .A(A[354]), .B(B[354]), .Z(n3871) );
  AND U6354 ( .A(B[355]), .B(A[355]), .Z(n3868) );
  NAND U6355 ( .A(n6756), .B(n6757), .Z(n3835) );
  AND U6356 ( .A(n3861), .B(n3857), .Z(n6757) );
  OR U6357 ( .A(A[356]), .B(B[356]), .Z(n3861) );
  AND U6358 ( .A(n3852), .B(n3848), .Z(n6756) );
  NANDN U6359 ( .A(n3847), .B(n6758), .Z(n3833) );
  NAND U6360 ( .A(n6759), .B(n3848), .Z(n6758) );
  OR U6361 ( .A(B[359]), .B(A[359]), .Z(n3848) );
  NANDN U6362 ( .A(n3850), .B(n6760), .Z(n6759) );
  NAND U6363 ( .A(n6761), .B(n3852), .Z(n6760) );
  OR U6364 ( .A(A[358]), .B(B[358]), .Z(n3852) );
  NANDN U6365 ( .A(n3854), .B(n6762), .Z(n6761) );
  NAND U6366 ( .A(n3857), .B(n3859), .Z(n6762) );
  AND U6367 ( .A(A[356]), .B(B[356]), .Z(n3859) );
  OR U6368 ( .A(A[357]), .B(B[357]), .Z(n3857) );
  AND U6369 ( .A(A[357]), .B(B[357]), .Z(n3854) );
  AND U6370 ( .A(A[358]), .B(B[358]), .Z(n3850) );
  AND U6371 ( .A(B[359]), .B(A[359]), .Z(n3847) );
  NAND U6372 ( .A(n6763), .B(n6764), .Z(n3813) );
  AND U6373 ( .A(n3831), .B(n3827), .Z(n6764) );
  OR U6374 ( .A(A[360]), .B(B[360]), .Z(n3831) );
  AND U6375 ( .A(n3822), .B(n3818), .Z(n6763) );
  NANDN U6376 ( .A(n3817), .B(n6765), .Z(n3811) );
  NAND U6377 ( .A(n6766), .B(n3818), .Z(n6765) );
  OR U6378 ( .A(B[363]), .B(A[363]), .Z(n3818) );
  NANDN U6379 ( .A(n3820), .B(n6767), .Z(n6766) );
  NAND U6380 ( .A(n6768), .B(n3822), .Z(n6767) );
  OR U6381 ( .A(A[362]), .B(B[362]), .Z(n3822) );
  NANDN U6382 ( .A(n3824), .B(n6769), .Z(n6768) );
  NAND U6383 ( .A(n3827), .B(n3829), .Z(n6769) );
  AND U6384 ( .A(A[360]), .B(B[360]), .Z(n3829) );
  OR U6385 ( .A(A[361]), .B(B[361]), .Z(n3827) );
  AND U6386 ( .A(A[361]), .B(B[361]), .Z(n3824) );
  AND U6387 ( .A(A[362]), .B(B[362]), .Z(n3820) );
  AND U6388 ( .A(B[363]), .B(A[363]), .Z(n3817) );
  AND U6389 ( .A(A[364]), .B(B[364]), .Z(n3806) );
  AND U6390 ( .A(A[365]), .B(B[365]), .Z(n3801) );
  AND U6391 ( .A(A[366]), .B(B[366]), .Z(n3797) );
  AND U6392 ( .A(B[367]), .B(A[367]), .Z(n3794) );
  NAND U6393 ( .A(n6770), .B(n6771), .Z(n6626) );
  AND U6394 ( .A(n6772), .B(n6773), .Z(n6771) );
  AND U6395 ( .A(n3711), .B(n3706), .Z(n6773) );
  OR U6396 ( .A(A[381]), .B(B[381]), .Z(n3706) );
  OR U6397 ( .A(A[380]), .B(B[380]), .Z(n3711) );
  AND U6398 ( .A(n3701), .B(n3697), .Z(n6772) );
  OR U6399 ( .A(B[383]), .B(A[383]), .Z(n3697) );
  OR U6400 ( .A(A[382]), .B(B[382]), .Z(n3701) );
  ANDN U6401 ( .B(n6774), .A(n3741), .Z(n6770) );
  NAND U6402 ( .A(n6775), .B(n6776), .Z(n3741) );
  AND U6403 ( .A(n3759), .B(n3755), .Z(n6776) );
  OR U6404 ( .A(A[373]), .B(B[373]), .Z(n3755) );
  OR U6405 ( .A(A[372]), .B(B[372]), .Z(n3759) );
  AND U6406 ( .A(n3750), .B(n3746), .Z(n6775) );
  OR U6407 ( .A(B[375]), .B(A[375]), .Z(n3746) );
  OR U6408 ( .A(A[374]), .B(B[374]), .Z(n3750) );
  NOR U6409 ( .A(n3763), .B(n3715), .Z(n6774) );
  NAND U6410 ( .A(n6777), .B(n6778), .Z(n3715) );
  AND U6411 ( .A(n3737), .B(n3733), .Z(n6778) );
  OR U6412 ( .A(A[377]), .B(B[377]), .Z(n3733) );
  OR U6413 ( .A(A[376]), .B(B[376]), .Z(n3737) );
  AND U6414 ( .A(n3728), .B(n3724), .Z(n6777) );
  OR U6415 ( .A(B[379]), .B(A[379]), .Z(n3724) );
  OR U6416 ( .A(A[378]), .B(B[378]), .Z(n3728) );
  NAND U6417 ( .A(n6779), .B(n6780), .Z(n3763) );
  AND U6418 ( .A(n3786), .B(n3777), .Z(n6780) );
  OR U6419 ( .A(A[369]), .B(B[369]), .Z(n3777) );
  OR U6420 ( .A(A[368]), .B(B[368]), .Z(n3786) );
  AND U6421 ( .A(n3772), .B(n3768), .Z(n6779) );
  OR U6422 ( .A(B[371]), .B(A[371]), .Z(n3768) );
  OR U6423 ( .A(A[370]), .B(B[370]), .Z(n3772) );
  NAND U6424 ( .A(n6781), .B(n6782), .Z(n3303) );
  ANDN U6425 ( .B(n3400), .A(n3497), .Z(n6782) );
  NOR U6426 ( .A(n3590), .B(n6783), .Z(n6781) );
  NAND U6427 ( .A(n6784), .B(n6785), .Z(n3590) );
  AND U6428 ( .A(n6786), .B(n6787), .Z(n6785) );
  AND U6429 ( .A(n3618), .B(n3613), .Z(n6787) );
  AND U6430 ( .A(n3608), .B(n3604), .Z(n6786) );
  ANDN U6431 ( .B(n6788), .A(n3671), .Z(n6784) );
  NAND U6432 ( .A(n6789), .B(n6790), .Z(n3671) );
  AND U6433 ( .A(n3688), .B(n3684), .Z(n6790) );
  OR U6434 ( .A(B[384]), .B(A[384]), .Z(n3688) );
  AND U6435 ( .A(n3679), .B(n3675), .Z(n6789) );
  ANDN U6436 ( .B(n3622), .A(n3644), .Z(n6788) );
  NAND U6437 ( .A(n6791), .B(n6792), .Z(n3301) );
  NAND U6438 ( .A(n6793), .B(n3308), .Z(n6792) );
  NANDN U6439 ( .A(n3310), .B(n6794), .Z(n6793) );
  NAND U6440 ( .A(n6795), .B(n3312), .Z(n6794) );
  NANDN U6441 ( .A(n3314), .B(n6796), .Z(n6795) );
  NAND U6442 ( .A(n6797), .B(n3317), .Z(n6796) );
  NANDN U6443 ( .A(n3319), .B(n6798), .Z(n6797) );
  NAND U6444 ( .A(n6799), .B(n3322), .Z(n6798) );
  NANDN U6445 ( .A(n3324), .B(n6800), .Z(n6799) );
  NANDN U6446 ( .A(n3326), .B(n6801), .Z(n6800) );
  NANDN U6447 ( .A(n3346), .B(n6802), .Z(n6801) );
  NANDN U6448 ( .A(n3348), .B(n3377), .Z(n6802) );
  NANDN U6449 ( .A(n3382), .B(n6803), .Z(n3377) );
  NAND U6450 ( .A(n6804), .B(n3383), .Z(n6803) );
  NANDN U6451 ( .A(n3385), .B(n6805), .Z(n6804) );
  NAND U6452 ( .A(n6806), .B(n3387), .Z(n6805) );
  NANDN U6453 ( .A(n3389), .B(n6807), .Z(n6806) );
  NAND U6454 ( .A(n3392), .B(n3394), .Z(n6807) );
  AND U6455 ( .A(A[432]), .B(B[432]), .Z(n3394) );
  AND U6456 ( .A(A[433]), .B(B[433]), .Z(n3389) );
  AND U6457 ( .A(A[434]), .B(B[434]), .Z(n3385) );
  AND U6458 ( .A(B[435]), .B(A[435]), .Z(n3382) );
  NANDN U6459 ( .A(n3360), .B(n6808), .Z(n3346) );
  NAND U6460 ( .A(n6809), .B(n3361), .Z(n6808) );
  NANDN U6461 ( .A(n3363), .B(n6810), .Z(n6809) );
  NAND U6462 ( .A(n6811), .B(n3365), .Z(n6810) );
  NANDN U6463 ( .A(n3367), .B(n6812), .Z(n6811) );
  NAND U6464 ( .A(n3370), .B(n3372), .Z(n6812) );
  AND U6465 ( .A(A[436]), .B(B[436]), .Z(n3372) );
  AND U6466 ( .A(A[437]), .B(B[437]), .Z(n3367) );
  AND U6467 ( .A(A[438]), .B(B[438]), .Z(n3363) );
  AND U6468 ( .A(B[439]), .B(A[439]), .Z(n3360) );
  NANDN U6469 ( .A(n3330), .B(n6813), .Z(n3324) );
  NAND U6470 ( .A(n6814), .B(n3331), .Z(n6813) );
  NANDN U6471 ( .A(n3333), .B(n6815), .Z(n6814) );
  NAND U6472 ( .A(n6816), .B(n3335), .Z(n6815) );
  NANDN U6473 ( .A(n3337), .B(n6817), .Z(n6816) );
  NAND U6474 ( .A(n3340), .B(n3342), .Z(n6817) );
  AND U6475 ( .A(A[440]), .B(B[440]), .Z(n3342) );
  AND U6476 ( .A(A[441]), .B(B[441]), .Z(n3337) );
  AND U6477 ( .A(A[442]), .B(B[442]), .Z(n3333) );
  AND U6478 ( .A(B[443]), .B(A[443]), .Z(n3330) );
  AND U6479 ( .A(A[444]), .B(B[444]), .Z(n3319) );
  AND U6480 ( .A(A[445]), .B(B[445]), .Z(n3314) );
  AND U6481 ( .A(A[446]), .B(B[446]), .Z(n3310) );
  ANDN U6482 ( .B(n6818), .A(n3307), .Z(n6791) );
  AND U6483 ( .A(B[447]), .B(A[447]), .Z(n3307) );
  NANDN U6484 ( .A(n6783), .B(n6819), .Z(n6818) );
  NANDN U6485 ( .A(n3398), .B(n6820), .Z(n6819) );
  NAND U6486 ( .A(n6821), .B(n3400), .Z(n6820) );
  AND U6487 ( .A(n6822), .B(n6823), .Z(n3400) );
  AND U6488 ( .A(n6824), .B(n6825), .Z(n6823) );
  AND U6489 ( .A(n3424), .B(n3414), .Z(n6825) );
  AND U6490 ( .A(n3409), .B(n3405), .Z(n6824) );
  ANDN U6491 ( .B(n6826), .A(n3472), .Z(n6822) );
  NAND U6492 ( .A(n6827), .B(n6828), .Z(n3472) );
  AND U6493 ( .A(n3493), .B(n3489), .Z(n6828) );
  OR U6494 ( .A(B[416]), .B(A[416]), .Z(n3493) );
  AND U6495 ( .A(n3484), .B(n3480), .Z(n6827) );
  ANDN U6496 ( .B(n3428), .A(n3450), .Z(n6826) );
  NANDN U6497 ( .A(n3495), .B(n6829), .Z(n6821) );
  NANDN U6498 ( .A(n3497), .B(n3589), .Z(n6829) );
  NANDN U6499 ( .A(n3603), .B(n6830), .Z(n3589) );
  NAND U6500 ( .A(n6831), .B(n3604), .Z(n6830) );
  OR U6501 ( .A(B[399]), .B(A[399]), .Z(n3604) );
  NANDN U6502 ( .A(n3606), .B(n6832), .Z(n6831) );
  NAND U6503 ( .A(n6833), .B(n3608), .Z(n6832) );
  OR U6504 ( .A(B[398]), .B(A[398]), .Z(n3608) );
  NANDN U6505 ( .A(n3610), .B(n6834), .Z(n6833) );
  NAND U6506 ( .A(n6835), .B(n3613), .Z(n6834) );
  OR U6507 ( .A(B[397]), .B(A[397]), .Z(n3613) );
  NANDN U6508 ( .A(n3615), .B(n6836), .Z(n6835) );
  NAND U6509 ( .A(n6837), .B(n3618), .Z(n6836) );
  OR U6510 ( .A(B[396]), .B(A[396]), .Z(n3618) );
  NANDN U6511 ( .A(n3620), .B(n6838), .Z(n6837) );
  NAND U6512 ( .A(n6839), .B(n3622), .Z(n6838) );
  AND U6513 ( .A(n6840), .B(n6841), .Z(n3622) );
  AND U6514 ( .A(n3640), .B(n3636), .Z(n6841) );
  OR U6515 ( .A(B[392]), .B(A[392]), .Z(n3640) );
  AND U6516 ( .A(n3631), .B(n3627), .Z(n6840) );
  NANDN U6517 ( .A(n3642), .B(n6842), .Z(n6839) );
  NANDN U6518 ( .A(n3644), .B(n3670), .Z(n6842) );
  NANDN U6519 ( .A(n3674), .B(n6843), .Z(n3670) );
  NAND U6520 ( .A(n6844), .B(n3675), .Z(n6843) );
  OR U6521 ( .A(B[387]), .B(A[387]), .Z(n3675) );
  NANDN U6522 ( .A(n3677), .B(n6845), .Z(n6844) );
  NAND U6523 ( .A(n6846), .B(n3679), .Z(n6845) );
  OR U6524 ( .A(B[386]), .B(A[386]), .Z(n3679) );
  NANDN U6525 ( .A(n3681), .B(n6847), .Z(n6846) );
  NAND U6526 ( .A(n3684), .B(n3686), .Z(n6847) );
  AND U6527 ( .A(B[384]), .B(A[384]), .Z(n3686) );
  OR U6528 ( .A(B[385]), .B(A[385]), .Z(n3684) );
  AND U6529 ( .A(B[385]), .B(A[385]), .Z(n3681) );
  AND U6530 ( .A(B[386]), .B(A[386]), .Z(n3677) );
  AND U6531 ( .A(B[387]), .B(A[387]), .Z(n3674) );
  NAND U6532 ( .A(n6848), .B(n6849), .Z(n3644) );
  AND U6533 ( .A(n3667), .B(n3658), .Z(n6849) );
  OR U6534 ( .A(B[388]), .B(A[388]), .Z(n3667) );
  AND U6535 ( .A(n3653), .B(n3649), .Z(n6848) );
  NANDN U6536 ( .A(n3648), .B(n6850), .Z(n3642) );
  NAND U6537 ( .A(n6851), .B(n3649), .Z(n6850) );
  OR U6538 ( .A(B[391]), .B(A[391]), .Z(n3649) );
  NANDN U6539 ( .A(n3651), .B(n6852), .Z(n6851) );
  NAND U6540 ( .A(n6853), .B(n3653), .Z(n6852) );
  OR U6541 ( .A(B[390]), .B(A[390]), .Z(n3653) );
  NANDN U6542 ( .A(n3655), .B(n6854), .Z(n6853) );
  NAND U6543 ( .A(n3658), .B(n3665), .Z(n6854) );
  AND U6544 ( .A(B[388]), .B(A[388]), .Z(n3665) );
  OR U6545 ( .A(B[389]), .B(A[389]), .Z(n3658) );
  AND U6546 ( .A(B[389]), .B(A[389]), .Z(n3655) );
  AND U6547 ( .A(B[390]), .B(A[390]), .Z(n3651) );
  AND U6548 ( .A(B[391]), .B(A[391]), .Z(n3648) );
  NANDN U6549 ( .A(n3626), .B(n6855), .Z(n3620) );
  NAND U6550 ( .A(n6856), .B(n3627), .Z(n6855) );
  OR U6551 ( .A(B[395]), .B(A[395]), .Z(n3627) );
  NANDN U6552 ( .A(n3629), .B(n6857), .Z(n6856) );
  NAND U6553 ( .A(n6858), .B(n3631), .Z(n6857) );
  OR U6554 ( .A(B[394]), .B(A[394]), .Z(n3631) );
  NANDN U6555 ( .A(n3633), .B(n6859), .Z(n6858) );
  NAND U6556 ( .A(n3636), .B(n3638), .Z(n6859) );
  AND U6557 ( .A(B[392]), .B(A[392]), .Z(n3638) );
  OR U6558 ( .A(B[393]), .B(A[393]), .Z(n3636) );
  AND U6559 ( .A(B[393]), .B(A[393]), .Z(n3633) );
  AND U6560 ( .A(B[394]), .B(A[394]), .Z(n3629) );
  AND U6561 ( .A(B[395]), .B(A[395]), .Z(n3626) );
  AND U6562 ( .A(B[396]), .B(A[396]), .Z(n3615) );
  AND U6563 ( .A(B[397]), .B(A[397]), .Z(n3610) );
  AND U6564 ( .A(B[398]), .B(A[398]), .Z(n3606) );
  AND U6565 ( .A(B[399]), .B(A[399]), .Z(n3603) );
  NAND U6566 ( .A(n6860), .B(n6861), .Z(n3497) );
  AND U6567 ( .A(n6862), .B(n6863), .Z(n6861) );
  AND U6568 ( .A(n3516), .B(n3511), .Z(n6863) );
  AND U6569 ( .A(n3506), .B(n3502), .Z(n6862) );
  ANDN U6570 ( .B(n6864), .A(n3569), .Z(n6860) );
  NAND U6571 ( .A(n6865), .B(n6866), .Z(n3569) );
  AND U6572 ( .A(n3586), .B(n3582), .Z(n6866) );
  OR U6573 ( .A(B[400]), .B(A[400]), .Z(n3586) );
  AND U6574 ( .A(n3577), .B(n3573), .Z(n6865) );
  ANDN U6575 ( .B(n3520), .A(n3547), .Z(n6864) );
  NANDN U6576 ( .A(n3501), .B(n6867), .Z(n3495) );
  NAND U6577 ( .A(n6868), .B(n3502), .Z(n6867) );
  OR U6578 ( .A(B[415]), .B(A[415]), .Z(n3502) );
  NANDN U6579 ( .A(n3504), .B(n6869), .Z(n6868) );
  NAND U6580 ( .A(n6870), .B(n3506), .Z(n6869) );
  OR U6581 ( .A(B[414]), .B(A[414]), .Z(n3506) );
  NANDN U6582 ( .A(n3508), .B(n6871), .Z(n6870) );
  NAND U6583 ( .A(n6872), .B(n3511), .Z(n6871) );
  OR U6584 ( .A(B[413]), .B(A[413]), .Z(n3511) );
  NANDN U6585 ( .A(n3513), .B(n6873), .Z(n6872) );
  NAND U6586 ( .A(n6874), .B(n3516), .Z(n6873) );
  OR U6587 ( .A(B[412]), .B(A[412]), .Z(n3516) );
  NANDN U6588 ( .A(n3518), .B(n6875), .Z(n6874) );
  NAND U6589 ( .A(n6876), .B(n3520), .Z(n6875) );
  AND U6590 ( .A(n6877), .B(n6878), .Z(n3520) );
  AND U6591 ( .A(n3543), .B(n3534), .Z(n6878) );
  OR U6592 ( .A(B[408]), .B(A[408]), .Z(n3543) );
  AND U6593 ( .A(n3529), .B(n3525), .Z(n6877) );
  NANDN U6594 ( .A(n3545), .B(n6879), .Z(n6876) );
  NANDN U6595 ( .A(n3547), .B(n3568), .Z(n6879) );
  NANDN U6596 ( .A(n3572), .B(n6880), .Z(n3568) );
  NAND U6597 ( .A(n6881), .B(n3573), .Z(n6880) );
  OR U6598 ( .A(B[403]), .B(A[403]), .Z(n3573) );
  NANDN U6599 ( .A(n3575), .B(n6882), .Z(n6881) );
  NAND U6600 ( .A(n6883), .B(n3577), .Z(n6882) );
  OR U6601 ( .A(B[402]), .B(A[402]), .Z(n3577) );
  NANDN U6602 ( .A(n3579), .B(n6884), .Z(n6883) );
  NAND U6603 ( .A(n3582), .B(n3584), .Z(n6884) );
  AND U6604 ( .A(B[400]), .B(A[400]), .Z(n3584) );
  OR U6605 ( .A(B[401]), .B(A[401]), .Z(n3582) );
  AND U6606 ( .A(B[401]), .B(A[401]), .Z(n3579) );
  AND U6607 ( .A(B[402]), .B(A[402]), .Z(n3575) );
  AND U6608 ( .A(B[403]), .B(A[403]), .Z(n3572) );
  NAND U6609 ( .A(n6885), .B(n6886), .Z(n3547) );
  AND U6610 ( .A(n3565), .B(n3561), .Z(n6886) );
  OR U6611 ( .A(B[404]), .B(A[404]), .Z(n3565) );
  AND U6612 ( .A(n3556), .B(n3552), .Z(n6885) );
  NANDN U6613 ( .A(n3551), .B(n6887), .Z(n3545) );
  NAND U6614 ( .A(n6888), .B(n3552), .Z(n6887) );
  OR U6615 ( .A(B[407]), .B(A[407]), .Z(n3552) );
  NANDN U6616 ( .A(n3554), .B(n6889), .Z(n6888) );
  NAND U6617 ( .A(n6890), .B(n3556), .Z(n6889) );
  OR U6618 ( .A(B[406]), .B(A[406]), .Z(n3556) );
  NANDN U6619 ( .A(n3558), .B(n6891), .Z(n6890) );
  NAND U6620 ( .A(n3561), .B(n3563), .Z(n6891) );
  AND U6621 ( .A(B[404]), .B(A[404]), .Z(n3563) );
  OR U6622 ( .A(B[405]), .B(A[405]), .Z(n3561) );
  AND U6623 ( .A(B[405]), .B(A[405]), .Z(n3558) );
  AND U6624 ( .A(B[406]), .B(A[406]), .Z(n3554) );
  AND U6625 ( .A(B[407]), .B(A[407]), .Z(n3551) );
  NANDN U6626 ( .A(n3524), .B(n6892), .Z(n3518) );
  NAND U6627 ( .A(n6893), .B(n3525), .Z(n6892) );
  OR U6628 ( .A(B[411]), .B(A[411]), .Z(n3525) );
  NANDN U6629 ( .A(n3527), .B(n6894), .Z(n6893) );
  NAND U6630 ( .A(n6895), .B(n3529), .Z(n6894) );
  OR U6631 ( .A(B[410]), .B(A[410]), .Z(n3529) );
  NANDN U6632 ( .A(n3531), .B(n6896), .Z(n6895) );
  NAND U6633 ( .A(n3534), .B(n3541), .Z(n6896) );
  AND U6634 ( .A(B[408]), .B(A[408]), .Z(n3541) );
  OR U6635 ( .A(B[409]), .B(A[409]), .Z(n3534) );
  AND U6636 ( .A(B[409]), .B(A[409]), .Z(n3531) );
  AND U6637 ( .A(B[410]), .B(A[410]), .Z(n3527) );
  AND U6638 ( .A(B[411]), .B(A[411]), .Z(n3524) );
  AND U6639 ( .A(B[412]), .B(A[412]), .Z(n3513) );
  AND U6640 ( .A(B[413]), .B(A[413]), .Z(n3508) );
  AND U6641 ( .A(B[414]), .B(A[414]), .Z(n3504) );
  AND U6642 ( .A(B[415]), .B(A[415]), .Z(n3501) );
  NANDN U6643 ( .A(n3404), .B(n6897), .Z(n3398) );
  NAND U6644 ( .A(n6898), .B(n3405), .Z(n6897) );
  OR U6645 ( .A(B[431]), .B(A[431]), .Z(n3405) );
  NANDN U6646 ( .A(n3407), .B(n6899), .Z(n6898) );
  NAND U6647 ( .A(n6900), .B(n3409), .Z(n6899) );
  OR U6648 ( .A(B[430]), .B(A[430]), .Z(n3409) );
  NANDN U6649 ( .A(n3411), .B(n6901), .Z(n6900) );
  NAND U6650 ( .A(n6902), .B(n3414), .Z(n6901) );
  OR U6651 ( .A(B[429]), .B(A[429]), .Z(n3414) );
  NANDN U6652 ( .A(n3421), .B(n6903), .Z(n6902) );
  NAND U6653 ( .A(n6904), .B(n3424), .Z(n6903) );
  OR U6654 ( .A(B[428]), .B(A[428]), .Z(n3424) );
  NANDN U6655 ( .A(n3426), .B(n6905), .Z(n6904) );
  NAND U6656 ( .A(n6906), .B(n3428), .Z(n6905) );
  AND U6657 ( .A(n6907), .B(n6908), .Z(n3428) );
  AND U6658 ( .A(n3446), .B(n3442), .Z(n6908) );
  OR U6659 ( .A(B[424]), .B(A[424]), .Z(n3446) );
  AND U6660 ( .A(n3437), .B(n3433), .Z(n6907) );
  NANDN U6661 ( .A(n3448), .B(n6909), .Z(n6906) );
  NANDN U6662 ( .A(n3450), .B(n3471), .Z(n6909) );
  NANDN U6663 ( .A(n3479), .B(n6910), .Z(n3471) );
  NAND U6664 ( .A(n6911), .B(n3480), .Z(n6910) );
  OR U6665 ( .A(B[419]), .B(A[419]), .Z(n3480) );
  NANDN U6666 ( .A(n3482), .B(n6912), .Z(n6911) );
  NAND U6667 ( .A(n6913), .B(n3484), .Z(n6912) );
  OR U6668 ( .A(B[418]), .B(A[418]), .Z(n3484) );
  NANDN U6669 ( .A(n3486), .B(n6914), .Z(n6913) );
  NAND U6670 ( .A(n3489), .B(n3491), .Z(n6914) );
  AND U6671 ( .A(B[416]), .B(A[416]), .Z(n3491) );
  OR U6672 ( .A(B[417]), .B(A[417]), .Z(n3489) );
  AND U6673 ( .A(B[417]), .B(A[417]), .Z(n3486) );
  AND U6674 ( .A(B[418]), .B(A[418]), .Z(n3482) );
  AND U6675 ( .A(B[419]), .B(A[419]), .Z(n3479) );
  NAND U6676 ( .A(n6915), .B(n6916), .Z(n3450) );
  AND U6677 ( .A(n3468), .B(n3464), .Z(n6916) );
  OR U6678 ( .A(B[420]), .B(A[420]), .Z(n3468) );
  AND U6679 ( .A(n3459), .B(n3455), .Z(n6915) );
  NANDN U6680 ( .A(n3454), .B(n6917), .Z(n3448) );
  NAND U6681 ( .A(n6918), .B(n3455), .Z(n6917) );
  OR U6682 ( .A(B[423]), .B(A[423]), .Z(n3455) );
  NANDN U6683 ( .A(n3457), .B(n6919), .Z(n6918) );
  NAND U6684 ( .A(n6920), .B(n3459), .Z(n6919) );
  OR U6685 ( .A(B[422]), .B(A[422]), .Z(n3459) );
  NANDN U6686 ( .A(n3461), .B(n6921), .Z(n6920) );
  NAND U6687 ( .A(n3464), .B(n3466), .Z(n6921) );
  AND U6688 ( .A(B[420]), .B(A[420]), .Z(n3466) );
  OR U6689 ( .A(B[421]), .B(A[421]), .Z(n3464) );
  AND U6690 ( .A(B[421]), .B(A[421]), .Z(n3461) );
  AND U6691 ( .A(B[422]), .B(A[422]), .Z(n3457) );
  AND U6692 ( .A(B[423]), .B(A[423]), .Z(n3454) );
  NANDN U6693 ( .A(n3432), .B(n6922), .Z(n3426) );
  NAND U6694 ( .A(n6923), .B(n3433), .Z(n6922) );
  OR U6695 ( .A(B[427]), .B(A[427]), .Z(n3433) );
  NANDN U6696 ( .A(n3435), .B(n6924), .Z(n6923) );
  NAND U6697 ( .A(n6925), .B(n3437), .Z(n6924) );
  OR U6698 ( .A(B[426]), .B(A[426]), .Z(n3437) );
  NANDN U6699 ( .A(n3439), .B(n6926), .Z(n6925) );
  NAND U6700 ( .A(n3442), .B(n3444), .Z(n6926) );
  AND U6701 ( .A(B[424]), .B(A[424]), .Z(n3444) );
  OR U6702 ( .A(B[425]), .B(A[425]), .Z(n3442) );
  AND U6703 ( .A(B[425]), .B(A[425]), .Z(n3439) );
  AND U6704 ( .A(B[426]), .B(A[426]), .Z(n3435) );
  AND U6705 ( .A(B[427]), .B(A[427]), .Z(n3432) );
  AND U6706 ( .A(B[428]), .B(A[428]), .Z(n3421) );
  AND U6707 ( .A(B[429]), .B(A[429]), .Z(n3411) );
  AND U6708 ( .A(B[430]), .B(A[430]), .Z(n3407) );
  AND U6709 ( .A(B[431]), .B(A[431]), .Z(n3404) );
  NAND U6710 ( .A(n6927), .B(n6928), .Z(n6783) );
  AND U6711 ( .A(n6929), .B(n6930), .Z(n6928) );
  AND U6712 ( .A(n3322), .B(n3317), .Z(n6930) );
  OR U6713 ( .A(A[445]), .B(B[445]), .Z(n3317) );
  OR U6714 ( .A(A[444]), .B(B[444]), .Z(n3322) );
  AND U6715 ( .A(n3312), .B(n3308), .Z(n6929) );
  OR U6716 ( .A(B[447]), .B(A[447]), .Z(n3308) );
  OR U6717 ( .A(A[446]), .B(B[446]), .Z(n3312) );
  ANDN U6718 ( .B(n6931), .A(n3348), .Z(n6927) );
  NAND U6719 ( .A(n6932), .B(n6933), .Z(n3348) );
  AND U6720 ( .A(n3374), .B(n3370), .Z(n6933) );
  OR U6721 ( .A(A[437]), .B(B[437]), .Z(n3370) );
  OR U6722 ( .A(A[436]), .B(B[436]), .Z(n3374) );
  AND U6723 ( .A(n3365), .B(n3361), .Z(n6932) );
  OR U6724 ( .A(B[439]), .B(A[439]), .Z(n3361) );
  OR U6725 ( .A(A[438]), .B(B[438]), .Z(n3365) );
  NOR U6726 ( .A(n3378), .B(n3326), .Z(n6931) );
  NAND U6727 ( .A(n6934), .B(n6935), .Z(n3326) );
  AND U6728 ( .A(n3344), .B(n3340), .Z(n6935) );
  OR U6729 ( .A(A[441]), .B(B[441]), .Z(n3340) );
  OR U6730 ( .A(A[440]), .B(B[440]), .Z(n3344) );
  AND U6731 ( .A(n3335), .B(n3331), .Z(n6934) );
  OR U6732 ( .A(B[443]), .B(A[443]), .Z(n3331) );
  OR U6733 ( .A(A[442]), .B(B[442]), .Z(n3335) );
  NAND U6734 ( .A(n6936), .B(n6937), .Z(n3378) );
  AND U6735 ( .A(n3396), .B(n3392), .Z(n6937) );
  OR U6736 ( .A(A[433]), .B(B[433]), .Z(n3392) );
  OR U6737 ( .A(A[432]), .B(B[432]), .Z(n3396) );
  AND U6738 ( .A(n3387), .B(n3383), .Z(n6936) );
  OR U6739 ( .A(B[435]), .B(A[435]), .Z(n3383) );
  OR U6740 ( .A(A[434]), .B(B[434]), .Z(n3387) );
  NAND U6741 ( .A(n6938), .B(n6939), .Z(n3205) );
  AND U6742 ( .A(n6940), .B(n6941), .Z(n6939) );
  AND U6743 ( .A(n3224), .B(n3219), .Z(n6941) );
  AND U6744 ( .A(n3214), .B(n3210), .Z(n6940) );
  ANDN U6745 ( .B(n6942), .A(n3277), .Z(n6938) );
  NAND U6746 ( .A(n6943), .B(n6944), .Z(n3277) );
  AND U6747 ( .A(n3299), .B(n3290), .Z(n6944) );
  OR U6748 ( .A(B[448]), .B(A[448]), .Z(n3299) );
  AND U6749 ( .A(n3285), .B(n3281), .Z(n6943) );
  ANDN U6750 ( .B(n3228), .A(n3255), .Z(n6942) );
  NANDN U6751 ( .A(n3209), .B(n6945), .Z(n3203) );
  NAND U6752 ( .A(n6946), .B(n3210), .Z(n6945) );
  OR U6753 ( .A(B[463]), .B(A[463]), .Z(n3210) );
  NANDN U6754 ( .A(n3212), .B(n6947), .Z(n6946) );
  NAND U6755 ( .A(n6948), .B(n3214), .Z(n6947) );
  OR U6756 ( .A(B[462]), .B(A[462]), .Z(n3214) );
  NANDN U6757 ( .A(n3216), .B(n6949), .Z(n6948) );
  NAND U6758 ( .A(n6950), .B(n3219), .Z(n6949) );
  OR U6759 ( .A(B[461]), .B(A[461]), .Z(n3219) );
  NANDN U6760 ( .A(n3221), .B(n6951), .Z(n6950) );
  NAND U6761 ( .A(n6952), .B(n3224), .Z(n6951) );
  OR U6762 ( .A(B[460]), .B(A[460]), .Z(n3224) );
  NANDN U6763 ( .A(n3226), .B(n6953), .Z(n6952) );
  NAND U6764 ( .A(n6954), .B(n3228), .Z(n6953) );
  AND U6765 ( .A(n6955), .B(n6956), .Z(n3228) );
  AND U6766 ( .A(n3251), .B(n3247), .Z(n6956) );
  OR U6767 ( .A(B[456]), .B(A[456]), .Z(n3251) );
  AND U6768 ( .A(n3242), .B(n3238), .Z(n6955) );
  NANDN U6769 ( .A(n3253), .B(n6957), .Z(n6954) );
  NANDN U6770 ( .A(n3255), .B(n3276), .Z(n6957) );
  NANDN U6771 ( .A(n3280), .B(n6958), .Z(n3276) );
  NAND U6772 ( .A(n6959), .B(n3281), .Z(n6958) );
  OR U6773 ( .A(B[451]), .B(A[451]), .Z(n3281) );
  NANDN U6774 ( .A(n3283), .B(n6960), .Z(n6959) );
  NAND U6775 ( .A(n6961), .B(n3285), .Z(n6960) );
  OR U6776 ( .A(B[450]), .B(A[450]), .Z(n3285) );
  NANDN U6777 ( .A(n3287), .B(n6962), .Z(n6961) );
  NAND U6778 ( .A(n3290), .B(n3297), .Z(n6962) );
  AND U6779 ( .A(B[448]), .B(A[448]), .Z(n3297) );
  OR U6780 ( .A(B[449]), .B(A[449]), .Z(n3290) );
  AND U6781 ( .A(B[449]), .B(A[449]), .Z(n3287) );
  AND U6782 ( .A(B[450]), .B(A[450]), .Z(n3283) );
  AND U6783 ( .A(B[451]), .B(A[451]), .Z(n3280) );
  NAND U6784 ( .A(n6963), .B(n6964), .Z(n3255) );
  AND U6785 ( .A(n3273), .B(n3269), .Z(n6964) );
  OR U6786 ( .A(B[452]), .B(A[452]), .Z(n3273) );
  AND U6787 ( .A(n3264), .B(n3260), .Z(n6963) );
  NANDN U6788 ( .A(n3259), .B(n6965), .Z(n3253) );
  NAND U6789 ( .A(n6966), .B(n3260), .Z(n6965) );
  OR U6790 ( .A(B[455]), .B(A[455]), .Z(n3260) );
  NANDN U6791 ( .A(n3262), .B(n6967), .Z(n6966) );
  NAND U6792 ( .A(n6968), .B(n3264), .Z(n6967) );
  OR U6793 ( .A(B[454]), .B(A[454]), .Z(n3264) );
  NANDN U6794 ( .A(n3266), .B(n6969), .Z(n6968) );
  NAND U6795 ( .A(n3269), .B(n3271), .Z(n6969) );
  AND U6796 ( .A(B[452]), .B(A[452]), .Z(n3271) );
  OR U6797 ( .A(B[453]), .B(A[453]), .Z(n3269) );
  AND U6798 ( .A(B[453]), .B(A[453]), .Z(n3266) );
  AND U6799 ( .A(B[454]), .B(A[454]), .Z(n3262) );
  AND U6800 ( .A(B[455]), .B(A[455]), .Z(n3259) );
  NANDN U6801 ( .A(n3237), .B(n6970), .Z(n3226) );
  NAND U6802 ( .A(n6971), .B(n3238), .Z(n6970) );
  OR U6803 ( .A(B[459]), .B(A[459]), .Z(n3238) );
  NANDN U6804 ( .A(n3240), .B(n6972), .Z(n6971) );
  NAND U6805 ( .A(n6973), .B(n3242), .Z(n6972) );
  OR U6806 ( .A(B[458]), .B(A[458]), .Z(n3242) );
  NANDN U6807 ( .A(n3244), .B(n6974), .Z(n6973) );
  NAND U6808 ( .A(n3247), .B(n3249), .Z(n6974) );
  AND U6809 ( .A(B[456]), .B(A[456]), .Z(n3249) );
  OR U6810 ( .A(B[457]), .B(A[457]), .Z(n3247) );
  AND U6811 ( .A(B[457]), .B(A[457]), .Z(n3244) );
  AND U6812 ( .A(B[458]), .B(A[458]), .Z(n3240) );
  AND U6813 ( .A(B[459]), .B(A[459]), .Z(n3237) );
  AND U6814 ( .A(B[460]), .B(A[460]), .Z(n3221) );
  AND U6815 ( .A(B[461]), .B(A[461]), .Z(n3216) );
  AND U6816 ( .A(B[462]), .B(A[462]), .Z(n3212) );
  AND U6817 ( .A(B[463]), .B(A[463]), .Z(n3209) );
  NAND U6818 ( .A(n6975), .B(n6976), .Z(n3104) );
  AND U6819 ( .A(n6977), .B(n6978), .Z(n6976) );
  AND U6820 ( .A(n3131), .B(n3126), .Z(n6978) );
  AND U6821 ( .A(n3121), .B(n3117), .Z(n6977) );
  ANDN U6822 ( .B(n6979), .A(n3184), .Z(n6975) );
  NAND U6823 ( .A(n6980), .B(n6981), .Z(n3184) );
  AND U6824 ( .A(n3201), .B(n3197), .Z(n6981) );
  OR U6825 ( .A(B[464]), .B(A[464]), .Z(n3201) );
  AND U6826 ( .A(n3192), .B(n3188), .Z(n6980) );
  ANDN U6827 ( .B(n3135), .A(n3157), .Z(n6979) );
  NANDN U6828 ( .A(n3116), .B(n6982), .Z(n3102) );
  NAND U6829 ( .A(n6983), .B(n3117), .Z(n6982) );
  OR U6830 ( .A(B[479]), .B(A[479]), .Z(n3117) );
  NANDN U6831 ( .A(n3119), .B(n6984), .Z(n6983) );
  NAND U6832 ( .A(n6985), .B(n3121), .Z(n6984) );
  OR U6833 ( .A(B[478]), .B(A[478]), .Z(n3121) );
  NANDN U6834 ( .A(n3123), .B(n6986), .Z(n6985) );
  NAND U6835 ( .A(n6987), .B(n3126), .Z(n6986) );
  OR U6836 ( .A(B[477]), .B(A[477]), .Z(n3126) );
  NANDN U6837 ( .A(n3128), .B(n6988), .Z(n6987) );
  NAND U6838 ( .A(n6989), .B(n3131), .Z(n6988) );
  OR U6839 ( .A(B[476]), .B(A[476]), .Z(n3131) );
  NANDN U6840 ( .A(n3133), .B(n6990), .Z(n6989) );
  NAND U6841 ( .A(n6991), .B(n3135), .Z(n6990) );
  AND U6842 ( .A(n6992), .B(n6993), .Z(n3135) );
  AND U6843 ( .A(n3153), .B(n3149), .Z(n6993) );
  OR U6844 ( .A(B[472]), .B(A[472]), .Z(n3153) );
  AND U6845 ( .A(n3144), .B(n3140), .Z(n6992) );
  NANDN U6846 ( .A(n3155), .B(n6994), .Z(n6991) );
  NANDN U6847 ( .A(n3157), .B(n3183), .Z(n6994) );
  NANDN U6848 ( .A(n3187), .B(n6995), .Z(n3183) );
  NAND U6849 ( .A(n6996), .B(n3188), .Z(n6995) );
  OR U6850 ( .A(B[467]), .B(A[467]), .Z(n3188) );
  NANDN U6851 ( .A(n3190), .B(n6997), .Z(n6996) );
  NAND U6852 ( .A(n6998), .B(n3192), .Z(n6997) );
  OR U6853 ( .A(B[466]), .B(A[466]), .Z(n3192) );
  NANDN U6854 ( .A(n3194), .B(n6999), .Z(n6998) );
  NAND U6855 ( .A(n3197), .B(n3199), .Z(n6999) );
  AND U6856 ( .A(B[464]), .B(A[464]), .Z(n3199) );
  OR U6857 ( .A(B[465]), .B(A[465]), .Z(n3197) );
  AND U6858 ( .A(B[465]), .B(A[465]), .Z(n3194) );
  AND U6859 ( .A(B[466]), .B(A[466]), .Z(n3190) );
  AND U6860 ( .A(B[467]), .B(A[467]), .Z(n3187) );
  NAND U6861 ( .A(n7000), .B(n7001), .Z(n3157) );
  AND U6862 ( .A(n3180), .B(n3171), .Z(n7001) );
  OR U6863 ( .A(B[468]), .B(A[468]), .Z(n3180) );
  AND U6864 ( .A(n3166), .B(n3162), .Z(n7000) );
  NANDN U6865 ( .A(n3161), .B(n7002), .Z(n3155) );
  NAND U6866 ( .A(n7003), .B(n3162), .Z(n7002) );
  OR U6867 ( .A(B[471]), .B(A[471]), .Z(n3162) );
  NANDN U6868 ( .A(n3164), .B(n7004), .Z(n7003) );
  NAND U6869 ( .A(n7005), .B(n3166), .Z(n7004) );
  OR U6870 ( .A(B[470]), .B(A[470]), .Z(n3166) );
  NANDN U6871 ( .A(n3168), .B(n7006), .Z(n7005) );
  NAND U6872 ( .A(n3171), .B(n3178), .Z(n7006) );
  AND U6873 ( .A(B[468]), .B(A[468]), .Z(n3178) );
  OR U6874 ( .A(B[469]), .B(A[469]), .Z(n3171) );
  AND U6875 ( .A(B[469]), .B(A[469]), .Z(n3168) );
  AND U6876 ( .A(B[470]), .B(A[470]), .Z(n3164) );
  AND U6877 ( .A(B[471]), .B(A[471]), .Z(n3161) );
  NANDN U6878 ( .A(n3139), .B(n7007), .Z(n3133) );
  NAND U6879 ( .A(n7008), .B(n3140), .Z(n7007) );
  OR U6880 ( .A(B[475]), .B(A[475]), .Z(n3140) );
  NANDN U6881 ( .A(n3142), .B(n7009), .Z(n7008) );
  NAND U6882 ( .A(n7010), .B(n3144), .Z(n7009) );
  OR U6883 ( .A(B[474]), .B(A[474]), .Z(n3144) );
  NANDN U6884 ( .A(n3146), .B(n7011), .Z(n7010) );
  NAND U6885 ( .A(n3149), .B(n3151), .Z(n7011) );
  AND U6886 ( .A(B[472]), .B(A[472]), .Z(n3151) );
  OR U6887 ( .A(B[473]), .B(A[473]), .Z(n3149) );
  AND U6888 ( .A(B[473]), .B(A[473]), .Z(n3146) );
  AND U6889 ( .A(B[474]), .B(A[474]), .Z(n3142) );
  AND U6890 ( .A(B[475]), .B(A[475]), .Z(n3139) );
  AND U6891 ( .A(B[476]), .B(A[476]), .Z(n3128) );
  AND U6892 ( .A(B[477]), .B(A[477]), .Z(n3123) );
  AND U6893 ( .A(B[478]), .B(A[478]), .Z(n3119) );
  AND U6894 ( .A(B[479]), .B(A[479]), .Z(n3116) );
  NAND U6895 ( .A(n7012), .B(n7013), .Z(n3015) );
  AND U6896 ( .A(n7014), .B(n7015), .Z(n7013) );
  AND U6897 ( .A(n3034), .B(n3029), .Z(n7015) );
  AND U6898 ( .A(n3024), .B(n3020), .Z(n7014) );
  ANDN U6899 ( .B(n7016), .A(n3083), .Z(n7012) );
  NAND U6900 ( .A(n7017), .B(n7018), .Z(n3083) );
  AND U6901 ( .A(n3100), .B(n3096), .Z(n7018) );
  OR U6902 ( .A(B[480]), .B(A[480]), .Z(n3100) );
  AND U6903 ( .A(n3091), .B(n3087), .Z(n7017) );
  ANDN U6904 ( .B(n3038), .A(n3061), .Z(n7016) );
  NANDN U6905 ( .A(n3019), .B(n7019), .Z(n3013) );
  NAND U6906 ( .A(n7020), .B(n3020), .Z(n7019) );
  OR U6907 ( .A(B[495]), .B(A[495]), .Z(n3020) );
  NANDN U6908 ( .A(n3022), .B(n7021), .Z(n7020) );
  NAND U6909 ( .A(n7022), .B(n3024), .Z(n7021) );
  OR U6910 ( .A(B[494]), .B(A[494]), .Z(n3024) );
  NANDN U6911 ( .A(n3026), .B(n7023), .Z(n7022) );
  NAND U6912 ( .A(n7024), .B(n3029), .Z(n7023) );
  OR U6913 ( .A(B[493]), .B(A[493]), .Z(n3029) );
  NANDN U6914 ( .A(n3031), .B(n7025), .Z(n7024) );
  NAND U6915 ( .A(n7026), .B(n3034), .Z(n7025) );
  OR U6916 ( .A(B[492]), .B(A[492]), .Z(n3034) );
  NANDN U6917 ( .A(n3036), .B(n7027), .Z(n7026) );
  NAND U6918 ( .A(n7028), .B(n3038), .Z(n7027) );
  AND U6919 ( .A(n7029), .B(n7030), .Z(n3038) );
  AND U6920 ( .A(n3057), .B(n3052), .Z(n7030) );
  OR U6921 ( .A(B[488]), .B(A[488]), .Z(n3057) );
  AND U6922 ( .A(n3047), .B(n3043), .Z(n7029) );
  NANDN U6923 ( .A(n3059), .B(n7031), .Z(n7028) );
  NANDN U6924 ( .A(n3061), .B(n3082), .Z(n7031) );
  NANDN U6925 ( .A(n3086), .B(n7032), .Z(n3082) );
  NAND U6926 ( .A(n7033), .B(n3087), .Z(n7032) );
  OR U6927 ( .A(B[483]), .B(A[483]), .Z(n3087) );
  NANDN U6928 ( .A(n3089), .B(n7034), .Z(n7033) );
  NAND U6929 ( .A(n7035), .B(n3091), .Z(n7034) );
  OR U6930 ( .A(B[482]), .B(A[482]), .Z(n3091) );
  NANDN U6931 ( .A(n3093), .B(n7036), .Z(n7035) );
  NAND U6932 ( .A(n3096), .B(n3098), .Z(n7036) );
  AND U6933 ( .A(B[480]), .B(A[480]), .Z(n3098) );
  OR U6934 ( .A(B[481]), .B(A[481]), .Z(n3096) );
  AND U6935 ( .A(B[481]), .B(A[481]), .Z(n3093) );
  AND U6936 ( .A(B[482]), .B(A[482]), .Z(n3089) );
  AND U6937 ( .A(B[483]), .B(A[483]), .Z(n3086) );
  NAND U6938 ( .A(n7037), .B(n7038), .Z(n3061) );
  AND U6939 ( .A(n3079), .B(n3075), .Z(n7038) );
  OR U6940 ( .A(B[484]), .B(A[484]), .Z(n3079) );
  AND U6941 ( .A(n3070), .B(n3066), .Z(n7037) );
  NANDN U6942 ( .A(n3065), .B(n7039), .Z(n3059) );
  NAND U6943 ( .A(n7040), .B(n3066), .Z(n7039) );
  OR U6944 ( .A(B[487]), .B(A[487]), .Z(n3066) );
  NANDN U6945 ( .A(n3068), .B(n7041), .Z(n7040) );
  NAND U6946 ( .A(n7042), .B(n3070), .Z(n7041) );
  OR U6947 ( .A(B[486]), .B(A[486]), .Z(n3070) );
  NANDN U6948 ( .A(n3072), .B(n7043), .Z(n7042) );
  NAND U6949 ( .A(n3075), .B(n3077), .Z(n7043) );
  AND U6950 ( .A(B[484]), .B(A[484]), .Z(n3077) );
  OR U6951 ( .A(B[485]), .B(A[485]), .Z(n3075) );
  AND U6952 ( .A(B[485]), .B(A[485]), .Z(n3072) );
  AND U6953 ( .A(B[486]), .B(A[486]), .Z(n3068) );
  AND U6954 ( .A(B[487]), .B(A[487]), .Z(n3065) );
  NANDN U6955 ( .A(n3042), .B(n7044), .Z(n3036) );
  NAND U6956 ( .A(n7045), .B(n3043), .Z(n7044) );
  OR U6957 ( .A(B[491]), .B(A[491]), .Z(n3043) );
  NANDN U6958 ( .A(n3045), .B(n7046), .Z(n7045) );
  NAND U6959 ( .A(n7047), .B(n3047), .Z(n7046) );
  OR U6960 ( .A(B[490]), .B(A[490]), .Z(n3047) );
  NANDN U6961 ( .A(n3049), .B(n7048), .Z(n7047) );
  NAND U6962 ( .A(n3052), .B(n3055), .Z(n7048) );
  AND U6963 ( .A(B[488]), .B(A[488]), .Z(n3055) );
  OR U6964 ( .A(B[489]), .B(A[489]), .Z(n3052) );
  AND U6965 ( .A(B[489]), .B(A[489]), .Z(n3049) );
  AND U6966 ( .A(B[490]), .B(A[490]), .Z(n3045) );
  AND U6967 ( .A(B[491]), .B(A[491]), .Z(n3042) );
  AND U6968 ( .A(B[492]), .B(A[492]), .Z(n3031) );
  AND U6969 ( .A(B[493]), .B(A[493]), .Z(n3026) );
  AND U6970 ( .A(B[494]), .B(A[494]), .Z(n3022) );
  AND U6971 ( .A(B[495]), .B(A[495]), .Z(n3019) );
  ANDN U6972 ( .B(n7049), .A(n2984), .Z(n5859) );
  NAND U6973 ( .A(n7050), .B(n7051), .Z(n2984) );
  AND U6974 ( .A(n3011), .B(n3007), .Z(n7051) );
  OR U6975 ( .A(B[496]), .B(A[496]), .Z(n3011) );
  ANDN U6976 ( .B(n2998), .A(n3001), .Z(n7050) );
  ANDN U6977 ( .B(n2963), .A(n2940), .Z(n7049) );
  ANDN U6978 ( .B(n7052), .A(n2919), .Z(n5857) );
  AND U6979 ( .A(B[510]), .B(A[510]), .Z(n2919) );
  NAND U6980 ( .A(n7053), .B(n2921), .Z(n7052) );
  OR U6981 ( .A(A[510]), .B(B[510]), .Z(n2921) );
  NANDN U6982 ( .A(n2923), .B(n7054), .Z(n7053) );
  NAND U6983 ( .A(n7055), .B(n2926), .Z(n7054) );
  OR U6984 ( .A(B[509]), .B(A[509]), .Z(n2926) );
  NANDN U6985 ( .A(n2933), .B(n7056), .Z(n7055) );
  NANDN U6986 ( .A(n2935), .B(n7057), .Z(n7056) );
  NANDN U6987 ( .A(n2938), .B(n7058), .Z(n7057) );
  NANDN U6988 ( .A(n2940), .B(n7059), .Z(n7058) );
  NANDN U6989 ( .A(n2960), .B(n7060), .Z(n7059) );
  NAND U6990 ( .A(n2983), .B(n2963), .Z(n7060) );
  AND U6991 ( .A(n7061), .B(n7062), .Z(n2963) );
  AND U6992 ( .A(n2980), .B(n2976), .Z(n7062) );
  OR U6993 ( .A(B[500]), .B(A[500]), .Z(n2980) );
  AND U6994 ( .A(n2971), .B(n2967), .Z(n7061) );
  NANDN U6995 ( .A(n2997), .B(n7063), .Z(n2983) );
  NAND U6996 ( .A(n7064), .B(n2998), .Z(n7063) );
  OR U6997 ( .A(B[499]), .B(A[499]), .Z(n2998) );
  NANDN U6998 ( .A(n3000), .B(n7065), .Z(n7064) );
  NANDN U6999 ( .A(n3001), .B(n7066), .Z(n7065) );
  NANDN U7000 ( .A(n3004), .B(n7067), .Z(n7066) );
  NAND U7001 ( .A(n3007), .B(n3009), .Z(n7067) );
  AND U7002 ( .A(A[496]), .B(B[496]), .Z(n3009) );
  OR U7003 ( .A(B[497]), .B(A[497]), .Z(n3007) );
  AND U7004 ( .A(B[497]), .B(A[497]), .Z(n3004) );
  NOR U7005 ( .A(B[498]), .B(A[498]), .Z(n3001) );
  AND U7006 ( .A(B[498]), .B(A[498]), .Z(n3000) );
  AND U7007 ( .A(B[499]), .B(A[499]), .Z(n2997) );
  NANDN U7008 ( .A(n2966), .B(n7068), .Z(n2960) );
  NAND U7009 ( .A(n7069), .B(n2967), .Z(n7068) );
  OR U7010 ( .A(B[503]), .B(A[503]), .Z(n2967) );
  NANDN U7011 ( .A(n2969), .B(n7070), .Z(n7069) );
  NAND U7012 ( .A(n7071), .B(n2971), .Z(n7070) );
  OR U7013 ( .A(B[502]), .B(A[502]), .Z(n2971) );
  NANDN U7014 ( .A(n2973), .B(n7072), .Z(n7071) );
  NAND U7015 ( .A(n2976), .B(n2978), .Z(n7072) );
  AND U7016 ( .A(B[500]), .B(A[500]), .Z(n2978) );
  OR U7017 ( .A(B[501]), .B(A[501]), .Z(n2976) );
  AND U7018 ( .A(B[501]), .B(A[501]), .Z(n2973) );
  AND U7019 ( .A(B[502]), .B(A[502]), .Z(n2969) );
  AND U7020 ( .A(B[503]), .B(A[503]), .Z(n2966) );
  NAND U7021 ( .A(n7073), .B(n7074), .Z(n2940) );
  AND U7022 ( .A(n2958), .B(n2954), .Z(n7074) );
  OR U7023 ( .A(B[504]), .B(A[504]), .Z(n2958) );
  AND U7024 ( .A(n2949), .B(n2945), .Z(n7073) );
  NANDN U7025 ( .A(n2944), .B(n7075), .Z(n2938) );
  NAND U7026 ( .A(n7076), .B(n2945), .Z(n7075) );
  OR U7027 ( .A(B[507]), .B(A[507]), .Z(n2945) );
  NANDN U7028 ( .A(n2947), .B(n7077), .Z(n7076) );
  NAND U7029 ( .A(n7078), .B(n2949), .Z(n7077) );
  OR U7030 ( .A(B[506]), .B(A[506]), .Z(n2949) );
  NANDN U7031 ( .A(n2951), .B(n7079), .Z(n7078) );
  NAND U7032 ( .A(n2954), .B(n2956), .Z(n7079) );
  AND U7033 ( .A(B[504]), .B(A[504]), .Z(n2956) );
  OR U7034 ( .A(B[505]), .B(A[505]), .Z(n2954) );
  AND U7035 ( .A(B[505]), .B(A[505]), .Z(n2951) );
  AND U7036 ( .A(B[506]), .B(A[506]), .Z(n2947) );
  AND U7037 ( .A(B[507]), .B(A[507]), .Z(n2944) );
  NOR U7038 ( .A(B[508]), .B(A[508]), .Z(n2935) );
  AND U7039 ( .A(B[508]), .B(A[508]), .Z(n2933) );
  AND U7040 ( .A(B[509]), .B(A[509]), .Z(n2923) );
  NOR U7041 ( .A(B[511]), .B(A[511]), .Z(n2916) );
  NOR U7042 ( .A(n2820), .B(n5747), .Z(n5830) );
  NAND U7043 ( .A(n7080), .B(n7081), .Z(n5747) );
  AND U7044 ( .A(n7082), .B(n7083), .Z(n7081) );
  AND U7045 ( .A(n2549), .B(n2544), .Z(n7083) );
  OR U7046 ( .A(A[573]), .B(B[573]), .Z(n2544) );
  OR U7047 ( .A(A[572]), .B(B[572]), .Z(n2549) );
  AND U7048 ( .A(n2539), .B(n2535), .Z(n7082) );
  OR U7049 ( .A(B[575]), .B(A[575]), .Z(n2535) );
  OR U7050 ( .A(A[574]), .B(B[574]), .Z(n2539) );
  ANDN U7051 ( .B(n7084), .A(n2580), .Z(n7080) );
  NAND U7052 ( .A(n7085), .B(n7086), .Z(n2580) );
  AND U7053 ( .A(n2598), .B(n2594), .Z(n7086) );
  OR U7054 ( .A(A[565]), .B(B[565]), .Z(n2594) );
  OR U7055 ( .A(A[564]), .B(B[564]), .Z(n2598) );
  AND U7056 ( .A(n2589), .B(n2585), .Z(n7085) );
  OR U7057 ( .A(B[567]), .B(A[567]), .Z(n2585) );
  OR U7058 ( .A(A[566]), .B(B[566]), .Z(n2589) );
  NOR U7059 ( .A(n2602), .B(n2553), .Z(n7084) );
  NAND U7060 ( .A(n7087), .B(n7088), .Z(n2553) );
  AND U7061 ( .A(n2576), .B(n2567), .Z(n7088) );
  OR U7062 ( .A(A[569]), .B(B[569]), .Z(n2567) );
  OR U7063 ( .A(A[568]), .B(B[568]), .Z(n2576) );
  AND U7064 ( .A(n2562), .B(n2558), .Z(n7087) );
  OR U7065 ( .A(B[571]), .B(A[571]), .Z(n2558) );
  OR U7066 ( .A(A[570]), .B(B[570]), .Z(n2562) );
  NAND U7067 ( .A(n7089), .B(n7090), .Z(n2602) );
  AND U7068 ( .A(n2620), .B(n2616), .Z(n7090) );
  OR U7069 ( .A(A[561]), .B(B[561]), .Z(n2616) );
  OR U7070 ( .A(A[560]), .B(B[560]), .Z(n2620) );
  AND U7071 ( .A(n2611), .B(n2607), .Z(n7089) );
  OR U7072 ( .A(B[563]), .B(A[563]), .Z(n2607) );
  OR U7073 ( .A(A[562]), .B(B[562]), .Z(n2611) );
  NAND U7074 ( .A(n7091), .B(n7092), .Z(n2820) );
  AND U7075 ( .A(n7093), .B(n7094), .Z(n7092) );
  AND U7076 ( .A(n2839), .B(n2834), .Z(n7094) );
  OR U7077 ( .A(A[525]), .B(B[525]), .Z(n2834) );
  OR U7078 ( .A(A[524]), .B(B[524]), .Z(n2839) );
  AND U7079 ( .A(n2829), .B(n2825), .Z(n7093) );
  OR U7080 ( .A(B[527]), .B(A[527]), .Z(n2825) );
  OR U7081 ( .A(A[526]), .B(B[526]), .Z(n2829) );
  ANDN U7082 ( .B(n7095), .A(n2895), .Z(n7091) );
  NAND U7083 ( .A(n7096), .B(n7097), .Z(n2895) );
  AND U7084 ( .A(n2912), .B(n2908), .Z(n7097) );
  OR U7085 ( .A(A[513]), .B(B[513]), .Z(n2908) );
  OR U7086 ( .A(A[512]), .B(B[512]), .Z(n2912) );
  AND U7087 ( .A(n2903), .B(n2899), .Z(n7096) );
  OR U7088 ( .A(B[515]), .B(A[515]), .Z(n2899) );
  OR U7089 ( .A(A[514]), .B(B[514]), .Z(n2903) );
  NOR U7090 ( .A(n2865), .B(n2843), .Z(n7095) );
  NAND U7091 ( .A(n7098), .B(n7099), .Z(n2843) );
  AND U7092 ( .A(n2861), .B(n2857), .Z(n7099) );
  OR U7093 ( .A(A[521]), .B(B[521]), .Z(n2857) );
  OR U7094 ( .A(A[520]), .B(B[520]), .Z(n2861) );
  AND U7095 ( .A(n2852), .B(n2848), .Z(n7098) );
  OR U7096 ( .A(B[523]), .B(A[523]), .Z(n2848) );
  OR U7097 ( .A(A[522]), .B(B[522]), .Z(n2852) );
  NAND U7098 ( .A(n7100), .B(n7101), .Z(n2865) );
  AND U7099 ( .A(n2891), .B(n2887), .Z(n7101) );
  OR U7100 ( .A(A[517]), .B(B[517]), .Z(n2887) );
  OR U7101 ( .A(A[516]), .B(B[516]), .Z(n2891) );
  AND U7102 ( .A(n2882), .B(n2878), .Z(n7100) );
  OR U7103 ( .A(B[519]), .B(A[519]), .Z(n2878) );
  OR U7104 ( .A(A[518]), .B(B[518]), .Z(n2882) );
  NAND U7105 ( .A(n7102), .B(n7103), .Z(n2136) );
  NOR U7106 ( .A(n2336), .B(n2238), .Z(n7103) );
  NOR U7107 ( .A(n2436), .B(n7104), .Z(n7102) );
  NAND U7108 ( .A(n7105), .B(n7106), .Z(n2436) );
  AND U7109 ( .A(n7107), .B(n7108), .Z(n7106) );
  AND U7110 ( .A(n2459), .B(n2449), .Z(n7108) );
  AND U7111 ( .A(n2444), .B(n2440), .Z(n7107) );
  ANDN U7112 ( .B(n7109), .A(n2507), .Z(n7105) );
  NAND U7113 ( .A(n7110), .B(n7111), .Z(n2507) );
  AND U7114 ( .A(n2528), .B(n2524), .Z(n7111) );
  OR U7115 ( .A(A[576]), .B(B[576]), .Z(n2528) );
  AND U7116 ( .A(n2519), .B(n2515), .Z(n7110) );
  NOR U7117 ( .A(n2485), .B(n2463), .Z(n7109) );
  NAND U7118 ( .A(n7112), .B(n7113), .Z(n2134) );
  NAND U7119 ( .A(n7114), .B(n2149), .Z(n7113) );
  NANDN U7120 ( .A(n2151), .B(n7115), .Z(n7114) );
  NAND U7121 ( .A(n7116), .B(n2153), .Z(n7115) );
  NANDN U7122 ( .A(n2155), .B(n7117), .Z(n7116) );
  NAND U7123 ( .A(n7118), .B(n2158), .Z(n7117) );
  NANDN U7124 ( .A(n2160), .B(n7119), .Z(n7118) );
  NAND U7125 ( .A(n7120), .B(n2163), .Z(n7119) );
  NANDN U7126 ( .A(n2165), .B(n7121), .Z(n7120) );
  NANDN U7127 ( .A(n2167), .B(n7122), .Z(n7121) );
  NANDN U7128 ( .A(n2187), .B(n7123), .Z(n7122) );
  NANDN U7129 ( .A(n2189), .B(n2215), .Z(n7123) );
  NANDN U7130 ( .A(n2220), .B(n7124), .Z(n2215) );
  NAND U7131 ( .A(n7125), .B(n2221), .Z(n7124) );
  NANDN U7132 ( .A(n2223), .B(n7126), .Z(n7125) );
  NAND U7133 ( .A(n7127), .B(n2225), .Z(n7126) );
  NANDN U7134 ( .A(n2227), .B(n7128), .Z(n7127) );
  NAND U7135 ( .A(n2230), .B(n2232), .Z(n7128) );
  AND U7136 ( .A(A[624]), .B(B[624]), .Z(n2232) );
  AND U7137 ( .A(A[625]), .B(B[625]), .Z(n2227) );
  AND U7138 ( .A(A[626]), .B(B[626]), .Z(n2223) );
  AND U7139 ( .A(B[627]), .B(A[627]), .Z(n2220) );
  NANDN U7140 ( .A(n2193), .B(n7129), .Z(n2187) );
  NAND U7141 ( .A(n7130), .B(n2194), .Z(n7129) );
  NANDN U7142 ( .A(n2196), .B(n7131), .Z(n7130) );
  NAND U7143 ( .A(n7132), .B(n2198), .Z(n7131) );
  NANDN U7144 ( .A(n2200), .B(n7133), .Z(n7132) );
  NAND U7145 ( .A(n2203), .B(n2210), .Z(n7133) );
  AND U7146 ( .A(A[628]), .B(B[628]), .Z(n2210) );
  AND U7147 ( .A(A[629]), .B(B[629]), .Z(n2200) );
  AND U7148 ( .A(A[630]), .B(B[630]), .Z(n2196) );
  AND U7149 ( .A(B[631]), .B(A[631]), .Z(n2193) );
  NANDN U7150 ( .A(n2171), .B(n7134), .Z(n2165) );
  NAND U7151 ( .A(n7135), .B(n2172), .Z(n7134) );
  NANDN U7152 ( .A(n2174), .B(n7136), .Z(n7135) );
  NAND U7153 ( .A(n7137), .B(n2176), .Z(n7136) );
  NANDN U7154 ( .A(n2178), .B(n7138), .Z(n7137) );
  NAND U7155 ( .A(n2181), .B(n2183), .Z(n7138) );
  AND U7156 ( .A(A[632]), .B(B[632]), .Z(n2183) );
  AND U7157 ( .A(A[633]), .B(B[633]), .Z(n2178) );
  AND U7158 ( .A(A[634]), .B(B[634]), .Z(n2174) );
  AND U7159 ( .A(B[635]), .B(A[635]), .Z(n2171) );
  AND U7160 ( .A(A[636]), .B(B[636]), .Z(n2160) );
  AND U7161 ( .A(A[637]), .B(B[637]), .Z(n2155) );
  AND U7162 ( .A(A[638]), .B(B[638]), .Z(n2151) );
  ANDN U7163 ( .B(n7139), .A(n2148), .Z(n7112) );
  AND U7164 ( .A(B[639]), .B(A[639]), .Z(n2148) );
  NANDN U7165 ( .A(n7104), .B(n7140), .Z(n7139) );
  NANDN U7166 ( .A(n2236), .B(n7141), .Z(n7140) );
  NANDN U7167 ( .A(n2238), .B(n7142), .Z(n7141) );
  NANDN U7168 ( .A(n2334), .B(n7143), .Z(n7142) );
  NANDN U7169 ( .A(n2336), .B(n2435), .Z(n7143) );
  NANDN U7170 ( .A(n2439), .B(n7144), .Z(n2435) );
  NAND U7171 ( .A(n7145), .B(n2440), .Z(n7144) );
  OR U7172 ( .A(B[591]), .B(A[591]), .Z(n2440) );
  NANDN U7173 ( .A(n2442), .B(n7146), .Z(n7145) );
  NAND U7174 ( .A(n7147), .B(n2444), .Z(n7146) );
  OR U7175 ( .A(A[590]), .B(B[590]), .Z(n2444) );
  NANDN U7176 ( .A(n2446), .B(n7148), .Z(n7147) );
  NAND U7177 ( .A(n7149), .B(n2449), .Z(n7148) );
  OR U7178 ( .A(A[589]), .B(B[589]), .Z(n2449) );
  NANDN U7179 ( .A(n2456), .B(n7150), .Z(n7149) );
  NAND U7180 ( .A(n7151), .B(n2459), .Z(n7150) );
  OR U7181 ( .A(A[588]), .B(B[588]), .Z(n2459) );
  NANDN U7182 ( .A(n2461), .B(n7152), .Z(n7151) );
  NANDN U7183 ( .A(n2463), .B(n7153), .Z(n7152) );
  NANDN U7184 ( .A(n2483), .B(n7154), .Z(n7153) );
  NANDN U7185 ( .A(n2485), .B(n2506), .Z(n7154) );
  NANDN U7186 ( .A(n2514), .B(n7155), .Z(n2506) );
  NAND U7187 ( .A(n7156), .B(n2515), .Z(n7155) );
  OR U7188 ( .A(B[579]), .B(A[579]), .Z(n2515) );
  NANDN U7189 ( .A(n2517), .B(n7157), .Z(n7156) );
  NAND U7190 ( .A(n7158), .B(n2519), .Z(n7157) );
  OR U7191 ( .A(A[578]), .B(B[578]), .Z(n2519) );
  NANDN U7192 ( .A(n2521), .B(n7159), .Z(n7158) );
  NAND U7193 ( .A(n2524), .B(n2526), .Z(n7159) );
  AND U7194 ( .A(A[576]), .B(B[576]), .Z(n2526) );
  OR U7195 ( .A(A[577]), .B(B[577]), .Z(n2524) );
  AND U7196 ( .A(A[577]), .B(B[577]), .Z(n2521) );
  AND U7197 ( .A(A[578]), .B(B[578]), .Z(n2517) );
  AND U7198 ( .A(B[579]), .B(A[579]), .Z(n2514) );
  NAND U7199 ( .A(n7160), .B(n7161), .Z(n2485) );
  AND U7200 ( .A(n2503), .B(n2499), .Z(n7161) );
  OR U7201 ( .A(A[580]), .B(B[580]), .Z(n2503) );
  AND U7202 ( .A(n2494), .B(n2490), .Z(n7160) );
  NANDN U7203 ( .A(n2489), .B(n7162), .Z(n2483) );
  NAND U7204 ( .A(n7163), .B(n2490), .Z(n7162) );
  OR U7205 ( .A(B[583]), .B(A[583]), .Z(n2490) );
  NANDN U7206 ( .A(n2492), .B(n7164), .Z(n7163) );
  NAND U7207 ( .A(n7165), .B(n2494), .Z(n7164) );
  OR U7208 ( .A(A[582]), .B(B[582]), .Z(n2494) );
  NANDN U7209 ( .A(n2496), .B(n7166), .Z(n7165) );
  NAND U7210 ( .A(n2499), .B(n2501), .Z(n7166) );
  AND U7211 ( .A(A[580]), .B(B[580]), .Z(n2501) );
  OR U7212 ( .A(A[581]), .B(B[581]), .Z(n2499) );
  AND U7213 ( .A(A[581]), .B(B[581]), .Z(n2496) );
  AND U7214 ( .A(A[582]), .B(B[582]), .Z(n2492) );
  AND U7215 ( .A(B[583]), .B(A[583]), .Z(n2489) );
  NAND U7216 ( .A(n7167), .B(n7168), .Z(n2463) );
  AND U7217 ( .A(n2481), .B(n2477), .Z(n7168) );
  OR U7218 ( .A(A[584]), .B(B[584]), .Z(n2481) );
  AND U7219 ( .A(n2472), .B(n2468), .Z(n7167) );
  NANDN U7220 ( .A(n2467), .B(n7169), .Z(n2461) );
  NAND U7221 ( .A(n7170), .B(n2468), .Z(n7169) );
  OR U7222 ( .A(B[587]), .B(A[587]), .Z(n2468) );
  NANDN U7223 ( .A(n2470), .B(n7171), .Z(n7170) );
  NAND U7224 ( .A(n7172), .B(n2472), .Z(n7171) );
  OR U7225 ( .A(A[586]), .B(B[586]), .Z(n2472) );
  NANDN U7226 ( .A(n2474), .B(n7173), .Z(n7172) );
  NAND U7227 ( .A(n2477), .B(n2479), .Z(n7173) );
  AND U7228 ( .A(A[584]), .B(B[584]), .Z(n2479) );
  OR U7229 ( .A(A[585]), .B(B[585]), .Z(n2477) );
  AND U7230 ( .A(A[585]), .B(B[585]), .Z(n2474) );
  AND U7231 ( .A(A[586]), .B(B[586]), .Z(n2470) );
  AND U7232 ( .A(B[587]), .B(A[587]), .Z(n2467) );
  AND U7233 ( .A(A[588]), .B(B[588]), .Z(n2456) );
  AND U7234 ( .A(A[589]), .B(B[589]), .Z(n2446) );
  AND U7235 ( .A(A[590]), .B(B[590]), .Z(n2442) );
  AND U7236 ( .A(B[591]), .B(A[591]), .Z(n2439) );
  NAND U7237 ( .A(n7174), .B(n7175), .Z(n2336) );
  AND U7238 ( .A(n7176), .B(n7177), .Z(n7175) );
  AND U7239 ( .A(n2355), .B(n2350), .Z(n7177) );
  AND U7240 ( .A(n2345), .B(n2341), .Z(n7176) );
  ANDN U7241 ( .B(n7178), .A(n2415), .Z(n7174) );
  NAND U7242 ( .A(n7179), .B(n7180), .Z(n2415) );
  AND U7243 ( .A(n2432), .B(n2428), .Z(n7180) );
  OR U7244 ( .A(A[592]), .B(B[592]), .Z(n2432) );
  AND U7245 ( .A(n2423), .B(n2419), .Z(n7179) );
  NOR U7246 ( .A(n2381), .B(n2359), .Z(n7178) );
  NANDN U7247 ( .A(n2340), .B(n7181), .Z(n2334) );
  NAND U7248 ( .A(n7182), .B(n2341), .Z(n7181) );
  OR U7249 ( .A(B[607]), .B(A[607]), .Z(n2341) );
  NANDN U7250 ( .A(n2343), .B(n7183), .Z(n7182) );
  NAND U7251 ( .A(n7184), .B(n2345), .Z(n7183) );
  OR U7252 ( .A(A[606]), .B(B[606]), .Z(n2345) );
  NANDN U7253 ( .A(n2347), .B(n7185), .Z(n7184) );
  NAND U7254 ( .A(n7186), .B(n2350), .Z(n7185) );
  OR U7255 ( .A(A[605]), .B(B[605]), .Z(n2350) );
  NANDN U7256 ( .A(n2352), .B(n7187), .Z(n7186) );
  NAND U7257 ( .A(n7188), .B(n2355), .Z(n7187) );
  OR U7258 ( .A(A[604]), .B(B[604]), .Z(n2355) );
  NANDN U7259 ( .A(n2357), .B(n7189), .Z(n7188) );
  NANDN U7260 ( .A(n2359), .B(n7190), .Z(n7189) );
  NANDN U7261 ( .A(n2379), .B(n7191), .Z(n7190) );
  NANDN U7262 ( .A(n2381), .B(n2414), .Z(n7191) );
  NANDN U7263 ( .A(n2418), .B(n7192), .Z(n2414) );
  NAND U7264 ( .A(n7193), .B(n2419), .Z(n7192) );
  OR U7265 ( .A(B[595]), .B(A[595]), .Z(n2419) );
  NANDN U7266 ( .A(n2421), .B(n7194), .Z(n7193) );
  NAND U7267 ( .A(n7195), .B(n2423), .Z(n7194) );
  OR U7268 ( .A(A[594]), .B(B[594]), .Z(n2423) );
  NANDN U7269 ( .A(n2425), .B(n7196), .Z(n7195) );
  NAND U7270 ( .A(n2428), .B(n2430), .Z(n7196) );
  AND U7271 ( .A(A[592]), .B(B[592]), .Z(n2430) );
  OR U7272 ( .A(A[593]), .B(B[593]), .Z(n2428) );
  AND U7273 ( .A(A[593]), .B(B[593]), .Z(n2425) );
  AND U7274 ( .A(A[594]), .B(B[594]), .Z(n2421) );
  AND U7275 ( .A(B[595]), .B(A[595]), .Z(n2418) );
  NAND U7276 ( .A(n7197), .B(n7198), .Z(n2381) );
  AND U7277 ( .A(n2411), .B(n2407), .Z(n7198) );
  OR U7278 ( .A(A[596]), .B(B[596]), .Z(n2411) );
  AND U7279 ( .A(n2402), .B(n2398), .Z(n7197) );
  NANDN U7280 ( .A(n2397), .B(n7199), .Z(n2379) );
  NAND U7281 ( .A(n7200), .B(n2398), .Z(n7199) );
  OR U7282 ( .A(B[599]), .B(A[599]), .Z(n2398) );
  NANDN U7283 ( .A(n2400), .B(n7201), .Z(n7200) );
  NAND U7284 ( .A(n7202), .B(n2402), .Z(n7201) );
  OR U7285 ( .A(A[598]), .B(B[598]), .Z(n2402) );
  NANDN U7286 ( .A(n2404), .B(n7203), .Z(n7202) );
  NAND U7287 ( .A(n2407), .B(n2409), .Z(n7203) );
  AND U7288 ( .A(A[596]), .B(B[596]), .Z(n2409) );
  OR U7289 ( .A(A[597]), .B(B[597]), .Z(n2407) );
  AND U7290 ( .A(A[597]), .B(B[597]), .Z(n2404) );
  AND U7291 ( .A(A[598]), .B(B[598]), .Z(n2400) );
  AND U7292 ( .A(B[599]), .B(A[599]), .Z(n2397) );
  NAND U7293 ( .A(n7204), .B(n7205), .Z(n2359) );
  AND U7294 ( .A(n2377), .B(n2373), .Z(n7205) );
  OR U7295 ( .A(A[600]), .B(B[600]), .Z(n2377) );
  AND U7296 ( .A(n2368), .B(n2364), .Z(n7204) );
  NANDN U7297 ( .A(n2363), .B(n7206), .Z(n2357) );
  NAND U7298 ( .A(n7207), .B(n2364), .Z(n7206) );
  OR U7299 ( .A(B[603]), .B(A[603]), .Z(n2364) );
  NANDN U7300 ( .A(n2366), .B(n7208), .Z(n7207) );
  NAND U7301 ( .A(n7209), .B(n2368), .Z(n7208) );
  OR U7302 ( .A(A[602]), .B(B[602]), .Z(n2368) );
  NANDN U7303 ( .A(n2370), .B(n7210), .Z(n7209) );
  NAND U7304 ( .A(n2373), .B(n2375), .Z(n7210) );
  AND U7305 ( .A(A[600]), .B(B[600]), .Z(n2375) );
  OR U7306 ( .A(A[601]), .B(B[601]), .Z(n2373) );
  AND U7307 ( .A(A[601]), .B(B[601]), .Z(n2370) );
  AND U7308 ( .A(A[602]), .B(B[602]), .Z(n2366) );
  AND U7309 ( .A(B[603]), .B(A[603]), .Z(n2363) );
  AND U7310 ( .A(A[604]), .B(B[604]), .Z(n2352) );
  AND U7311 ( .A(A[605]), .B(B[605]), .Z(n2347) );
  AND U7312 ( .A(A[606]), .B(B[606]), .Z(n2343) );
  AND U7313 ( .A(B[607]), .B(A[607]), .Z(n2340) );
  NAND U7314 ( .A(n7211), .B(n7212), .Z(n2238) );
  AND U7315 ( .A(n7213), .B(n7214), .Z(n7212) );
  AND U7316 ( .A(n2257), .B(n2252), .Z(n7214) );
  AND U7317 ( .A(n2247), .B(n2243), .Z(n7213) );
  ANDN U7318 ( .B(n7215), .A(n2310), .Z(n7211) );
  NAND U7319 ( .A(n7216), .B(n7217), .Z(n2310) );
  AND U7320 ( .A(n2332), .B(n2323), .Z(n7217) );
  OR U7321 ( .A(A[608]), .B(B[608]), .Z(n2332) );
  AND U7322 ( .A(n2318), .B(n2314), .Z(n7216) );
  NOR U7323 ( .A(n2288), .B(n2261), .Z(n7215) );
  NANDN U7324 ( .A(n2242), .B(n7218), .Z(n2236) );
  NAND U7325 ( .A(n7219), .B(n2243), .Z(n7218) );
  OR U7326 ( .A(B[623]), .B(A[623]), .Z(n2243) );
  NANDN U7327 ( .A(n2245), .B(n7220), .Z(n7219) );
  NAND U7328 ( .A(n7221), .B(n2247), .Z(n7220) );
  OR U7329 ( .A(A[622]), .B(B[622]), .Z(n2247) );
  NANDN U7330 ( .A(n2249), .B(n7222), .Z(n7221) );
  NAND U7331 ( .A(n7223), .B(n2252), .Z(n7222) );
  OR U7332 ( .A(A[621]), .B(B[621]), .Z(n2252) );
  NANDN U7333 ( .A(n2254), .B(n7224), .Z(n7223) );
  NAND U7334 ( .A(n7225), .B(n2257), .Z(n7224) );
  OR U7335 ( .A(A[620]), .B(B[620]), .Z(n2257) );
  NANDN U7336 ( .A(n2259), .B(n7226), .Z(n7225) );
  NANDN U7337 ( .A(n2261), .B(n7227), .Z(n7226) );
  NANDN U7338 ( .A(n2286), .B(n7228), .Z(n7227) );
  NANDN U7339 ( .A(n2288), .B(n2309), .Z(n7228) );
  NANDN U7340 ( .A(n2313), .B(n7229), .Z(n2309) );
  NAND U7341 ( .A(n7230), .B(n2314), .Z(n7229) );
  OR U7342 ( .A(B[611]), .B(A[611]), .Z(n2314) );
  NANDN U7343 ( .A(n2316), .B(n7231), .Z(n7230) );
  NAND U7344 ( .A(n7232), .B(n2318), .Z(n7231) );
  OR U7345 ( .A(A[610]), .B(B[610]), .Z(n2318) );
  NANDN U7346 ( .A(n2320), .B(n7233), .Z(n7232) );
  NAND U7347 ( .A(n2323), .B(n2330), .Z(n7233) );
  AND U7348 ( .A(A[608]), .B(B[608]), .Z(n2330) );
  OR U7349 ( .A(A[609]), .B(B[609]), .Z(n2323) );
  AND U7350 ( .A(A[609]), .B(B[609]), .Z(n2320) );
  AND U7351 ( .A(A[610]), .B(B[610]), .Z(n2316) );
  AND U7352 ( .A(B[611]), .B(A[611]), .Z(n2313) );
  NAND U7353 ( .A(n7234), .B(n7235), .Z(n2288) );
  AND U7354 ( .A(n2306), .B(n2302), .Z(n7235) );
  OR U7355 ( .A(A[612]), .B(B[612]), .Z(n2306) );
  AND U7356 ( .A(n2297), .B(n2293), .Z(n7234) );
  NANDN U7357 ( .A(n2292), .B(n7236), .Z(n2286) );
  NAND U7358 ( .A(n7237), .B(n2293), .Z(n7236) );
  OR U7359 ( .A(B[615]), .B(A[615]), .Z(n2293) );
  NANDN U7360 ( .A(n2295), .B(n7238), .Z(n7237) );
  NAND U7361 ( .A(n7239), .B(n2297), .Z(n7238) );
  OR U7362 ( .A(A[614]), .B(B[614]), .Z(n2297) );
  NANDN U7363 ( .A(n2299), .B(n7240), .Z(n7239) );
  NAND U7364 ( .A(n2302), .B(n2304), .Z(n7240) );
  AND U7365 ( .A(A[612]), .B(B[612]), .Z(n2304) );
  OR U7366 ( .A(A[613]), .B(B[613]), .Z(n2302) );
  AND U7367 ( .A(A[613]), .B(B[613]), .Z(n2299) );
  AND U7368 ( .A(A[614]), .B(B[614]), .Z(n2295) );
  AND U7369 ( .A(B[615]), .B(A[615]), .Z(n2292) );
  NAND U7370 ( .A(n7241), .B(n7242), .Z(n2261) );
  AND U7371 ( .A(n2284), .B(n2280), .Z(n7242) );
  OR U7372 ( .A(A[616]), .B(B[616]), .Z(n2284) );
  AND U7373 ( .A(n2275), .B(n2271), .Z(n7241) );
  NANDN U7374 ( .A(n2270), .B(n7243), .Z(n2259) );
  NAND U7375 ( .A(n7244), .B(n2271), .Z(n7243) );
  OR U7376 ( .A(B[619]), .B(A[619]), .Z(n2271) );
  NANDN U7377 ( .A(n2273), .B(n7245), .Z(n7244) );
  NAND U7378 ( .A(n7246), .B(n2275), .Z(n7245) );
  OR U7379 ( .A(A[618]), .B(B[618]), .Z(n2275) );
  NANDN U7380 ( .A(n2277), .B(n7247), .Z(n7246) );
  NAND U7381 ( .A(n2280), .B(n2282), .Z(n7247) );
  AND U7382 ( .A(A[616]), .B(B[616]), .Z(n2282) );
  OR U7383 ( .A(A[617]), .B(B[617]), .Z(n2280) );
  AND U7384 ( .A(A[617]), .B(B[617]), .Z(n2277) );
  AND U7385 ( .A(A[618]), .B(B[618]), .Z(n2273) );
  AND U7386 ( .A(B[619]), .B(A[619]), .Z(n2270) );
  AND U7387 ( .A(A[620]), .B(B[620]), .Z(n2254) );
  AND U7388 ( .A(A[621]), .B(B[621]), .Z(n2249) );
  AND U7389 ( .A(A[622]), .B(B[622]), .Z(n2245) );
  AND U7390 ( .A(B[623]), .B(A[623]), .Z(n2242) );
  NAND U7391 ( .A(n7248), .B(n7249), .Z(n7104) );
  AND U7392 ( .A(n7250), .B(n7251), .Z(n7249) );
  AND U7393 ( .A(n2163), .B(n2158), .Z(n7251) );
  OR U7394 ( .A(A[637]), .B(B[637]), .Z(n2158) );
  OR U7395 ( .A(A[636]), .B(B[636]), .Z(n2163) );
  AND U7396 ( .A(n2153), .B(n2149), .Z(n7250) );
  OR U7397 ( .A(B[639]), .B(A[639]), .Z(n2149) );
  OR U7398 ( .A(A[638]), .B(B[638]), .Z(n2153) );
  ANDN U7399 ( .B(n7252), .A(n2189), .Z(n7248) );
  NAND U7400 ( .A(n7253), .B(n7254), .Z(n2189) );
  AND U7401 ( .A(n2212), .B(n2203), .Z(n7254) );
  OR U7402 ( .A(A[629]), .B(B[629]), .Z(n2203) );
  OR U7403 ( .A(A[628]), .B(B[628]), .Z(n2212) );
  AND U7404 ( .A(n2198), .B(n2194), .Z(n7253) );
  OR U7405 ( .A(B[631]), .B(A[631]), .Z(n2194) );
  OR U7406 ( .A(A[630]), .B(B[630]), .Z(n2198) );
  NOR U7407 ( .A(n2216), .B(n2167), .Z(n7252) );
  NAND U7408 ( .A(n7255), .B(n7256), .Z(n2167) );
  AND U7409 ( .A(n2185), .B(n2181), .Z(n7256) );
  OR U7410 ( .A(A[633]), .B(B[633]), .Z(n2181) );
  OR U7411 ( .A(A[632]), .B(B[632]), .Z(n2185) );
  AND U7412 ( .A(n2176), .B(n2172), .Z(n7255) );
  OR U7413 ( .A(B[635]), .B(A[635]), .Z(n2172) );
  OR U7414 ( .A(A[634]), .B(B[634]), .Z(n2176) );
  NAND U7415 ( .A(n7257), .B(n7258), .Z(n2216) );
  AND U7416 ( .A(n2234), .B(n2230), .Z(n7258) );
  OR U7417 ( .A(A[625]), .B(B[625]), .Z(n2230) );
  OR U7418 ( .A(A[624]), .B(B[624]), .Z(n2234) );
  AND U7419 ( .A(n2225), .B(n2221), .Z(n7257) );
  OR U7420 ( .A(B[627]), .B(A[627]), .Z(n2221) );
  OR U7421 ( .A(A[626]), .B(B[626]), .Z(n2225) );
  NAND U7422 ( .A(n7259), .B(n7260), .Z(n1754) );
  ANDN U7423 ( .B(n1855), .A(n1951), .Z(n7260) );
  NOR U7424 ( .A(n2048), .B(n7261), .Z(n7259) );
  NAND U7425 ( .A(n7262), .B(n7263), .Z(n2048) );
  AND U7426 ( .A(n7264), .B(n7265), .Z(n7263) );
  AND U7427 ( .A(n2066), .B(n2061), .Z(n7265) );
  AND U7428 ( .A(n2056), .B(n2052), .Z(n7264) );
  ANDN U7429 ( .B(n7266), .A(n2115), .Z(n7262) );
  NAND U7430 ( .A(n7267), .B(n7268), .Z(n2115) );
  AND U7431 ( .A(n2132), .B(n2128), .Z(n7268) );
  OR U7432 ( .A(B[640]), .B(A[640]), .Z(n2132) );
  AND U7433 ( .A(n2123), .B(n2119), .Z(n7267) );
  ANDN U7434 ( .B(n2070), .A(n2093), .Z(n7266) );
  NAND U7435 ( .A(n7269), .B(n7270), .Z(n1752) );
  NAND U7436 ( .A(n7271), .B(n1759), .Z(n7270) );
  NANDN U7437 ( .A(n1761), .B(n7272), .Z(n7271) );
  NAND U7438 ( .A(n7273), .B(n1763), .Z(n7272) );
  NANDN U7439 ( .A(n1765), .B(n7274), .Z(n7273) );
  NAND U7440 ( .A(n7275), .B(n1768), .Z(n7274) );
  NANDN U7441 ( .A(n1770), .B(n7276), .Z(n7275) );
  NAND U7442 ( .A(n7277), .B(n1773), .Z(n7276) );
  NANDN U7443 ( .A(n1775), .B(n7278), .Z(n7277) );
  NANDN U7444 ( .A(n1777), .B(n7279), .Z(n7278) );
  NANDN U7445 ( .A(n1804), .B(n7280), .Z(n7279) );
  NANDN U7446 ( .A(n1806), .B(n1827), .Z(n7280) );
  NANDN U7447 ( .A(n1832), .B(n7281), .Z(n1827) );
  NAND U7448 ( .A(n7282), .B(n1833), .Z(n7281) );
  NANDN U7449 ( .A(n1835), .B(n7283), .Z(n7282) );
  NAND U7450 ( .A(n7284), .B(n1837), .Z(n7283) );
  NANDN U7451 ( .A(n1839), .B(n7285), .Z(n7284) );
  NAND U7452 ( .A(n1842), .B(n1849), .Z(n7285) );
  AND U7453 ( .A(A[688]), .B(B[688]), .Z(n1849) );
  AND U7454 ( .A(A[689]), .B(B[689]), .Z(n1839) );
  AND U7455 ( .A(A[690]), .B(B[690]), .Z(n1835) );
  AND U7456 ( .A(B[691]), .B(A[691]), .Z(n1832) );
  NANDN U7457 ( .A(n1810), .B(n7286), .Z(n1804) );
  NAND U7458 ( .A(n7287), .B(n1811), .Z(n7286) );
  NANDN U7459 ( .A(n1813), .B(n7288), .Z(n7287) );
  NAND U7460 ( .A(n7289), .B(n1815), .Z(n7288) );
  NANDN U7461 ( .A(n1817), .B(n7290), .Z(n7289) );
  NAND U7462 ( .A(n1820), .B(n1822), .Z(n7290) );
  AND U7463 ( .A(A[692]), .B(B[692]), .Z(n1822) );
  AND U7464 ( .A(A[693]), .B(B[693]), .Z(n1817) );
  AND U7465 ( .A(A[694]), .B(B[694]), .Z(n1813) );
  AND U7466 ( .A(B[695]), .B(A[695]), .Z(n1810) );
  NANDN U7467 ( .A(n1788), .B(n7291), .Z(n1775) );
  NAND U7468 ( .A(n7292), .B(n1789), .Z(n7291) );
  NANDN U7469 ( .A(n1791), .B(n7293), .Z(n7292) );
  NAND U7470 ( .A(n7294), .B(n1793), .Z(n7293) );
  NANDN U7471 ( .A(n1795), .B(n7295), .Z(n7294) );
  NAND U7472 ( .A(n1798), .B(n1800), .Z(n7295) );
  AND U7473 ( .A(A[696]), .B(B[696]), .Z(n1800) );
  AND U7474 ( .A(A[697]), .B(B[697]), .Z(n1795) );
  AND U7475 ( .A(A[698]), .B(B[698]), .Z(n1791) );
  AND U7476 ( .A(B[699]), .B(A[699]), .Z(n1788) );
  AND U7477 ( .A(A[700]), .B(B[700]), .Z(n1770) );
  AND U7478 ( .A(A[701]), .B(B[701]), .Z(n1765) );
  AND U7479 ( .A(A[702]), .B(B[702]), .Z(n1761) );
  ANDN U7480 ( .B(n7296), .A(n1758), .Z(n7269) );
  AND U7481 ( .A(B[703]), .B(A[703]), .Z(n1758) );
  NANDN U7482 ( .A(n7261), .B(n7297), .Z(n7296) );
  NANDN U7483 ( .A(n1853), .B(n7298), .Z(n7297) );
  NAND U7484 ( .A(n7299), .B(n1855), .Z(n7298) );
  AND U7485 ( .A(n7300), .B(n7301), .Z(n1855) );
  AND U7486 ( .A(n7302), .B(n7303), .Z(n7301) );
  AND U7487 ( .A(n1874), .B(n1869), .Z(n7303) );
  AND U7488 ( .A(n1864), .B(n1860), .Z(n7302) );
  ANDN U7489 ( .B(n7304), .A(n1930), .Z(n7300) );
  NAND U7490 ( .A(n7305), .B(n7306), .Z(n1930) );
  AND U7491 ( .A(n1947), .B(n1943), .Z(n7306) );
  OR U7492 ( .A(B[672]), .B(A[672]), .Z(n1947) );
  AND U7493 ( .A(n1938), .B(n1934), .Z(n7305) );
  ANDN U7494 ( .B(n1878), .A(n1900), .Z(n7304) );
  NANDN U7495 ( .A(n1949), .B(n7307), .Z(n7299) );
  NANDN U7496 ( .A(n1951), .B(n2047), .Z(n7307) );
  NANDN U7497 ( .A(n2051), .B(n7308), .Z(n2047) );
  NAND U7498 ( .A(n7309), .B(n2052), .Z(n7308) );
  OR U7499 ( .A(B[655]), .B(A[655]), .Z(n2052) );
  NANDN U7500 ( .A(n2054), .B(n7310), .Z(n7309) );
  NAND U7501 ( .A(n7311), .B(n2056), .Z(n7310) );
  OR U7502 ( .A(B[654]), .B(A[654]), .Z(n2056) );
  NANDN U7503 ( .A(n2058), .B(n7312), .Z(n7311) );
  NAND U7504 ( .A(n7313), .B(n2061), .Z(n7312) );
  OR U7505 ( .A(B[653]), .B(A[653]), .Z(n2061) );
  NANDN U7506 ( .A(n2063), .B(n7314), .Z(n7313) );
  NAND U7507 ( .A(n7315), .B(n2066), .Z(n7314) );
  OR U7508 ( .A(B[652]), .B(A[652]), .Z(n2066) );
  NANDN U7509 ( .A(n2068), .B(n7316), .Z(n7315) );
  NAND U7510 ( .A(n7317), .B(n2070), .Z(n7316) );
  AND U7511 ( .A(n7318), .B(n7319), .Z(n2070) );
  AND U7512 ( .A(n2089), .B(n2084), .Z(n7319) );
  OR U7513 ( .A(B[648]), .B(A[648]), .Z(n2089) );
  AND U7514 ( .A(n2079), .B(n2075), .Z(n7318) );
  NANDN U7515 ( .A(n2091), .B(n7320), .Z(n7317) );
  NANDN U7516 ( .A(n2093), .B(n2114), .Z(n7320) );
  NANDN U7517 ( .A(n2118), .B(n7321), .Z(n2114) );
  NAND U7518 ( .A(n7322), .B(n2119), .Z(n7321) );
  OR U7519 ( .A(B[643]), .B(A[643]), .Z(n2119) );
  NANDN U7520 ( .A(n2121), .B(n7323), .Z(n7322) );
  NAND U7521 ( .A(n7324), .B(n2123), .Z(n7323) );
  OR U7522 ( .A(B[642]), .B(A[642]), .Z(n2123) );
  NANDN U7523 ( .A(n2125), .B(n7325), .Z(n7324) );
  NAND U7524 ( .A(n2128), .B(n2130), .Z(n7325) );
  AND U7525 ( .A(B[640]), .B(A[640]), .Z(n2130) );
  OR U7526 ( .A(B[641]), .B(A[641]), .Z(n2128) );
  AND U7527 ( .A(B[641]), .B(A[641]), .Z(n2125) );
  AND U7528 ( .A(B[642]), .B(A[642]), .Z(n2121) );
  AND U7529 ( .A(B[643]), .B(A[643]), .Z(n2118) );
  NAND U7530 ( .A(n7326), .B(n7327), .Z(n2093) );
  AND U7531 ( .A(n2111), .B(n2107), .Z(n7327) );
  OR U7532 ( .A(B[644]), .B(A[644]), .Z(n2111) );
  AND U7533 ( .A(n2102), .B(n2098), .Z(n7326) );
  NANDN U7534 ( .A(n2097), .B(n7328), .Z(n2091) );
  NAND U7535 ( .A(n7329), .B(n2098), .Z(n7328) );
  OR U7536 ( .A(B[647]), .B(A[647]), .Z(n2098) );
  NANDN U7537 ( .A(n2100), .B(n7330), .Z(n7329) );
  NAND U7538 ( .A(n7331), .B(n2102), .Z(n7330) );
  OR U7539 ( .A(B[646]), .B(A[646]), .Z(n2102) );
  NANDN U7540 ( .A(n2104), .B(n7332), .Z(n7331) );
  NAND U7541 ( .A(n2107), .B(n2109), .Z(n7332) );
  AND U7542 ( .A(B[644]), .B(A[644]), .Z(n2109) );
  OR U7543 ( .A(B[645]), .B(A[645]), .Z(n2107) );
  AND U7544 ( .A(B[645]), .B(A[645]), .Z(n2104) );
  AND U7545 ( .A(B[646]), .B(A[646]), .Z(n2100) );
  AND U7546 ( .A(B[647]), .B(A[647]), .Z(n2097) );
  NANDN U7547 ( .A(n2074), .B(n7333), .Z(n2068) );
  NAND U7548 ( .A(n7334), .B(n2075), .Z(n7333) );
  OR U7549 ( .A(B[651]), .B(A[651]), .Z(n2075) );
  NANDN U7550 ( .A(n2077), .B(n7335), .Z(n7334) );
  NAND U7551 ( .A(n7336), .B(n2079), .Z(n7335) );
  OR U7552 ( .A(B[650]), .B(A[650]), .Z(n2079) );
  NANDN U7553 ( .A(n2081), .B(n7337), .Z(n7336) );
  NAND U7554 ( .A(n2084), .B(n2087), .Z(n7337) );
  AND U7555 ( .A(B[648]), .B(A[648]), .Z(n2087) );
  OR U7556 ( .A(B[649]), .B(A[649]), .Z(n2084) );
  AND U7557 ( .A(B[649]), .B(A[649]), .Z(n2081) );
  AND U7558 ( .A(B[650]), .B(A[650]), .Z(n2077) );
  AND U7559 ( .A(B[651]), .B(A[651]), .Z(n2074) );
  AND U7560 ( .A(B[652]), .B(A[652]), .Z(n2063) );
  AND U7561 ( .A(B[653]), .B(A[653]), .Z(n2058) );
  AND U7562 ( .A(B[654]), .B(A[654]), .Z(n2054) );
  AND U7563 ( .A(B[655]), .B(A[655]), .Z(n2051) );
  NAND U7564 ( .A(n7338), .B(n7339), .Z(n1951) );
  AND U7565 ( .A(n7340), .B(n7341), .Z(n7339) );
  AND U7566 ( .A(n1975), .B(n1965), .Z(n7341) );
  AND U7567 ( .A(n1960), .B(n1956), .Z(n7340) );
  ANDN U7568 ( .B(n7342), .A(n2023), .Z(n7338) );
  NAND U7569 ( .A(n7343), .B(n7344), .Z(n2023) );
  AND U7570 ( .A(n2044), .B(n2040), .Z(n7344) );
  OR U7571 ( .A(B[656]), .B(A[656]), .Z(n2044) );
  AND U7572 ( .A(n2035), .B(n2031), .Z(n7343) );
  ANDN U7573 ( .B(n1979), .A(n2001), .Z(n7342) );
  NANDN U7574 ( .A(n1955), .B(n7345), .Z(n1949) );
  NAND U7575 ( .A(n7346), .B(n1956), .Z(n7345) );
  OR U7576 ( .A(B[671]), .B(A[671]), .Z(n1956) );
  NANDN U7577 ( .A(n1958), .B(n7347), .Z(n7346) );
  NAND U7578 ( .A(n7348), .B(n1960), .Z(n7347) );
  OR U7579 ( .A(B[670]), .B(A[670]), .Z(n1960) );
  NANDN U7580 ( .A(n1962), .B(n7349), .Z(n7348) );
  NAND U7581 ( .A(n7350), .B(n1965), .Z(n7349) );
  OR U7582 ( .A(B[669]), .B(A[669]), .Z(n1965) );
  NANDN U7583 ( .A(n1972), .B(n7351), .Z(n7350) );
  NAND U7584 ( .A(n7352), .B(n1975), .Z(n7351) );
  OR U7585 ( .A(B[668]), .B(A[668]), .Z(n1975) );
  NANDN U7586 ( .A(n1977), .B(n7353), .Z(n7352) );
  NAND U7587 ( .A(n7354), .B(n1979), .Z(n7353) );
  AND U7588 ( .A(n7355), .B(n7356), .Z(n1979) );
  AND U7589 ( .A(n1997), .B(n1993), .Z(n7356) );
  OR U7590 ( .A(B[664]), .B(A[664]), .Z(n1997) );
  AND U7591 ( .A(n1988), .B(n1984), .Z(n7355) );
  NANDN U7592 ( .A(n1999), .B(n7357), .Z(n7354) );
  NANDN U7593 ( .A(n2001), .B(n2022), .Z(n7357) );
  NANDN U7594 ( .A(n2030), .B(n7358), .Z(n2022) );
  NAND U7595 ( .A(n7359), .B(n2031), .Z(n7358) );
  OR U7596 ( .A(B[659]), .B(A[659]), .Z(n2031) );
  NANDN U7597 ( .A(n2033), .B(n7360), .Z(n7359) );
  NAND U7598 ( .A(n7361), .B(n2035), .Z(n7360) );
  OR U7599 ( .A(B[658]), .B(A[658]), .Z(n2035) );
  NANDN U7600 ( .A(n2037), .B(n7362), .Z(n7361) );
  NAND U7601 ( .A(n2040), .B(n2042), .Z(n7362) );
  AND U7602 ( .A(B[656]), .B(A[656]), .Z(n2042) );
  OR U7603 ( .A(B[657]), .B(A[657]), .Z(n2040) );
  AND U7604 ( .A(B[657]), .B(A[657]), .Z(n2037) );
  AND U7605 ( .A(B[658]), .B(A[658]), .Z(n2033) );
  AND U7606 ( .A(B[659]), .B(A[659]), .Z(n2030) );
  NAND U7607 ( .A(n7363), .B(n7364), .Z(n2001) );
  AND U7608 ( .A(n2019), .B(n2015), .Z(n7364) );
  OR U7609 ( .A(B[660]), .B(A[660]), .Z(n2019) );
  AND U7610 ( .A(n2010), .B(n2006), .Z(n7363) );
  NANDN U7611 ( .A(n2005), .B(n7365), .Z(n1999) );
  NAND U7612 ( .A(n7366), .B(n2006), .Z(n7365) );
  OR U7613 ( .A(B[663]), .B(A[663]), .Z(n2006) );
  NANDN U7614 ( .A(n2008), .B(n7367), .Z(n7366) );
  NAND U7615 ( .A(n7368), .B(n2010), .Z(n7367) );
  OR U7616 ( .A(B[662]), .B(A[662]), .Z(n2010) );
  NANDN U7617 ( .A(n2012), .B(n7369), .Z(n7368) );
  NAND U7618 ( .A(n2015), .B(n2017), .Z(n7369) );
  AND U7619 ( .A(B[660]), .B(A[660]), .Z(n2017) );
  OR U7620 ( .A(B[661]), .B(A[661]), .Z(n2015) );
  AND U7621 ( .A(B[661]), .B(A[661]), .Z(n2012) );
  AND U7622 ( .A(B[662]), .B(A[662]), .Z(n2008) );
  AND U7623 ( .A(B[663]), .B(A[663]), .Z(n2005) );
  NANDN U7624 ( .A(n1983), .B(n7370), .Z(n1977) );
  NAND U7625 ( .A(n7371), .B(n1984), .Z(n7370) );
  OR U7626 ( .A(B[667]), .B(A[667]), .Z(n1984) );
  NANDN U7627 ( .A(n1986), .B(n7372), .Z(n7371) );
  NAND U7628 ( .A(n7373), .B(n1988), .Z(n7372) );
  OR U7629 ( .A(B[666]), .B(A[666]), .Z(n1988) );
  NANDN U7630 ( .A(n1990), .B(n7374), .Z(n7373) );
  NAND U7631 ( .A(n1993), .B(n1995), .Z(n7374) );
  AND U7632 ( .A(B[664]), .B(A[664]), .Z(n1995) );
  OR U7633 ( .A(B[665]), .B(A[665]), .Z(n1993) );
  AND U7634 ( .A(B[665]), .B(A[665]), .Z(n1990) );
  AND U7635 ( .A(B[666]), .B(A[666]), .Z(n1986) );
  AND U7636 ( .A(B[667]), .B(A[667]), .Z(n1983) );
  AND U7637 ( .A(B[668]), .B(A[668]), .Z(n1972) );
  AND U7638 ( .A(B[669]), .B(A[669]), .Z(n1962) );
  AND U7639 ( .A(B[670]), .B(A[670]), .Z(n1958) );
  AND U7640 ( .A(B[671]), .B(A[671]), .Z(n1955) );
  NANDN U7641 ( .A(n1859), .B(n7375), .Z(n1853) );
  NAND U7642 ( .A(n7376), .B(n1860), .Z(n7375) );
  OR U7643 ( .A(B[687]), .B(A[687]), .Z(n1860) );
  NANDN U7644 ( .A(n1862), .B(n7377), .Z(n7376) );
  NAND U7645 ( .A(n7378), .B(n1864), .Z(n7377) );
  OR U7646 ( .A(B[686]), .B(A[686]), .Z(n1864) );
  NANDN U7647 ( .A(n1866), .B(n7379), .Z(n7378) );
  NAND U7648 ( .A(n7380), .B(n1869), .Z(n7379) );
  OR U7649 ( .A(B[685]), .B(A[685]), .Z(n1869) );
  NANDN U7650 ( .A(n1871), .B(n7381), .Z(n7380) );
  NAND U7651 ( .A(n7382), .B(n1874), .Z(n7381) );
  OR U7652 ( .A(B[684]), .B(A[684]), .Z(n1874) );
  NANDN U7653 ( .A(n1876), .B(n7383), .Z(n7382) );
  NAND U7654 ( .A(n7384), .B(n1878), .Z(n7383) );
  AND U7655 ( .A(n7385), .B(n7386), .Z(n1878) );
  AND U7656 ( .A(n1896), .B(n1892), .Z(n7386) );
  OR U7657 ( .A(B[680]), .B(A[680]), .Z(n1896) );
  AND U7658 ( .A(n1887), .B(n1883), .Z(n7385) );
  NANDN U7659 ( .A(n1898), .B(n7387), .Z(n7384) );
  NANDN U7660 ( .A(n1900), .B(n1929), .Z(n7387) );
  NANDN U7661 ( .A(n1933), .B(n7388), .Z(n1929) );
  NAND U7662 ( .A(n7389), .B(n1934), .Z(n7388) );
  OR U7663 ( .A(B[675]), .B(A[675]), .Z(n1934) );
  NANDN U7664 ( .A(n1936), .B(n7390), .Z(n7389) );
  NAND U7665 ( .A(n7391), .B(n1938), .Z(n7390) );
  OR U7666 ( .A(B[674]), .B(A[674]), .Z(n1938) );
  NANDN U7667 ( .A(n1940), .B(n7392), .Z(n7391) );
  NAND U7668 ( .A(n1943), .B(n1945), .Z(n7392) );
  AND U7669 ( .A(B[672]), .B(A[672]), .Z(n1945) );
  OR U7670 ( .A(B[673]), .B(A[673]), .Z(n1943) );
  AND U7671 ( .A(B[673]), .B(A[673]), .Z(n1940) );
  AND U7672 ( .A(B[674]), .B(A[674]), .Z(n1936) );
  AND U7673 ( .A(B[675]), .B(A[675]), .Z(n1933) );
  NAND U7674 ( .A(n7393), .B(n7394), .Z(n1900) );
  AND U7675 ( .A(n1926), .B(n1922), .Z(n7394) );
  OR U7676 ( .A(B[676]), .B(A[676]), .Z(n1926) );
  AND U7677 ( .A(n1917), .B(n1913), .Z(n7393) );
  NANDN U7678 ( .A(n1912), .B(n7395), .Z(n1898) );
  NAND U7679 ( .A(n7396), .B(n1913), .Z(n7395) );
  OR U7680 ( .A(B[679]), .B(A[679]), .Z(n1913) );
  NANDN U7681 ( .A(n1915), .B(n7397), .Z(n7396) );
  NAND U7682 ( .A(n7398), .B(n1917), .Z(n7397) );
  OR U7683 ( .A(B[678]), .B(A[678]), .Z(n1917) );
  NANDN U7684 ( .A(n1919), .B(n7399), .Z(n7398) );
  NAND U7685 ( .A(n1922), .B(n1924), .Z(n7399) );
  AND U7686 ( .A(B[676]), .B(A[676]), .Z(n1924) );
  OR U7687 ( .A(B[677]), .B(A[677]), .Z(n1922) );
  AND U7688 ( .A(B[677]), .B(A[677]), .Z(n1919) );
  AND U7689 ( .A(B[678]), .B(A[678]), .Z(n1915) );
  AND U7690 ( .A(B[679]), .B(A[679]), .Z(n1912) );
  NANDN U7691 ( .A(n1882), .B(n7400), .Z(n1876) );
  NAND U7692 ( .A(n7401), .B(n1883), .Z(n7400) );
  OR U7693 ( .A(B[683]), .B(A[683]), .Z(n1883) );
  NANDN U7694 ( .A(n1885), .B(n7402), .Z(n7401) );
  NAND U7695 ( .A(n7403), .B(n1887), .Z(n7402) );
  OR U7696 ( .A(B[682]), .B(A[682]), .Z(n1887) );
  NANDN U7697 ( .A(n1889), .B(n7404), .Z(n7403) );
  NAND U7698 ( .A(n1892), .B(n1894), .Z(n7404) );
  AND U7699 ( .A(B[680]), .B(A[680]), .Z(n1894) );
  OR U7700 ( .A(B[681]), .B(A[681]), .Z(n1892) );
  AND U7701 ( .A(B[681]), .B(A[681]), .Z(n1889) );
  AND U7702 ( .A(B[682]), .B(A[682]), .Z(n1885) );
  AND U7703 ( .A(B[683]), .B(A[683]), .Z(n1882) );
  AND U7704 ( .A(B[684]), .B(A[684]), .Z(n1871) );
  AND U7705 ( .A(B[685]), .B(A[685]), .Z(n1866) );
  AND U7706 ( .A(B[686]), .B(A[686]), .Z(n1862) );
  AND U7707 ( .A(B[687]), .B(A[687]), .Z(n1859) );
  NAND U7708 ( .A(n7405), .B(n7406), .Z(n7261) );
  AND U7709 ( .A(n7407), .B(n7408), .Z(n7406) );
  AND U7710 ( .A(n1773), .B(n1768), .Z(n7408) );
  OR U7711 ( .A(A[701]), .B(B[701]), .Z(n1768) );
  OR U7712 ( .A(A[700]), .B(B[700]), .Z(n1773) );
  AND U7713 ( .A(n1763), .B(n1759), .Z(n7407) );
  OR U7714 ( .A(B[703]), .B(A[703]), .Z(n1759) );
  OR U7715 ( .A(A[702]), .B(B[702]), .Z(n1763) );
  ANDN U7716 ( .B(n7409), .A(n1806), .Z(n7405) );
  NAND U7717 ( .A(n7410), .B(n7411), .Z(n1806) );
  AND U7718 ( .A(n1824), .B(n1820), .Z(n7411) );
  OR U7719 ( .A(A[693]), .B(B[693]), .Z(n1820) );
  OR U7720 ( .A(A[692]), .B(B[692]), .Z(n1824) );
  AND U7721 ( .A(n1815), .B(n1811), .Z(n7410) );
  OR U7722 ( .A(B[695]), .B(A[695]), .Z(n1811) );
  OR U7723 ( .A(A[694]), .B(B[694]), .Z(n1815) );
  NOR U7724 ( .A(n1828), .B(n1777), .Z(n7409) );
  NAND U7725 ( .A(n7412), .B(n7413), .Z(n1777) );
  AND U7726 ( .A(n1802), .B(n1798), .Z(n7413) );
  OR U7727 ( .A(A[697]), .B(B[697]), .Z(n1798) );
  OR U7728 ( .A(A[696]), .B(B[696]), .Z(n1802) );
  AND U7729 ( .A(n1793), .B(n1789), .Z(n7412) );
  OR U7730 ( .A(B[699]), .B(A[699]), .Z(n1789) );
  OR U7731 ( .A(A[698]), .B(B[698]), .Z(n1793) );
  NAND U7732 ( .A(n7414), .B(n7415), .Z(n1828) );
  AND U7733 ( .A(n1851), .B(n1842), .Z(n7415) );
  OR U7734 ( .A(A[689]), .B(B[689]), .Z(n1842) );
  OR U7735 ( .A(A[688]), .B(B[688]), .Z(n1851) );
  AND U7736 ( .A(n1837), .B(n1833), .Z(n7414) );
  OR U7737 ( .A(B[691]), .B(A[691]), .Z(n1833) );
  OR U7738 ( .A(A[690]), .B(B[690]), .Z(n1837) );
  NAND U7739 ( .A(n7416), .B(n7417), .Z(n1653) );
  AND U7740 ( .A(n7418), .B(n7419), .Z(n7417) );
  AND U7741 ( .A(n1680), .B(n1675), .Z(n7419) );
  AND U7742 ( .A(n1670), .B(n1666), .Z(n7418) );
  ANDN U7743 ( .B(n7420), .A(n1733), .Z(n7416) );
  NAND U7744 ( .A(n7421), .B(n7422), .Z(n1733) );
  AND U7745 ( .A(n1750), .B(n1746), .Z(n7422) );
  OR U7746 ( .A(B[704]), .B(A[704]), .Z(n1750) );
  AND U7747 ( .A(n1741), .B(n1737), .Z(n7421) );
  ANDN U7748 ( .B(n1684), .A(n1706), .Z(n7420) );
  NANDN U7749 ( .A(n1665), .B(n7423), .Z(n1651) );
  NAND U7750 ( .A(n7424), .B(n1666), .Z(n7423) );
  OR U7751 ( .A(B[719]), .B(A[719]), .Z(n1666) );
  NANDN U7752 ( .A(n1668), .B(n7425), .Z(n7424) );
  NAND U7753 ( .A(n7426), .B(n1670), .Z(n7425) );
  OR U7754 ( .A(B[718]), .B(A[718]), .Z(n1670) );
  NANDN U7755 ( .A(n1672), .B(n7427), .Z(n7426) );
  NAND U7756 ( .A(n7428), .B(n1675), .Z(n7427) );
  OR U7757 ( .A(B[717]), .B(A[717]), .Z(n1675) );
  NANDN U7758 ( .A(n1677), .B(n7429), .Z(n7428) );
  NAND U7759 ( .A(n7430), .B(n1680), .Z(n7429) );
  OR U7760 ( .A(B[716]), .B(A[716]), .Z(n1680) );
  NANDN U7761 ( .A(n1682), .B(n7431), .Z(n7430) );
  NAND U7762 ( .A(n7432), .B(n1684), .Z(n7431) );
  AND U7763 ( .A(n7433), .B(n7434), .Z(n1684) );
  AND U7764 ( .A(n1702), .B(n1698), .Z(n7434) );
  OR U7765 ( .A(B[712]), .B(A[712]), .Z(n1702) );
  AND U7766 ( .A(n1693), .B(n1689), .Z(n7433) );
  NANDN U7767 ( .A(n1704), .B(n7435), .Z(n7432) );
  NANDN U7768 ( .A(n1706), .B(n1732), .Z(n7435) );
  NANDN U7769 ( .A(n1736), .B(n7436), .Z(n1732) );
  NAND U7770 ( .A(n7437), .B(n1737), .Z(n7436) );
  OR U7771 ( .A(B[707]), .B(A[707]), .Z(n1737) );
  NANDN U7772 ( .A(n1739), .B(n7438), .Z(n7437) );
  NAND U7773 ( .A(n7439), .B(n1741), .Z(n7438) );
  OR U7774 ( .A(B[706]), .B(A[706]), .Z(n1741) );
  NANDN U7775 ( .A(n1743), .B(n7440), .Z(n7439) );
  NAND U7776 ( .A(n1746), .B(n1748), .Z(n7440) );
  AND U7777 ( .A(B[704]), .B(A[704]), .Z(n1748) );
  OR U7778 ( .A(B[705]), .B(A[705]), .Z(n1746) );
  AND U7779 ( .A(B[705]), .B(A[705]), .Z(n1743) );
  AND U7780 ( .A(B[706]), .B(A[706]), .Z(n1739) );
  AND U7781 ( .A(B[707]), .B(A[707]), .Z(n1736) );
  NAND U7782 ( .A(n7441), .B(n7442), .Z(n1706) );
  AND U7783 ( .A(n1729), .B(n1720), .Z(n7442) );
  OR U7784 ( .A(B[708]), .B(A[708]), .Z(n1729) );
  AND U7785 ( .A(n1715), .B(n1711), .Z(n7441) );
  NANDN U7786 ( .A(n1710), .B(n7443), .Z(n1704) );
  NAND U7787 ( .A(n7444), .B(n1711), .Z(n7443) );
  OR U7788 ( .A(B[711]), .B(A[711]), .Z(n1711) );
  NANDN U7789 ( .A(n1713), .B(n7445), .Z(n7444) );
  NAND U7790 ( .A(n7446), .B(n1715), .Z(n7445) );
  OR U7791 ( .A(B[710]), .B(A[710]), .Z(n1715) );
  NANDN U7792 ( .A(n1717), .B(n7447), .Z(n7446) );
  NAND U7793 ( .A(n1720), .B(n1727), .Z(n7447) );
  AND U7794 ( .A(B[708]), .B(A[708]), .Z(n1727) );
  OR U7795 ( .A(B[709]), .B(A[709]), .Z(n1720) );
  AND U7796 ( .A(B[709]), .B(A[709]), .Z(n1717) );
  AND U7797 ( .A(B[710]), .B(A[710]), .Z(n1713) );
  AND U7798 ( .A(B[711]), .B(A[711]), .Z(n1710) );
  NANDN U7799 ( .A(n1688), .B(n7448), .Z(n1682) );
  NAND U7800 ( .A(n7449), .B(n1689), .Z(n7448) );
  OR U7801 ( .A(B[715]), .B(A[715]), .Z(n1689) );
  NANDN U7802 ( .A(n1691), .B(n7450), .Z(n7449) );
  NAND U7803 ( .A(n7451), .B(n1693), .Z(n7450) );
  OR U7804 ( .A(B[714]), .B(A[714]), .Z(n1693) );
  NANDN U7805 ( .A(n1695), .B(n7452), .Z(n7451) );
  NAND U7806 ( .A(n1698), .B(n1700), .Z(n7452) );
  AND U7807 ( .A(B[712]), .B(A[712]), .Z(n1700) );
  OR U7808 ( .A(B[713]), .B(A[713]), .Z(n1698) );
  AND U7809 ( .A(B[713]), .B(A[713]), .Z(n1695) );
  AND U7810 ( .A(B[714]), .B(A[714]), .Z(n1691) );
  AND U7811 ( .A(B[715]), .B(A[715]), .Z(n1688) );
  AND U7812 ( .A(B[716]), .B(A[716]), .Z(n1677) );
  AND U7813 ( .A(B[717]), .B(A[717]), .Z(n1672) );
  AND U7814 ( .A(B[718]), .B(A[718]), .Z(n1668) );
  AND U7815 ( .A(B[719]), .B(A[719]), .Z(n1665) );
  NAND U7816 ( .A(n7453), .B(n7454), .Z(n1560) );
  AND U7817 ( .A(n7455), .B(n7456), .Z(n7454) );
  AND U7818 ( .A(n1579), .B(n1574), .Z(n7456) );
  AND U7819 ( .A(n1569), .B(n1565), .Z(n7455) );
  ANDN U7820 ( .B(n7457), .A(n1632), .Z(n7453) );
  NAND U7821 ( .A(n7458), .B(n7459), .Z(n1632) );
  AND U7822 ( .A(n1649), .B(n1645), .Z(n7459) );
  OR U7823 ( .A(B[720]), .B(A[720]), .Z(n1649) );
  AND U7824 ( .A(n1640), .B(n1636), .Z(n7458) );
  ANDN U7825 ( .B(n1583), .A(n1610), .Z(n7457) );
  NANDN U7826 ( .A(n1564), .B(n7460), .Z(n1558) );
  NAND U7827 ( .A(n7461), .B(n1565), .Z(n7460) );
  OR U7828 ( .A(B[735]), .B(A[735]), .Z(n1565) );
  NANDN U7829 ( .A(n1567), .B(n7462), .Z(n7461) );
  NAND U7830 ( .A(n7463), .B(n1569), .Z(n7462) );
  OR U7831 ( .A(B[734]), .B(A[734]), .Z(n1569) );
  NANDN U7832 ( .A(n1571), .B(n7464), .Z(n7463) );
  NAND U7833 ( .A(n7465), .B(n1574), .Z(n7464) );
  OR U7834 ( .A(B[733]), .B(A[733]), .Z(n1574) );
  NANDN U7835 ( .A(n1576), .B(n7466), .Z(n7465) );
  NAND U7836 ( .A(n7467), .B(n1579), .Z(n7466) );
  OR U7837 ( .A(B[732]), .B(A[732]), .Z(n1579) );
  NANDN U7838 ( .A(n1581), .B(n7468), .Z(n7467) );
  NAND U7839 ( .A(n7469), .B(n1583), .Z(n7468) );
  AND U7840 ( .A(n7470), .B(n7471), .Z(n1583) );
  AND U7841 ( .A(n1606), .B(n1597), .Z(n7471) );
  OR U7842 ( .A(B[728]), .B(A[728]), .Z(n1606) );
  AND U7843 ( .A(n1592), .B(n1588), .Z(n7470) );
  NANDN U7844 ( .A(n1608), .B(n7472), .Z(n7469) );
  NANDN U7845 ( .A(n1610), .B(n1631), .Z(n7472) );
  NANDN U7846 ( .A(n1635), .B(n7473), .Z(n1631) );
  NAND U7847 ( .A(n7474), .B(n1636), .Z(n7473) );
  OR U7848 ( .A(B[723]), .B(A[723]), .Z(n1636) );
  NANDN U7849 ( .A(n1638), .B(n7475), .Z(n7474) );
  NAND U7850 ( .A(n7476), .B(n1640), .Z(n7475) );
  OR U7851 ( .A(B[722]), .B(A[722]), .Z(n1640) );
  NANDN U7852 ( .A(n1642), .B(n7477), .Z(n7476) );
  NAND U7853 ( .A(n1645), .B(n1647), .Z(n7477) );
  AND U7854 ( .A(B[720]), .B(A[720]), .Z(n1647) );
  OR U7855 ( .A(B[721]), .B(A[721]), .Z(n1645) );
  AND U7856 ( .A(B[721]), .B(A[721]), .Z(n1642) );
  AND U7857 ( .A(B[722]), .B(A[722]), .Z(n1638) );
  AND U7858 ( .A(B[723]), .B(A[723]), .Z(n1635) );
  NAND U7859 ( .A(n7478), .B(n7479), .Z(n1610) );
  AND U7860 ( .A(n1628), .B(n1624), .Z(n7479) );
  OR U7861 ( .A(B[724]), .B(A[724]), .Z(n1628) );
  AND U7862 ( .A(n1619), .B(n1615), .Z(n7478) );
  NANDN U7863 ( .A(n1614), .B(n7480), .Z(n1608) );
  NAND U7864 ( .A(n7481), .B(n1615), .Z(n7480) );
  OR U7865 ( .A(B[727]), .B(A[727]), .Z(n1615) );
  NANDN U7866 ( .A(n1617), .B(n7482), .Z(n7481) );
  NAND U7867 ( .A(n7483), .B(n1619), .Z(n7482) );
  OR U7868 ( .A(B[726]), .B(A[726]), .Z(n1619) );
  NANDN U7869 ( .A(n1621), .B(n7484), .Z(n7483) );
  NAND U7870 ( .A(n1624), .B(n1626), .Z(n7484) );
  AND U7871 ( .A(B[724]), .B(A[724]), .Z(n1626) );
  OR U7872 ( .A(B[725]), .B(A[725]), .Z(n1624) );
  AND U7873 ( .A(B[725]), .B(A[725]), .Z(n1621) );
  AND U7874 ( .A(B[726]), .B(A[726]), .Z(n1617) );
  AND U7875 ( .A(B[727]), .B(A[727]), .Z(n1614) );
  NANDN U7876 ( .A(n1587), .B(n7485), .Z(n1581) );
  NAND U7877 ( .A(n7486), .B(n1588), .Z(n7485) );
  OR U7878 ( .A(B[731]), .B(A[731]), .Z(n1588) );
  NANDN U7879 ( .A(n1590), .B(n7487), .Z(n7486) );
  NAND U7880 ( .A(n7488), .B(n1592), .Z(n7487) );
  OR U7881 ( .A(B[730]), .B(A[730]), .Z(n1592) );
  NANDN U7882 ( .A(n1594), .B(n7489), .Z(n7488) );
  NAND U7883 ( .A(n1597), .B(n1604), .Z(n7489) );
  AND U7884 ( .A(B[728]), .B(A[728]), .Z(n1604) );
  OR U7885 ( .A(B[729]), .B(A[729]), .Z(n1597) );
  AND U7886 ( .A(B[729]), .B(A[729]), .Z(n1594) );
  AND U7887 ( .A(B[730]), .B(A[730]), .Z(n1590) );
  AND U7888 ( .A(B[731]), .B(A[731]), .Z(n1587) );
  AND U7889 ( .A(B[732]), .B(A[732]), .Z(n1576) );
  AND U7890 ( .A(B[733]), .B(A[733]), .Z(n1571) );
  AND U7891 ( .A(B[734]), .B(A[734]), .Z(n1567) );
  AND U7892 ( .A(B[735]), .B(A[735]), .Z(n1564) );
  NAND U7893 ( .A(n7490), .B(n7491), .Z(n1463) );
  AND U7894 ( .A(n7492), .B(n7493), .Z(n7491) );
  AND U7895 ( .A(n1487), .B(n1477), .Z(n7493) );
  AND U7896 ( .A(n1472), .B(n1468), .Z(n7492) );
  ANDN U7897 ( .B(n7494), .A(n1535), .Z(n7490) );
  NAND U7898 ( .A(n7495), .B(n7496), .Z(n1535) );
  AND U7899 ( .A(n1556), .B(n1552), .Z(n7496) );
  OR U7900 ( .A(B[736]), .B(A[736]), .Z(n1556) );
  AND U7901 ( .A(n1547), .B(n1543), .Z(n7495) );
  ANDN U7902 ( .B(n1491), .A(n1513), .Z(n7494) );
  NANDN U7903 ( .A(n1467), .B(n7497), .Z(n1461) );
  NAND U7904 ( .A(n7498), .B(n1468), .Z(n7497) );
  OR U7905 ( .A(B[751]), .B(A[751]), .Z(n1468) );
  NANDN U7906 ( .A(n1470), .B(n7499), .Z(n7498) );
  NAND U7907 ( .A(n7500), .B(n1472), .Z(n7499) );
  OR U7908 ( .A(B[750]), .B(A[750]), .Z(n1472) );
  NANDN U7909 ( .A(n1474), .B(n7501), .Z(n7500) );
  NAND U7910 ( .A(n7502), .B(n1477), .Z(n7501) );
  OR U7911 ( .A(B[749]), .B(A[749]), .Z(n1477) );
  NANDN U7912 ( .A(n1484), .B(n7503), .Z(n7502) );
  NAND U7913 ( .A(n7504), .B(n1487), .Z(n7503) );
  OR U7914 ( .A(B[748]), .B(A[748]), .Z(n1487) );
  NANDN U7915 ( .A(n1489), .B(n7505), .Z(n7504) );
  NAND U7916 ( .A(n7506), .B(n1491), .Z(n7505) );
  AND U7917 ( .A(n7507), .B(n7508), .Z(n1491) );
  AND U7918 ( .A(n1509), .B(n1505), .Z(n7508) );
  OR U7919 ( .A(B[744]), .B(A[744]), .Z(n1509) );
  AND U7920 ( .A(n1500), .B(n1496), .Z(n7507) );
  NANDN U7921 ( .A(n1511), .B(n7509), .Z(n7506) );
  NANDN U7922 ( .A(n1513), .B(n1534), .Z(n7509) );
  NANDN U7923 ( .A(n1542), .B(n7510), .Z(n1534) );
  NAND U7924 ( .A(n7511), .B(n1543), .Z(n7510) );
  OR U7925 ( .A(B[739]), .B(A[739]), .Z(n1543) );
  NANDN U7926 ( .A(n1545), .B(n7512), .Z(n7511) );
  NAND U7927 ( .A(n7513), .B(n1547), .Z(n7512) );
  OR U7928 ( .A(B[738]), .B(A[738]), .Z(n1547) );
  NANDN U7929 ( .A(n1549), .B(n7514), .Z(n7513) );
  NAND U7930 ( .A(n1552), .B(n1554), .Z(n7514) );
  AND U7931 ( .A(B[736]), .B(A[736]), .Z(n1554) );
  OR U7932 ( .A(B[737]), .B(A[737]), .Z(n1552) );
  AND U7933 ( .A(B[737]), .B(A[737]), .Z(n1549) );
  AND U7934 ( .A(B[738]), .B(A[738]), .Z(n1545) );
  AND U7935 ( .A(B[739]), .B(A[739]), .Z(n1542) );
  NAND U7936 ( .A(n7515), .B(n7516), .Z(n1513) );
  AND U7937 ( .A(n1531), .B(n1527), .Z(n7516) );
  OR U7938 ( .A(B[740]), .B(A[740]), .Z(n1531) );
  AND U7939 ( .A(n1522), .B(n1518), .Z(n7515) );
  NANDN U7940 ( .A(n1517), .B(n7517), .Z(n1511) );
  NAND U7941 ( .A(n7518), .B(n1518), .Z(n7517) );
  OR U7942 ( .A(B[743]), .B(A[743]), .Z(n1518) );
  NANDN U7943 ( .A(n1520), .B(n7519), .Z(n7518) );
  NAND U7944 ( .A(n7520), .B(n1522), .Z(n7519) );
  OR U7945 ( .A(B[742]), .B(A[742]), .Z(n1522) );
  NANDN U7946 ( .A(n1524), .B(n7521), .Z(n7520) );
  NAND U7947 ( .A(n1527), .B(n1529), .Z(n7521) );
  AND U7948 ( .A(B[740]), .B(A[740]), .Z(n1529) );
  OR U7949 ( .A(B[741]), .B(A[741]), .Z(n1527) );
  AND U7950 ( .A(B[741]), .B(A[741]), .Z(n1524) );
  AND U7951 ( .A(B[742]), .B(A[742]), .Z(n1520) );
  AND U7952 ( .A(B[743]), .B(A[743]), .Z(n1517) );
  NANDN U7953 ( .A(n1495), .B(n7522), .Z(n1489) );
  NAND U7954 ( .A(n7523), .B(n1496), .Z(n7522) );
  OR U7955 ( .A(B[747]), .B(A[747]), .Z(n1496) );
  NANDN U7956 ( .A(n1498), .B(n7524), .Z(n7523) );
  NAND U7957 ( .A(n7525), .B(n1500), .Z(n7524) );
  OR U7958 ( .A(B[746]), .B(A[746]), .Z(n1500) );
  NANDN U7959 ( .A(n1502), .B(n7526), .Z(n7525) );
  NAND U7960 ( .A(n1505), .B(n1507), .Z(n7526) );
  AND U7961 ( .A(B[744]), .B(A[744]), .Z(n1507) );
  OR U7962 ( .A(B[745]), .B(A[745]), .Z(n1505) );
  AND U7963 ( .A(B[745]), .B(A[745]), .Z(n1502) );
  AND U7964 ( .A(B[746]), .B(A[746]), .Z(n1498) );
  AND U7965 ( .A(B[747]), .B(A[747]), .Z(n1495) );
  AND U7966 ( .A(B[748]), .B(A[748]), .Z(n1484) );
  AND U7967 ( .A(B[749]), .B(A[749]), .Z(n1474) );
  AND U7968 ( .A(B[750]), .B(A[750]), .Z(n1470) );
  AND U7969 ( .A(B[751]), .B(A[751]), .Z(n1467) );
  ANDN U7970 ( .B(n7527), .A(n1441), .Z(n5703) );
  NAND U7971 ( .A(n7528), .B(n7529), .Z(n1441) );
  AND U7972 ( .A(n1459), .B(n1455), .Z(n7529) );
  OR U7973 ( .A(B[752]), .B(A[752]), .Z(n1459) );
  ANDN U7974 ( .B(n1446), .A(n1449), .Z(n7528) );
  ANDN U7975 ( .B(n1412), .A(n1389), .Z(n7527) );
  ANDN U7976 ( .B(n7530), .A(n1373), .Z(n5701) );
  AND U7977 ( .A(B[766]), .B(A[766]), .Z(n1373) );
  NAND U7978 ( .A(n7531), .B(n1375), .Z(n7530) );
  OR U7979 ( .A(A[766]), .B(B[766]), .Z(n1375) );
  NANDN U7980 ( .A(n1377), .B(n7532), .Z(n7531) );
  NAND U7981 ( .A(n7533), .B(n1380), .Z(n7532) );
  OR U7982 ( .A(B[765]), .B(A[765]), .Z(n1380) );
  NANDN U7983 ( .A(n1382), .B(n7534), .Z(n7533) );
  NANDN U7984 ( .A(n1384), .B(n7535), .Z(n7534) );
  NANDN U7985 ( .A(n1387), .B(n7536), .Z(n7535) );
  NANDN U7986 ( .A(n1389), .B(n7537), .Z(n7536) );
  NANDN U7987 ( .A(n1409), .B(n7538), .Z(n7537) );
  NAND U7988 ( .A(n1440), .B(n1412), .Z(n7538) );
  AND U7989 ( .A(n7539), .B(n7540), .Z(n1412) );
  AND U7990 ( .A(n1437), .B(n1433), .Z(n7540) );
  OR U7991 ( .A(B[756]), .B(A[756]), .Z(n1437) );
  AND U7992 ( .A(n1428), .B(n1424), .Z(n7539) );
  NANDN U7993 ( .A(n1445), .B(n7541), .Z(n1440) );
  NAND U7994 ( .A(n7542), .B(n1446), .Z(n7541) );
  OR U7995 ( .A(B[755]), .B(A[755]), .Z(n1446) );
  NANDN U7996 ( .A(n1448), .B(n7543), .Z(n7542) );
  NANDN U7997 ( .A(n1449), .B(n7544), .Z(n7543) );
  NANDN U7998 ( .A(n1452), .B(n7545), .Z(n7544) );
  NAND U7999 ( .A(n1455), .B(n1457), .Z(n7545) );
  AND U8000 ( .A(A[752]), .B(B[752]), .Z(n1457) );
  OR U8001 ( .A(B[753]), .B(A[753]), .Z(n1455) );
  AND U8002 ( .A(B[753]), .B(A[753]), .Z(n1452) );
  NOR U8003 ( .A(B[754]), .B(A[754]), .Z(n1449) );
  AND U8004 ( .A(B[754]), .B(A[754]), .Z(n1448) );
  AND U8005 ( .A(B[755]), .B(A[755]), .Z(n1445) );
  NANDN U8006 ( .A(n1423), .B(n7546), .Z(n1409) );
  NAND U8007 ( .A(n7547), .B(n1424), .Z(n7546) );
  OR U8008 ( .A(B[759]), .B(A[759]), .Z(n1424) );
  NANDN U8009 ( .A(n1426), .B(n7548), .Z(n7547) );
  NAND U8010 ( .A(n7549), .B(n1428), .Z(n7548) );
  OR U8011 ( .A(B[758]), .B(A[758]), .Z(n1428) );
  NANDN U8012 ( .A(n1430), .B(n7550), .Z(n7549) );
  NAND U8013 ( .A(n1433), .B(n1435), .Z(n7550) );
  AND U8014 ( .A(B[756]), .B(A[756]), .Z(n1435) );
  OR U8015 ( .A(B[757]), .B(A[757]), .Z(n1433) );
  AND U8016 ( .A(B[757]), .B(A[757]), .Z(n1430) );
  AND U8017 ( .A(B[758]), .B(A[758]), .Z(n1426) );
  AND U8018 ( .A(B[759]), .B(A[759]), .Z(n1423) );
  NAND U8019 ( .A(n7551), .B(n7552), .Z(n1389) );
  AND U8020 ( .A(n1407), .B(n1403), .Z(n7552) );
  OR U8021 ( .A(B[760]), .B(A[760]), .Z(n1407) );
  AND U8022 ( .A(n1398), .B(n1394), .Z(n7551) );
  NANDN U8023 ( .A(n1393), .B(n7553), .Z(n1387) );
  NAND U8024 ( .A(n7554), .B(n1394), .Z(n7553) );
  OR U8025 ( .A(B[763]), .B(A[763]), .Z(n1394) );
  NANDN U8026 ( .A(n1396), .B(n7555), .Z(n7554) );
  NAND U8027 ( .A(n7556), .B(n1398), .Z(n7555) );
  OR U8028 ( .A(B[762]), .B(A[762]), .Z(n1398) );
  NANDN U8029 ( .A(n1400), .B(n7557), .Z(n7556) );
  NAND U8030 ( .A(n1403), .B(n1405), .Z(n7557) );
  AND U8031 ( .A(B[760]), .B(A[760]), .Z(n1405) );
  OR U8032 ( .A(B[761]), .B(A[761]), .Z(n1403) );
  AND U8033 ( .A(B[761]), .B(A[761]), .Z(n1400) );
  AND U8034 ( .A(B[762]), .B(A[762]), .Z(n1396) );
  AND U8035 ( .A(B[763]), .B(A[763]), .Z(n1393) );
  NOR U8036 ( .A(B[764]), .B(A[764]), .Z(n1384) );
  AND U8037 ( .A(B[764]), .B(A[764]), .Z(n1382) );
  AND U8038 ( .A(B[765]), .B(A[765]), .Z(n1377) );
  NOR U8039 ( .A(B[767]), .B(A[767]), .Z(n1370) );
  NOR U8040 ( .A(n1343), .B(n1294), .Z(n5696) );
  NAND U8041 ( .A(n7558), .B(n7559), .Z(n1343) );
  AND U8042 ( .A(n1366), .B(n1357), .Z(n7559) );
  OR U8043 ( .A(B[768]), .B(A[768]), .Z(n1366) );
  ANDN U8044 ( .B(n1348), .A(n1351), .Z(n7558) );
  ANDN U8045 ( .B(n7560), .A(n1287), .Z(n5694) );
  AND U8046 ( .A(B[780]), .B(A[780]), .Z(n1287) );
  NAND U8047 ( .A(n7561), .B(n1290), .Z(n7560) );
  OR U8048 ( .A(A[780]), .B(B[780]), .Z(n1290) );
  NANDN U8049 ( .A(n1292), .B(n7562), .Z(n7561) );
  NANDN U8050 ( .A(n1294), .B(n7563), .Z(n7562) );
  NANDN U8051 ( .A(n1319), .B(n7564), .Z(n7563) );
  NAND U8052 ( .A(n1342), .B(n1322), .Z(n7564) );
  AND U8053 ( .A(n7565), .B(n7566), .Z(n1322) );
  AND U8054 ( .A(n1339), .B(n1335), .Z(n7566) );
  OR U8055 ( .A(B[772]), .B(A[772]), .Z(n1339) );
  AND U8056 ( .A(n1330), .B(n1326), .Z(n7565) );
  NANDN U8057 ( .A(n1347), .B(n7567), .Z(n1342) );
  NAND U8058 ( .A(n7568), .B(n1348), .Z(n7567) );
  OR U8059 ( .A(B[771]), .B(A[771]), .Z(n1348) );
  NANDN U8060 ( .A(n1350), .B(n7569), .Z(n7568) );
  NANDN U8061 ( .A(n1351), .B(n7570), .Z(n7569) );
  NANDN U8062 ( .A(n1354), .B(n7571), .Z(n7570) );
  NAND U8063 ( .A(n1357), .B(n1364), .Z(n7571) );
  AND U8064 ( .A(A[768]), .B(B[768]), .Z(n1364) );
  OR U8065 ( .A(B[769]), .B(A[769]), .Z(n1357) );
  AND U8066 ( .A(B[769]), .B(A[769]), .Z(n1354) );
  NOR U8067 ( .A(B[770]), .B(A[770]), .Z(n1351) );
  AND U8068 ( .A(B[770]), .B(A[770]), .Z(n1350) );
  AND U8069 ( .A(B[771]), .B(A[771]), .Z(n1347) );
  NANDN U8070 ( .A(n1325), .B(n7572), .Z(n1319) );
  NAND U8071 ( .A(n7573), .B(n1326), .Z(n7572) );
  OR U8072 ( .A(B[775]), .B(A[775]), .Z(n1326) );
  NANDN U8073 ( .A(n1328), .B(n7574), .Z(n7573) );
  NAND U8074 ( .A(n7575), .B(n1330), .Z(n7574) );
  OR U8075 ( .A(B[774]), .B(A[774]), .Z(n1330) );
  NANDN U8076 ( .A(n1332), .B(n7576), .Z(n7575) );
  NAND U8077 ( .A(n1335), .B(n1337), .Z(n7576) );
  AND U8078 ( .A(B[772]), .B(A[772]), .Z(n1337) );
  OR U8079 ( .A(B[773]), .B(A[773]), .Z(n1335) );
  AND U8080 ( .A(B[773]), .B(A[773]), .Z(n1332) );
  AND U8081 ( .A(B[774]), .B(A[774]), .Z(n1328) );
  AND U8082 ( .A(B[775]), .B(A[775]), .Z(n1325) );
  NAND U8083 ( .A(n7577), .B(n7578), .Z(n1294) );
  AND U8084 ( .A(n1317), .B(n1313), .Z(n7578) );
  OR U8085 ( .A(B[776]), .B(A[776]), .Z(n1317) );
  AND U8086 ( .A(n1308), .B(n1304), .Z(n7577) );
  NANDN U8087 ( .A(n1303), .B(n7579), .Z(n1292) );
  NAND U8088 ( .A(n7580), .B(n1304), .Z(n7579) );
  OR U8089 ( .A(B[779]), .B(A[779]), .Z(n1304) );
  NANDN U8090 ( .A(n1306), .B(n7581), .Z(n7580) );
  NAND U8091 ( .A(n7582), .B(n1308), .Z(n7581) );
  OR U8092 ( .A(B[778]), .B(A[778]), .Z(n1308) );
  NANDN U8093 ( .A(n1310), .B(n7583), .Z(n7582) );
  NAND U8094 ( .A(n1313), .B(n1315), .Z(n7583) );
  AND U8095 ( .A(B[776]), .B(A[776]), .Z(n1315) );
  OR U8096 ( .A(B[777]), .B(A[777]), .Z(n1313) );
  AND U8097 ( .A(B[777]), .B(A[777]), .Z(n1310) );
  AND U8098 ( .A(B[778]), .B(A[778]), .Z(n1306) );
  AND U8099 ( .A(B[779]), .B(A[779]), .Z(n1303) );
  NOR U8100 ( .A(B[781]), .B(A[781]), .Z(n1284) );
  AND U8101 ( .A(B[781]), .B(A[781]), .Z(n1282) );
  NOR U8102 ( .A(B[782]), .B(A[782]), .Z(n1279) );
  AND U8103 ( .A(B[782]), .B(A[782]), .Z(n1278) );
  NOR U8104 ( .A(B[783]), .B(A[783]), .Z(n1275) );
  NOR U8105 ( .A(n1253), .B(n1204), .Z(n5685) );
  NAND U8106 ( .A(n7584), .B(n7585), .Z(n1253) );
  AND U8107 ( .A(n1271), .B(n1267), .Z(n7585) );
  OR U8108 ( .A(B[784]), .B(A[784]), .Z(n1271) );
  ANDN U8109 ( .B(n1258), .A(n1261), .Z(n7584) );
  ANDN U8110 ( .B(n7586), .A(n1197), .Z(n5683) );
  AND U8111 ( .A(B[796]), .B(A[796]), .Z(n1197) );
  NAND U8112 ( .A(n7587), .B(n1200), .Z(n7586) );
  OR U8113 ( .A(A[796]), .B(B[796]), .Z(n1200) );
  NANDN U8114 ( .A(n1202), .B(n7588), .Z(n7587) );
  NANDN U8115 ( .A(n1204), .B(n7589), .Z(n7588) );
  NANDN U8116 ( .A(n1224), .B(n7590), .Z(n7589) );
  NAND U8117 ( .A(n1252), .B(n1227), .Z(n7590) );
  AND U8118 ( .A(n7591), .B(n7592), .Z(n1227) );
  AND U8119 ( .A(n1249), .B(n1240), .Z(n7592) );
  OR U8120 ( .A(B[788]), .B(A[788]), .Z(n1249) );
  AND U8121 ( .A(n1235), .B(n1231), .Z(n7591) );
  NANDN U8122 ( .A(n1257), .B(n7593), .Z(n1252) );
  NAND U8123 ( .A(n7594), .B(n1258), .Z(n7593) );
  OR U8124 ( .A(B[787]), .B(A[787]), .Z(n1258) );
  NANDN U8125 ( .A(n1260), .B(n7595), .Z(n7594) );
  NANDN U8126 ( .A(n1261), .B(n7596), .Z(n7595) );
  NANDN U8127 ( .A(n1264), .B(n7597), .Z(n7596) );
  NAND U8128 ( .A(n1267), .B(n1269), .Z(n7597) );
  AND U8129 ( .A(A[784]), .B(B[784]), .Z(n1269) );
  OR U8130 ( .A(B[785]), .B(A[785]), .Z(n1267) );
  AND U8131 ( .A(B[785]), .B(A[785]), .Z(n1264) );
  NOR U8132 ( .A(B[786]), .B(A[786]), .Z(n1261) );
  AND U8133 ( .A(B[786]), .B(A[786]), .Z(n1260) );
  AND U8134 ( .A(B[787]), .B(A[787]), .Z(n1257) );
  NANDN U8135 ( .A(n1230), .B(n7598), .Z(n1224) );
  NAND U8136 ( .A(n7599), .B(n1231), .Z(n7598) );
  OR U8137 ( .A(B[791]), .B(A[791]), .Z(n1231) );
  NANDN U8138 ( .A(n1233), .B(n7600), .Z(n7599) );
  NAND U8139 ( .A(n7601), .B(n1235), .Z(n7600) );
  OR U8140 ( .A(B[790]), .B(A[790]), .Z(n1235) );
  NANDN U8141 ( .A(n1237), .B(n7602), .Z(n7601) );
  NAND U8142 ( .A(n1240), .B(n1247), .Z(n7602) );
  AND U8143 ( .A(B[788]), .B(A[788]), .Z(n1247) );
  OR U8144 ( .A(B[789]), .B(A[789]), .Z(n1240) );
  AND U8145 ( .A(B[789]), .B(A[789]), .Z(n1237) );
  AND U8146 ( .A(B[790]), .B(A[790]), .Z(n1233) );
  AND U8147 ( .A(B[791]), .B(A[791]), .Z(n1230) );
  NAND U8148 ( .A(n7603), .B(n7604), .Z(n1204) );
  AND U8149 ( .A(n1222), .B(n1218), .Z(n7604) );
  OR U8150 ( .A(B[792]), .B(A[792]), .Z(n1222) );
  AND U8151 ( .A(n1213), .B(n1209), .Z(n7603) );
  NANDN U8152 ( .A(n1208), .B(n7605), .Z(n1202) );
  NAND U8153 ( .A(n7606), .B(n1209), .Z(n7605) );
  OR U8154 ( .A(B[795]), .B(A[795]), .Z(n1209) );
  NANDN U8155 ( .A(n1211), .B(n7607), .Z(n7606) );
  NAND U8156 ( .A(n7608), .B(n1213), .Z(n7607) );
  OR U8157 ( .A(B[794]), .B(A[794]), .Z(n1213) );
  NANDN U8158 ( .A(n1215), .B(n7609), .Z(n7608) );
  NAND U8159 ( .A(n1218), .B(n1220), .Z(n7609) );
  AND U8160 ( .A(B[792]), .B(A[792]), .Z(n1220) );
  OR U8161 ( .A(B[793]), .B(A[793]), .Z(n1218) );
  AND U8162 ( .A(B[793]), .B(A[793]), .Z(n1215) );
  AND U8163 ( .A(B[794]), .B(A[794]), .Z(n1211) );
  AND U8164 ( .A(B[795]), .B(A[795]), .Z(n1208) );
  NOR U8165 ( .A(B[797]), .B(A[797]), .Z(n1194) );
  AND U8166 ( .A(B[797]), .B(A[797]), .Z(n1192) );
  NOR U8167 ( .A(B[798]), .B(A[798]), .Z(n1189) );
  AND U8168 ( .A(B[798]), .B(A[798]), .Z(n1188) );
  NOR U8169 ( .A(B[799]), .B(A[799]), .Z(n1185) );
  NOR U8170 ( .A(n1149), .B(n1104), .Z(n5674) );
  NAND U8171 ( .A(n7610), .B(n7611), .Z(n1149) );
  AND U8172 ( .A(n1167), .B(n1163), .Z(n7611) );
  OR U8173 ( .A(B[800]), .B(A[800]), .Z(n1167) );
  ANDN U8174 ( .B(n1154), .A(n1157), .Z(n7610) );
  ANDN U8175 ( .B(n7612), .A(n1097), .Z(n5672) );
  AND U8176 ( .A(B[812]), .B(A[812]), .Z(n1097) );
  NAND U8177 ( .A(n7613), .B(n1100), .Z(n7612) );
  OR U8178 ( .A(A[812]), .B(B[812]), .Z(n1100) );
  NANDN U8179 ( .A(n1102), .B(n7614), .Z(n7613) );
  NANDN U8180 ( .A(n1104), .B(n7615), .Z(n7614) );
  NANDN U8181 ( .A(n1125), .B(n7616), .Z(n7615) );
  NAND U8182 ( .A(n1148), .B(n1128), .Z(n7616) );
  AND U8183 ( .A(n7617), .B(n7618), .Z(n1128) );
  AND U8184 ( .A(n1145), .B(n1141), .Z(n7618) );
  OR U8185 ( .A(B[804]), .B(A[804]), .Z(n1145) );
  AND U8186 ( .A(n1136), .B(n1132), .Z(n7617) );
  NANDN U8187 ( .A(n1153), .B(n7619), .Z(n1148) );
  NAND U8188 ( .A(n7620), .B(n1154), .Z(n7619) );
  OR U8189 ( .A(B[803]), .B(A[803]), .Z(n1154) );
  NANDN U8190 ( .A(n1156), .B(n7621), .Z(n7620) );
  NANDN U8191 ( .A(n1157), .B(n7622), .Z(n7621) );
  NANDN U8192 ( .A(n1160), .B(n7623), .Z(n7622) );
  NAND U8193 ( .A(n1163), .B(n1165), .Z(n7623) );
  AND U8194 ( .A(A[800]), .B(B[800]), .Z(n1165) );
  OR U8195 ( .A(B[801]), .B(A[801]), .Z(n1163) );
  AND U8196 ( .A(B[801]), .B(A[801]), .Z(n1160) );
  NOR U8197 ( .A(B[802]), .B(A[802]), .Z(n1157) );
  AND U8198 ( .A(B[802]), .B(A[802]), .Z(n1156) );
  AND U8199 ( .A(B[803]), .B(A[803]), .Z(n1153) );
  NANDN U8200 ( .A(n1131), .B(n7624), .Z(n1125) );
  NAND U8201 ( .A(n7625), .B(n1132), .Z(n7624) );
  OR U8202 ( .A(B[807]), .B(A[807]), .Z(n1132) );
  NANDN U8203 ( .A(n1134), .B(n7626), .Z(n7625) );
  NAND U8204 ( .A(n7627), .B(n1136), .Z(n7626) );
  OR U8205 ( .A(B[806]), .B(A[806]), .Z(n1136) );
  NANDN U8206 ( .A(n1138), .B(n7628), .Z(n7627) );
  NAND U8207 ( .A(n1141), .B(n1143), .Z(n7628) );
  AND U8208 ( .A(B[804]), .B(A[804]), .Z(n1143) );
  OR U8209 ( .A(B[805]), .B(A[805]), .Z(n1141) );
  AND U8210 ( .A(B[805]), .B(A[805]), .Z(n1138) );
  AND U8211 ( .A(B[806]), .B(A[806]), .Z(n1134) );
  AND U8212 ( .A(B[807]), .B(A[807]), .Z(n1131) );
  NAND U8213 ( .A(n7629), .B(n7630), .Z(n1104) );
  AND U8214 ( .A(n1123), .B(n1118), .Z(n7630) );
  OR U8215 ( .A(B[808]), .B(A[808]), .Z(n1123) );
  AND U8216 ( .A(n1113), .B(n1109), .Z(n7629) );
  NANDN U8217 ( .A(n1108), .B(n7631), .Z(n1102) );
  NAND U8218 ( .A(n7632), .B(n1109), .Z(n7631) );
  OR U8219 ( .A(B[811]), .B(A[811]), .Z(n1109) );
  NANDN U8220 ( .A(n1111), .B(n7633), .Z(n7632) );
  NAND U8221 ( .A(n7634), .B(n1113), .Z(n7633) );
  OR U8222 ( .A(B[810]), .B(A[810]), .Z(n1113) );
  NANDN U8223 ( .A(n1115), .B(n7635), .Z(n7634) );
  NAND U8224 ( .A(n1118), .B(n1121), .Z(n7635) );
  AND U8225 ( .A(B[808]), .B(A[808]), .Z(n1121) );
  OR U8226 ( .A(B[809]), .B(A[809]), .Z(n1118) );
  AND U8227 ( .A(B[809]), .B(A[809]), .Z(n1115) );
  AND U8228 ( .A(B[810]), .B(A[810]), .Z(n1111) );
  AND U8229 ( .A(B[811]), .B(A[811]), .Z(n1108) );
  NOR U8230 ( .A(B[813]), .B(A[813]), .Z(n1094) );
  AND U8231 ( .A(B[813]), .B(A[813]), .Z(n1092) );
  NOR U8232 ( .A(B[814]), .B(A[814]), .Z(n1089) );
  AND U8233 ( .A(B[814]), .B(A[814]), .Z(n1088) );
  NOR U8234 ( .A(B[815]), .B(A[815]), .Z(n1085) );
  NOR U8235 ( .A(n1059), .B(n1015), .Z(n5663) );
  NAND U8236 ( .A(n7636), .B(n7637), .Z(n1059) );
  AND U8237 ( .A(n1081), .B(n1077), .Z(n7637) );
  OR U8238 ( .A(B[816]), .B(A[816]), .Z(n1081) );
  ANDN U8239 ( .B(n1068), .A(n1071), .Z(n7636) );
  ANDN U8240 ( .B(n7638), .A(n1008), .Z(n5661) );
  AND U8241 ( .A(B[828]), .B(A[828]), .Z(n1008) );
  NAND U8242 ( .A(n7639), .B(n1011), .Z(n7638) );
  OR U8243 ( .A(A[828]), .B(B[828]), .Z(n1011) );
  NANDN U8244 ( .A(n1013), .B(n7640), .Z(n7639) );
  NANDN U8245 ( .A(n1015), .B(n7641), .Z(n7640) );
  NANDN U8246 ( .A(n1035), .B(n7642), .Z(n7641) );
  NAND U8247 ( .A(n1058), .B(n1038), .Z(n7642) );
  AND U8248 ( .A(n7643), .B(n7644), .Z(n1038) );
  AND U8249 ( .A(n1055), .B(n1051), .Z(n7644) );
  OR U8250 ( .A(B[820]), .B(A[820]), .Z(n1055) );
  AND U8251 ( .A(n1046), .B(n1042), .Z(n7643) );
  NANDN U8252 ( .A(n1067), .B(n7645), .Z(n1058) );
  NAND U8253 ( .A(n7646), .B(n1068), .Z(n7645) );
  OR U8254 ( .A(B[819]), .B(A[819]), .Z(n1068) );
  NANDN U8255 ( .A(n1070), .B(n7647), .Z(n7646) );
  NANDN U8256 ( .A(n1071), .B(n7648), .Z(n7647) );
  NANDN U8257 ( .A(n1074), .B(n7649), .Z(n7648) );
  NAND U8258 ( .A(n1077), .B(n1079), .Z(n7649) );
  AND U8259 ( .A(A[816]), .B(B[816]), .Z(n1079) );
  OR U8260 ( .A(B[817]), .B(A[817]), .Z(n1077) );
  AND U8261 ( .A(B[817]), .B(A[817]), .Z(n1074) );
  NOR U8262 ( .A(B[818]), .B(A[818]), .Z(n1071) );
  AND U8263 ( .A(B[818]), .B(A[818]), .Z(n1070) );
  AND U8264 ( .A(B[819]), .B(A[819]), .Z(n1067) );
  NANDN U8265 ( .A(n1041), .B(n7650), .Z(n1035) );
  NAND U8266 ( .A(n7651), .B(n1042), .Z(n7650) );
  OR U8267 ( .A(B[823]), .B(A[823]), .Z(n1042) );
  NANDN U8268 ( .A(n1044), .B(n7652), .Z(n7651) );
  NAND U8269 ( .A(n7653), .B(n1046), .Z(n7652) );
  OR U8270 ( .A(B[822]), .B(A[822]), .Z(n1046) );
  NANDN U8271 ( .A(n1048), .B(n7654), .Z(n7653) );
  NAND U8272 ( .A(n1051), .B(n1053), .Z(n7654) );
  AND U8273 ( .A(B[820]), .B(A[820]), .Z(n1053) );
  OR U8274 ( .A(B[821]), .B(A[821]), .Z(n1051) );
  AND U8275 ( .A(B[821]), .B(A[821]), .Z(n1048) );
  AND U8276 ( .A(B[822]), .B(A[822]), .Z(n1044) );
  AND U8277 ( .A(B[823]), .B(A[823]), .Z(n1041) );
  NAND U8278 ( .A(n7655), .B(n7656), .Z(n1015) );
  AND U8279 ( .A(n1033), .B(n1029), .Z(n7656) );
  OR U8280 ( .A(B[824]), .B(A[824]), .Z(n1033) );
  AND U8281 ( .A(n1024), .B(n1020), .Z(n7655) );
  NANDN U8282 ( .A(n1019), .B(n7657), .Z(n1013) );
  NAND U8283 ( .A(n7658), .B(n1020), .Z(n7657) );
  OR U8284 ( .A(B[827]), .B(A[827]), .Z(n1020) );
  NANDN U8285 ( .A(n1022), .B(n7659), .Z(n7658) );
  NAND U8286 ( .A(n7660), .B(n1024), .Z(n7659) );
  OR U8287 ( .A(B[826]), .B(A[826]), .Z(n1024) );
  NANDN U8288 ( .A(n1026), .B(n7661), .Z(n7660) );
  NAND U8289 ( .A(n1029), .B(n1031), .Z(n7661) );
  AND U8290 ( .A(B[824]), .B(A[824]), .Z(n1031) );
  OR U8291 ( .A(B[825]), .B(A[825]), .Z(n1029) );
  AND U8292 ( .A(B[825]), .B(A[825]), .Z(n1026) );
  AND U8293 ( .A(B[826]), .B(A[826]), .Z(n1022) );
  AND U8294 ( .A(B[827]), .B(A[827]), .Z(n1019) );
  NOR U8295 ( .A(B[829]), .B(A[829]), .Z(n1000) );
  AND U8296 ( .A(B[829]), .B(A[829]), .Z(n998) );
  NOR U8297 ( .A(B[830]), .B(A[830]), .Z(n995) );
  AND U8298 ( .A(B[830]), .B(A[830]), .Z(n994) );
  NOR U8299 ( .A(B[831]), .B(A[831]), .Z(n991) );
  NOR U8300 ( .A(n969), .B(n917), .Z(n5652) );
  NAND U8301 ( .A(n7662), .B(n7663), .Z(n969) );
  AND U8302 ( .A(n987), .B(n983), .Z(n7663) );
  OR U8303 ( .A(B[832]), .B(A[832]), .Z(n987) );
  ANDN U8304 ( .B(n974), .A(n977), .Z(n7662) );
  ANDN U8305 ( .B(n7664), .A(n910), .Z(n5650) );
  AND U8306 ( .A(B[844]), .B(A[844]), .Z(n910) );
  NAND U8307 ( .A(n7665), .B(n913), .Z(n7664) );
  OR U8308 ( .A(A[844]), .B(B[844]), .Z(n913) );
  NANDN U8309 ( .A(n915), .B(n7666), .Z(n7665) );
  NANDN U8310 ( .A(n917), .B(n7667), .Z(n7666) );
  NANDN U8311 ( .A(n937), .B(n7668), .Z(n7667) );
  NAND U8312 ( .A(n968), .B(n940), .Z(n7668) );
  AND U8313 ( .A(n7669), .B(n7670), .Z(n940) );
  AND U8314 ( .A(n965), .B(n961), .Z(n7670) );
  OR U8315 ( .A(B[836]), .B(A[836]), .Z(n965) );
  AND U8316 ( .A(n956), .B(n952), .Z(n7669) );
  NANDN U8317 ( .A(n973), .B(n7671), .Z(n968) );
  NAND U8318 ( .A(n7672), .B(n974), .Z(n7671) );
  OR U8319 ( .A(B[835]), .B(A[835]), .Z(n974) );
  NANDN U8320 ( .A(n976), .B(n7673), .Z(n7672) );
  NANDN U8321 ( .A(n977), .B(n7674), .Z(n7673) );
  NANDN U8322 ( .A(n980), .B(n7675), .Z(n7674) );
  NAND U8323 ( .A(n983), .B(n985), .Z(n7675) );
  AND U8324 ( .A(A[832]), .B(B[832]), .Z(n985) );
  OR U8325 ( .A(B[833]), .B(A[833]), .Z(n983) );
  AND U8326 ( .A(B[833]), .B(A[833]), .Z(n980) );
  NOR U8327 ( .A(B[834]), .B(A[834]), .Z(n977) );
  AND U8328 ( .A(B[834]), .B(A[834]), .Z(n976) );
  AND U8329 ( .A(B[835]), .B(A[835]), .Z(n973) );
  NANDN U8330 ( .A(n951), .B(n7676), .Z(n937) );
  NAND U8331 ( .A(n7677), .B(n952), .Z(n7676) );
  OR U8332 ( .A(B[839]), .B(A[839]), .Z(n952) );
  NANDN U8333 ( .A(n954), .B(n7678), .Z(n7677) );
  NAND U8334 ( .A(n7679), .B(n956), .Z(n7678) );
  OR U8335 ( .A(B[838]), .B(A[838]), .Z(n956) );
  NANDN U8336 ( .A(n958), .B(n7680), .Z(n7679) );
  NAND U8337 ( .A(n961), .B(n963), .Z(n7680) );
  AND U8338 ( .A(B[836]), .B(A[836]), .Z(n963) );
  OR U8339 ( .A(B[837]), .B(A[837]), .Z(n961) );
  AND U8340 ( .A(B[837]), .B(A[837]), .Z(n958) );
  AND U8341 ( .A(B[838]), .B(A[838]), .Z(n954) );
  AND U8342 ( .A(B[839]), .B(A[839]), .Z(n951) );
  NAND U8343 ( .A(n7681), .B(n7682), .Z(n917) );
  AND U8344 ( .A(n935), .B(n931), .Z(n7682) );
  OR U8345 ( .A(B[840]), .B(A[840]), .Z(n935) );
  AND U8346 ( .A(n926), .B(n922), .Z(n7681) );
  NANDN U8347 ( .A(n921), .B(n7683), .Z(n915) );
  NAND U8348 ( .A(n7684), .B(n922), .Z(n7683) );
  OR U8349 ( .A(B[843]), .B(A[843]), .Z(n922) );
  NANDN U8350 ( .A(n924), .B(n7685), .Z(n7684) );
  NAND U8351 ( .A(n7686), .B(n926), .Z(n7685) );
  OR U8352 ( .A(B[842]), .B(A[842]), .Z(n926) );
  NANDN U8353 ( .A(n928), .B(n7687), .Z(n7686) );
  NAND U8354 ( .A(n931), .B(n933), .Z(n7687) );
  AND U8355 ( .A(B[840]), .B(A[840]), .Z(n933) );
  OR U8356 ( .A(B[841]), .B(A[841]), .Z(n931) );
  AND U8357 ( .A(B[841]), .B(A[841]), .Z(n928) );
  AND U8358 ( .A(B[842]), .B(A[842]), .Z(n924) );
  AND U8359 ( .A(B[843]), .B(A[843]), .Z(n921) );
  NOR U8360 ( .A(B[845]), .B(A[845]), .Z(n907) );
  AND U8361 ( .A(B[845]), .B(A[845]), .Z(n905) );
  NOR U8362 ( .A(B[846]), .B(A[846]), .Z(n902) );
  AND U8363 ( .A(B[846]), .B(A[846]), .Z(n901) );
  NOR U8364 ( .A(B[847]), .B(A[847]), .Z(n898) );
  NOR U8365 ( .A(n871), .B(n823), .Z(n5641) );
  NAND U8366 ( .A(n7688), .B(n7689), .Z(n871) );
  AND U8367 ( .A(n894), .B(n885), .Z(n7689) );
  OR U8368 ( .A(B[848]), .B(A[848]), .Z(n894) );
  ANDN U8369 ( .B(n876), .A(n879), .Z(n7688) );
  ANDN U8370 ( .B(n7690), .A(n816), .Z(n5639) );
  AND U8371 ( .A(B[860]), .B(A[860]), .Z(n816) );
  NAND U8372 ( .A(n7691), .B(n819), .Z(n7690) );
  OR U8373 ( .A(A[860]), .B(B[860]), .Z(n819) );
  NANDN U8374 ( .A(n821), .B(n7692), .Z(n7691) );
  NANDN U8375 ( .A(n823), .B(n7693), .Z(n7692) );
  NANDN U8376 ( .A(n847), .B(n7694), .Z(n7693) );
  NAND U8377 ( .A(n870), .B(n850), .Z(n7694) );
  AND U8378 ( .A(n7695), .B(n7696), .Z(n850) );
  AND U8379 ( .A(n867), .B(n863), .Z(n7696) );
  OR U8380 ( .A(B[852]), .B(A[852]), .Z(n867) );
  AND U8381 ( .A(n858), .B(n854), .Z(n7695) );
  NANDN U8382 ( .A(n875), .B(n7697), .Z(n870) );
  NAND U8383 ( .A(n7698), .B(n876), .Z(n7697) );
  OR U8384 ( .A(B[851]), .B(A[851]), .Z(n876) );
  NANDN U8385 ( .A(n878), .B(n7699), .Z(n7698) );
  NANDN U8386 ( .A(n879), .B(n7700), .Z(n7699) );
  NANDN U8387 ( .A(n882), .B(n7701), .Z(n7700) );
  NAND U8388 ( .A(n885), .B(n892), .Z(n7701) );
  AND U8389 ( .A(A[848]), .B(B[848]), .Z(n892) );
  OR U8390 ( .A(B[849]), .B(A[849]), .Z(n885) );
  AND U8391 ( .A(B[849]), .B(A[849]), .Z(n882) );
  NOR U8392 ( .A(B[850]), .B(A[850]), .Z(n879) );
  AND U8393 ( .A(B[850]), .B(A[850]), .Z(n878) );
  AND U8394 ( .A(B[851]), .B(A[851]), .Z(n875) );
  NANDN U8395 ( .A(n853), .B(n7702), .Z(n847) );
  NAND U8396 ( .A(n7703), .B(n854), .Z(n7702) );
  OR U8397 ( .A(B[855]), .B(A[855]), .Z(n854) );
  NANDN U8398 ( .A(n856), .B(n7704), .Z(n7703) );
  NAND U8399 ( .A(n7705), .B(n858), .Z(n7704) );
  OR U8400 ( .A(B[854]), .B(A[854]), .Z(n858) );
  NANDN U8401 ( .A(n860), .B(n7706), .Z(n7705) );
  NAND U8402 ( .A(n863), .B(n865), .Z(n7706) );
  AND U8403 ( .A(B[852]), .B(A[852]), .Z(n865) );
  OR U8404 ( .A(B[853]), .B(A[853]), .Z(n863) );
  AND U8405 ( .A(B[853]), .B(A[853]), .Z(n860) );
  AND U8406 ( .A(B[854]), .B(A[854]), .Z(n856) );
  AND U8407 ( .A(B[855]), .B(A[855]), .Z(n853) );
  NAND U8408 ( .A(n7707), .B(n7708), .Z(n823) );
  AND U8409 ( .A(n845), .B(n841), .Z(n7708) );
  OR U8410 ( .A(B[856]), .B(A[856]), .Z(n845) );
  AND U8411 ( .A(n836), .B(n832), .Z(n7707) );
  NANDN U8412 ( .A(n831), .B(n7709), .Z(n821) );
  NAND U8413 ( .A(n7710), .B(n832), .Z(n7709) );
  OR U8414 ( .A(B[859]), .B(A[859]), .Z(n832) );
  NANDN U8415 ( .A(n834), .B(n7711), .Z(n7710) );
  NAND U8416 ( .A(n7712), .B(n836), .Z(n7711) );
  OR U8417 ( .A(B[858]), .B(A[858]), .Z(n836) );
  NANDN U8418 ( .A(n838), .B(n7713), .Z(n7712) );
  NAND U8419 ( .A(n841), .B(n843), .Z(n7713) );
  AND U8420 ( .A(B[856]), .B(A[856]), .Z(n843) );
  OR U8421 ( .A(B[857]), .B(A[857]), .Z(n841) );
  AND U8422 ( .A(B[857]), .B(A[857]), .Z(n838) );
  AND U8423 ( .A(B[858]), .B(A[858]), .Z(n834) );
  AND U8424 ( .A(B[859]), .B(A[859]), .Z(n831) );
  NOR U8425 ( .A(B[861]), .B(A[861]), .Z(n813) );
  AND U8426 ( .A(B[861]), .B(A[861]), .Z(n811) );
  NOR U8427 ( .A(B[862]), .B(A[862]), .Z(n808) );
  AND U8428 ( .A(B[862]), .B(A[862]), .Z(n807) );
  NOR U8429 ( .A(B[863]), .B(A[863]), .Z(n804) );
  NOR U8430 ( .A(n782), .B(n733), .Z(n5630) );
  NAND U8431 ( .A(n7714), .B(n7715), .Z(n782) );
  AND U8432 ( .A(n800), .B(n796), .Z(n7715) );
  OR U8433 ( .A(B[864]), .B(A[864]), .Z(n800) );
  ANDN U8434 ( .B(n787), .A(n790), .Z(n7714) );
  ANDN U8435 ( .B(n7716), .A(n726), .Z(n5628) );
  AND U8436 ( .A(B[876]), .B(A[876]), .Z(n726) );
  NAND U8437 ( .A(n7717), .B(n729), .Z(n7716) );
  OR U8438 ( .A(A[876]), .B(B[876]), .Z(n729) );
  NANDN U8439 ( .A(n731), .B(n7718), .Z(n7717) );
  NANDN U8440 ( .A(n733), .B(n7719), .Z(n7718) );
  NANDN U8441 ( .A(n753), .B(n7720), .Z(n7719) );
  NAND U8442 ( .A(n781), .B(n756), .Z(n7720) );
  AND U8443 ( .A(n7721), .B(n7722), .Z(n756) );
  AND U8444 ( .A(n778), .B(n769), .Z(n7722) );
  OR U8445 ( .A(B[868]), .B(A[868]), .Z(n778) );
  AND U8446 ( .A(n764), .B(n760), .Z(n7721) );
  NANDN U8447 ( .A(n786), .B(n7723), .Z(n781) );
  NAND U8448 ( .A(n7724), .B(n787), .Z(n7723) );
  OR U8449 ( .A(B[867]), .B(A[867]), .Z(n787) );
  NANDN U8450 ( .A(n789), .B(n7725), .Z(n7724) );
  NANDN U8451 ( .A(n790), .B(n7726), .Z(n7725) );
  NANDN U8452 ( .A(n793), .B(n7727), .Z(n7726) );
  NAND U8453 ( .A(n796), .B(n798), .Z(n7727) );
  AND U8454 ( .A(A[864]), .B(B[864]), .Z(n798) );
  OR U8455 ( .A(B[865]), .B(A[865]), .Z(n796) );
  AND U8456 ( .A(B[865]), .B(A[865]), .Z(n793) );
  NOR U8457 ( .A(B[866]), .B(A[866]), .Z(n790) );
  AND U8458 ( .A(B[866]), .B(A[866]), .Z(n789) );
  AND U8459 ( .A(B[867]), .B(A[867]), .Z(n786) );
  NANDN U8460 ( .A(n759), .B(n7728), .Z(n753) );
  NAND U8461 ( .A(n7729), .B(n760), .Z(n7728) );
  OR U8462 ( .A(B[871]), .B(A[871]), .Z(n760) );
  NANDN U8463 ( .A(n762), .B(n7730), .Z(n7729) );
  NAND U8464 ( .A(n7731), .B(n764), .Z(n7730) );
  OR U8465 ( .A(B[870]), .B(A[870]), .Z(n764) );
  NANDN U8466 ( .A(n766), .B(n7732), .Z(n7731) );
  NAND U8467 ( .A(n769), .B(n776), .Z(n7732) );
  AND U8468 ( .A(B[868]), .B(A[868]), .Z(n776) );
  OR U8469 ( .A(B[869]), .B(A[869]), .Z(n769) );
  AND U8470 ( .A(B[869]), .B(A[869]), .Z(n766) );
  AND U8471 ( .A(B[870]), .B(A[870]), .Z(n762) );
  AND U8472 ( .A(B[871]), .B(A[871]), .Z(n759) );
  NAND U8473 ( .A(n7733), .B(n7734), .Z(n733) );
  AND U8474 ( .A(n751), .B(n747), .Z(n7734) );
  OR U8475 ( .A(B[872]), .B(A[872]), .Z(n751) );
  AND U8476 ( .A(n742), .B(n738), .Z(n7733) );
  NANDN U8477 ( .A(n737), .B(n7735), .Z(n731) );
  NAND U8478 ( .A(n7736), .B(n738), .Z(n7735) );
  OR U8479 ( .A(B[875]), .B(A[875]), .Z(n738) );
  NANDN U8480 ( .A(n740), .B(n7737), .Z(n7736) );
  NAND U8481 ( .A(n7738), .B(n742), .Z(n7737) );
  OR U8482 ( .A(B[874]), .B(A[874]), .Z(n742) );
  NANDN U8483 ( .A(n744), .B(n7739), .Z(n7738) );
  NAND U8484 ( .A(n747), .B(n749), .Z(n7739) );
  AND U8485 ( .A(B[872]), .B(A[872]), .Z(n749) );
  OR U8486 ( .A(B[873]), .B(A[873]), .Z(n747) );
  AND U8487 ( .A(B[873]), .B(A[873]), .Z(n744) );
  AND U8488 ( .A(B[874]), .B(A[874]), .Z(n740) );
  AND U8489 ( .A(B[875]), .B(A[875]), .Z(n737) );
  NOR U8490 ( .A(B[877]), .B(A[877]), .Z(n723) );
  AND U8491 ( .A(B[877]), .B(A[877]), .Z(n721) );
  NOR U8492 ( .A(B[878]), .B(A[878]), .Z(n718) );
  AND U8493 ( .A(B[878]), .B(A[878]), .Z(n717) );
  NOR U8494 ( .A(B[879]), .B(A[879]), .Z(n714) );
  NOR U8495 ( .A(n684), .B(n635), .Z(n5619) );
  NAND U8496 ( .A(n7740), .B(n7741), .Z(n684) );
  AND U8497 ( .A(n702), .B(n698), .Z(n7741) );
  OR U8498 ( .A(B[880]), .B(A[880]), .Z(n702) );
  ANDN U8499 ( .B(n689), .A(n692), .Z(n7740) );
  ANDN U8500 ( .B(n7742), .A(n628), .Z(n5617) );
  AND U8501 ( .A(B[892]), .B(A[892]), .Z(n628) );
  NAND U8502 ( .A(n7743), .B(n631), .Z(n7742) );
  OR U8503 ( .A(A[892]), .B(B[892]), .Z(n631) );
  NANDN U8504 ( .A(n633), .B(n7744), .Z(n7743) );
  NANDN U8505 ( .A(n635), .B(n7745), .Z(n7744) );
  NANDN U8506 ( .A(n660), .B(n7746), .Z(n7745) );
  NAND U8507 ( .A(n683), .B(n663), .Z(n7746) );
  AND U8508 ( .A(n7747), .B(n7748), .Z(n663) );
  AND U8509 ( .A(n680), .B(n676), .Z(n7748) );
  OR U8510 ( .A(B[884]), .B(A[884]), .Z(n680) );
  AND U8511 ( .A(n671), .B(n667), .Z(n7747) );
  NANDN U8512 ( .A(n688), .B(n7749), .Z(n683) );
  NAND U8513 ( .A(n7750), .B(n689), .Z(n7749) );
  OR U8514 ( .A(B[883]), .B(A[883]), .Z(n689) );
  NANDN U8515 ( .A(n691), .B(n7751), .Z(n7750) );
  NANDN U8516 ( .A(n692), .B(n7752), .Z(n7751) );
  NANDN U8517 ( .A(n695), .B(n7753), .Z(n7752) );
  NAND U8518 ( .A(n698), .B(n700), .Z(n7753) );
  AND U8519 ( .A(A[880]), .B(B[880]), .Z(n700) );
  OR U8520 ( .A(B[881]), .B(A[881]), .Z(n698) );
  AND U8521 ( .A(B[881]), .B(A[881]), .Z(n695) );
  NOR U8522 ( .A(B[882]), .B(A[882]), .Z(n692) );
  AND U8523 ( .A(B[882]), .B(A[882]), .Z(n691) );
  AND U8524 ( .A(B[883]), .B(A[883]), .Z(n688) );
  NANDN U8525 ( .A(n666), .B(n7754), .Z(n660) );
  NAND U8526 ( .A(n7755), .B(n667), .Z(n7754) );
  OR U8527 ( .A(B[887]), .B(A[887]), .Z(n667) );
  NANDN U8528 ( .A(n669), .B(n7756), .Z(n7755) );
  NAND U8529 ( .A(n7757), .B(n671), .Z(n7756) );
  OR U8530 ( .A(B[886]), .B(A[886]), .Z(n671) );
  NANDN U8531 ( .A(n673), .B(n7758), .Z(n7757) );
  NAND U8532 ( .A(n676), .B(n678), .Z(n7758) );
  AND U8533 ( .A(B[884]), .B(A[884]), .Z(n678) );
  OR U8534 ( .A(B[885]), .B(A[885]), .Z(n676) );
  AND U8535 ( .A(B[885]), .B(A[885]), .Z(n673) );
  AND U8536 ( .A(B[886]), .B(A[886]), .Z(n669) );
  AND U8537 ( .A(B[887]), .B(A[887]), .Z(n666) );
  NAND U8538 ( .A(n7759), .B(n7760), .Z(n635) );
  AND U8539 ( .A(n658), .B(n649), .Z(n7760) );
  OR U8540 ( .A(B[888]), .B(A[888]), .Z(n658) );
  AND U8541 ( .A(n644), .B(n640), .Z(n7759) );
  NANDN U8542 ( .A(n639), .B(n7761), .Z(n633) );
  NAND U8543 ( .A(n7762), .B(n640), .Z(n7761) );
  OR U8544 ( .A(B[891]), .B(A[891]), .Z(n640) );
  NANDN U8545 ( .A(n642), .B(n7763), .Z(n7762) );
  NAND U8546 ( .A(n7764), .B(n644), .Z(n7763) );
  OR U8547 ( .A(B[890]), .B(A[890]), .Z(n644) );
  NANDN U8548 ( .A(n646), .B(n7765), .Z(n7764) );
  NAND U8549 ( .A(n649), .B(n656), .Z(n7765) );
  AND U8550 ( .A(B[888]), .B(A[888]), .Z(n656) );
  OR U8551 ( .A(B[889]), .B(A[889]), .Z(n649) );
  AND U8552 ( .A(B[889]), .B(A[889]), .Z(n646) );
  AND U8553 ( .A(B[890]), .B(A[890]), .Z(n642) );
  AND U8554 ( .A(B[891]), .B(A[891]), .Z(n639) );
  NOR U8555 ( .A(B[893]), .B(A[893]), .Z(n625) );
  AND U8556 ( .A(B[893]), .B(A[893]), .Z(n623) );
  NOR U8557 ( .A(B[894]), .B(A[894]), .Z(n620) );
  AND U8558 ( .A(B[894]), .B(A[894]), .Z(n619) );
  NOR U8559 ( .A(B[895]), .B(A[895]), .Z(n616) );
  NOR U8560 ( .A(n586), .B(n542), .Z(n5608) );
  NAND U8561 ( .A(n7766), .B(n7767), .Z(n586) );
  AND U8562 ( .A(n612), .B(n608), .Z(n7767) );
  OR U8563 ( .A(B[896]), .B(A[896]), .Z(n612) );
  ANDN U8564 ( .B(n599), .A(n602), .Z(n7766) );
  ANDN U8565 ( .B(n7768), .A(n535), .Z(n5606) );
  AND U8566 ( .A(B[908]), .B(A[908]), .Z(n535) );
  NAND U8567 ( .A(n7769), .B(n538), .Z(n7768) );
  OR U8568 ( .A(A[908]), .B(B[908]), .Z(n538) );
  NANDN U8569 ( .A(n540), .B(n7770), .Z(n7769) );
  NANDN U8570 ( .A(n542), .B(n7771), .Z(n7770) );
  NANDN U8571 ( .A(n562), .B(n7772), .Z(n7771) );
  NAND U8572 ( .A(n585), .B(n565), .Z(n7772) );
  AND U8573 ( .A(n7773), .B(n7774), .Z(n565) );
  AND U8574 ( .A(n582), .B(n578), .Z(n7774) );
  OR U8575 ( .A(B[900]), .B(A[900]), .Z(n582) );
  AND U8576 ( .A(n573), .B(n569), .Z(n7773) );
  NANDN U8577 ( .A(n598), .B(n7775), .Z(n585) );
  NAND U8578 ( .A(n7776), .B(n599), .Z(n7775) );
  OR U8579 ( .A(B[899]), .B(A[899]), .Z(n599) );
  NANDN U8580 ( .A(n601), .B(n7777), .Z(n7776) );
  NANDN U8581 ( .A(n602), .B(n7778), .Z(n7777) );
  NANDN U8582 ( .A(n605), .B(n7779), .Z(n7778) );
  NAND U8583 ( .A(n608), .B(n610), .Z(n7779) );
  AND U8584 ( .A(A[896]), .B(B[896]), .Z(n610) );
  OR U8585 ( .A(B[897]), .B(A[897]), .Z(n608) );
  AND U8586 ( .A(B[897]), .B(A[897]), .Z(n605) );
  NOR U8587 ( .A(B[898]), .B(A[898]), .Z(n602) );
  AND U8588 ( .A(B[898]), .B(A[898]), .Z(n601) );
  AND U8589 ( .A(B[899]), .B(A[899]), .Z(n598) );
  NANDN U8590 ( .A(n568), .B(n7780), .Z(n562) );
  NAND U8591 ( .A(n7781), .B(n569), .Z(n7780) );
  OR U8592 ( .A(B[903]), .B(A[903]), .Z(n569) );
  NANDN U8593 ( .A(n571), .B(n7782), .Z(n7781) );
  NAND U8594 ( .A(n7783), .B(n573), .Z(n7782) );
  OR U8595 ( .A(B[902]), .B(A[902]), .Z(n573) );
  NANDN U8596 ( .A(n575), .B(n7784), .Z(n7783) );
  NAND U8597 ( .A(n578), .B(n580), .Z(n7784) );
  AND U8598 ( .A(B[900]), .B(A[900]), .Z(n580) );
  OR U8599 ( .A(B[901]), .B(A[901]), .Z(n578) );
  AND U8600 ( .A(B[901]), .B(A[901]), .Z(n575) );
  AND U8601 ( .A(B[902]), .B(A[902]), .Z(n571) );
  AND U8602 ( .A(B[903]), .B(A[903]), .Z(n568) );
  NAND U8603 ( .A(n7785), .B(n7786), .Z(n542) );
  AND U8604 ( .A(n560), .B(n556), .Z(n7786) );
  OR U8605 ( .A(B[904]), .B(A[904]), .Z(n560) );
  AND U8606 ( .A(n551), .B(n547), .Z(n7785) );
  NANDN U8607 ( .A(n546), .B(n7787), .Z(n540) );
  NAND U8608 ( .A(n7788), .B(n547), .Z(n7787) );
  OR U8609 ( .A(B[907]), .B(A[907]), .Z(n547) );
  NANDN U8610 ( .A(n549), .B(n7789), .Z(n7788) );
  NAND U8611 ( .A(n7790), .B(n551), .Z(n7789) );
  OR U8612 ( .A(B[906]), .B(A[906]), .Z(n551) );
  NANDN U8613 ( .A(n553), .B(n7791), .Z(n7790) );
  NAND U8614 ( .A(n556), .B(n558), .Z(n7791) );
  AND U8615 ( .A(B[904]), .B(A[904]), .Z(n558) );
  OR U8616 ( .A(B[905]), .B(A[905]), .Z(n556) );
  AND U8617 ( .A(B[905]), .B(A[905]), .Z(n553) );
  AND U8618 ( .A(B[906]), .B(A[906]), .Z(n549) );
  AND U8619 ( .A(B[907]), .B(A[907]), .Z(n546) );
  NOR U8620 ( .A(B[909]), .B(A[909]), .Z(n527) );
  AND U8621 ( .A(B[909]), .B(A[909]), .Z(n525) );
  NOR U8622 ( .A(B[910]), .B(A[910]), .Z(n522) );
  AND U8623 ( .A(B[910]), .B(A[910]), .Z(n521) );
  NOR U8624 ( .A(B[911]), .B(A[911]), .Z(n518) );
  NOR U8625 ( .A(n496), .B(n444), .Z(n5597) );
  NAND U8626 ( .A(n7792), .B(n7793), .Z(n496) );
  AND U8627 ( .A(n514), .B(n510), .Z(n7793) );
  OR U8628 ( .A(B[912]), .B(A[912]), .Z(n514) );
  ANDN U8629 ( .B(n501), .A(n504), .Z(n7792) );
  ANDN U8630 ( .B(n7794), .A(n437), .Z(n5595) );
  AND U8631 ( .A(B[924]), .B(A[924]), .Z(n437) );
  NAND U8632 ( .A(n7795), .B(n440), .Z(n7794) );
  OR U8633 ( .A(A[924]), .B(B[924]), .Z(n440) );
  NANDN U8634 ( .A(n442), .B(n7796), .Z(n7795) );
  NANDN U8635 ( .A(n444), .B(n7797), .Z(n7796) );
  NANDN U8636 ( .A(n464), .B(n7798), .Z(n7797) );
  NAND U8637 ( .A(n495), .B(n467), .Z(n7798) );
  AND U8638 ( .A(n7799), .B(n7800), .Z(n467) );
  AND U8639 ( .A(n492), .B(n488), .Z(n7800) );
  OR U8640 ( .A(B[916]), .B(A[916]), .Z(n492) );
  AND U8641 ( .A(n483), .B(n479), .Z(n7799) );
  NANDN U8642 ( .A(n500), .B(n7801), .Z(n495) );
  NAND U8643 ( .A(n7802), .B(n501), .Z(n7801) );
  OR U8644 ( .A(B[915]), .B(A[915]), .Z(n501) );
  NANDN U8645 ( .A(n503), .B(n7803), .Z(n7802) );
  NANDN U8646 ( .A(n504), .B(n7804), .Z(n7803) );
  NANDN U8647 ( .A(n507), .B(n7805), .Z(n7804) );
  NAND U8648 ( .A(n510), .B(n512), .Z(n7805) );
  AND U8649 ( .A(A[912]), .B(B[912]), .Z(n512) );
  OR U8650 ( .A(B[913]), .B(A[913]), .Z(n510) );
  AND U8651 ( .A(B[913]), .B(A[913]), .Z(n507) );
  NOR U8652 ( .A(B[914]), .B(A[914]), .Z(n504) );
  AND U8653 ( .A(B[914]), .B(A[914]), .Z(n503) );
  AND U8654 ( .A(B[915]), .B(A[915]), .Z(n500) );
  NANDN U8655 ( .A(n478), .B(n7806), .Z(n464) );
  NAND U8656 ( .A(n7807), .B(n479), .Z(n7806) );
  OR U8657 ( .A(B[919]), .B(A[919]), .Z(n479) );
  NANDN U8658 ( .A(n481), .B(n7808), .Z(n7807) );
  NAND U8659 ( .A(n7809), .B(n483), .Z(n7808) );
  OR U8660 ( .A(B[918]), .B(A[918]), .Z(n483) );
  NANDN U8661 ( .A(n485), .B(n7810), .Z(n7809) );
  NAND U8662 ( .A(n488), .B(n490), .Z(n7810) );
  AND U8663 ( .A(B[916]), .B(A[916]), .Z(n490) );
  OR U8664 ( .A(B[917]), .B(A[917]), .Z(n488) );
  AND U8665 ( .A(B[917]), .B(A[917]), .Z(n485) );
  AND U8666 ( .A(B[918]), .B(A[918]), .Z(n481) );
  AND U8667 ( .A(B[919]), .B(A[919]), .Z(n478) );
  NAND U8668 ( .A(n7811), .B(n7812), .Z(n444) );
  AND U8669 ( .A(n462), .B(n458), .Z(n7812) );
  OR U8670 ( .A(B[920]), .B(A[920]), .Z(n462) );
  AND U8671 ( .A(n453), .B(n449), .Z(n7811) );
  NANDN U8672 ( .A(n448), .B(n7813), .Z(n442) );
  NAND U8673 ( .A(n7814), .B(n449), .Z(n7813) );
  OR U8674 ( .A(B[923]), .B(A[923]), .Z(n449) );
  NANDN U8675 ( .A(n451), .B(n7815), .Z(n7814) );
  NAND U8676 ( .A(n7816), .B(n453), .Z(n7815) );
  OR U8677 ( .A(B[922]), .B(A[922]), .Z(n453) );
  NANDN U8678 ( .A(n455), .B(n7817), .Z(n7816) );
  NAND U8679 ( .A(n458), .B(n460), .Z(n7817) );
  AND U8680 ( .A(B[920]), .B(A[920]), .Z(n460) );
  OR U8681 ( .A(B[921]), .B(A[921]), .Z(n458) );
  AND U8682 ( .A(B[921]), .B(A[921]), .Z(n455) );
  AND U8683 ( .A(B[922]), .B(A[922]), .Z(n451) );
  AND U8684 ( .A(B[923]), .B(A[923]), .Z(n448) );
  NOR U8685 ( .A(B[925]), .B(A[925]), .Z(n434) );
  AND U8686 ( .A(B[925]), .B(A[925]), .Z(n432) );
  NOR U8687 ( .A(B[926]), .B(A[926]), .Z(n429) );
  AND U8688 ( .A(B[926]), .B(A[926]), .Z(n428) );
  NOR U8689 ( .A(B[927]), .B(A[927]), .Z(n425) );
  NOR U8690 ( .A(n398), .B(n349), .Z(n5586) );
  NAND U8691 ( .A(n7818), .B(n7819), .Z(n398) );
  AND U8692 ( .A(n421), .B(n412), .Z(n7819) );
  OR U8693 ( .A(B[928]), .B(A[928]), .Z(n421) );
  ANDN U8694 ( .B(n403), .A(n406), .Z(n7818) );
  ANDN U8695 ( .B(n7820), .A(n342), .Z(n5584) );
  AND U8696 ( .A(B[940]), .B(A[940]), .Z(n342) );
  NAND U8697 ( .A(n7821), .B(n345), .Z(n7820) );
  OR U8698 ( .A(A[940]), .B(B[940]), .Z(n345) );
  NANDN U8699 ( .A(n347), .B(n7822), .Z(n7821) );
  NANDN U8700 ( .A(n349), .B(n7823), .Z(n7822) );
  NANDN U8701 ( .A(n374), .B(n7824), .Z(n7823) );
  NAND U8702 ( .A(n397), .B(n377), .Z(n7824) );
  AND U8703 ( .A(n7825), .B(n7826), .Z(n377) );
  AND U8704 ( .A(n394), .B(n390), .Z(n7826) );
  OR U8705 ( .A(B[932]), .B(A[932]), .Z(n394) );
  AND U8706 ( .A(n385), .B(n381), .Z(n7825) );
  NANDN U8707 ( .A(n402), .B(n7827), .Z(n397) );
  NAND U8708 ( .A(n7828), .B(n403), .Z(n7827) );
  OR U8709 ( .A(B[931]), .B(A[931]), .Z(n403) );
  NANDN U8710 ( .A(n405), .B(n7829), .Z(n7828) );
  NANDN U8711 ( .A(n406), .B(n7830), .Z(n7829) );
  NANDN U8712 ( .A(n409), .B(n7831), .Z(n7830) );
  NAND U8713 ( .A(n412), .B(n419), .Z(n7831) );
  AND U8714 ( .A(A[928]), .B(B[928]), .Z(n419) );
  OR U8715 ( .A(B[929]), .B(A[929]), .Z(n412) );
  AND U8716 ( .A(B[929]), .B(A[929]), .Z(n409) );
  NOR U8717 ( .A(B[930]), .B(A[930]), .Z(n406) );
  AND U8718 ( .A(B[930]), .B(A[930]), .Z(n405) );
  AND U8719 ( .A(B[931]), .B(A[931]), .Z(n402) );
  NANDN U8720 ( .A(n380), .B(n7832), .Z(n374) );
  NAND U8721 ( .A(n7833), .B(n381), .Z(n7832) );
  OR U8722 ( .A(B[935]), .B(A[935]), .Z(n381) );
  NANDN U8723 ( .A(n383), .B(n7834), .Z(n7833) );
  NAND U8724 ( .A(n7835), .B(n385), .Z(n7834) );
  OR U8725 ( .A(B[934]), .B(A[934]), .Z(n385) );
  NANDN U8726 ( .A(n387), .B(n7836), .Z(n7835) );
  NAND U8727 ( .A(n390), .B(n392), .Z(n7836) );
  AND U8728 ( .A(B[932]), .B(A[932]), .Z(n392) );
  OR U8729 ( .A(B[933]), .B(A[933]), .Z(n390) );
  AND U8730 ( .A(B[933]), .B(A[933]), .Z(n387) );
  AND U8731 ( .A(B[934]), .B(A[934]), .Z(n383) );
  AND U8732 ( .A(B[935]), .B(A[935]), .Z(n380) );
  NAND U8733 ( .A(n7837), .B(n7838), .Z(n349) );
  AND U8734 ( .A(n372), .B(n368), .Z(n7838) );
  OR U8735 ( .A(B[936]), .B(A[936]), .Z(n372) );
  AND U8736 ( .A(n363), .B(n359), .Z(n7837) );
  NANDN U8737 ( .A(n358), .B(n7839), .Z(n347) );
  NAND U8738 ( .A(n7840), .B(n359), .Z(n7839) );
  OR U8739 ( .A(B[939]), .B(A[939]), .Z(n359) );
  NANDN U8740 ( .A(n361), .B(n7841), .Z(n7840) );
  NAND U8741 ( .A(n7842), .B(n363), .Z(n7841) );
  OR U8742 ( .A(B[938]), .B(A[938]), .Z(n363) );
  NANDN U8743 ( .A(n365), .B(n7843), .Z(n7842) );
  NAND U8744 ( .A(n368), .B(n370), .Z(n7843) );
  AND U8745 ( .A(B[936]), .B(A[936]), .Z(n370) );
  OR U8746 ( .A(B[937]), .B(A[937]), .Z(n368) );
  AND U8747 ( .A(B[937]), .B(A[937]), .Z(n365) );
  AND U8748 ( .A(B[938]), .B(A[938]), .Z(n361) );
  AND U8749 ( .A(B[939]), .B(A[939]), .Z(n358) );
  NOR U8750 ( .A(B[941]), .B(A[941]), .Z(n339) );
  AND U8751 ( .A(B[941]), .B(A[941]), .Z(n337) );
  NOR U8752 ( .A(B[942]), .B(A[942]), .Z(n334) );
  AND U8753 ( .A(B[942]), .B(A[942]), .Z(n333) );
  NOR U8754 ( .A(B[943]), .B(A[943]), .Z(n330) );
  NOR U8755 ( .A(n308), .B(n259), .Z(n5575) );
  NAND U8756 ( .A(n7844), .B(n7845), .Z(n308) );
  AND U8757 ( .A(n326), .B(n322), .Z(n7845) );
  OR U8758 ( .A(B[944]), .B(A[944]), .Z(n326) );
  ANDN U8759 ( .B(n313), .A(n316), .Z(n7844) );
  ANDN U8760 ( .B(n7846), .A(n252), .Z(n5573) );
  AND U8761 ( .A(B[956]), .B(A[956]), .Z(n252) );
  NAND U8762 ( .A(n7847), .B(n255), .Z(n7846) );
  OR U8763 ( .A(A[956]), .B(B[956]), .Z(n255) );
  NANDN U8764 ( .A(n257), .B(n7848), .Z(n7847) );
  NANDN U8765 ( .A(n259), .B(n7849), .Z(n7848) );
  NANDN U8766 ( .A(n279), .B(n7850), .Z(n7849) );
  NAND U8767 ( .A(n307), .B(n282), .Z(n7850) );
  AND U8768 ( .A(n7851), .B(n7852), .Z(n282) );
  AND U8769 ( .A(n304), .B(n295), .Z(n7852) );
  OR U8770 ( .A(B[948]), .B(A[948]), .Z(n304) );
  AND U8771 ( .A(n290), .B(n286), .Z(n7851) );
  NANDN U8772 ( .A(n312), .B(n7853), .Z(n307) );
  NAND U8773 ( .A(n7854), .B(n313), .Z(n7853) );
  OR U8774 ( .A(B[947]), .B(A[947]), .Z(n313) );
  NANDN U8775 ( .A(n315), .B(n7855), .Z(n7854) );
  NANDN U8776 ( .A(n316), .B(n7856), .Z(n7855) );
  NANDN U8777 ( .A(n319), .B(n7857), .Z(n7856) );
  NAND U8778 ( .A(n322), .B(n324), .Z(n7857) );
  AND U8779 ( .A(A[944]), .B(B[944]), .Z(n324) );
  OR U8780 ( .A(B[945]), .B(A[945]), .Z(n322) );
  AND U8781 ( .A(B[945]), .B(A[945]), .Z(n319) );
  NOR U8782 ( .A(B[946]), .B(A[946]), .Z(n316) );
  AND U8783 ( .A(B[946]), .B(A[946]), .Z(n315) );
  AND U8784 ( .A(B[947]), .B(A[947]), .Z(n312) );
  NANDN U8785 ( .A(n285), .B(n7858), .Z(n279) );
  NAND U8786 ( .A(n7859), .B(n286), .Z(n7858) );
  OR U8787 ( .A(B[951]), .B(A[951]), .Z(n286) );
  NANDN U8788 ( .A(n288), .B(n7860), .Z(n7859) );
  NAND U8789 ( .A(n7861), .B(n290), .Z(n7860) );
  OR U8790 ( .A(B[950]), .B(A[950]), .Z(n290) );
  NANDN U8791 ( .A(n292), .B(n7862), .Z(n7861) );
  NAND U8792 ( .A(n295), .B(n302), .Z(n7862) );
  AND U8793 ( .A(B[948]), .B(A[948]), .Z(n302) );
  OR U8794 ( .A(B[949]), .B(A[949]), .Z(n295) );
  AND U8795 ( .A(B[949]), .B(A[949]), .Z(n292) );
  AND U8796 ( .A(B[950]), .B(A[950]), .Z(n288) );
  AND U8797 ( .A(B[951]), .B(A[951]), .Z(n285) );
  NAND U8798 ( .A(n7863), .B(n7864), .Z(n259) );
  AND U8799 ( .A(n277), .B(n273), .Z(n7864) );
  OR U8800 ( .A(B[952]), .B(A[952]), .Z(n277) );
  AND U8801 ( .A(n268), .B(n264), .Z(n7863) );
  NANDN U8802 ( .A(n263), .B(n7865), .Z(n257) );
  NAND U8803 ( .A(n7866), .B(n264), .Z(n7865) );
  OR U8804 ( .A(B[955]), .B(A[955]), .Z(n264) );
  NANDN U8805 ( .A(n266), .B(n7867), .Z(n7866) );
  NAND U8806 ( .A(n7868), .B(n268), .Z(n7867) );
  OR U8807 ( .A(B[954]), .B(A[954]), .Z(n268) );
  NANDN U8808 ( .A(n270), .B(n7869), .Z(n7868) );
  NAND U8809 ( .A(n273), .B(n275), .Z(n7869) );
  AND U8810 ( .A(B[952]), .B(A[952]), .Z(n275) );
  OR U8811 ( .A(B[953]), .B(A[953]), .Z(n273) );
  AND U8812 ( .A(B[953]), .B(A[953]), .Z(n270) );
  AND U8813 ( .A(B[954]), .B(A[954]), .Z(n266) );
  AND U8814 ( .A(B[955]), .B(A[955]), .Z(n263) );
  NOR U8815 ( .A(B[957]), .B(A[957]), .Z(n249) );
  AND U8816 ( .A(B[957]), .B(A[957]), .Z(n247) );
  NOR U8817 ( .A(B[958]), .B(A[958]), .Z(n244) );
  AND U8818 ( .A(B[958]), .B(A[958]), .Z(n243) );
  NOR U8819 ( .A(B[959]), .B(A[959]), .Z(n240) );
  OR U8820 ( .A(A[961]), .B(B[961]), .Z(n223) );
  AND U8821 ( .A(n218), .B(n214), .Z(n5564) );
  OR U8822 ( .A(B[963]), .B(A[963]), .Z(n214) );
  OR U8823 ( .A(A[962]), .B(B[962]), .Z(n218) );
  NAND U8824 ( .A(n7870), .B(n7871), .Z(n189) );
  AND U8825 ( .A(n207), .B(n203), .Z(n7871) );
  OR U8826 ( .A(A[964]), .B(B[964]), .Z(n207) );
  AND U8827 ( .A(n198), .B(n194), .Z(n7870) );
  NANDN U8828 ( .A(n193), .B(n7872), .Z(n187) );
  NAND U8829 ( .A(n7873), .B(n194), .Z(n7872) );
  OR U8830 ( .A(B[967]), .B(A[967]), .Z(n194) );
  NANDN U8831 ( .A(n196), .B(n7874), .Z(n7873) );
  NAND U8832 ( .A(n7875), .B(n198), .Z(n7874) );
  OR U8833 ( .A(A[966]), .B(B[966]), .Z(n198) );
  NANDN U8834 ( .A(n200), .B(n7876), .Z(n7875) );
  NAND U8835 ( .A(n203), .B(n205), .Z(n7876) );
  AND U8836 ( .A(A[964]), .B(B[964]), .Z(n205) );
  OR U8837 ( .A(A[965]), .B(B[965]), .Z(n203) );
  AND U8838 ( .A(A[965]), .B(B[965]), .Z(n200) );
  AND U8839 ( .A(A[966]), .B(B[966]), .Z(n196) );
  AND U8840 ( .A(B[967]), .B(A[967]), .Z(n193) );
  NAND U8841 ( .A(n7877), .B(n7878), .Z(n166) );
  AND U8842 ( .A(n185), .B(n180), .Z(n7878) );
  OR U8843 ( .A(B[968]), .B(A[968]), .Z(n185) );
  AND U8844 ( .A(n175), .B(n171), .Z(n7877) );
  NANDN U8845 ( .A(n170), .B(n7879), .Z(n164) );
  NAND U8846 ( .A(n7880), .B(n171), .Z(n7879) );
  OR U8847 ( .A(B[971]), .B(A[971]), .Z(n171) );
  NANDN U8848 ( .A(n173), .B(n7881), .Z(n7880) );
  NAND U8849 ( .A(n7882), .B(n175), .Z(n7881) );
  OR U8850 ( .A(B[970]), .B(A[970]), .Z(n175) );
  NANDN U8851 ( .A(n177), .B(n7883), .Z(n7882) );
  NAND U8852 ( .A(n180), .B(n183), .Z(n7883) );
  AND U8853 ( .A(B[968]), .B(A[968]), .Z(n183) );
  OR U8854 ( .A(B[969]), .B(A[969]), .Z(n180) );
  AND U8855 ( .A(B[969]), .B(A[969]), .Z(n177) );
  AND U8856 ( .A(B[970]), .B(A[970]), .Z(n173) );
  AND U8857 ( .A(B[971]), .B(A[971]), .Z(n170) );
  NOR U8858 ( .A(B[972]), .B(A[972]), .Z(n161) );
  AND U8859 ( .A(B[972]), .B(A[972]), .Z(n159) );
  NOR U8860 ( .A(B[973]), .B(A[973]), .Z(n156) );
  AND U8861 ( .A(B[973]), .B(A[973]), .Z(n154) );
  NOR U8862 ( .A(B[974]), .B(A[974]), .Z(n151) );
  AND U8863 ( .A(B[974]), .B(A[974]), .Z(n150) );
  NOR U8864 ( .A(B[975]), .B(A[975]), .Z(n147) );
  OR U8865 ( .A(A[977]), .B(B[977]), .Z(n138) );
  AND U8866 ( .A(n133), .B(n129), .Z(n5543) );
  OR U8867 ( .A(B[979]), .B(A[979]), .Z(n129) );
  OR U8868 ( .A(A[978]), .B(B[978]), .Z(n133) );
  NAND U8869 ( .A(n7884), .B(n7885), .Z(n99) );
  AND U8870 ( .A(n117), .B(n113), .Z(n7885) );
  OR U8871 ( .A(A[980]), .B(B[980]), .Z(n117) );
  AND U8872 ( .A(n108), .B(n104), .Z(n7884) );
  NANDN U8873 ( .A(n103), .B(n7886), .Z(n97) );
  NAND U8874 ( .A(n7887), .B(n104), .Z(n7886) );
  OR U8875 ( .A(B[983]), .B(A[983]), .Z(n104) );
  NANDN U8876 ( .A(n106), .B(n7888), .Z(n7887) );
  NAND U8877 ( .A(n7889), .B(n108), .Z(n7888) );
  OR U8878 ( .A(A[982]), .B(B[982]), .Z(n108) );
  NANDN U8879 ( .A(n110), .B(n7890), .Z(n7889) );
  NAND U8880 ( .A(n113), .B(n115), .Z(n7890) );
  AND U8881 ( .A(A[980]), .B(B[980]), .Z(n115) );
  OR U8882 ( .A(A[981]), .B(B[981]), .Z(n113) );
  AND U8883 ( .A(A[981]), .B(B[981]), .Z(n110) );
  AND U8884 ( .A(A[982]), .B(B[982]), .Z(n106) );
  AND U8885 ( .A(B[983]), .B(A[983]), .Z(n103) );
  NAND U8886 ( .A(n7891), .B(n7892), .Z(n77) );
  AND U8887 ( .A(n95), .B(n91), .Z(n7892) );
  OR U8888 ( .A(B[984]), .B(A[984]), .Z(n95) );
  AND U8889 ( .A(n86), .B(n82), .Z(n7891) );
  NANDN U8890 ( .A(n81), .B(n7893), .Z(n75) );
  NAND U8891 ( .A(n7894), .B(n82), .Z(n7893) );
  OR U8892 ( .A(B[987]), .B(A[987]), .Z(n82) );
  NANDN U8893 ( .A(n84), .B(n7895), .Z(n7894) );
  NAND U8894 ( .A(n7896), .B(n86), .Z(n7895) );
  OR U8895 ( .A(B[986]), .B(A[986]), .Z(n86) );
  NANDN U8896 ( .A(n88), .B(n7897), .Z(n7896) );
  NAND U8897 ( .A(n91), .B(n93), .Z(n7897) );
  AND U8898 ( .A(B[984]), .B(A[984]), .Z(n93) );
  OR U8899 ( .A(B[985]), .B(A[985]), .Z(n91) );
  AND U8900 ( .A(B[985]), .B(A[985]), .Z(n88) );
  AND U8901 ( .A(B[986]), .B(A[986]), .Z(n84) );
  AND U8902 ( .A(B[987]), .B(A[987]), .Z(n81) );
  NOR U8903 ( .A(B[988]), .B(A[988]), .Z(n72) );
  AND U8904 ( .A(B[988]), .B(A[988]), .Z(n70) );
  NOR U8905 ( .A(B[989]), .B(A[989]), .Z(n62) );
  AND U8906 ( .A(B[989]), .B(A[989]), .Z(n60) );
  NOR U8907 ( .A(B[990]), .B(A[990]), .Z(n57) );
  AND U8908 ( .A(B[990]), .B(A[990]), .Z(n56) );
  NOR U8909 ( .A(B[991]), .B(A[991]), .Z(n53) );
  NAND U8910 ( .A(n7898), .B(n7899), .Z(n5475) );
  AND U8911 ( .A(n20), .B(n25), .Z(n7899) );
  AND U8912 ( .A(n16), .B(n30), .Z(n7898) );
  OR U8913 ( .A(B[996]), .B(A[996]), .Z(n30) );
  NANDN U8914 ( .A(n15), .B(n7900), .Z(n5471) );
  NAND U8915 ( .A(n7901), .B(n16), .Z(n7900) );
  OR U8916 ( .A(B[999]), .B(A[999]), .Z(n16) );
  NANDN U8917 ( .A(n18), .B(n7902), .Z(n7901) );
  NAND U8918 ( .A(n7903), .B(n20), .Z(n7902) );
  OR U8919 ( .A(B[998]), .B(A[998]), .Z(n20) );
  NANDN U8920 ( .A(n22), .B(n7904), .Z(n7903) );
  NANDN U8921 ( .A(n27), .B(n25), .Z(n7904) );
  OR U8922 ( .A(B[997]), .B(A[997]), .Z(n25) );
  NAND U8923 ( .A(B[996]), .B(A[996]), .Z(n27) );
  AND U8924 ( .A(B[997]), .B(A[997]), .Z(n22) );
  AND U8925 ( .A(A[998]), .B(B[998]), .Z(n18) );
  AND U8926 ( .A(B[999]), .B(A[999]), .Z(n15) );
  ANDN U8927 ( .B(n7905), .A(n4791), .Z(SUM[0]) );
  AND U8928 ( .A(A[0]), .B(B[0]), .Z(n4791) );
  OR U8929 ( .A(A[0]), .B(B[0]), .Z(n7905) );
endmodule


module mult_N1024_CC512_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [1023:0] A;
  input [1:0] B;
  output [1025:0] PRODUCT;
  input TC;
  wire   \P1[512] , \P1[511] , \P1[510] , \P1[509] , \P1[508] , \P1[507] ,
         \P1[506] , \P1[505] , \P1[504] , \P1[503] , \P1[502] , \P1[501] ,
         \P1[500] , \P1[499] , \P1[498] , \P1[497] , \P1[496] , \P1[495] ,
         \P1[494] , \P1[493] , \P1[492] , \P1[491] , \P1[490] , \P1[489] ,
         \P1[488] , \P1[487] , \P1[486] , \P1[485] , \P1[484] , \P1[483] ,
         \P1[482] , \P1[481] , \P1[480] , \P1[479] , \P1[478] , \P1[477] ,
         \P1[476] , \P1[475] , \P1[474] , \P1[473] , \P1[472] , \P1[471] ,
         \P1[470] , \P1[469] , \P1[468] , \P1[467] , \P1[466] , \P1[465] ,
         \P1[464] , \P1[463] , \P1[462] , \P1[461] , \P1[460] , \P1[459] ,
         \P1[458] , \P1[457] , \P1[456] , \P1[455] , \P1[454] , \P1[453] ,
         \P1[452] , \P1[451] , \P1[450] , \P1[449] , \P1[448] , \P1[447] ,
         \P1[446] , \P1[445] , \P1[444] , \P1[443] , \P1[442] , \P1[441] ,
         \P1[440] , \P1[439] , \P1[438] , \P1[437] , \P1[436] , \P1[435] ,
         \P1[434] , \P1[433] , \P1[432] , \P1[431] , \P1[430] , \P1[429] ,
         \P1[428] , \P1[427] , \P1[426] , \P1[425] , \P1[424] , \P1[423] ,
         \P1[422] , \P1[421] , \P1[420] , \P1[419] , \P1[418] , \P1[417] ,
         \P1[416] , \P1[415] , \P1[414] , \P1[413] , \P1[412] , \P1[411] ,
         \P1[410] , \P1[409] , \P1[408] , \P1[407] , \P1[406] , \P1[405] ,
         \P1[404] , \P1[403] , \P1[402] , \P1[401] , \P1[400] , \P1[399] ,
         \P1[398] , \P1[397] , \P1[396] , \P1[395] , \P1[394] , \P1[393] ,
         \P1[392] , \P1[391] , \P1[390] , \P1[389] , \P1[388] , \P1[387] ,
         \P1[386] , \P1[385] , \P1[384] , \P1[383] , \P1[382] , \P1[381] ,
         \P1[380] , \P1[379] , \P1[378] , \P1[377] , \P1[376] , \P1[375] ,
         \P1[374] , \P1[373] , \P1[372] , \P1[371] , \P1[370] , \P1[369] ,
         \P1[368] , \P1[367] , \P1[366] , \P1[365] , \P1[364] , \P1[363] ,
         \P1[362] , \P1[361] , \P1[360] , \P1[359] , \P1[358] , \P1[357] ,
         \P1[356] , \P1[355] , \P1[354] , \P1[353] , \P1[352] , \P1[351] ,
         \P1[350] , \P1[349] , \P1[348] , \P1[347] , \P1[346] , \P1[345] ,
         \P1[344] , \P1[343] , \P1[342] , \P1[341] , \P1[340] , \P1[339] ,
         \P1[338] , \P1[337] , \P1[336] , \P1[335] , \P1[334] , \P1[333] ,
         \P1[332] , \P1[331] , \P1[330] , \P1[329] , \P1[328] , \P1[327] ,
         \P1[326] , \P1[325] , \P1[324] , \P1[323] , \P1[322] , \P1[321] ,
         \P1[320] , \P1[319] , \P1[318] , \P1[317] , \P1[316] , \P1[315] ,
         \P1[314] , \P1[313] , \P1[312] , \P1[311] , \P1[310] , \P1[309] ,
         \P1[308] , \P1[307] , \P1[306] , \P1[305] , \P1[304] , \P1[303] ,
         \P1[302] , \P1[301] , \P1[300] , \P1[299] , \P1[298] , \P1[297] ,
         \P1[296] , \P1[295] , \P1[294] , \P1[293] , \P1[292] , \P1[291] ,
         \P1[290] , \P1[289] , \P1[288] , \P1[287] , \P1[286] , \P1[285] ,
         \P1[284] , \P1[283] , \P1[282] , \P1[281] , \P1[280] , \P1[279] ,
         \P1[278] , \P1[277] , \P1[276] , \P1[275] , \P1[274] , \P1[273] ,
         \P1[272] , \P1[271] , \P1[270] , \P1[269] , \P1[268] , \P1[267] ,
         \P1[266] , \P1[265] , \P1[264] , \P1[263] , \P1[262] , \P1[261] ,
         \P1[260] , \P1[259] , \P1[258] , \P1[257] , \P1[256] , \P1[255] ,
         \P1[254] , \P1[253] , \P1[252] , \P1[251] , \P1[250] , \P1[249] ,
         \P1[248] , \P1[247] , \P1[246] , \P1[245] , \P1[244] , \P1[243] ,
         \P1[242] , \P1[241] , \P1[240] , \P1[239] , \P1[238] , \P1[237] ,
         \P1[236] , \P1[235] , \P1[234] , \P1[233] , \P1[232] , \P1[231] ,
         \P1[230] , \P1[229] , \P1[228] , \P1[227] , \P1[226] , \P1[225] ,
         \P1[224] , \P1[223] , \P1[222] , \P1[221] , \P1[220] , \P1[219] ,
         \P1[218] , \P1[217] , \P1[216] , \P1[215] , \P1[214] , \P1[213] ,
         \P1[212] , \P1[211] , \P1[210] , \P1[209] , \P1[208] , \P1[207] ,
         \P1[206] , \P1[205] , \P1[204] , \P1[203] , \P1[202] , \P1[201] ,
         \P1[200] , \P1[199] , \P1[198] , \P1[197] , \P1[196] , \P1[195] ,
         \P1[194] , \P1[193] , \P1[192] , \P1[191] , \P1[190] , \P1[189] ,
         \P1[188] , \P1[187] , \P1[186] , \P1[185] , \P1[184] , \P1[183] ,
         \P1[182] , \P1[181] , \P1[180] , \P1[179] , \P1[178] , \P1[177] ,
         \P1[176] , \P1[175] , \P1[174] , \P1[173] , \P1[172] , \P1[171] ,
         \P1[170] , \P1[169] , \P1[168] , \P1[167] , \P1[166] , \P1[165] ,
         \P1[164] , \P1[163] , \P1[162] , \P1[161] , \P1[160] , \P1[159] ,
         \P1[158] , \P1[157] , \P1[156] , \P1[155] , \P1[154] , \P1[153] ,
         \P1[152] , \P1[151] , \P1[150] , \P1[149] , \P1[148] , \P1[147] ,
         \P1[146] , \P1[145] , \P1[144] , \P1[143] , \P1[142] , \P1[141] ,
         \P1[140] , \P1[139] , \P1[138] , \P1[137] , \P1[136] , \P1[135] ,
         \P1[134] , \P1[133] , \P1[132] , \P1[131] , \P1[130] , \P1[129] ,
         \P1[128] , \P1[127] , \P1[126] , \P1[125] , \P1[124] , \P1[123] ,
         \P1[122] , \P1[121] , \P1[120] , \P1[119] , \P1[118] , \P1[117] ,
         \P1[116] , \P1[115] , \P1[114] , \P1[113] , \P1[112] , \P1[111] ,
         \P1[110] , \P1[109] , \P1[108] , \P1[107] , \P1[106] , \P1[105] ,
         \P1[104] , \P1[103] , \P1[102] , \P1[101] , \P1[100] , \P1[99] ,
         \P1[98] , \P1[97] , \P1[96] , \P1[95] , \P1[94] , \P1[93] , \P1[92] ,
         \P1[91] , \P1[90] , \P1[89] , \P1[88] , \P1[87] , \P1[86] , \P1[85] ,
         \P1[84] , \P1[83] , \P1[82] , \P1[81] , \P1[80] , \P1[79] , \P1[78] ,
         \P1[77] , \P1[76] , \P1[75] , \P1[74] , \P1[73] , \P1[72] , \P1[71] ,
         \P1[70] , \P1[69] , \P1[68] , \P1[67] , \P1[66] , \P1[65] , \P1[64] ,
         \P1[63] , \P1[62] , \P1[61] , \P1[60] , \P1[59] , \P1[58] , \P1[57] ,
         \P1[56] , \P1[55] , \P1[54] , \P1[53] , \P1[52] , \P1[51] , \P1[50] ,
         \P1[49] , \P1[48] , \P1[47] , \P1[46] , \P1[45] , \P1[44] , \P1[43] ,
         \P1[42] , \P1[41] , \P1[40] , \P1[39] , \P1[38] , \P1[37] , \P1[36] ,
         \P1[35] , \P1[34] , \P1[33] , \P1[32] , \P1[31] , \P1[30] , \P1[29] ,
         \P1[28] , \P1[27] , \P1[26] , \P1[25] , \P1[24] , \P1[23] , \P1[22] ,
         \P1[21] , \P1[20] , \P1[19] , \P1[18] , \P1[17] , \P1[16] , \P1[15] ,
         \P1[14] , \P1[13] , \P1[12] , \P1[11] , \P1[10] , \P1[9] , \P1[8] ,
         \P1[7] , \P1[6] , \P1[5] , \P1[4] , \P1[3] , \P1[2] , \P1[1] ,
         \P0[512] , \P0[511] , \P0[510] , \P0[509] , \P0[508] , \P0[507] ,
         \P0[506] , \P0[505] , \P0[504] , \P0[503] , \P0[502] , \P0[501] ,
         \P0[500] , \P0[499] , \P0[498] , \P0[497] , \P0[496] , \P0[495] ,
         \P0[494] , \P0[493] , \P0[492] , \P0[491] , \P0[490] , \P0[489] ,
         \P0[488] , \P0[487] , \P0[486] , \P0[485] , \P0[484] , \P0[483] ,
         \P0[482] , \P0[481] , \P0[480] , \P0[479] , \P0[478] , \P0[477] ,
         \P0[476] , \P0[475] , \P0[474] , \P0[473] , \P0[472] , \P0[471] ,
         \P0[470] , \P0[469] , \P0[468] , \P0[467] , \P0[466] , \P0[465] ,
         \P0[464] , \P0[463] , \P0[462] , \P0[461] , \P0[460] , \P0[459] ,
         \P0[458] , \P0[457] , \P0[456] , \P0[455] , \P0[454] , \P0[453] ,
         \P0[452] , \P0[451] , \P0[450] , \P0[449] , \P0[448] , \P0[447] ,
         \P0[446] , \P0[445] , \P0[444] , \P0[443] , \P0[442] , \P0[441] ,
         \P0[440] , \P0[439] , \P0[438] , \P0[437] , \P0[436] , \P0[435] ,
         \P0[434] , \P0[433] , \P0[432] , \P0[431] , \P0[430] , \P0[429] ,
         \P0[428] , \P0[427] , \P0[426] , \P0[425] , \P0[424] , \P0[423] ,
         \P0[422] , \P0[421] , \P0[420] , \P0[419] , \P0[418] , \P0[417] ,
         \P0[416] , \P0[415] , \P0[414] , \P0[413] , \P0[412] , \P0[411] ,
         \P0[410] , \P0[409] , \P0[408] , \P0[407] , \P0[406] , \P0[405] ,
         \P0[404] , \P0[403] , \P0[402] , \P0[401] , \P0[400] , \P0[399] ,
         \P0[398] , \P0[397] , \P0[396] , \P0[395] , \P0[394] , \P0[393] ,
         \P0[392] , \P0[391] , \P0[390] , \P0[389] , \P0[388] , \P0[387] ,
         \P0[386] , \P0[385] , \P0[384] , \P0[383] , \P0[382] , \P0[381] ,
         \P0[380] , \P0[379] , \P0[378] , \P0[377] , \P0[376] , \P0[375] ,
         \P0[374] , \P0[373] , \P0[372] , \P0[371] , \P0[370] , \P0[369] ,
         \P0[368] , \P0[367] , \P0[366] , \P0[365] , \P0[364] , \P0[363] ,
         \P0[362] , \P0[361] , \P0[360] , \P0[359] , \P0[358] , \P0[357] ,
         \P0[356] , \P0[355] , \P0[354] , \P0[353] , \P0[352] , \P0[351] ,
         \P0[350] , \P0[349] , \P0[348] , \P0[347] , \P0[346] , \P0[345] ,
         \P0[344] , \P0[343] , \P0[342] , \P0[341] , \P0[340] , \P0[339] ,
         \P0[338] , \P0[337] , \P0[336] , \P0[335] , \P0[334] , \P0[333] ,
         \P0[332] , \P0[331] , \P0[330] , \P0[329] , \P0[328] , \P0[327] ,
         \P0[326] , \P0[325] , \P0[324] , \P0[323] , \P0[322] , \P0[321] ,
         \P0[320] , \P0[319] , \P0[318] , \P0[317] , \P0[316] , \P0[315] ,
         \P0[314] , \P0[313] , \P0[312] , \P0[311] , \P0[310] , \P0[309] ,
         \P0[308] , \P0[307] , \P0[306] , \P0[305] , \P0[304] , \P0[303] ,
         \P0[302] , \P0[301] , \P0[300] , \P0[299] , \P0[298] , \P0[297] ,
         \P0[296] , \P0[295] , \P0[294] , \P0[293] , \P0[292] , \P0[291] ,
         \P0[290] , \P0[289] , \P0[288] , \P0[287] , \P0[286] , \P0[285] ,
         \P0[284] , \P0[283] , \P0[282] , \P0[281] , \P0[280] , \P0[279] ,
         \P0[278] , \P0[277] , \P0[276] , \P0[275] , \P0[274] , \P0[273] ,
         \P0[272] , \P0[271] , \P0[270] , \P0[269] , \P0[268] , \P0[267] ,
         \P0[266] , \P0[265] , \P0[264] , \P0[263] , \P0[262] , \P0[261] ,
         \P0[260] , \P0[259] , \P0[258] , \P0[257] , \P0[256] , \P0[255] ,
         \P0[254] , \P0[253] , \P0[252] , \P0[251] , \P0[250] , \P0[249] ,
         \P0[248] , \P0[247] , \P0[246] , \P0[245] , \P0[244] , \P0[243] ,
         \P0[242] , \P0[241] , \P0[240] , \P0[239] , \P0[238] , \P0[237] ,
         \P0[236] , \P0[235] , \P0[234] , \P0[233] , \P0[232] , \P0[231] ,
         \P0[230] , \P0[229] , \P0[228] , \P0[227] , \P0[226] , \P0[225] ,
         \P0[224] , \P0[223] , \P0[222] , \P0[221] , \P0[220] , \P0[219] ,
         \P0[218] , \P0[217] , \P0[216] , \P0[215] , \P0[214] , \P0[213] ,
         \P0[212] , \P0[211] , \P0[210] , \P0[209] , \P0[208] , \P0[207] ,
         \P0[206] , \P0[205] , \P0[204] , \P0[203] , \P0[202] , \P0[201] ,
         \P0[200] , \P0[199] , \P0[198] , \P0[197] , \P0[196] , \P0[195] ,
         \P0[194] , \P0[193] , \P0[192] , \P0[191] , \P0[190] , \P0[189] ,
         \P0[188] , \P0[187] , \P0[186] , \P0[185] , \P0[184] , \P0[183] ,
         \P0[182] , \P0[181] , \P0[180] , \P0[179] , \P0[178] , \P0[177] ,
         \P0[176] , \P0[175] , \P0[174] , \P0[173] , \P0[172] , \P0[171] ,
         \P0[170] , \P0[169] , \P0[168] , \P0[167] , \P0[166] , \P0[165] ,
         \P0[164] , \P0[163] , \P0[162] , \P0[161] , \P0[160] , \P0[159] ,
         \P0[158] , \P0[157] , \P0[156] , \P0[155] , \P0[154] , \P0[153] ,
         \P0[152] , \P0[151] , \P0[150] , \P0[149] , \P0[148] , \P0[147] ,
         \P0[146] , \P0[145] , \P0[144] , \P0[143] , \P0[142] , \P0[141] ,
         \P0[140] , \P0[139] , \P0[138] , \P0[137] , \P0[136] , \P0[135] ,
         \P0[134] , \P0[133] , \P0[132] , \P0[131] , \P0[130] , \P0[129] ,
         \P0[128] , \P0[127] , \P0[126] , \P0[125] , \P0[124] , \P0[123] ,
         \P0[122] , \P0[121] , \P0[120] , \P0[119] , \P0[118] , \P0[117] ,
         \P0[116] , \P0[115] , \P0[114] , \P0[113] , \P0[112] , \P0[111] ,
         \P0[110] , \P0[109] , \P0[108] , \P0[107] , \P0[106] , \P0[105] ,
         \P0[104] , \P0[103] , \P0[102] , \P0[101] , \P0[100] , \P0[99] ,
         \P0[98] , \P0[97] , \P0[96] , \P0[95] , \P0[94] , \P0[93] , \P0[92] ,
         \P0[91] , \P0[90] , \P0[89] , \P0[88] , \P0[87] , \P0[86] , \P0[85] ,
         \P0[84] , \P0[83] , \P0[82] , \P0[81] , \P0[80] , \P0[79] , \P0[78] ,
         \P0[77] , \P0[76] , \P0[75] , \P0[74] , \P0[73] , \P0[72] , \P0[71] ,
         \P0[70] , \P0[69] , \P0[68] , \P0[67] , \P0[66] , \P0[65] , \P0[64] ,
         \P0[63] , \P0[62] , \P0[61] , \P0[60] , \P0[59] , \P0[58] , \P0[57] ,
         \P0[56] , \P0[55] , \P0[54] , \P0[53] , \P0[52] , \P0[51] , \P0[50] ,
         \P0[49] , \P0[48] , \P0[47] , \P0[46] , \P0[45] , \P0[44] , \P0[43] ,
         \P0[42] , \P0[41] , \P0[40] , \P0[39] , \P0[38] , \P0[37] , \P0[36] ,
         \P0[35] , \P0[34] , \P0[33] , \P0[32] , \P0[31] , \P0[30] , \P0[29] ,
         \P0[28] , \P0[27] , \P0[26] , \P0[25] , \P0[24] , \P0[23] , \P0[22] ,
         \P0[21] , \P0[20] , \P0[19] , \P0[18] , \P0[17] , \P0[16] , \P0[15] ,
         \P0[14] , \P0[13] , \P0[12] , \P0[11] , \P0[10] , \P0[9] , \P0[8] ,
         \P0[7] , \P0[6] , \P0[5] , \P0[4] , \P0[3] , \P0[2] , \P0[1] ,
         \P1[1024] , \P1[1023] , \P1[1022] , \P1[1021] , \P1[1020] ,
         \P1[1019] , \P1[1018] , \P1[1017] , \P1[1016] , \P1[1015] ,
         \P1[1014] , \P1[1013] , \P1[1012] , \P1[1011] , \P1[1010] ,
         \P1[1009] , \P1[1008] , \P1[1007] , \P1[1006] , \P1[1005] ,
         \P1[1004] , \P1[1003] , \P1[1002] , \P1[1001] , \P1[1000] , \P1[999] ,
         \P1[998] , \P1[997] , \P1[996] , \P1[995] , \P1[994] , \P1[993] ,
         \P1[992] , \P1[991] , \P1[990] , \P1[989] , \P1[988] , \P1[987] ,
         \P1[986] , \P1[985] , \P1[984] , \P1[983] , \P1[982] , \P1[981] ,
         \P1[980] , \P1[979] , \P1[978] , \P1[977] , \P1[976] , \P1[975] ,
         \P1[974] , \P1[973] , \P1[972] , \P1[971] , \P1[970] , \P1[969] ,
         \P1[968] , \P1[967] , \P1[966] , \P1[965] , \P1[964] , \P1[963] ,
         \P1[962] , \P1[961] , \P1[960] , \P1[959] , \P1[958] , \P1[957] ,
         \P1[956] , \P1[955] , \P1[954] , \P1[953] , \P1[952] , \P1[951] ,
         \P1[950] , \P1[949] , \P1[948] , \P1[947] , \P1[946] , \P1[945] ,
         \P1[944] , \P1[943] , \P1[942] , \P1[941] , \P1[940] , \P1[939] ,
         \P1[938] , \P1[937] , \P1[936] , \P1[935] , \P1[934] , \P1[933] ,
         \P1[932] , \P1[931] , \P1[930] , \P1[929] , \P1[928] , \P1[927] ,
         \P1[926] , \P1[925] , \P1[924] , \P1[923] , \P1[922] , \P1[921] ,
         \P1[920] , \P1[919] , \P1[918] , \P1[917] , \P1[916] , \P1[915] ,
         \P1[914] , \P1[913] , \P1[912] , \P1[911] , \P1[910] , \P1[909] ,
         \P1[908] , \P1[907] , \P1[906] , \P1[905] , \P1[904] , \P1[903] ,
         \P1[902] , \P1[901] , \P1[900] , \P1[899] , \P1[898] , \P1[897] ,
         \P1[896] , \P1[895] , \P1[894] , \P1[893] , \P1[892] , \P1[891] ,
         \P1[890] , \P1[889] , \P1[888] , \P1[887] , \P1[886] , \P1[885] ,
         \P1[884] , \P1[883] , \P1[882] , \P1[881] , \P1[880] , \P1[879] ,
         \P1[878] , \P1[877] , \P1[876] , \P1[875] , \P1[874] , \P1[873] ,
         \P1[872] , \P1[871] , \P1[870] , \P1[869] , \P1[868] , \P1[867] ,
         \P1[866] , \P1[865] , \P1[864] , \P1[863] , \P1[862] , \P1[861] ,
         \P1[860] , \P1[859] , \P1[858] , \P1[857] , \P1[856] , \P1[855] ,
         \P1[854] , \P1[853] , \P1[852] , \P1[851] , \P1[850] , \P1[849] ,
         \P1[848] , \P1[847] , \P1[846] , \P1[845] , \P1[844] , \P1[843] ,
         \P1[842] , \P1[841] , \P1[840] , \P1[839] , \P1[838] , \P1[837] ,
         \P1[836] , \P1[835] , \P1[834] , \P1[833] , \P1[832] , \P1[831] ,
         \P1[830] , \P1[829] , \P1[828] , \P1[827] , \P1[826] , \P1[825] ,
         \P1[824] , \P1[823] , \P1[822] , \P1[821] , \P1[820] , \P1[819] ,
         \P1[818] , \P1[817] , \P1[816] , \P1[815] , \P1[814] , \P1[813] ,
         \P1[812] , \P1[811] , \P1[810] , \P1[809] , \P1[808] , \P1[807] ,
         \P1[806] , \P1[805] , \P1[804] , \P1[803] , \P1[802] , \P1[801] ,
         \P1[800] , \P1[799] , \P1[798] , \P1[797] , \P1[796] , \P1[795] ,
         \P1[794] , \P1[793] , \P1[792] , \P1[791] , \P1[790] , \P1[789] ,
         \P1[788] , \P1[787] , \P1[786] , \P1[785] , \P1[784] , \P1[783] ,
         \P1[782] , \P1[781] , \P1[780] , \P1[779] , \P1[778] , \P1[777] ,
         \P1[776] , \P1[775] , \P1[774] , \P1[773] , \P1[772] , \P1[771] ,
         \P1[770] , \P1[769] , \P1[768] , \P1[767] , \P1[766] , \P1[765] ,
         \P1[764] , \P1[763] , \P1[762] , \P1[761] , \P1[760] , \P1[759] ,
         \P1[758] , \P1[757] , \P1[756] , \P1[755] , \P1[754] , \P1[753] ,
         \P1[752] , \P1[751] , \P1[750] , \P1[749] , \P1[748] , \P1[747] ,
         \P1[746] , \P1[745] , \P1[744] , \P1[743] , \P1[742] , \P1[741] ,
         \P1[740] , \P1[739] , \P1[738] , \P1[737] , \P1[736] , \P1[735] ,
         \P1[734] , \P1[733] , \P1[732] , \P1[731] , \P1[730] , \P1[729] ,
         \P1[728] , \P1[727] , \P1[726] , \P1[725] , \P1[724] , \P1[723] ,
         \P1[722] , \P1[721] , \P1[720] , \P1[719] , \P1[718] , \P1[717] ,
         \P1[716] , \P1[715] , \P1[714] , \P1[713] , \P1[712] , \P1[711] ,
         \P1[710] , \P1[709] , \P1[708] , \P1[707] , \P1[706] , \P1[705] ,
         \P1[704] , \P1[703] , \P1[702] , \P1[701] , \P1[700] , \P1[699] ,
         \P1[698] , \P1[697] , \P1[696] , \P1[695] , \P1[694] , \P1[693] ,
         \P1[692] , \P1[691] , \P1[690] , \P1[689] , \P1[688] , \P1[687] ,
         \P1[686] , \P1[685] , \P1[684] , \P1[683] , \P1[682] , \P1[681] ,
         \P1[680] , \P1[679] , \P1[678] , \P1[677] , \P1[676] , \P1[675] ,
         \P1[674] , \P1[673] , \P1[672] , \P1[671] , \P1[670] , \P1[669] ,
         \P1[668] , \P1[667] , \P1[666] , \P1[665] , \P1[664] , \P1[663] ,
         \P1[662] , \P1[661] , \P1[660] , \P1[659] , \P1[658] , \P1[657] ,
         \P1[656] , \P1[655] , \P1[654] , \P1[653] , \P1[652] , \P1[651] ,
         \P1[650] , \P1[649] , \P1[648] , \P1[647] , \P1[646] , \P1[645] ,
         \P1[644] , \P1[643] , \P1[642] , \P1[641] , \P1[640] , \P1[639] ,
         \P1[638] , \P1[637] , \P1[636] , \P1[635] , \P1[634] , \P1[633] ,
         \P1[632] , \P1[631] , \P1[630] , \P1[629] , \P1[628] , \P1[627] ,
         \P1[626] , \P1[625] , \P1[624] , \P1[623] , \P1[622] , \P1[621] ,
         \P1[620] , \P1[619] , \P1[618] , \P1[617] , \P1[616] , \P1[615] ,
         \P1[614] , \P1[613] , \P1[612] , \P1[611] , \P1[610] , \P1[609] ,
         \P1[608] , \P1[607] , \P1[606] , \P1[605] , \P1[604] , \P1[603] ,
         \P1[602] , \P1[601] , \P1[600] , \P1[599] , \P1[598] , \P1[597] ,
         \P1[596] , \P1[595] , \P1[594] , \P1[593] , \P1[592] , \P1[591] ,
         \P1[590] , \P1[589] , \P1[588] , \P1[587] , \P1[586] , \P1[585] ,
         \P1[584] , \P1[583] , \P1[582] , \P1[581] , \P1[580] , \P1[579] ,
         \P1[578] , \P1[577] , \P1[576] , \P1[575] , \P1[574] , \P1[573] ,
         \P1[572] , \P1[571] , \P1[570] , \P1[569] , \P1[568] , \P1[567] ,
         \P1[566] , \P1[565] , \P1[564] , \P1[563] , \P1[562] , \P1[561] ,
         \P1[560] , \P1[559] , \P1[558] , \P1[557] , \P1[556] , \P1[555] ,
         \P1[554] , \P1[553] , \P1[552] , \P1[551] , \P1[550] , \P1[549] ,
         \P1[548] , \P1[547] , \P1[546] , \P1[545] , \P1[544] , \P1[543] ,
         \P1[542] , \P1[541] , \P1[540] , \P1[539] , \P1[538] , \P1[537] ,
         \P1[536] , \P1[535] , \P1[534] , \P1[533] , \P1[532] , \P1[531] ,
         \P1[530] , \P1[529] , \P1[528] , \P1[527] , \P1[526] , \P1[525] ,
         \P1[524] , \P1[523] , \P1[522] , \P1[521] , \P1[520] , \P1[519] ,
         \P1[518] , \P1[517] , \P1[516] , \P1[515] , \P1[514] , \P1[513] ,
         \P0[1023] , \P0[1022] , \P0[1021] , \P0[1020] , \P0[1019] ,
         \P0[1018] , \P0[1017] , \P0[1016] , \P0[1015] , \P0[1014] ,
         \P0[1013] , \P0[1012] , \P0[1011] , \P0[1010] , \P0[1009] ,
         \P0[1008] , \P0[1007] , \P0[1006] , \P0[1005] , \P0[1004] ,
         \P0[1003] , \P0[1002] , \P0[1001] , \P0[1000] , \P0[999] , \P0[998] ,
         \P0[997] , \P0[996] , \P0[995] , \P0[994] , \P0[993] , \P0[992] ,
         \P0[991] , \P0[990] , \P0[989] , \P0[988] , \P0[987] , \P0[986] ,
         \P0[985] , \P0[984] , \P0[983] , \P0[982] , \P0[981] , \P0[980] ,
         \P0[979] , \P0[978] , \P0[977] , \P0[976] , \P0[975] , \P0[974] ,
         \P0[973] , \P0[972] , \P0[971] , \P0[970] , \P0[969] , \P0[968] ,
         \P0[967] , \P0[966] , \P0[965] , \P0[964] , \P0[963] , \P0[962] ,
         \P0[961] , \P0[960] , \P0[959] , \P0[958] , \P0[957] , \P0[956] ,
         \P0[955] , \P0[954] , \P0[953] , \P0[952] , \P0[951] , \P0[950] ,
         \P0[949] , \P0[948] , \P0[947] , \P0[946] , \P0[945] , \P0[944] ,
         \P0[943] , \P0[942] , \P0[941] , \P0[940] , \P0[939] , \P0[938] ,
         \P0[937] , \P0[936] , \P0[935] , \P0[934] , \P0[933] , \P0[932] ,
         \P0[931] , \P0[930] , \P0[929] , \P0[928] , \P0[927] , \P0[926] ,
         \P0[925] , \P0[924] , \P0[923] , \P0[922] , \P0[921] , \P0[920] ,
         \P0[919] , \P0[918] , \P0[917] , \P0[916] , \P0[915] , \P0[914] ,
         \P0[913] , \P0[912] , \P0[911] , \P0[910] , \P0[909] , \P0[908] ,
         \P0[907] , \P0[906] , \P0[905] , \P0[904] , \P0[903] , \P0[902] ,
         \P0[901] , \P0[900] , \P0[899] , \P0[898] , \P0[897] , \P0[896] ,
         \P0[895] , \P0[894] , \P0[893] , \P0[892] , \P0[891] , \P0[890] ,
         \P0[889] , \P0[888] , \P0[887] , \P0[886] , \P0[885] , \P0[884] ,
         \P0[883] , \P0[882] , \P0[881] , \P0[880] , \P0[879] , \P0[878] ,
         \P0[877] , \P0[876] , \P0[875] , \P0[874] , \P0[873] , \P0[872] ,
         \P0[871] , \P0[870] , \P0[869] , \P0[868] , \P0[867] , \P0[866] ,
         \P0[865] , \P0[864] , \P0[863] , \P0[862] , \P0[861] , \P0[860] ,
         \P0[859] , \P0[858] , \P0[857] , \P0[856] , \P0[855] , \P0[854] ,
         \P0[853] , \P0[852] , \P0[851] , \P0[850] , \P0[849] , \P0[848] ,
         \P0[847] , \P0[846] , \P0[845] , \P0[844] , \P0[843] , \P0[842] ,
         \P0[841] , \P0[840] , \P0[839] , \P0[838] , \P0[837] , \P0[836] ,
         \P0[835] , \P0[834] , \P0[833] , \P0[832] , \P0[831] , \P0[830] ,
         \P0[829] , \P0[828] , \P0[827] , \P0[826] , \P0[825] , \P0[824] ,
         \P0[823] , \P0[822] , \P0[821] , \P0[820] , \P0[819] , \P0[818] ,
         \P0[817] , \P0[816] , \P0[815] , \P0[814] , \P0[813] , \P0[812] ,
         \P0[811] , \P0[810] , \P0[809] , \P0[808] , \P0[807] , \P0[806] ,
         \P0[805] , \P0[804] , \P0[803] , \P0[802] , \P0[801] , \P0[800] ,
         \P0[799] , \P0[798] , \P0[797] , \P0[796] , \P0[795] , \P0[794] ,
         \P0[793] , \P0[792] , \P0[791] , \P0[790] , \P0[789] , \P0[788] ,
         \P0[787] , \P0[786] , \P0[785] , \P0[784] , \P0[783] , \P0[782] ,
         \P0[781] , \P0[780] , \P0[779] , \P0[778] , \P0[777] , \P0[776] ,
         \P0[775] , \P0[774] , \P0[773] , \P0[772] , \P0[771] , \P0[770] ,
         \P0[769] , \P0[768] , \P0[767] , \P0[766] , \P0[765] , \P0[764] ,
         \P0[763] , \P0[762] , \P0[761] , \P0[760] , \P0[759] , \P0[758] ,
         \P0[757] , \P0[756] , \P0[755] , \P0[754] , \P0[753] , \P0[752] ,
         \P0[751] , \P0[750] , \P0[749] , \P0[748] , \P0[747] , \P0[746] ,
         \P0[745] , \P0[744] , \P0[743] , \P0[742] , \P0[741] , \P0[740] ,
         \P0[739] , \P0[738] , \P0[737] , \P0[736] , \P0[735] , \P0[734] ,
         \P0[733] , \P0[732] , \P0[731] , \P0[730] , \P0[729] , \P0[728] ,
         \P0[727] , \P0[726] , \P0[725] , \P0[724] , \P0[723] , \P0[722] ,
         \P0[721] , \P0[720] , \P0[719] , \P0[718] , \P0[717] , \P0[716] ,
         \P0[715] , \P0[714] , \P0[713] , \P0[712] , \P0[711] , \P0[710] ,
         \P0[709] , \P0[708] , \P0[707] , \P0[706] , \P0[705] , \P0[704] ,
         \P0[703] , \P0[702] , \P0[701] , \P0[700] , \P0[699] , \P0[698] ,
         \P0[697] , \P0[696] , \P0[695] , \P0[694] , \P0[693] , \P0[692] ,
         \P0[691] , \P0[690] , \P0[689] , \P0[688] , \P0[687] , \P0[686] ,
         \P0[685] , \P0[684] , \P0[683] , \P0[682] , \P0[681] , \P0[680] ,
         \P0[679] , \P0[678] , \P0[677] , \P0[676] , \P0[675] , \P0[674] ,
         \P0[673] , \P0[672] , \P0[671] , \P0[670] , \P0[669] , \P0[668] ,
         \P0[667] , \P0[666] , \P0[665] , \P0[664] , \P0[663] , \P0[662] ,
         \P0[661] , \P0[660] , \P0[659] , \P0[658] , \P0[657] , \P0[656] ,
         \P0[655] , \P0[654] , \P0[653] , \P0[652] , \P0[651] , \P0[650] ,
         \P0[649] , \P0[648] , \P0[647] , \P0[646] , \P0[645] , \P0[644] ,
         \P0[643] , \P0[642] , \P0[641] , \P0[640] , \P0[639] , \P0[638] ,
         \P0[637] , \P0[636] , \P0[635] , \P0[634] , \P0[633] , \P0[632] ,
         \P0[631] , \P0[630] , \P0[629] , \P0[628] , \P0[627] , \P0[626] ,
         \P0[625] , \P0[624] , \P0[623] , \P0[622] , \P0[621] , \P0[620] ,
         \P0[619] , \P0[618] , \P0[617] , \P0[616] , \P0[615] , \P0[614] ,
         \P0[613] , \P0[612] , \P0[611] , \P0[610] , \P0[609] , \P0[608] ,
         \P0[607] , \P0[606] , \P0[605] , \P0[604] , \P0[603] , \P0[602] ,
         \P0[601] , \P0[600] , \P0[599] , \P0[598] , \P0[597] , \P0[596] ,
         \P0[595] , \P0[594] , \P0[593] , \P0[592] , \P0[591] , \P0[590] ,
         \P0[589] , \P0[588] , \P0[587] , \P0[586] , \P0[585] , \P0[584] ,
         \P0[583] , \P0[582] , \P0[581] , \P0[580] , \P0[579] , \P0[578] ,
         \P0[577] , \P0[576] , \P0[575] , \P0[574] , \P0[573] , \P0[572] ,
         \P0[571] , \P0[570] , \P0[569] , \P0[568] , \P0[567] , \P0[566] ,
         \P0[565] , \P0[564] , \P0[563] , \P0[562] , \P0[561] , \P0[560] ,
         \P0[559] , \P0[558] , \P0[557] , \P0[556] , \P0[555] , \P0[554] ,
         \P0[553] , \P0[552] , \P0[551] , \P0[550] , \P0[549] , \P0[548] ,
         \P0[547] , \P0[546] , \P0[545] , \P0[544] , \P0[543] , \P0[542] ,
         \P0[541] , \P0[540] , \P0[539] , \P0[538] , \P0[537] , \P0[536] ,
         \P0[535] , \P0[534] , \P0[533] , \P0[532] , \P0[531] , \P0[530] ,
         \P0[529] , \P0[528] , \P0[527] , \P0[526] , \P0[525] , \P0[524] ,
         \P0[523] , \P0[522] , \P0[521] , \P0[520] , \P0[519] , \P0[518] ,
         \P0[517] , \P0[516] , \P0[515] , \P0[514] , \P0[513] ;
  wire   SYNOPSYS_UNCONNECTED__0;

  mult_N1024_CC512_DW01_add_0 FS_3 ( .A({1'b0, \P0[1023] , \P0[1022] , 
        \P0[1021] , \P0[1020] , \P0[1019] , \P0[1018] , \P0[1017] , \P0[1016] , 
        \P0[1015] , \P0[1014] , \P0[1013] , \P0[1012] , \P0[1011] , \P0[1010] , 
        \P0[1009] , \P0[1008] , \P0[1007] , \P0[1006] , \P0[1005] , \P0[1004] , 
        \P0[1003] , \P0[1002] , \P0[1001] , \P0[1000] , \P0[999] , \P0[998] , 
        \P0[997] , \P0[996] , \P0[995] , \P0[994] , \P0[993] , \P0[992] , 
        \P0[991] , \P0[990] , \P0[989] , \P0[988] , \P0[987] , \P0[986] , 
        \P0[985] , \P0[984] , \P0[983] , \P0[982] , \P0[981] , \P0[980] , 
        \P0[979] , \P0[978] , \P0[977] , \P0[976] , \P0[975] , \P0[974] , 
        \P0[973] , \P0[972] , \P0[971] , \P0[970] , \P0[969] , \P0[968] , 
        \P0[967] , \P0[966] , \P0[965] , \P0[964] , \P0[963] , \P0[962] , 
        \P0[961] , \P0[960] , \P0[959] , \P0[958] , \P0[957] , \P0[956] , 
        \P0[955] , \P0[954] , \P0[953] , \P0[952] , \P0[951] , \P0[950] , 
        \P0[949] , \P0[948] , \P0[947] , \P0[946] , \P0[945] , \P0[944] , 
        \P0[943] , \P0[942] , \P0[941] , \P0[940] , \P0[939] , \P0[938] , 
        \P0[937] , \P0[936] , \P0[935] , \P0[934] , \P0[933] , \P0[932] , 
        \P0[931] , \P0[930] , \P0[929] , \P0[928] , \P0[927] , \P0[926] , 
        \P0[925] , \P0[924] , \P0[923] , \P0[922] , \P0[921] , \P0[920] , 
        \P0[919] , \P0[918] , \P0[917] , \P0[916] , \P0[915] , \P0[914] , 
        \P0[913] , \P0[912] , \P0[911] , \P0[910] , \P0[909] , \P0[908] , 
        \P0[907] , \P0[906] , \P0[905] , \P0[904] , \P0[903] , \P0[902] , 
        \P0[901] , \P0[900] , \P0[899] , \P0[898] , \P0[897] , \P0[896] , 
        \P0[895] , \P0[894] , \P0[893] , \P0[892] , \P0[891] , \P0[890] , 
        \P0[889] , \P0[888] , \P0[887] , \P0[886] , \P0[885] , \P0[884] , 
        \P0[883] , \P0[882] , \P0[881] , \P0[880] , \P0[879] , \P0[878] , 
        \P0[877] , \P0[876] , \P0[875] , \P0[874] , \P0[873] , \P0[872] , 
        \P0[871] , \P0[870] , \P0[869] , \P0[868] , \P0[867] , \P0[866] , 
        \P0[865] , \P0[864] , \P0[863] , \P0[862] , \P0[861] , \P0[860] , 
        \P0[859] , \P0[858] , \P0[857] , \P0[856] , \P0[855] , \P0[854] , 
        \P0[853] , \P0[852] , \P0[851] , \P0[850] , \P0[849] , \P0[848] , 
        \P0[847] , \P0[846] , \P0[845] , \P0[844] , \P0[843] , \P0[842] , 
        \P0[841] , \P0[840] , \P0[839] , \P0[838] , \P0[837] , \P0[836] , 
        \P0[835] , \P0[834] , \P0[833] , \P0[832] , \P0[831] , \P0[830] , 
        \P0[829] , \P0[828] , \P0[827] , \P0[826] , \P0[825] , \P0[824] , 
        \P0[823] , \P0[822] , \P0[821] , \P0[820] , \P0[819] , \P0[818] , 
        \P0[817] , \P0[816] , \P0[815] , \P0[814] , \P0[813] , \P0[812] , 
        \P0[811] , \P0[810] , \P0[809] , \P0[808] , \P0[807] , \P0[806] , 
        \P0[805] , \P0[804] , \P0[803] , \P0[802] , \P0[801] , \P0[800] , 
        \P0[799] , \P0[798] , \P0[797] , \P0[796] , \P0[795] , \P0[794] , 
        \P0[793] , \P0[792] , \P0[791] , \P0[790] , \P0[789] , \P0[788] , 
        \P0[787] , \P0[786] , \P0[785] , \P0[784] , \P0[783] , \P0[782] , 
        \P0[781] , \P0[780] , \P0[779] , \P0[778] , \P0[777] , \P0[776] , 
        \P0[775] , \P0[774] , \P0[773] , \P0[772] , \P0[771] , \P0[770] , 
        \P0[769] , \P0[768] , \P0[767] , \P0[766] , \P0[765] , \P0[764] , 
        \P0[763] , \P0[762] , \P0[761] , \P0[760] , \P0[759] , \P0[758] , 
        \P0[757] , \P0[756] , \P0[755] , \P0[754] , \P0[753] , \P0[752] , 
        \P0[751] , \P0[750] , \P0[749] , \P0[748] , \P0[747] , \P0[746] , 
        \P0[745] , \P0[744] , \P0[743] , \P0[742] , \P0[741] , \P0[740] , 
        \P0[739] , \P0[738] , \P0[737] , \P0[736] , \P0[735] , \P0[734] , 
        \P0[733] , \P0[732] , \P0[731] , \P0[730] , \P0[729] , \P0[728] , 
        \P0[727] , \P0[726] , \P0[725] , \P0[724] , \P0[723] , \P0[722] , 
        \P0[721] , \P0[720] , \P0[719] , \P0[718] , \P0[717] , \P0[716] , 
        \P0[715] , \P0[714] , \P0[713] , \P0[712] , \P0[711] , \P0[710] , 
        \P0[709] , \P0[708] , \P0[707] , \P0[706] , \P0[705] , \P0[704] , 
        \P0[703] , \P0[702] , \P0[701] , \P0[700] , \P0[699] , \P0[698] , 
        \P0[697] , \P0[696] , \P0[695] , \P0[694] , \P0[693] , \P0[692] , 
        \P0[691] , \P0[690] , \P0[689] , \P0[688] , \P0[687] , \P0[686] , 
        \P0[685] , \P0[684] , \P0[683] , \P0[682] , \P0[681] , \P0[680] , 
        \P0[679] , \P0[678] , \P0[677] , \P0[676] , \P0[675] , \P0[674] , 
        \P0[673] , \P0[672] , \P0[671] , \P0[670] , \P0[669] , \P0[668] , 
        \P0[667] , \P0[666] , \P0[665] , \P0[664] , \P0[663] , \P0[662] , 
        \P0[661] , \P0[660] , \P0[659] , \P0[658] , \P0[657] , \P0[656] , 
        \P0[655] , \P0[654] , \P0[653] , \P0[652] , \P0[651] , \P0[650] , 
        \P0[649] , \P0[648] , \P0[647] , \P0[646] , \P0[645] , \P0[644] , 
        \P0[643] , \P0[642] , \P0[641] , \P0[640] , \P0[639] , \P0[638] , 
        \P0[637] , \P0[636] , \P0[635] , \P0[634] , \P0[633] , \P0[632] , 
        \P0[631] , \P0[630] , \P0[629] , \P0[628] , \P0[627] , \P0[626] , 
        \P0[625] , \P0[624] , \P0[623] , \P0[622] , \P0[621] , \P0[620] , 
        \P0[619] , \P0[618] , \P0[617] , \P0[616] , \P0[615] , \P0[614] , 
        \P0[613] , \P0[612] , \P0[611] , \P0[610] , \P0[609] , \P0[608] , 
        \P0[607] , \P0[606] , \P0[605] , \P0[604] , \P0[603] , \P0[602] , 
        \P0[601] , \P0[600] , \P0[599] , \P0[598] , \P0[597] , \P0[596] , 
        \P0[595] , \P0[594] , \P0[593] , \P0[592] , \P0[591] , \P0[590] , 
        \P0[589] , \P0[588] , \P0[587] , \P0[586] , \P0[585] , \P0[584] , 
        \P0[583] , \P0[582] , \P0[581] , \P0[580] , \P0[579] , \P0[578] , 
        \P0[577] , \P0[576] , \P0[575] , \P0[574] , \P0[573] , \P0[572] , 
        \P0[571] , \P0[570] , \P0[569] , \P0[568] , \P0[567] , \P0[566] , 
        \P0[565] , \P0[564] , \P0[563] , \P0[562] , \P0[561] , \P0[560] , 
        \P0[559] , \P0[558] , \P0[557] , \P0[556] , \P0[555] , \P0[554] , 
        \P0[553] , \P0[552] , \P0[551] , \P0[550] , \P0[549] , \P0[548] , 
        \P0[547] , \P0[546] , \P0[545] , \P0[544] , \P0[543] , \P0[542] , 
        \P0[541] , \P0[540] , \P0[539] , \P0[538] , \P0[537] , \P0[536] , 
        \P0[535] , \P0[534] , \P0[533] , \P0[532] , \P0[531] , \P0[530] , 
        \P0[529] , \P0[528] , \P0[527] , \P0[526] , \P0[525] , \P0[524] , 
        \P0[523] , \P0[522] , \P0[521] , \P0[520] , \P0[519] , \P0[518] , 
        \P0[517] , \P0[516] , \P0[515] , \P0[514] , \P0[513] , \P0[512] , 
        \P0[511] , \P0[510] , \P0[509] , \P0[508] , \P0[507] , \P0[506] , 
        \P0[505] , \P0[504] , \P0[503] , \P0[502] , \P0[501] , \P0[500] , 
        \P0[499] , \P0[498] , \P0[497] , \P0[496] , \P0[495] , \P0[494] , 
        \P0[493] , \P0[492] , \P0[491] , \P0[490] , \P0[489] , \P0[488] , 
        \P0[487] , \P0[486] , \P0[485] , \P0[484] , \P0[483] , \P0[482] , 
        \P0[481] , \P0[480] , \P0[479] , \P0[478] , \P0[477] , \P0[476] , 
        \P0[475] , \P0[474] , \P0[473] , \P0[472] , \P0[471] , \P0[470] , 
        \P0[469] , \P0[468] , \P0[467] , \P0[466] , \P0[465] , \P0[464] , 
        \P0[463] , \P0[462] , \P0[461] , \P0[460] , \P0[459] , \P0[458] , 
        \P0[457] , \P0[456] , \P0[455] , \P0[454] , \P0[453] , \P0[452] , 
        \P0[451] , \P0[450] , \P0[449] , \P0[448] , \P0[447] , \P0[446] , 
        \P0[445] , \P0[444] , \P0[443] , \P0[442] , \P0[441] , \P0[440] , 
        \P0[439] , \P0[438] , \P0[437] , \P0[436] , \P0[435] , \P0[434] , 
        \P0[433] , \P0[432] , \P0[431] , \P0[430] , \P0[429] , \P0[428] , 
        \P0[427] , \P0[426] , \P0[425] , \P0[424] , \P0[423] , \P0[422] , 
        \P0[421] , \P0[420] , \P0[419] , \P0[418] , \P0[417] , \P0[416] , 
        \P0[415] , \P0[414] , \P0[413] , \P0[412] , \P0[411] , \P0[410] , 
        \P0[409] , \P0[408] , \P0[407] , \P0[406] , \P0[405] , \P0[404] , 
        \P0[403] , \P0[402] , \P0[401] , \P0[400] , \P0[399] , \P0[398] , 
        \P0[397] , \P0[396] , \P0[395] , \P0[394] , \P0[393] , \P0[392] , 
        \P0[391] , \P0[390] , \P0[389] , \P0[388] , \P0[387] , \P0[386] , 
        \P0[385] , \P0[384] , \P0[383] , \P0[382] , \P0[381] , \P0[380] , 
        \P0[379] , \P0[378] , \P0[377] , \P0[376] , \P0[375] , \P0[374] , 
        \P0[373] , \P0[372] , \P0[371] , \P0[370] , \P0[369] , \P0[368] , 
        \P0[367] , \P0[366] , \P0[365] , \P0[364] , \P0[363] , \P0[362] , 
        \P0[361] , \P0[360] , \P0[359] , \P0[358] , \P0[357] , \P0[356] , 
        \P0[355] , \P0[354] , \P0[353] , \P0[352] , \P0[351] , \P0[350] , 
        \P0[349] , \P0[348] , \P0[347] , \P0[346] , \P0[345] , \P0[344] , 
        \P0[343] , \P0[342] , \P0[341] , \P0[340] , \P0[339] , \P0[338] , 
        \P0[337] , \P0[336] , \P0[335] , \P0[334] , \P0[333] , \P0[332] , 
        \P0[331] , \P0[330] , \P0[329] , \P0[328] , \P0[327] , \P0[326] , 
        \P0[325] , \P0[324] , \P0[323] , \P0[322] , \P0[321] , \P0[320] , 
        \P0[319] , \P0[318] , \P0[317] , \P0[316] , \P0[315] , \P0[314] , 
        \P0[313] , \P0[312] , \P0[311] , \P0[310] , \P0[309] , \P0[308] , 
        \P0[307] , \P0[306] , \P0[305] , \P0[304] , \P0[303] , \P0[302] , 
        \P0[301] , \P0[300] , \P0[299] , \P0[298] , \P0[297] , \P0[296] , 
        \P0[295] , \P0[294] , \P0[293] , \P0[292] , \P0[291] , \P0[290] , 
        \P0[289] , \P0[288] , \P0[287] , \P0[286] , \P0[285] , \P0[284] , 
        \P0[283] , \P0[282] , \P0[281] , \P0[280] , \P0[279] , \P0[278] , 
        \P0[277] , \P0[276] , \P0[275] , \P0[274] , \P0[273] , \P0[272] , 
        \P0[271] , \P0[270] , \P0[269] , \P0[268] , \P0[267] , \P0[266] , 
        \P0[265] , \P0[264] , \P0[263] , \P0[262] , \P0[261] , \P0[260] , 
        \P0[259] , \P0[258] , \P0[257] , \P0[256] , \P0[255] , \P0[254] , 
        \P0[253] , \P0[252] , \P0[251] , \P0[250] , \P0[249] , \P0[248] , 
        \P0[247] , \P0[246] , \P0[245] , \P0[244] , \P0[243] , \P0[242] , 
        \P0[241] , \P0[240] , \P0[239] , \P0[238] , \P0[237] , \P0[236] , 
        \P0[235] , \P0[234] , \P0[233] , \P0[232] , \P0[231] , \P0[230] , 
        \P0[229] , \P0[228] , \P0[227] , \P0[226] , \P0[225] , \P0[224] , 
        \P0[223] , \P0[222] , \P0[221] , \P0[220] , \P0[219] , \P0[218] , 
        \P0[217] , \P0[216] , \P0[215] , \P0[214] , \P0[213] , \P0[212] , 
        \P0[211] , \P0[210] , \P0[209] , \P0[208] , \P0[207] , \P0[206] , 
        \P0[205] , \P0[204] , \P0[203] , \P0[202] , \P0[201] , \P0[200] , 
        \P0[199] , \P0[198] , \P0[197] , \P0[196] , \P0[195] , \P0[194] , 
        \P0[193] , \P0[192] , \P0[191] , \P0[190] , \P0[189] , \P0[188] , 
        \P0[187] , \P0[186] , \P0[185] , \P0[184] , \P0[183] , \P0[182] , 
        \P0[181] , \P0[180] , \P0[179] , \P0[178] , \P0[177] , \P0[176] , 
        \P0[175] , \P0[174] , \P0[173] , \P0[172] , \P0[171] , \P0[170] , 
        \P0[169] , \P0[168] , \P0[167] , \P0[166] , \P0[165] , \P0[164] , 
        \P0[163] , \P0[162] , \P0[161] , \P0[160] , \P0[159] , \P0[158] , 
        \P0[157] , \P0[156] , \P0[155] , \P0[154] , \P0[153] , \P0[152] , 
        \P0[151] , \P0[150] , \P0[149] , \P0[148] , \P0[147] , \P0[146] , 
        \P0[145] , \P0[144] , \P0[143] , \P0[142] , \P0[141] , \P0[140] , 
        \P0[139] , \P0[138] , \P0[137] , \P0[136] , \P0[135] , \P0[134] , 
        \P0[133] , \P0[132] , \P0[131] , \P0[130] , \P0[129] , \P0[128] , 
        \P0[127] , \P0[126] , \P0[125] , \P0[124] , \P0[123] , \P0[122] , 
        \P0[121] , \P0[120] , \P0[119] , \P0[118] , \P0[117] , \P0[116] , 
        \P0[115] , \P0[114] , \P0[113] , \P0[112] , \P0[111] , \P0[110] , 
        \P0[109] , \P0[108] , \P0[107] , \P0[106] , \P0[105] , \P0[104] , 
        \P0[103] , \P0[102] , \P0[101] , \P0[100] , \P0[99] , \P0[98] , 
        \P0[97] , \P0[96] , \P0[95] , \P0[94] , \P0[93] , \P0[92] , \P0[91] , 
        \P0[90] , \P0[89] , \P0[88] , \P0[87] , \P0[86] , \P0[85] , \P0[84] , 
        \P0[83] , \P0[82] , \P0[81] , \P0[80] , \P0[79] , \P0[78] , \P0[77] , 
        \P0[76] , \P0[75] , \P0[74] , \P0[73] , \P0[72] , \P0[71] , \P0[70] , 
        \P0[69] , \P0[68] , \P0[67] , \P0[66] , \P0[65] , \P0[64] , \P0[63] , 
        \P0[62] , \P0[61] , \P0[60] , \P0[59] , \P0[58] , \P0[57] , \P0[56] , 
        \P0[55] , \P0[54] , \P0[53] , \P0[52] , \P0[51] , \P0[50] , \P0[49] , 
        \P0[48] , \P0[47] , \P0[46] , \P0[45] , \P0[44] , \P0[43] , \P0[42] , 
        \P0[41] , \P0[40] , \P0[39] , \P0[38] , \P0[37] , \P0[36] , \P0[35] , 
        \P0[34] , \P0[33] , \P0[32] , \P0[31] , \P0[30] , \P0[29] , \P0[28] , 
        \P0[27] , \P0[26] , \P0[25] , \P0[24] , \P0[23] , \P0[22] , \P0[21] , 
        \P0[20] , \P0[19] , \P0[18] , \P0[17] , \P0[16] , \P0[15] , \P0[14] , 
        \P0[13] , \P0[12] , \P0[11] , \P0[10] , \P0[9] , \P0[8] , \P0[7] , 
        \P0[6] , \P0[5] , \P0[4] , \P0[3] , \P0[2] , \P0[1] }), .B({\P1[1024] , 
        \P1[1023] , \P1[1022] , \P1[1021] , \P1[1020] , \P1[1019] , \P1[1018] , 
        \P1[1017] , \P1[1016] , \P1[1015] , \P1[1014] , \P1[1013] , \P1[1012] , 
        \P1[1011] , \P1[1010] , \P1[1009] , \P1[1008] , \P1[1007] , \P1[1006] , 
        \P1[1005] , \P1[1004] , \P1[1003] , \P1[1002] , \P1[1001] , \P1[1000] , 
        \P1[999] , \P1[998] , \P1[997] , \P1[996] , \P1[995] , \P1[994] , 
        \P1[993] , \P1[992] , \P1[991] , \P1[990] , \P1[989] , \P1[988] , 
        \P1[987] , \P1[986] , \P1[985] , \P1[984] , \P1[983] , \P1[982] , 
        \P1[981] , \P1[980] , \P1[979] , \P1[978] , \P1[977] , \P1[976] , 
        \P1[975] , \P1[974] , \P1[973] , \P1[972] , \P1[971] , \P1[970] , 
        \P1[969] , \P1[968] , \P1[967] , \P1[966] , \P1[965] , \P1[964] , 
        \P1[963] , \P1[962] , \P1[961] , \P1[960] , \P1[959] , \P1[958] , 
        \P1[957] , \P1[956] , \P1[955] , \P1[954] , \P1[953] , \P1[952] , 
        \P1[951] , \P1[950] , \P1[949] , \P1[948] , \P1[947] , \P1[946] , 
        \P1[945] , \P1[944] , \P1[943] , \P1[942] , \P1[941] , \P1[940] , 
        \P1[939] , \P1[938] , \P1[937] , \P1[936] , \P1[935] , \P1[934] , 
        \P1[933] , \P1[932] , \P1[931] , \P1[930] , \P1[929] , \P1[928] , 
        \P1[927] , \P1[926] , \P1[925] , \P1[924] , \P1[923] , \P1[922] , 
        \P1[921] , \P1[920] , \P1[919] , \P1[918] , \P1[917] , \P1[916] , 
        \P1[915] , \P1[914] , \P1[913] , \P1[912] , \P1[911] , \P1[910] , 
        \P1[909] , \P1[908] , \P1[907] , \P1[906] , \P1[905] , \P1[904] , 
        \P1[903] , \P1[902] , \P1[901] , \P1[900] , \P1[899] , \P1[898] , 
        \P1[897] , \P1[896] , \P1[895] , \P1[894] , \P1[893] , \P1[892] , 
        \P1[891] , \P1[890] , \P1[889] , \P1[888] , \P1[887] , \P1[886] , 
        \P1[885] , \P1[884] , \P1[883] , \P1[882] , \P1[881] , \P1[880] , 
        \P1[879] , \P1[878] , \P1[877] , \P1[876] , \P1[875] , \P1[874] , 
        \P1[873] , \P1[872] , \P1[871] , \P1[870] , \P1[869] , \P1[868] , 
        \P1[867] , \P1[866] , \P1[865] , \P1[864] , \P1[863] , \P1[862] , 
        \P1[861] , \P1[860] , \P1[859] , \P1[858] , \P1[857] , \P1[856] , 
        \P1[855] , \P1[854] , \P1[853] , \P1[852] , \P1[851] , \P1[850] , 
        \P1[849] , \P1[848] , \P1[847] , \P1[846] , \P1[845] , \P1[844] , 
        \P1[843] , \P1[842] , \P1[841] , \P1[840] , \P1[839] , \P1[838] , 
        \P1[837] , \P1[836] , \P1[835] , \P1[834] , \P1[833] , \P1[832] , 
        \P1[831] , \P1[830] , \P1[829] , \P1[828] , \P1[827] , \P1[826] , 
        \P1[825] , \P1[824] , \P1[823] , \P1[822] , \P1[821] , \P1[820] , 
        \P1[819] , \P1[818] , \P1[817] , \P1[816] , \P1[815] , \P1[814] , 
        \P1[813] , \P1[812] , \P1[811] , \P1[810] , \P1[809] , \P1[808] , 
        \P1[807] , \P1[806] , \P1[805] , \P1[804] , \P1[803] , \P1[802] , 
        \P1[801] , \P1[800] , \P1[799] , \P1[798] , \P1[797] , \P1[796] , 
        \P1[795] , \P1[794] , \P1[793] , \P1[792] , \P1[791] , \P1[790] , 
        \P1[789] , \P1[788] , \P1[787] , \P1[786] , \P1[785] , \P1[784] , 
        \P1[783] , \P1[782] , \P1[781] , \P1[780] , \P1[779] , \P1[778] , 
        \P1[777] , \P1[776] , \P1[775] , \P1[774] , \P1[773] , \P1[772] , 
        \P1[771] , \P1[770] , \P1[769] , \P1[768] , \P1[767] , \P1[766] , 
        \P1[765] , \P1[764] , \P1[763] , \P1[762] , \P1[761] , \P1[760] , 
        \P1[759] , \P1[758] , \P1[757] , \P1[756] , \P1[755] , \P1[754] , 
        \P1[753] , \P1[752] , \P1[751] , \P1[750] , \P1[749] , \P1[748] , 
        \P1[747] , \P1[746] , \P1[745] , \P1[744] , \P1[743] , \P1[742] , 
        \P1[741] , \P1[740] , \P1[739] , \P1[738] , \P1[737] , \P1[736] , 
        \P1[735] , \P1[734] , \P1[733] , \P1[732] , \P1[731] , \P1[730] , 
        \P1[729] , \P1[728] , \P1[727] , \P1[726] , \P1[725] , \P1[724] , 
        \P1[723] , \P1[722] , \P1[721] , \P1[720] , \P1[719] , \P1[718] , 
        \P1[717] , \P1[716] , \P1[715] , \P1[714] , \P1[713] , \P1[712] , 
        \P1[711] , \P1[710] , \P1[709] , \P1[708] , \P1[707] , \P1[706] , 
        \P1[705] , \P1[704] , \P1[703] , \P1[702] , \P1[701] , \P1[700] , 
        \P1[699] , \P1[698] , \P1[697] , \P1[696] , \P1[695] , \P1[694] , 
        \P1[693] , \P1[692] , \P1[691] , \P1[690] , \P1[689] , \P1[688] , 
        \P1[687] , \P1[686] , \P1[685] , \P1[684] , \P1[683] , \P1[682] , 
        \P1[681] , \P1[680] , \P1[679] , \P1[678] , \P1[677] , \P1[676] , 
        \P1[675] , \P1[674] , \P1[673] , \P1[672] , \P1[671] , \P1[670] , 
        \P1[669] , \P1[668] , \P1[667] , \P1[666] , \P1[665] , \P1[664] , 
        \P1[663] , \P1[662] , \P1[661] , \P1[660] , \P1[659] , \P1[658] , 
        \P1[657] , \P1[656] , \P1[655] , \P1[654] , \P1[653] , \P1[652] , 
        \P1[651] , \P1[650] , \P1[649] , \P1[648] , \P1[647] , \P1[646] , 
        \P1[645] , \P1[644] , \P1[643] , \P1[642] , \P1[641] , \P1[640] , 
        \P1[639] , \P1[638] , \P1[637] , \P1[636] , \P1[635] , \P1[634] , 
        \P1[633] , \P1[632] , \P1[631] , \P1[630] , \P1[629] , \P1[628] , 
        \P1[627] , \P1[626] , \P1[625] , \P1[624] , \P1[623] , \P1[622] , 
        \P1[621] , \P1[620] , \P1[619] , \P1[618] , \P1[617] , \P1[616] , 
        \P1[615] , \P1[614] , \P1[613] , \P1[612] , \P1[611] , \P1[610] , 
        \P1[609] , \P1[608] , \P1[607] , \P1[606] , \P1[605] , \P1[604] , 
        \P1[603] , \P1[602] , \P1[601] , \P1[600] , \P1[599] , \P1[598] , 
        \P1[597] , \P1[596] , \P1[595] , \P1[594] , \P1[593] , \P1[592] , 
        \P1[591] , \P1[590] , \P1[589] , \P1[588] , \P1[587] , \P1[586] , 
        \P1[585] , \P1[584] , \P1[583] , \P1[582] , \P1[581] , \P1[580] , 
        \P1[579] , \P1[578] , \P1[577] , \P1[576] , \P1[575] , \P1[574] , 
        \P1[573] , \P1[572] , \P1[571] , \P1[570] , \P1[569] , \P1[568] , 
        \P1[567] , \P1[566] , \P1[565] , \P1[564] , \P1[563] , \P1[562] , 
        \P1[561] , \P1[560] , \P1[559] , \P1[558] , \P1[557] , \P1[556] , 
        \P1[555] , \P1[554] , \P1[553] , \P1[552] , \P1[551] , \P1[550] , 
        \P1[549] , \P1[548] , \P1[547] , \P1[546] , \P1[545] , \P1[544] , 
        \P1[543] , \P1[542] , \P1[541] , \P1[540] , \P1[539] , \P1[538] , 
        \P1[537] , \P1[536] , \P1[535] , \P1[534] , \P1[533] , \P1[532] , 
        \P1[531] , \P1[530] , \P1[529] , \P1[528] , \P1[527] , \P1[526] , 
        \P1[525] , \P1[524] , \P1[523] , \P1[522] , \P1[521] , \P1[520] , 
        \P1[519] , \P1[518] , \P1[517] , \P1[516] , \P1[515] , \P1[514] , 
        \P1[513] , \P1[512] , \P1[511] , \P1[510] , \P1[509] , \P1[508] , 
        \P1[507] , \P1[506] , \P1[505] , \P1[504] , \P1[503] , \P1[502] , 
        \P1[501] , \P1[500] , \P1[499] , \P1[498] , \P1[497] , \P1[496] , 
        \P1[495] , \P1[494] , \P1[493] , \P1[492] , \P1[491] , \P1[490] , 
        \P1[489] , \P1[488] , \P1[487] , \P1[486] , \P1[485] , \P1[484] , 
        \P1[483] , \P1[482] , \P1[481] , \P1[480] , \P1[479] , \P1[478] , 
        \P1[477] , \P1[476] , \P1[475] , \P1[474] , \P1[473] , \P1[472] , 
        \P1[471] , \P1[470] , \P1[469] , \P1[468] , \P1[467] , \P1[466] , 
        \P1[465] , \P1[464] , \P1[463] , \P1[462] , \P1[461] , \P1[460] , 
        \P1[459] , \P1[458] , \P1[457] , \P1[456] , \P1[455] , \P1[454] , 
        \P1[453] , \P1[452] , \P1[451] , \P1[450] , \P1[449] , \P1[448] , 
        \P1[447] , \P1[446] , \P1[445] , \P1[444] , \P1[443] , \P1[442] , 
        \P1[441] , \P1[440] , \P1[439] , \P1[438] , \P1[437] , \P1[436] , 
        \P1[435] , \P1[434] , \P1[433] , \P1[432] , \P1[431] , \P1[430] , 
        \P1[429] , \P1[428] , \P1[427] , \P1[426] , \P1[425] , \P1[424] , 
        \P1[423] , \P1[422] , \P1[421] , \P1[420] , \P1[419] , \P1[418] , 
        \P1[417] , \P1[416] , \P1[415] , \P1[414] , \P1[413] , \P1[412] , 
        \P1[411] , \P1[410] , \P1[409] , \P1[408] , \P1[407] , \P1[406] , 
        \P1[405] , \P1[404] , \P1[403] , \P1[402] , \P1[401] , \P1[400] , 
        \P1[399] , \P1[398] , \P1[397] , \P1[396] , \P1[395] , \P1[394] , 
        \P1[393] , \P1[392] , \P1[391] , \P1[390] , \P1[389] , \P1[388] , 
        \P1[387] , \P1[386] , \P1[385] , \P1[384] , \P1[383] , \P1[382] , 
        \P1[381] , \P1[380] , \P1[379] , \P1[378] , \P1[377] , \P1[376] , 
        \P1[375] , \P1[374] , \P1[373] , \P1[372] , \P1[371] , \P1[370] , 
        \P1[369] , \P1[368] , \P1[367] , \P1[366] , \P1[365] , \P1[364] , 
        \P1[363] , \P1[362] , \P1[361] , \P1[360] , \P1[359] , \P1[358] , 
        \P1[357] , \P1[356] , \P1[355] , \P1[354] , \P1[353] , \P1[352] , 
        \P1[351] , \P1[350] , \P1[349] , \P1[348] , \P1[347] , \P1[346] , 
        \P1[345] , \P1[344] , \P1[343] , \P1[342] , \P1[341] , \P1[340] , 
        \P1[339] , \P1[338] , \P1[337] , \P1[336] , \P1[335] , \P1[334] , 
        \P1[333] , \P1[332] , \P1[331] , \P1[330] , \P1[329] , \P1[328] , 
        \P1[327] , \P1[326] , \P1[325] , \P1[324] , \P1[323] , \P1[322] , 
        \P1[321] , \P1[320] , \P1[319] , \P1[318] , \P1[317] , \P1[316] , 
        \P1[315] , \P1[314] , \P1[313] , \P1[312] , \P1[311] , \P1[310] , 
        \P1[309] , \P1[308] , \P1[307] , \P1[306] , \P1[305] , \P1[304] , 
        \P1[303] , \P1[302] , \P1[301] , \P1[300] , \P1[299] , \P1[298] , 
        \P1[297] , \P1[296] , \P1[295] , \P1[294] , \P1[293] , \P1[292] , 
        \P1[291] , \P1[290] , \P1[289] , \P1[288] , \P1[287] , \P1[286] , 
        \P1[285] , \P1[284] , \P1[283] , \P1[282] , \P1[281] , \P1[280] , 
        \P1[279] , \P1[278] , \P1[277] , \P1[276] , \P1[275] , \P1[274] , 
        \P1[273] , \P1[272] , \P1[271] , \P1[270] , \P1[269] , \P1[268] , 
        \P1[267] , \P1[266] , \P1[265] , \P1[264] , \P1[263] , \P1[262] , 
        \P1[261] , \P1[260] , \P1[259] , \P1[258] , \P1[257] , \P1[256] , 
        \P1[255] , \P1[254] , \P1[253] , \P1[252] , \P1[251] , \P1[250] , 
        \P1[249] , \P1[248] , \P1[247] , \P1[246] , \P1[245] , \P1[244] , 
        \P1[243] , \P1[242] , \P1[241] , \P1[240] , \P1[239] , \P1[238] , 
        \P1[237] , \P1[236] , \P1[235] , \P1[234] , \P1[233] , \P1[232] , 
        \P1[231] , \P1[230] , \P1[229] , \P1[228] , \P1[227] , \P1[226] , 
        \P1[225] , \P1[224] , \P1[223] , \P1[222] , \P1[221] , \P1[220] , 
        \P1[219] , \P1[218] , \P1[217] , \P1[216] , \P1[215] , \P1[214] , 
        \P1[213] , \P1[212] , \P1[211] , \P1[210] , \P1[209] , \P1[208] , 
        \P1[207] , \P1[206] , \P1[205] , \P1[204] , \P1[203] , \P1[202] , 
        \P1[201] , \P1[200] , \P1[199] , \P1[198] , \P1[197] , \P1[196] , 
        \P1[195] , \P1[194] , \P1[193] , \P1[192] , \P1[191] , \P1[190] , 
        \P1[189] , \P1[188] , \P1[187] , \P1[186] , \P1[185] , \P1[184] , 
        \P1[183] , \P1[182] , \P1[181] , \P1[180] , \P1[179] , \P1[178] , 
        \P1[177] , \P1[176] , \P1[175] , \P1[174] , \P1[173] , \P1[172] , 
        \P1[171] , \P1[170] , \P1[169] , \P1[168] , \P1[167] , \P1[166] , 
        \P1[165] , \P1[164] , \P1[163] , \P1[162] , \P1[161] , \P1[160] , 
        \P1[159] , \P1[158] , \P1[157] , \P1[156] , \P1[155] , \P1[154] , 
        \P1[153] , \P1[152] , \P1[151] , \P1[150] , \P1[149] , \P1[148] , 
        \P1[147] , \P1[146] , \P1[145] , \P1[144] , \P1[143] , \P1[142] , 
        \P1[141] , \P1[140] , \P1[139] , \P1[138] , \P1[137] , \P1[136] , 
        \P1[135] , \P1[134] , \P1[133] , \P1[132] , \P1[131] , \P1[130] , 
        \P1[129] , \P1[128] , \P1[127] , \P1[126] , \P1[125] , \P1[124] , 
        \P1[123] , \P1[122] , \P1[121] , \P1[120] , \P1[119] , \P1[118] , 
        \P1[117] , \P1[116] , \P1[115] , \P1[114] , \P1[113] , \P1[112] , 
        \P1[111] , \P1[110] , \P1[109] , \P1[108] , \P1[107] , \P1[106] , 
        \P1[105] , \P1[104] , \P1[103] , \P1[102] , \P1[101] , \P1[100] , 
        \P1[99] , \P1[98] , \P1[97] , \P1[96] , \P1[95] , \P1[94] , \P1[93] , 
        \P1[92] , \P1[91] , \P1[90] , \P1[89] , \P1[88] , \P1[87] , \P1[86] , 
        \P1[85] , \P1[84] , \P1[83] , \P1[82] , \P1[81] , \P1[80] , \P1[79] , 
        \P1[78] , \P1[77] , \P1[76] , \P1[75] , \P1[74] , \P1[73] , \P1[72] , 
        \P1[71] , \P1[70] , \P1[69] , \P1[68] , \P1[67] , \P1[66] , \P1[65] , 
        \P1[64] , \P1[63] , \P1[62] , \P1[61] , \P1[60] , \P1[59] , \P1[58] , 
        \P1[57] , \P1[56] , \P1[55] , \P1[54] , \P1[53] , \P1[52] , \P1[51] , 
        \P1[50] , \P1[49] , \P1[48] , \P1[47] , \P1[46] , \P1[45] , \P1[44] , 
        \P1[43] , \P1[42] , \P1[41] , \P1[40] , \P1[39] , \P1[38] , \P1[37] , 
        \P1[36] , \P1[35] , \P1[34] , \P1[33] , \P1[32] , \P1[31] , \P1[30] , 
        \P1[29] , \P1[28] , \P1[27] , \P1[26] , \P1[25] , \P1[24] , \P1[23] , 
        \P1[22] , \P1[21] , \P1[20] , \P1[19] , \P1[18] , \P1[17] , \P1[16] , 
        \P1[15] , \P1[14] , \P1[13] , \P1[12] , \P1[11] , \P1[10] , \P1[9] , 
        \P1[8] , \P1[7] , \P1[6] , \P1[5] , \P1[4] , \P1[3] , \P1[2] , \P1[1] }), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__0, PRODUCT[1023:1]}) );
  AND U2 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
  AND U3 ( .A(A[8]), .B(B[1]), .Z(\P1[9] ) );
  AND U4 ( .A(B[1]), .B(A[98]), .Z(\P1[99] ) );
  AND U5 ( .A(B[1]), .B(A[998]), .Z(\P1[999] ) );
  AND U6 ( .A(B[1]), .B(A[997]), .Z(\P1[998] ) );
  AND U7 ( .A(B[1]), .B(A[996]), .Z(\P1[997] ) );
  AND U8 ( .A(B[1]), .B(A[995]), .Z(\P1[996] ) );
  AND U9 ( .A(B[1]), .B(A[994]), .Z(\P1[995] ) );
  AND U10 ( .A(B[1]), .B(A[993]), .Z(\P1[994] ) );
  AND U11 ( .A(B[1]), .B(A[992]), .Z(\P1[993] ) );
  AND U12 ( .A(B[1]), .B(A[991]), .Z(\P1[992] ) );
  AND U13 ( .A(B[1]), .B(A[990]), .Z(\P1[991] ) );
  AND U14 ( .A(B[1]), .B(A[989]), .Z(\P1[990] ) );
  AND U15 ( .A(B[1]), .B(A[97]), .Z(\P1[98] ) );
  AND U16 ( .A(B[1]), .B(A[988]), .Z(\P1[989] ) );
  AND U17 ( .A(B[1]), .B(A[987]), .Z(\P1[988] ) );
  AND U18 ( .A(B[1]), .B(A[986]), .Z(\P1[987] ) );
  AND U19 ( .A(B[1]), .B(A[985]), .Z(\P1[986] ) );
  AND U20 ( .A(B[1]), .B(A[984]), .Z(\P1[985] ) );
  AND U21 ( .A(B[1]), .B(A[983]), .Z(\P1[984] ) );
  AND U22 ( .A(B[1]), .B(A[982]), .Z(\P1[983] ) );
  AND U23 ( .A(B[1]), .B(A[981]), .Z(\P1[982] ) );
  AND U24 ( .A(B[1]), .B(A[980]), .Z(\P1[981] ) );
  AND U25 ( .A(B[1]), .B(A[979]), .Z(\P1[980] ) );
  AND U26 ( .A(B[1]), .B(A[96]), .Z(\P1[97] ) );
  AND U27 ( .A(B[1]), .B(A[978]), .Z(\P1[979] ) );
  AND U28 ( .A(B[1]), .B(A[977]), .Z(\P1[978] ) );
  AND U29 ( .A(B[1]), .B(A[976]), .Z(\P1[977] ) );
  AND U30 ( .A(B[1]), .B(A[975]), .Z(\P1[976] ) );
  AND U31 ( .A(B[1]), .B(A[974]), .Z(\P1[975] ) );
  AND U32 ( .A(B[1]), .B(A[973]), .Z(\P1[974] ) );
  AND U33 ( .A(B[1]), .B(A[972]), .Z(\P1[973] ) );
  AND U34 ( .A(B[1]), .B(A[971]), .Z(\P1[972] ) );
  AND U35 ( .A(B[1]), .B(A[970]), .Z(\P1[971] ) );
  AND U36 ( .A(B[1]), .B(A[969]), .Z(\P1[970] ) );
  AND U37 ( .A(B[1]), .B(A[95]), .Z(\P1[96] ) );
  AND U38 ( .A(B[1]), .B(A[968]), .Z(\P1[969] ) );
  AND U39 ( .A(B[1]), .B(A[967]), .Z(\P1[968] ) );
  AND U40 ( .A(B[1]), .B(A[966]), .Z(\P1[967] ) );
  AND U41 ( .A(B[1]), .B(A[965]), .Z(\P1[966] ) );
  AND U42 ( .A(B[1]), .B(A[964]), .Z(\P1[965] ) );
  AND U43 ( .A(B[1]), .B(A[963]), .Z(\P1[964] ) );
  AND U44 ( .A(B[1]), .B(A[962]), .Z(\P1[963] ) );
  AND U45 ( .A(B[1]), .B(A[961]), .Z(\P1[962] ) );
  AND U46 ( .A(B[1]), .B(A[960]), .Z(\P1[961] ) );
  AND U47 ( .A(B[1]), .B(A[959]), .Z(\P1[960] ) );
  AND U48 ( .A(B[1]), .B(A[94]), .Z(\P1[95] ) );
  AND U49 ( .A(B[1]), .B(A[958]), .Z(\P1[959] ) );
  AND U50 ( .A(B[1]), .B(A[957]), .Z(\P1[958] ) );
  AND U51 ( .A(B[1]), .B(A[956]), .Z(\P1[957] ) );
  AND U52 ( .A(B[1]), .B(A[955]), .Z(\P1[956] ) );
  AND U53 ( .A(B[1]), .B(A[954]), .Z(\P1[955] ) );
  AND U54 ( .A(B[1]), .B(A[953]), .Z(\P1[954] ) );
  AND U55 ( .A(B[1]), .B(A[952]), .Z(\P1[953] ) );
  AND U56 ( .A(B[1]), .B(A[951]), .Z(\P1[952] ) );
  AND U57 ( .A(B[1]), .B(A[950]), .Z(\P1[951] ) );
  AND U58 ( .A(B[1]), .B(A[949]), .Z(\P1[950] ) );
  AND U59 ( .A(B[1]), .B(A[93]), .Z(\P1[94] ) );
  AND U60 ( .A(B[1]), .B(A[948]), .Z(\P1[949] ) );
  AND U61 ( .A(B[1]), .B(A[947]), .Z(\P1[948] ) );
  AND U62 ( .A(B[1]), .B(A[946]), .Z(\P1[947] ) );
  AND U63 ( .A(B[1]), .B(A[945]), .Z(\P1[946] ) );
  AND U64 ( .A(B[1]), .B(A[944]), .Z(\P1[945] ) );
  AND U65 ( .A(B[1]), .B(A[943]), .Z(\P1[944] ) );
  AND U66 ( .A(B[1]), .B(A[942]), .Z(\P1[943] ) );
  AND U67 ( .A(B[1]), .B(A[941]), .Z(\P1[942] ) );
  AND U68 ( .A(B[1]), .B(A[940]), .Z(\P1[941] ) );
  AND U69 ( .A(B[1]), .B(A[939]), .Z(\P1[940] ) );
  AND U70 ( .A(B[1]), .B(A[92]), .Z(\P1[93] ) );
  AND U71 ( .A(B[1]), .B(A[938]), .Z(\P1[939] ) );
  AND U72 ( .A(B[1]), .B(A[937]), .Z(\P1[938] ) );
  AND U73 ( .A(B[1]), .B(A[936]), .Z(\P1[937] ) );
  AND U74 ( .A(B[1]), .B(A[935]), .Z(\P1[936] ) );
  AND U75 ( .A(B[1]), .B(A[934]), .Z(\P1[935] ) );
  AND U76 ( .A(B[1]), .B(A[933]), .Z(\P1[934] ) );
  AND U77 ( .A(B[1]), .B(A[932]), .Z(\P1[933] ) );
  AND U78 ( .A(B[1]), .B(A[931]), .Z(\P1[932] ) );
  AND U79 ( .A(B[1]), .B(A[930]), .Z(\P1[931] ) );
  AND U80 ( .A(B[1]), .B(A[929]), .Z(\P1[930] ) );
  AND U81 ( .A(B[1]), .B(A[91]), .Z(\P1[92] ) );
  AND U82 ( .A(B[1]), .B(A[928]), .Z(\P1[929] ) );
  AND U83 ( .A(B[1]), .B(A[927]), .Z(\P1[928] ) );
  AND U84 ( .A(B[1]), .B(A[926]), .Z(\P1[927] ) );
  AND U85 ( .A(B[1]), .B(A[925]), .Z(\P1[926] ) );
  AND U86 ( .A(B[1]), .B(A[924]), .Z(\P1[925] ) );
  AND U87 ( .A(B[1]), .B(A[923]), .Z(\P1[924] ) );
  AND U88 ( .A(B[1]), .B(A[922]), .Z(\P1[923] ) );
  AND U89 ( .A(B[1]), .B(A[921]), .Z(\P1[922] ) );
  AND U90 ( .A(B[1]), .B(A[920]), .Z(\P1[921] ) );
  AND U91 ( .A(B[1]), .B(A[919]), .Z(\P1[920] ) );
  AND U92 ( .A(B[1]), .B(A[90]), .Z(\P1[91] ) );
  AND U93 ( .A(B[1]), .B(A[918]), .Z(\P1[919] ) );
  AND U94 ( .A(B[1]), .B(A[917]), .Z(\P1[918] ) );
  AND U95 ( .A(B[1]), .B(A[916]), .Z(\P1[917] ) );
  AND U96 ( .A(B[1]), .B(A[915]), .Z(\P1[916] ) );
  AND U97 ( .A(B[1]), .B(A[914]), .Z(\P1[915] ) );
  AND U98 ( .A(B[1]), .B(A[913]), .Z(\P1[914] ) );
  AND U99 ( .A(B[1]), .B(A[912]), .Z(\P1[913] ) );
  AND U100 ( .A(B[1]), .B(A[911]), .Z(\P1[912] ) );
  AND U101 ( .A(B[1]), .B(A[910]), .Z(\P1[911] ) );
  AND U102 ( .A(B[1]), .B(A[909]), .Z(\P1[910] ) );
  AND U103 ( .A(B[1]), .B(A[89]), .Z(\P1[90] ) );
  AND U104 ( .A(B[1]), .B(A[908]), .Z(\P1[909] ) );
  AND U105 ( .A(B[1]), .B(A[907]), .Z(\P1[908] ) );
  AND U106 ( .A(B[1]), .B(A[906]), .Z(\P1[907] ) );
  AND U107 ( .A(B[1]), .B(A[905]), .Z(\P1[906] ) );
  AND U108 ( .A(B[1]), .B(A[904]), .Z(\P1[905] ) );
  AND U109 ( .A(B[1]), .B(A[903]), .Z(\P1[904] ) );
  AND U110 ( .A(B[1]), .B(A[902]), .Z(\P1[903] ) );
  AND U111 ( .A(B[1]), .B(A[901]), .Z(\P1[902] ) );
  AND U112 ( .A(B[1]), .B(A[900]), .Z(\P1[901] ) );
  AND U113 ( .A(B[1]), .B(A[899]), .Z(\P1[900] ) );
  AND U114 ( .A(B[1]), .B(A[7]), .Z(\P1[8] ) );
  AND U115 ( .A(B[1]), .B(A[88]), .Z(\P1[89] ) );
  AND U116 ( .A(B[1]), .B(A[898]), .Z(\P1[899] ) );
  AND U117 ( .A(B[1]), .B(A[897]), .Z(\P1[898] ) );
  AND U118 ( .A(B[1]), .B(A[896]), .Z(\P1[897] ) );
  AND U119 ( .A(B[1]), .B(A[895]), .Z(\P1[896] ) );
  AND U120 ( .A(B[1]), .B(A[894]), .Z(\P1[895] ) );
  AND U121 ( .A(B[1]), .B(A[893]), .Z(\P1[894] ) );
  AND U122 ( .A(B[1]), .B(A[892]), .Z(\P1[893] ) );
  AND U123 ( .A(B[1]), .B(A[891]), .Z(\P1[892] ) );
  AND U124 ( .A(B[1]), .B(A[890]), .Z(\P1[891] ) );
  AND U125 ( .A(B[1]), .B(A[889]), .Z(\P1[890] ) );
  AND U126 ( .A(B[1]), .B(A[87]), .Z(\P1[88] ) );
  AND U127 ( .A(B[1]), .B(A[888]), .Z(\P1[889] ) );
  AND U128 ( .A(B[1]), .B(A[887]), .Z(\P1[888] ) );
  AND U129 ( .A(B[1]), .B(A[886]), .Z(\P1[887] ) );
  AND U130 ( .A(B[1]), .B(A[885]), .Z(\P1[886] ) );
  AND U131 ( .A(B[1]), .B(A[884]), .Z(\P1[885] ) );
  AND U132 ( .A(B[1]), .B(A[883]), .Z(\P1[884] ) );
  AND U133 ( .A(B[1]), .B(A[882]), .Z(\P1[883] ) );
  AND U134 ( .A(B[1]), .B(A[881]), .Z(\P1[882] ) );
  AND U135 ( .A(B[1]), .B(A[880]), .Z(\P1[881] ) );
  AND U136 ( .A(B[1]), .B(A[879]), .Z(\P1[880] ) );
  AND U137 ( .A(B[1]), .B(A[86]), .Z(\P1[87] ) );
  AND U138 ( .A(B[1]), .B(A[878]), .Z(\P1[879] ) );
  AND U139 ( .A(B[1]), .B(A[877]), .Z(\P1[878] ) );
  AND U140 ( .A(B[1]), .B(A[876]), .Z(\P1[877] ) );
  AND U141 ( .A(B[1]), .B(A[875]), .Z(\P1[876] ) );
  AND U142 ( .A(B[1]), .B(A[874]), .Z(\P1[875] ) );
  AND U143 ( .A(B[1]), .B(A[873]), .Z(\P1[874] ) );
  AND U144 ( .A(B[1]), .B(A[872]), .Z(\P1[873] ) );
  AND U145 ( .A(B[1]), .B(A[871]), .Z(\P1[872] ) );
  AND U146 ( .A(B[1]), .B(A[870]), .Z(\P1[871] ) );
  AND U147 ( .A(B[1]), .B(A[869]), .Z(\P1[870] ) );
  AND U148 ( .A(B[1]), .B(A[85]), .Z(\P1[86] ) );
  AND U149 ( .A(B[1]), .B(A[868]), .Z(\P1[869] ) );
  AND U150 ( .A(B[1]), .B(A[867]), .Z(\P1[868] ) );
  AND U151 ( .A(B[1]), .B(A[866]), .Z(\P1[867] ) );
  AND U152 ( .A(B[1]), .B(A[865]), .Z(\P1[866] ) );
  AND U153 ( .A(B[1]), .B(A[864]), .Z(\P1[865] ) );
  AND U154 ( .A(B[1]), .B(A[863]), .Z(\P1[864] ) );
  AND U155 ( .A(B[1]), .B(A[862]), .Z(\P1[863] ) );
  AND U156 ( .A(B[1]), .B(A[861]), .Z(\P1[862] ) );
  AND U157 ( .A(B[1]), .B(A[860]), .Z(\P1[861] ) );
  AND U158 ( .A(B[1]), .B(A[859]), .Z(\P1[860] ) );
  AND U159 ( .A(B[1]), .B(A[84]), .Z(\P1[85] ) );
  AND U160 ( .A(B[1]), .B(A[858]), .Z(\P1[859] ) );
  AND U161 ( .A(B[1]), .B(A[857]), .Z(\P1[858] ) );
  AND U162 ( .A(B[1]), .B(A[856]), .Z(\P1[857] ) );
  AND U163 ( .A(B[1]), .B(A[855]), .Z(\P1[856] ) );
  AND U164 ( .A(B[1]), .B(A[854]), .Z(\P1[855] ) );
  AND U165 ( .A(B[1]), .B(A[853]), .Z(\P1[854] ) );
  AND U166 ( .A(B[1]), .B(A[852]), .Z(\P1[853] ) );
  AND U167 ( .A(B[1]), .B(A[851]), .Z(\P1[852] ) );
  AND U168 ( .A(B[1]), .B(A[850]), .Z(\P1[851] ) );
  AND U169 ( .A(B[1]), .B(A[849]), .Z(\P1[850] ) );
  AND U170 ( .A(B[1]), .B(A[83]), .Z(\P1[84] ) );
  AND U171 ( .A(B[1]), .B(A[848]), .Z(\P1[849] ) );
  AND U172 ( .A(B[1]), .B(A[847]), .Z(\P1[848] ) );
  AND U173 ( .A(B[1]), .B(A[846]), .Z(\P1[847] ) );
  AND U174 ( .A(B[1]), .B(A[845]), .Z(\P1[846] ) );
  AND U175 ( .A(B[1]), .B(A[844]), .Z(\P1[845] ) );
  AND U176 ( .A(B[1]), .B(A[843]), .Z(\P1[844] ) );
  AND U177 ( .A(B[1]), .B(A[842]), .Z(\P1[843] ) );
  AND U178 ( .A(B[1]), .B(A[841]), .Z(\P1[842] ) );
  AND U179 ( .A(B[1]), .B(A[840]), .Z(\P1[841] ) );
  AND U180 ( .A(B[1]), .B(A[839]), .Z(\P1[840] ) );
  AND U181 ( .A(B[1]), .B(A[82]), .Z(\P1[83] ) );
  AND U182 ( .A(B[1]), .B(A[838]), .Z(\P1[839] ) );
  AND U183 ( .A(B[1]), .B(A[837]), .Z(\P1[838] ) );
  AND U184 ( .A(B[1]), .B(A[836]), .Z(\P1[837] ) );
  AND U185 ( .A(B[1]), .B(A[835]), .Z(\P1[836] ) );
  AND U186 ( .A(B[1]), .B(A[834]), .Z(\P1[835] ) );
  AND U187 ( .A(B[1]), .B(A[833]), .Z(\P1[834] ) );
  AND U188 ( .A(B[1]), .B(A[832]), .Z(\P1[833] ) );
  AND U189 ( .A(B[1]), .B(A[831]), .Z(\P1[832] ) );
  AND U190 ( .A(B[1]), .B(A[830]), .Z(\P1[831] ) );
  AND U191 ( .A(B[1]), .B(A[829]), .Z(\P1[830] ) );
  AND U192 ( .A(B[1]), .B(A[81]), .Z(\P1[82] ) );
  AND U193 ( .A(B[1]), .B(A[828]), .Z(\P1[829] ) );
  AND U194 ( .A(B[1]), .B(A[827]), .Z(\P1[828] ) );
  AND U195 ( .A(B[1]), .B(A[826]), .Z(\P1[827] ) );
  AND U196 ( .A(B[1]), .B(A[825]), .Z(\P1[826] ) );
  AND U197 ( .A(B[1]), .B(A[824]), .Z(\P1[825] ) );
  AND U198 ( .A(B[1]), .B(A[823]), .Z(\P1[824] ) );
  AND U199 ( .A(B[1]), .B(A[822]), .Z(\P1[823] ) );
  AND U200 ( .A(B[1]), .B(A[821]), .Z(\P1[822] ) );
  AND U201 ( .A(B[1]), .B(A[820]), .Z(\P1[821] ) );
  AND U202 ( .A(B[1]), .B(A[819]), .Z(\P1[820] ) );
  AND U203 ( .A(B[1]), .B(A[80]), .Z(\P1[81] ) );
  AND U204 ( .A(B[1]), .B(A[818]), .Z(\P1[819] ) );
  AND U205 ( .A(B[1]), .B(A[817]), .Z(\P1[818] ) );
  AND U206 ( .A(B[1]), .B(A[816]), .Z(\P1[817] ) );
  AND U207 ( .A(B[1]), .B(A[815]), .Z(\P1[816] ) );
  AND U208 ( .A(B[1]), .B(A[814]), .Z(\P1[815] ) );
  AND U209 ( .A(B[1]), .B(A[813]), .Z(\P1[814] ) );
  AND U210 ( .A(B[1]), .B(A[812]), .Z(\P1[813] ) );
  AND U211 ( .A(B[1]), .B(A[811]), .Z(\P1[812] ) );
  AND U212 ( .A(B[1]), .B(A[810]), .Z(\P1[811] ) );
  AND U213 ( .A(B[1]), .B(A[809]), .Z(\P1[810] ) );
  AND U214 ( .A(B[1]), .B(A[79]), .Z(\P1[80] ) );
  AND U215 ( .A(B[1]), .B(A[808]), .Z(\P1[809] ) );
  AND U216 ( .A(B[1]), .B(A[807]), .Z(\P1[808] ) );
  AND U217 ( .A(B[1]), .B(A[806]), .Z(\P1[807] ) );
  AND U218 ( .A(B[1]), .B(A[805]), .Z(\P1[806] ) );
  AND U219 ( .A(B[1]), .B(A[804]), .Z(\P1[805] ) );
  AND U220 ( .A(B[1]), .B(A[803]), .Z(\P1[804] ) );
  AND U221 ( .A(B[1]), .B(A[802]), .Z(\P1[803] ) );
  AND U222 ( .A(B[1]), .B(A[801]), .Z(\P1[802] ) );
  AND U223 ( .A(B[1]), .B(A[800]), .Z(\P1[801] ) );
  AND U224 ( .A(B[1]), .B(A[799]), .Z(\P1[800] ) );
  AND U225 ( .A(B[1]), .B(A[6]), .Z(\P1[7] ) );
  AND U226 ( .A(B[1]), .B(A[78]), .Z(\P1[79] ) );
  AND U227 ( .A(B[1]), .B(A[798]), .Z(\P1[799] ) );
  AND U228 ( .A(B[1]), .B(A[797]), .Z(\P1[798] ) );
  AND U229 ( .A(B[1]), .B(A[796]), .Z(\P1[797] ) );
  AND U230 ( .A(B[1]), .B(A[795]), .Z(\P1[796] ) );
  AND U231 ( .A(B[1]), .B(A[794]), .Z(\P1[795] ) );
  AND U232 ( .A(B[1]), .B(A[793]), .Z(\P1[794] ) );
  AND U233 ( .A(B[1]), .B(A[792]), .Z(\P1[793] ) );
  AND U234 ( .A(B[1]), .B(A[791]), .Z(\P1[792] ) );
  AND U235 ( .A(B[1]), .B(A[790]), .Z(\P1[791] ) );
  AND U236 ( .A(B[1]), .B(A[789]), .Z(\P1[790] ) );
  AND U237 ( .A(B[1]), .B(A[77]), .Z(\P1[78] ) );
  AND U238 ( .A(B[1]), .B(A[788]), .Z(\P1[789] ) );
  AND U239 ( .A(B[1]), .B(A[787]), .Z(\P1[788] ) );
  AND U240 ( .A(B[1]), .B(A[786]), .Z(\P1[787] ) );
  AND U241 ( .A(B[1]), .B(A[785]), .Z(\P1[786] ) );
  AND U242 ( .A(B[1]), .B(A[784]), .Z(\P1[785] ) );
  AND U243 ( .A(B[1]), .B(A[783]), .Z(\P1[784] ) );
  AND U244 ( .A(B[1]), .B(A[782]), .Z(\P1[783] ) );
  AND U245 ( .A(B[1]), .B(A[781]), .Z(\P1[782] ) );
  AND U246 ( .A(B[1]), .B(A[780]), .Z(\P1[781] ) );
  AND U247 ( .A(B[1]), .B(A[779]), .Z(\P1[780] ) );
  AND U248 ( .A(B[1]), .B(A[76]), .Z(\P1[77] ) );
  AND U249 ( .A(B[1]), .B(A[778]), .Z(\P1[779] ) );
  AND U250 ( .A(B[1]), .B(A[777]), .Z(\P1[778] ) );
  AND U251 ( .A(B[1]), .B(A[776]), .Z(\P1[777] ) );
  AND U252 ( .A(B[1]), .B(A[775]), .Z(\P1[776] ) );
  AND U253 ( .A(B[1]), .B(A[774]), .Z(\P1[775] ) );
  AND U254 ( .A(B[1]), .B(A[773]), .Z(\P1[774] ) );
  AND U255 ( .A(B[1]), .B(A[772]), .Z(\P1[773] ) );
  AND U256 ( .A(B[1]), .B(A[771]), .Z(\P1[772] ) );
  AND U257 ( .A(B[1]), .B(A[770]), .Z(\P1[771] ) );
  AND U258 ( .A(B[1]), .B(A[769]), .Z(\P1[770] ) );
  AND U259 ( .A(B[1]), .B(A[75]), .Z(\P1[76] ) );
  AND U260 ( .A(B[1]), .B(A[768]), .Z(\P1[769] ) );
  AND U261 ( .A(B[1]), .B(A[767]), .Z(\P1[768] ) );
  AND U262 ( .A(B[1]), .B(A[766]), .Z(\P1[767] ) );
  AND U263 ( .A(B[1]), .B(A[765]), .Z(\P1[766] ) );
  AND U264 ( .A(B[1]), .B(A[764]), .Z(\P1[765] ) );
  AND U265 ( .A(B[1]), .B(A[763]), .Z(\P1[764] ) );
  AND U266 ( .A(B[1]), .B(A[762]), .Z(\P1[763] ) );
  AND U267 ( .A(B[1]), .B(A[761]), .Z(\P1[762] ) );
  AND U268 ( .A(B[1]), .B(A[760]), .Z(\P1[761] ) );
  AND U269 ( .A(B[1]), .B(A[759]), .Z(\P1[760] ) );
  AND U270 ( .A(B[1]), .B(A[74]), .Z(\P1[75] ) );
  AND U271 ( .A(B[1]), .B(A[758]), .Z(\P1[759] ) );
  AND U272 ( .A(B[1]), .B(A[757]), .Z(\P1[758] ) );
  AND U273 ( .A(B[1]), .B(A[756]), .Z(\P1[757] ) );
  AND U274 ( .A(B[1]), .B(A[755]), .Z(\P1[756] ) );
  AND U275 ( .A(B[1]), .B(A[754]), .Z(\P1[755] ) );
  AND U276 ( .A(B[1]), .B(A[753]), .Z(\P1[754] ) );
  AND U277 ( .A(B[1]), .B(A[752]), .Z(\P1[753] ) );
  AND U278 ( .A(B[1]), .B(A[751]), .Z(\P1[752] ) );
  AND U279 ( .A(B[1]), .B(A[750]), .Z(\P1[751] ) );
  AND U280 ( .A(B[1]), .B(A[749]), .Z(\P1[750] ) );
  AND U281 ( .A(B[1]), .B(A[73]), .Z(\P1[74] ) );
  AND U282 ( .A(B[1]), .B(A[748]), .Z(\P1[749] ) );
  AND U283 ( .A(B[1]), .B(A[747]), .Z(\P1[748] ) );
  AND U284 ( .A(B[1]), .B(A[746]), .Z(\P1[747] ) );
  AND U285 ( .A(B[1]), .B(A[745]), .Z(\P1[746] ) );
  AND U286 ( .A(B[1]), .B(A[744]), .Z(\P1[745] ) );
  AND U287 ( .A(B[1]), .B(A[743]), .Z(\P1[744] ) );
  AND U288 ( .A(B[1]), .B(A[742]), .Z(\P1[743] ) );
  AND U289 ( .A(B[1]), .B(A[741]), .Z(\P1[742] ) );
  AND U290 ( .A(B[1]), .B(A[740]), .Z(\P1[741] ) );
  AND U291 ( .A(B[1]), .B(A[739]), .Z(\P1[740] ) );
  AND U292 ( .A(B[1]), .B(A[72]), .Z(\P1[73] ) );
  AND U293 ( .A(B[1]), .B(A[738]), .Z(\P1[739] ) );
  AND U294 ( .A(B[1]), .B(A[737]), .Z(\P1[738] ) );
  AND U295 ( .A(B[1]), .B(A[736]), .Z(\P1[737] ) );
  AND U296 ( .A(B[1]), .B(A[735]), .Z(\P1[736] ) );
  AND U297 ( .A(B[1]), .B(A[734]), .Z(\P1[735] ) );
  AND U298 ( .A(B[1]), .B(A[733]), .Z(\P1[734] ) );
  AND U299 ( .A(B[1]), .B(A[732]), .Z(\P1[733] ) );
  AND U300 ( .A(B[1]), .B(A[731]), .Z(\P1[732] ) );
  AND U301 ( .A(B[1]), .B(A[730]), .Z(\P1[731] ) );
  AND U302 ( .A(B[1]), .B(A[729]), .Z(\P1[730] ) );
  AND U303 ( .A(B[1]), .B(A[71]), .Z(\P1[72] ) );
  AND U304 ( .A(B[1]), .B(A[728]), .Z(\P1[729] ) );
  AND U305 ( .A(B[1]), .B(A[727]), .Z(\P1[728] ) );
  AND U306 ( .A(B[1]), .B(A[726]), .Z(\P1[727] ) );
  AND U307 ( .A(B[1]), .B(A[725]), .Z(\P1[726] ) );
  AND U308 ( .A(B[1]), .B(A[724]), .Z(\P1[725] ) );
  AND U309 ( .A(B[1]), .B(A[723]), .Z(\P1[724] ) );
  AND U310 ( .A(B[1]), .B(A[722]), .Z(\P1[723] ) );
  AND U311 ( .A(B[1]), .B(A[721]), .Z(\P1[722] ) );
  AND U312 ( .A(B[1]), .B(A[720]), .Z(\P1[721] ) );
  AND U313 ( .A(B[1]), .B(A[719]), .Z(\P1[720] ) );
  AND U314 ( .A(B[1]), .B(A[70]), .Z(\P1[71] ) );
  AND U315 ( .A(B[1]), .B(A[718]), .Z(\P1[719] ) );
  AND U316 ( .A(B[1]), .B(A[717]), .Z(\P1[718] ) );
  AND U317 ( .A(B[1]), .B(A[716]), .Z(\P1[717] ) );
  AND U318 ( .A(B[1]), .B(A[715]), .Z(\P1[716] ) );
  AND U319 ( .A(B[1]), .B(A[714]), .Z(\P1[715] ) );
  AND U320 ( .A(B[1]), .B(A[713]), .Z(\P1[714] ) );
  AND U321 ( .A(B[1]), .B(A[712]), .Z(\P1[713] ) );
  AND U322 ( .A(B[1]), .B(A[711]), .Z(\P1[712] ) );
  AND U323 ( .A(B[1]), .B(A[710]), .Z(\P1[711] ) );
  AND U324 ( .A(B[1]), .B(A[709]), .Z(\P1[710] ) );
  AND U325 ( .A(B[1]), .B(A[69]), .Z(\P1[70] ) );
  AND U326 ( .A(B[1]), .B(A[708]), .Z(\P1[709] ) );
  AND U327 ( .A(B[1]), .B(A[707]), .Z(\P1[708] ) );
  AND U328 ( .A(B[1]), .B(A[706]), .Z(\P1[707] ) );
  AND U329 ( .A(B[1]), .B(A[705]), .Z(\P1[706] ) );
  AND U330 ( .A(B[1]), .B(A[704]), .Z(\P1[705] ) );
  AND U331 ( .A(B[1]), .B(A[703]), .Z(\P1[704] ) );
  AND U332 ( .A(B[1]), .B(A[702]), .Z(\P1[703] ) );
  AND U333 ( .A(B[1]), .B(A[701]), .Z(\P1[702] ) );
  AND U334 ( .A(B[1]), .B(A[700]), .Z(\P1[701] ) );
  AND U335 ( .A(B[1]), .B(A[699]), .Z(\P1[700] ) );
  AND U336 ( .A(B[1]), .B(A[5]), .Z(\P1[6] ) );
  AND U337 ( .A(B[1]), .B(A[68]), .Z(\P1[69] ) );
  AND U338 ( .A(B[1]), .B(A[698]), .Z(\P1[699] ) );
  AND U339 ( .A(B[1]), .B(A[697]), .Z(\P1[698] ) );
  AND U340 ( .A(B[1]), .B(A[696]), .Z(\P1[697] ) );
  AND U341 ( .A(B[1]), .B(A[695]), .Z(\P1[696] ) );
  AND U342 ( .A(B[1]), .B(A[694]), .Z(\P1[695] ) );
  AND U343 ( .A(B[1]), .B(A[693]), .Z(\P1[694] ) );
  AND U344 ( .A(B[1]), .B(A[692]), .Z(\P1[693] ) );
  AND U345 ( .A(B[1]), .B(A[691]), .Z(\P1[692] ) );
  AND U346 ( .A(B[1]), .B(A[690]), .Z(\P1[691] ) );
  AND U347 ( .A(B[1]), .B(A[689]), .Z(\P1[690] ) );
  AND U348 ( .A(B[1]), .B(A[67]), .Z(\P1[68] ) );
  AND U349 ( .A(B[1]), .B(A[688]), .Z(\P1[689] ) );
  AND U350 ( .A(B[1]), .B(A[687]), .Z(\P1[688] ) );
  AND U351 ( .A(B[1]), .B(A[686]), .Z(\P1[687] ) );
  AND U352 ( .A(B[1]), .B(A[685]), .Z(\P1[686] ) );
  AND U353 ( .A(B[1]), .B(A[684]), .Z(\P1[685] ) );
  AND U354 ( .A(B[1]), .B(A[683]), .Z(\P1[684] ) );
  AND U355 ( .A(B[1]), .B(A[682]), .Z(\P1[683] ) );
  AND U356 ( .A(B[1]), .B(A[681]), .Z(\P1[682] ) );
  AND U357 ( .A(B[1]), .B(A[680]), .Z(\P1[681] ) );
  AND U358 ( .A(B[1]), .B(A[679]), .Z(\P1[680] ) );
  AND U359 ( .A(B[1]), .B(A[66]), .Z(\P1[67] ) );
  AND U360 ( .A(B[1]), .B(A[678]), .Z(\P1[679] ) );
  AND U361 ( .A(B[1]), .B(A[677]), .Z(\P1[678] ) );
  AND U362 ( .A(B[1]), .B(A[676]), .Z(\P1[677] ) );
  AND U363 ( .A(B[1]), .B(A[675]), .Z(\P1[676] ) );
  AND U364 ( .A(B[1]), .B(A[674]), .Z(\P1[675] ) );
  AND U365 ( .A(B[1]), .B(A[673]), .Z(\P1[674] ) );
  AND U366 ( .A(B[1]), .B(A[672]), .Z(\P1[673] ) );
  AND U367 ( .A(B[1]), .B(A[671]), .Z(\P1[672] ) );
  AND U368 ( .A(B[1]), .B(A[670]), .Z(\P1[671] ) );
  AND U369 ( .A(B[1]), .B(A[669]), .Z(\P1[670] ) );
  AND U370 ( .A(B[1]), .B(A[65]), .Z(\P1[66] ) );
  AND U371 ( .A(B[1]), .B(A[668]), .Z(\P1[669] ) );
  AND U372 ( .A(B[1]), .B(A[667]), .Z(\P1[668] ) );
  AND U373 ( .A(B[1]), .B(A[666]), .Z(\P1[667] ) );
  AND U374 ( .A(B[1]), .B(A[665]), .Z(\P1[666] ) );
  AND U375 ( .A(B[1]), .B(A[664]), .Z(\P1[665] ) );
  AND U376 ( .A(B[1]), .B(A[663]), .Z(\P1[664] ) );
  AND U377 ( .A(B[1]), .B(A[662]), .Z(\P1[663] ) );
  AND U378 ( .A(B[1]), .B(A[661]), .Z(\P1[662] ) );
  AND U379 ( .A(B[1]), .B(A[660]), .Z(\P1[661] ) );
  AND U380 ( .A(B[1]), .B(A[659]), .Z(\P1[660] ) );
  AND U381 ( .A(B[1]), .B(A[64]), .Z(\P1[65] ) );
  AND U382 ( .A(B[1]), .B(A[658]), .Z(\P1[659] ) );
  AND U383 ( .A(B[1]), .B(A[657]), .Z(\P1[658] ) );
  AND U384 ( .A(B[1]), .B(A[656]), .Z(\P1[657] ) );
  AND U385 ( .A(B[1]), .B(A[655]), .Z(\P1[656] ) );
  AND U386 ( .A(B[1]), .B(A[654]), .Z(\P1[655] ) );
  AND U387 ( .A(B[1]), .B(A[653]), .Z(\P1[654] ) );
  AND U388 ( .A(B[1]), .B(A[652]), .Z(\P1[653] ) );
  AND U389 ( .A(B[1]), .B(A[651]), .Z(\P1[652] ) );
  AND U390 ( .A(B[1]), .B(A[650]), .Z(\P1[651] ) );
  AND U391 ( .A(B[1]), .B(A[649]), .Z(\P1[650] ) );
  AND U392 ( .A(B[1]), .B(A[63]), .Z(\P1[64] ) );
  AND U393 ( .A(B[1]), .B(A[648]), .Z(\P1[649] ) );
  AND U394 ( .A(B[1]), .B(A[647]), .Z(\P1[648] ) );
  AND U395 ( .A(B[1]), .B(A[646]), .Z(\P1[647] ) );
  AND U396 ( .A(B[1]), .B(A[645]), .Z(\P1[646] ) );
  AND U397 ( .A(B[1]), .B(A[644]), .Z(\P1[645] ) );
  AND U398 ( .A(B[1]), .B(A[643]), .Z(\P1[644] ) );
  AND U399 ( .A(B[1]), .B(A[642]), .Z(\P1[643] ) );
  AND U400 ( .A(B[1]), .B(A[641]), .Z(\P1[642] ) );
  AND U401 ( .A(B[1]), .B(A[640]), .Z(\P1[641] ) );
  AND U402 ( .A(B[1]), .B(A[639]), .Z(\P1[640] ) );
  AND U403 ( .A(B[1]), .B(A[62]), .Z(\P1[63] ) );
  AND U404 ( .A(B[1]), .B(A[638]), .Z(\P1[639] ) );
  AND U405 ( .A(B[1]), .B(A[637]), .Z(\P1[638] ) );
  AND U406 ( .A(B[1]), .B(A[636]), .Z(\P1[637] ) );
  AND U407 ( .A(B[1]), .B(A[635]), .Z(\P1[636] ) );
  AND U408 ( .A(B[1]), .B(A[634]), .Z(\P1[635] ) );
  AND U409 ( .A(B[1]), .B(A[633]), .Z(\P1[634] ) );
  AND U410 ( .A(B[1]), .B(A[632]), .Z(\P1[633] ) );
  AND U411 ( .A(B[1]), .B(A[631]), .Z(\P1[632] ) );
  AND U412 ( .A(B[1]), .B(A[630]), .Z(\P1[631] ) );
  AND U413 ( .A(B[1]), .B(A[629]), .Z(\P1[630] ) );
  AND U414 ( .A(B[1]), .B(A[61]), .Z(\P1[62] ) );
  AND U415 ( .A(B[1]), .B(A[628]), .Z(\P1[629] ) );
  AND U416 ( .A(B[1]), .B(A[627]), .Z(\P1[628] ) );
  AND U417 ( .A(B[1]), .B(A[626]), .Z(\P1[627] ) );
  AND U418 ( .A(B[1]), .B(A[625]), .Z(\P1[626] ) );
  AND U419 ( .A(B[1]), .B(A[624]), .Z(\P1[625] ) );
  AND U420 ( .A(B[1]), .B(A[623]), .Z(\P1[624] ) );
  AND U421 ( .A(B[1]), .B(A[622]), .Z(\P1[623] ) );
  AND U422 ( .A(B[1]), .B(A[621]), .Z(\P1[622] ) );
  AND U423 ( .A(B[1]), .B(A[620]), .Z(\P1[621] ) );
  AND U424 ( .A(B[1]), .B(A[619]), .Z(\P1[620] ) );
  AND U425 ( .A(B[1]), .B(A[60]), .Z(\P1[61] ) );
  AND U426 ( .A(B[1]), .B(A[618]), .Z(\P1[619] ) );
  AND U427 ( .A(B[1]), .B(A[617]), .Z(\P1[618] ) );
  AND U428 ( .A(B[1]), .B(A[616]), .Z(\P1[617] ) );
  AND U429 ( .A(B[1]), .B(A[615]), .Z(\P1[616] ) );
  AND U430 ( .A(B[1]), .B(A[614]), .Z(\P1[615] ) );
  AND U431 ( .A(B[1]), .B(A[613]), .Z(\P1[614] ) );
  AND U432 ( .A(B[1]), .B(A[612]), .Z(\P1[613] ) );
  AND U433 ( .A(B[1]), .B(A[611]), .Z(\P1[612] ) );
  AND U434 ( .A(B[1]), .B(A[610]), .Z(\P1[611] ) );
  AND U435 ( .A(B[1]), .B(A[609]), .Z(\P1[610] ) );
  AND U436 ( .A(B[1]), .B(A[59]), .Z(\P1[60] ) );
  AND U437 ( .A(B[1]), .B(A[608]), .Z(\P1[609] ) );
  AND U438 ( .A(B[1]), .B(A[607]), .Z(\P1[608] ) );
  AND U439 ( .A(B[1]), .B(A[606]), .Z(\P1[607] ) );
  AND U440 ( .A(B[1]), .B(A[605]), .Z(\P1[606] ) );
  AND U441 ( .A(B[1]), .B(A[604]), .Z(\P1[605] ) );
  AND U442 ( .A(B[1]), .B(A[603]), .Z(\P1[604] ) );
  AND U443 ( .A(B[1]), .B(A[602]), .Z(\P1[603] ) );
  AND U444 ( .A(B[1]), .B(A[601]), .Z(\P1[602] ) );
  AND U445 ( .A(B[1]), .B(A[600]), .Z(\P1[601] ) );
  AND U446 ( .A(B[1]), .B(A[599]), .Z(\P1[600] ) );
  AND U447 ( .A(B[1]), .B(A[4]), .Z(\P1[5] ) );
  AND U448 ( .A(B[1]), .B(A[58]), .Z(\P1[59] ) );
  AND U449 ( .A(B[1]), .B(A[598]), .Z(\P1[599] ) );
  AND U450 ( .A(B[1]), .B(A[597]), .Z(\P1[598] ) );
  AND U451 ( .A(B[1]), .B(A[596]), .Z(\P1[597] ) );
  AND U452 ( .A(B[1]), .B(A[595]), .Z(\P1[596] ) );
  AND U453 ( .A(B[1]), .B(A[594]), .Z(\P1[595] ) );
  AND U454 ( .A(B[1]), .B(A[593]), .Z(\P1[594] ) );
  AND U455 ( .A(B[1]), .B(A[592]), .Z(\P1[593] ) );
  AND U456 ( .A(B[1]), .B(A[591]), .Z(\P1[592] ) );
  AND U457 ( .A(B[1]), .B(A[590]), .Z(\P1[591] ) );
  AND U458 ( .A(B[1]), .B(A[589]), .Z(\P1[590] ) );
  AND U459 ( .A(B[1]), .B(A[57]), .Z(\P1[58] ) );
  AND U460 ( .A(B[1]), .B(A[588]), .Z(\P1[589] ) );
  AND U461 ( .A(B[1]), .B(A[587]), .Z(\P1[588] ) );
  AND U462 ( .A(B[1]), .B(A[586]), .Z(\P1[587] ) );
  AND U463 ( .A(B[1]), .B(A[585]), .Z(\P1[586] ) );
  AND U464 ( .A(B[1]), .B(A[584]), .Z(\P1[585] ) );
  AND U465 ( .A(B[1]), .B(A[583]), .Z(\P1[584] ) );
  AND U466 ( .A(B[1]), .B(A[582]), .Z(\P1[583] ) );
  AND U467 ( .A(B[1]), .B(A[581]), .Z(\P1[582] ) );
  AND U468 ( .A(B[1]), .B(A[580]), .Z(\P1[581] ) );
  AND U469 ( .A(B[1]), .B(A[579]), .Z(\P1[580] ) );
  AND U470 ( .A(B[1]), .B(A[56]), .Z(\P1[57] ) );
  AND U471 ( .A(B[1]), .B(A[578]), .Z(\P1[579] ) );
  AND U472 ( .A(B[1]), .B(A[577]), .Z(\P1[578] ) );
  AND U473 ( .A(B[1]), .B(A[576]), .Z(\P1[577] ) );
  AND U474 ( .A(B[1]), .B(A[575]), .Z(\P1[576] ) );
  AND U475 ( .A(B[1]), .B(A[574]), .Z(\P1[575] ) );
  AND U476 ( .A(B[1]), .B(A[573]), .Z(\P1[574] ) );
  AND U477 ( .A(B[1]), .B(A[572]), .Z(\P1[573] ) );
  AND U478 ( .A(B[1]), .B(A[571]), .Z(\P1[572] ) );
  AND U479 ( .A(B[1]), .B(A[570]), .Z(\P1[571] ) );
  AND U480 ( .A(B[1]), .B(A[569]), .Z(\P1[570] ) );
  AND U481 ( .A(B[1]), .B(A[55]), .Z(\P1[56] ) );
  AND U482 ( .A(B[1]), .B(A[568]), .Z(\P1[569] ) );
  AND U483 ( .A(B[1]), .B(A[567]), .Z(\P1[568] ) );
  AND U484 ( .A(B[1]), .B(A[566]), .Z(\P1[567] ) );
  AND U485 ( .A(B[1]), .B(A[565]), .Z(\P1[566] ) );
  AND U486 ( .A(B[1]), .B(A[564]), .Z(\P1[565] ) );
  AND U487 ( .A(B[1]), .B(A[563]), .Z(\P1[564] ) );
  AND U488 ( .A(B[1]), .B(A[562]), .Z(\P1[563] ) );
  AND U489 ( .A(B[1]), .B(A[561]), .Z(\P1[562] ) );
  AND U490 ( .A(B[1]), .B(A[560]), .Z(\P1[561] ) );
  AND U491 ( .A(B[1]), .B(A[559]), .Z(\P1[560] ) );
  AND U492 ( .A(B[1]), .B(A[54]), .Z(\P1[55] ) );
  AND U493 ( .A(B[1]), .B(A[558]), .Z(\P1[559] ) );
  AND U494 ( .A(B[1]), .B(A[557]), .Z(\P1[558] ) );
  AND U495 ( .A(B[1]), .B(A[556]), .Z(\P1[557] ) );
  AND U496 ( .A(B[1]), .B(A[555]), .Z(\P1[556] ) );
  AND U497 ( .A(B[1]), .B(A[554]), .Z(\P1[555] ) );
  AND U498 ( .A(B[1]), .B(A[553]), .Z(\P1[554] ) );
  AND U499 ( .A(B[1]), .B(A[552]), .Z(\P1[553] ) );
  AND U500 ( .A(B[1]), .B(A[551]), .Z(\P1[552] ) );
  AND U501 ( .A(B[1]), .B(A[550]), .Z(\P1[551] ) );
  AND U502 ( .A(B[1]), .B(A[549]), .Z(\P1[550] ) );
  AND U503 ( .A(B[1]), .B(A[53]), .Z(\P1[54] ) );
  AND U504 ( .A(B[1]), .B(A[548]), .Z(\P1[549] ) );
  AND U505 ( .A(B[1]), .B(A[547]), .Z(\P1[548] ) );
  AND U506 ( .A(B[1]), .B(A[546]), .Z(\P1[547] ) );
  AND U507 ( .A(B[1]), .B(A[545]), .Z(\P1[546] ) );
  AND U508 ( .A(B[1]), .B(A[544]), .Z(\P1[545] ) );
  AND U509 ( .A(B[1]), .B(A[543]), .Z(\P1[544] ) );
  AND U510 ( .A(B[1]), .B(A[542]), .Z(\P1[543] ) );
  AND U511 ( .A(B[1]), .B(A[541]), .Z(\P1[542] ) );
  AND U512 ( .A(B[1]), .B(A[540]), .Z(\P1[541] ) );
  AND U513 ( .A(B[1]), .B(A[539]), .Z(\P1[540] ) );
  AND U514 ( .A(B[1]), .B(A[52]), .Z(\P1[53] ) );
  AND U515 ( .A(B[1]), .B(A[538]), .Z(\P1[539] ) );
  AND U516 ( .A(B[1]), .B(A[537]), .Z(\P1[538] ) );
  AND U517 ( .A(B[1]), .B(A[536]), .Z(\P1[537] ) );
  AND U518 ( .A(B[1]), .B(A[535]), .Z(\P1[536] ) );
  AND U519 ( .A(B[1]), .B(A[534]), .Z(\P1[535] ) );
  AND U520 ( .A(B[1]), .B(A[533]), .Z(\P1[534] ) );
  AND U521 ( .A(B[1]), .B(A[532]), .Z(\P1[533] ) );
  AND U522 ( .A(B[1]), .B(A[531]), .Z(\P1[532] ) );
  AND U523 ( .A(B[1]), .B(A[530]), .Z(\P1[531] ) );
  AND U524 ( .A(B[1]), .B(A[529]), .Z(\P1[530] ) );
  AND U525 ( .A(B[1]), .B(A[51]), .Z(\P1[52] ) );
  AND U526 ( .A(B[1]), .B(A[528]), .Z(\P1[529] ) );
  AND U527 ( .A(B[1]), .B(A[527]), .Z(\P1[528] ) );
  AND U528 ( .A(B[1]), .B(A[526]), .Z(\P1[527] ) );
  AND U529 ( .A(B[1]), .B(A[525]), .Z(\P1[526] ) );
  AND U530 ( .A(B[1]), .B(A[524]), .Z(\P1[525] ) );
  AND U531 ( .A(B[1]), .B(A[523]), .Z(\P1[524] ) );
  AND U532 ( .A(B[1]), .B(A[522]), .Z(\P1[523] ) );
  AND U533 ( .A(B[1]), .B(A[521]), .Z(\P1[522] ) );
  AND U534 ( .A(B[1]), .B(A[520]), .Z(\P1[521] ) );
  AND U535 ( .A(B[1]), .B(A[519]), .Z(\P1[520] ) );
  AND U536 ( .A(B[1]), .B(A[50]), .Z(\P1[51] ) );
  AND U537 ( .A(B[1]), .B(A[518]), .Z(\P1[519] ) );
  AND U538 ( .A(B[1]), .B(A[517]), .Z(\P1[518] ) );
  AND U539 ( .A(B[1]), .B(A[516]), .Z(\P1[517] ) );
  AND U540 ( .A(B[1]), .B(A[515]), .Z(\P1[516] ) );
  AND U541 ( .A(B[1]), .B(A[514]), .Z(\P1[515] ) );
  AND U542 ( .A(B[1]), .B(A[513]), .Z(\P1[514] ) );
  AND U543 ( .A(B[1]), .B(A[512]), .Z(\P1[513] ) );
  AND U544 ( .A(B[1]), .B(A[511]), .Z(\P1[512] ) );
  AND U545 ( .A(B[1]), .B(A[510]), .Z(\P1[511] ) );
  AND U546 ( .A(B[1]), .B(A[509]), .Z(\P1[510] ) );
  AND U547 ( .A(B[1]), .B(A[49]), .Z(\P1[50] ) );
  AND U548 ( .A(B[1]), .B(A[508]), .Z(\P1[509] ) );
  AND U549 ( .A(B[1]), .B(A[507]), .Z(\P1[508] ) );
  AND U550 ( .A(B[1]), .B(A[506]), .Z(\P1[507] ) );
  AND U551 ( .A(B[1]), .B(A[505]), .Z(\P1[506] ) );
  AND U552 ( .A(B[1]), .B(A[504]), .Z(\P1[505] ) );
  AND U553 ( .A(B[1]), .B(A[503]), .Z(\P1[504] ) );
  AND U554 ( .A(B[1]), .B(A[502]), .Z(\P1[503] ) );
  AND U555 ( .A(B[1]), .B(A[501]), .Z(\P1[502] ) );
  AND U556 ( .A(B[1]), .B(A[500]), .Z(\P1[501] ) );
  AND U557 ( .A(B[1]), .B(A[499]), .Z(\P1[500] ) );
  AND U558 ( .A(B[1]), .B(A[3]), .Z(\P1[4] ) );
  AND U559 ( .A(B[1]), .B(A[48]), .Z(\P1[49] ) );
  AND U560 ( .A(B[1]), .B(A[498]), .Z(\P1[499] ) );
  AND U561 ( .A(B[1]), .B(A[497]), .Z(\P1[498] ) );
  AND U562 ( .A(B[1]), .B(A[496]), .Z(\P1[497] ) );
  AND U563 ( .A(B[1]), .B(A[495]), .Z(\P1[496] ) );
  AND U564 ( .A(B[1]), .B(A[494]), .Z(\P1[495] ) );
  AND U565 ( .A(B[1]), .B(A[493]), .Z(\P1[494] ) );
  AND U566 ( .A(B[1]), .B(A[492]), .Z(\P1[493] ) );
  AND U567 ( .A(B[1]), .B(A[491]), .Z(\P1[492] ) );
  AND U568 ( .A(B[1]), .B(A[490]), .Z(\P1[491] ) );
  AND U569 ( .A(B[1]), .B(A[489]), .Z(\P1[490] ) );
  AND U570 ( .A(B[1]), .B(A[47]), .Z(\P1[48] ) );
  AND U571 ( .A(B[1]), .B(A[488]), .Z(\P1[489] ) );
  AND U572 ( .A(B[1]), .B(A[487]), .Z(\P1[488] ) );
  AND U573 ( .A(B[1]), .B(A[486]), .Z(\P1[487] ) );
  AND U574 ( .A(B[1]), .B(A[485]), .Z(\P1[486] ) );
  AND U575 ( .A(B[1]), .B(A[484]), .Z(\P1[485] ) );
  AND U576 ( .A(B[1]), .B(A[483]), .Z(\P1[484] ) );
  AND U577 ( .A(B[1]), .B(A[482]), .Z(\P1[483] ) );
  AND U578 ( .A(B[1]), .B(A[481]), .Z(\P1[482] ) );
  AND U579 ( .A(B[1]), .B(A[480]), .Z(\P1[481] ) );
  AND U580 ( .A(B[1]), .B(A[479]), .Z(\P1[480] ) );
  AND U581 ( .A(B[1]), .B(A[46]), .Z(\P1[47] ) );
  AND U582 ( .A(B[1]), .B(A[478]), .Z(\P1[479] ) );
  AND U583 ( .A(B[1]), .B(A[477]), .Z(\P1[478] ) );
  AND U584 ( .A(B[1]), .B(A[476]), .Z(\P1[477] ) );
  AND U585 ( .A(B[1]), .B(A[475]), .Z(\P1[476] ) );
  AND U586 ( .A(B[1]), .B(A[474]), .Z(\P1[475] ) );
  AND U587 ( .A(B[1]), .B(A[473]), .Z(\P1[474] ) );
  AND U588 ( .A(B[1]), .B(A[472]), .Z(\P1[473] ) );
  AND U589 ( .A(B[1]), .B(A[471]), .Z(\P1[472] ) );
  AND U590 ( .A(B[1]), .B(A[470]), .Z(\P1[471] ) );
  AND U591 ( .A(B[1]), .B(A[469]), .Z(\P1[470] ) );
  AND U592 ( .A(B[1]), .B(A[45]), .Z(\P1[46] ) );
  AND U593 ( .A(B[1]), .B(A[468]), .Z(\P1[469] ) );
  AND U594 ( .A(B[1]), .B(A[467]), .Z(\P1[468] ) );
  AND U595 ( .A(B[1]), .B(A[466]), .Z(\P1[467] ) );
  AND U596 ( .A(B[1]), .B(A[465]), .Z(\P1[466] ) );
  AND U597 ( .A(B[1]), .B(A[464]), .Z(\P1[465] ) );
  AND U598 ( .A(B[1]), .B(A[463]), .Z(\P1[464] ) );
  AND U599 ( .A(B[1]), .B(A[462]), .Z(\P1[463] ) );
  AND U600 ( .A(B[1]), .B(A[461]), .Z(\P1[462] ) );
  AND U601 ( .A(B[1]), .B(A[460]), .Z(\P1[461] ) );
  AND U602 ( .A(B[1]), .B(A[459]), .Z(\P1[460] ) );
  AND U603 ( .A(B[1]), .B(A[44]), .Z(\P1[45] ) );
  AND U604 ( .A(B[1]), .B(A[458]), .Z(\P1[459] ) );
  AND U605 ( .A(B[1]), .B(A[457]), .Z(\P1[458] ) );
  AND U606 ( .A(B[1]), .B(A[456]), .Z(\P1[457] ) );
  AND U607 ( .A(B[1]), .B(A[455]), .Z(\P1[456] ) );
  AND U608 ( .A(B[1]), .B(A[454]), .Z(\P1[455] ) );
  AND U609 ( .A(B[1]), .B(A[453]), .Z(\P1[454] ) );
  AND U610 ( .A(B[1]), .B(A[452]), .Z(\P1[453] ) );
  AND U611 ( .A(B[1]), .B(A[451]), .Z(\P1[452] ) );
  AND U612 ( .A(B[1]), .B(A[450]), .Z(\P1[451] ) );
  AND U613 ( .A(B[1]), .B(A[449]), .Z(\P1[450] ) );
  AND U614 ( .A(B[1]), .B(A[43]), .Z(\P1[44] ) );
  AND U615 ( .A(B[1]), .B(A[448]), .Z(\P1[449] ) );
  AND U616 ( .A(B[1]), .B(A[447]), .Z(\P1[448] ) );
  AND U617 ( .A(B[1]), .B(A[446]), .Z(\P1[447] ) );
  AND U618 ( .A(B[1]), .B(A[445]), .Z(\P1[446] ) );
  AND U619 ( .A(B[1]), .B(A[444]), .Z(\P1[445] ) );
  AND U620 ( .A(B[1]), .B(A[443]), .Z(\P1[444] ) );
  AND U621 ( .A(B[1]), .B(A[442]), .Z(\P1[443] ) );
  AND U622 ( .A(B[1]), .B(A[441]), .Z(\P1[442] ) );
  AND U623 ( .A(B[1]), .B(A[440]), .Z(\P1[441] ) );
  AND U624 ( .A(B[1]), .B(A[439]), .Z(\P1[440] ) );
  AND U625 ( .A(B[1]), .B(A[42]), .Z(\P1[43] ) );
  AND U626 ( .A(B[1]), .B(A[438]), .Z(\P1[439] ) );
  AND U627 ( .A(B[1]), .B(A[437]), .Z(\P1[438] ) );
  AND U628 ( .A(B[1]), .B(A[436]), .Z(\P1[437] ) );
  AND U629 ( .A(B[1]), .B(A[435]), .Z(\P1[436] ) );
  AND U630 ( .A(B[1]), .B(A[434]), .Z(\P1[435] ) );
  AND U631 ( .A(B[1]), .B(A[433]), .Z(\P1[434] ) );
  AND U632 ( .A(B[1]), .B(A[432]), .Z(\P1[433] ) );
  AND U633 ( .A(B[1]), .B(A[431]), .Z(\P1[432] ) );
  AND U634 ( .A(B[1]), .B(A[430]), .Z(\P1[431] ) );
  AND U635 ( .A(B[1]), .B(A[429]), .Z(\P1[430] ) );
  AND U636 ( .A(B[1]), .B(A[41]), .Z(\P1[42] ) );
  AND U637 ( .A(B[1]), .B(A[428]), .Z(\P1[429] ) );
  AND U638 ( .A(B[1]), .B(A[427]), .Z(\P1[428] ) );
  AND U639 ( .A(B[1]), .B(A[426]), .Z(\P1[427] ) );
  AND U640 ( .A(B[1]), .B(A[425]), .Z(\P1[426] ) );
  AND U641 ( .A(B[1]), .B(A[424]), .Z(\P1[425] ) );
  AND U642 ( .A(B[1]), .B(A[423]), .Z(\P1[424] ) );
  AND U643 ( .A(B[1]), .B(A[422]), .Z(\P1[423] ) );
  AND U644 ( .A(B[1]), .B(A[421]), .Z(\P1[422] ) );
  AND U645 ( .A(B[1]), .B(A[420]), .Z(\P1[421] ) );
  AND U646 ( .A(B[1]), .B(A[419]), .Z(\P1[420] ) );
  AND U647 ( .A(B[1]), .B(A[40]), .Z(\P1[41] ) );
  AND U648 ( .A(B[1]), .B(A[418]), .Z(\P1[419] ) );
  AND U649 ( .A(B[1]), .B(A[417]), .Z(\P1[418] ) );
  AND U650 ( .A(B[1]), .B(A[416]), .Z(\P1[417] ) );
  AND U651 ( .A(B[1]), .B(A[415]), .Z(\P1[416] ) );
  AND U652 ( .A(B[1]), .B(A[414]), .Z(\P1[415] ) );
  AND U653 ( .A(B[1]), .B(A[413]), .Z(\P1[414] ) );
  AND U654 ( .A(B[1]), .B(A[412]), .Z(\P1[413] ) );
  AND U655 ( .A(B[1]), .B(A[411]), .Z(\P1[412] ) );
  AND U656 ( .A(B[1]), .B(A[410]), .Z(\P1[411] ) );
  AND U657 ( .A(B[1]), .B(A[409]), .Z(\P1[410] ) );
  AND U658 ( .A(B[1]), .B(A[39]), .Z(\P1[40] ) );
  AND U659 ( .A(B[1]), .B(A[408]), .Z(\P1[409] ) );
  AND U660 ( .A(B[1]), .B(A[407]), .Z(\P1[408] ) );
  AND U661 ( .A(B[1]), .B(A[406]), .Z(\P1[407] ) );
  AND U662 ( .A(B[1]), .B(A[405]), .Z(\P1[406] ) );
  AND U663 ( .A(B[1]), .B(A[404]), .Z(\P1[405] ) );
  AND U664 ( .A(B[1]), .B(A[403]), .Z(\P1[404] ) );
  AND U665 ( .A(B[1]), .B(A[402]), .Z(\P1[403] ) );
  AND U666 ( .A(B[1]), .B(A[401]), .Z(\P1[402] ) );
  AND U667 ( .A(B[1]), .B(A[400]), .Z(\P1[401] ) );
  AND U668 ( .A(B[1]), .B(A[399]), .Z(\P1[400] ) );
  AND U669 ( .A(B[1]), .B(A[2]), .Z(\P1[3] ) );
  AND U670 ( .A(B[1]), .B(A[38]), .Z(\P1[39] ) );
  AND U671 ( .A(B[1]), .B(A[398]), .Z(\P1[399] ) );
  AND U672 ( .A(B[1]), .B(A[397]), .Z(\P1[398] ) );
  AND U673 ( .A(B[1]), .B(A[396]), .Z(\P1[397] ) );
  AND U674 ( .A(B[1]), .B(A[395]), .Z(\P1[396] ) );
  AND U675 ( .A(B[1]), .B(A[394]), .Z(\P1[395] ) );
  AND U676 ( .A(B[1]), .B(A[393]), .Z(\P1[394] ) );
  AND U677 ( .A(B[1]), .B(A[392]), .Z(\P1[393] ) );
  AND U678 ( .A(B[1]), .B(A[391]), .Z(\P1[392] ) );
  AND U679 ( .A(B[1]), .B(A[390]), .Z(\P1[391] ) );
  AND U680 ( .A(B[1]), .B(A[389]), .Z(\P1[390] ) );
  AND U681 ( .A(B[1]), .B(A[37]), .Z(\P1[38] ) );
  AND U682 ( .A(B[1]), .B(A[388]), .Z(\P1[389] ) );
  AND U683 ( .A(B[1]), .B(A[387]), .Z(\P1[388] ) );
  AND U684 ( .A(B[1]), .B(A[386]), .Z(\P1[387] ) );
  AND U685 ( .A(B[1]), .B(A[385]), .Z(\P1[386] ) );
  AND U686 ( .A(B[1]), .B(A[384]), .Z(\P1[385] ) );
  AND U687 ( .A(B[1]), .B(A[383]), .Z(\P1[384] ) );
  AND U688 ( .A(B[1]), .B(A[382]), .Z(\P1[383] ) );
  AND U689 ( .A(B[1]), .B(A[381]), .Z(\P1[382] ) );
  AND U690 ( .A(B[1]), .B(A[380]), .Z(\P1[381] ) );
  AND U691 ( .A(B[1]), .B(A[379]), .Z(\P1[380] ) );
  AND U692 ( .A(B[1]), .B(A[36]), .Z(\P1[37] ) );
  AND U693 ( .A(B[1]), .B(A[378]), .Z(\P1[379] ) );
  AND U694 ( .A(B[1]), .B(A[377]), .Z(\P1[378] ) );
  AND U695 ( .A(B[1]), .B(A[376]), .Z(\P1[377] ) );
  AND U696 ( .A(B[1]), .B(A[375]), .Z(\P1[376] ) );
  AND U697 ( .A(B[1]), .B(A[374]), .Z(\P1[375] ) );
  AND U698 ( .A(B[1]), .B(A[373]), .Z(\P1[374] ) );
  AND U699 ( .A(B[1]), .B(A[372]), .Z(\P1[373] ) );
  AND U700 ( .A(B[1]), .B(A[371]), .Z(\P1[372] ) );
  AND U701 ( .A(B[1]), .B(A[370]), .Z(\P1[371] ) );
  AND U702 ( .A(B[1]), .B(A[369]), .Z(\P1[370] ) );
  AND U703 ( .A(B[1]), .B(A[35]), .Z(\P1[36] ) );
  AND U704 ( .A(B[1]), .B(A[368]), .Z(\P1[369] ) );
  AND U705 ( .A(B[1]), .B(A[367]), .Z(\P1[368] ) );
  AND U706 ( .A(B[1]), .B(A[366]), .Z(\P1[367] ) );
  AND U707 ( .A(B[1]), .B(A[365]), .Z(\P1[366] ) );
  AND U708 ( .A(B[1]), .B(A[364]), .Z(\P1[365] ) );
  AND U709 ( .A(B[1]), .B(A[363]), .Z(\P1[364] ) );
  AND U710 ( .A(B[1]), .B(A[362]), .Z(\P1[363] ) );
  AND U711 ( .A(B[1]), .B(A[361]), .Z(\P1[362] ) );
  AND U712 ( .A(B[1]), .B(A[360]), .Z(\P1[361] ) );
  AND U713 ( .A(B[1]), .B(A[359]), .Z(\P1[360] ) );
  AND U714 ( .A(B[1]), .B(A[34]), .Z(\P1[35] ) );
  AND U715 ( .A(B[1]), .B(A[358]), .Z(\P1[359] ) );
  AND U716 ( .A(B[1]), .B(A[357]), .Z(\P1[358] ) );
  AND U717 ( .A(B[1]), .B(A[356]), .Z(\P1[357] ) );
  AND U718 ( .A(B[1]), .B(A[355]), .Z(\P1[356] ) );
  AND U719 ( .A(B[1]), .B(A[354]), .Z(\P1[355] ) );
  AND U720 ( .A(B[1]), .B(A[353]), .Z(\P1[354] ) );
  AND U721 ( .A(B[1]), .B(A[352]), .Z(\P1[353] ) );
  AND U722 ( .A(B[1]), .B(A[351]), .Z(\P1[352] ) );
  AND U723 ( .A(B[1]), .B(A[350]), .Z(\P1[351] ) );
  AND U724 ( .A(B[1]), .B(A[349]), .Z(\P1[350] ) );
  AND U725 ( .A(B[1]), .B(A[33]), .Z(\P1[34] ) );
  AND U726 ( .A(B[1]), .B(A[348]), .Z(\P1[349] ) );
  AND U727 ( .A(B[1]), .B(A[347]), .Z(\P1[348] ) );
  AND U728 ( .A(B[1]), .B(A[346]), .Z(\P1[347] ) );
  AND U729 ( .A(B[1]), .B(A[345]), .Z(\P1[346] ) );
  AND U730 ( .A(B[1]), .B(A[344]), .Z(\P1[345] ) );
  AND U731 ( .A(B[1]), .B(A[343]), .Z(\P1[344] ) );
  AND U732 ( .A(B[1]), .B(A[342]), .Z(\P1[343] ) );
  AND U733 ( .A(B[1]), .B(A[341]), .Z(\P1[342] ) );
  AND U734 ( .A(B[1]), .B(A[340]), .Z(\P1[341] ) );
  AND U735 ( .A(B[1]), .B(A[339]), .Z(\P1[340] ) );
  AND U736 ( .A(B[1]), .B(A[32]), .Z(\P1[33] ) );
  AND U737 ( .A(B[1]), .B(A[338]), .Z(\P1[339] ) );
  AND U738 ( .A(B[1]), .B(A[337]), .Z(\P1[338] ) );
  AND U739 ( .A(B[1]), .B(A[336]), .Z(\P1[337] ) );
  AND U740 ( .A(B[1]), .B(A[335]), .Z(\P1[336] ) );
  AND U741 ( .A(B[1]), .B(A[334]), .Z(\P1[335] ) );
  AND U742 ( .A(B[1]), .B(A[333]), .Z(\P1[334] ) );
  AND U743 ( .A(B[1]), .B(A[332]), .Z(\P1[333] ) );
  AND U744 ( .A(B[1]), .B(A[331]), .Z(\P1[332] ) );
  AND U745 ( .A(B[1]), .B(A[330]), .Z(\P1[331] ) );
  AND U746 ( .A(B[1]), .B(A[329]), .Z(\P1[330] ) );
  AND U747 ( .A(B[1]), .B(A[31]), .Z(\P1[32] ) );
  AND U748 ( .A(B[1]), .B(A[328]), .Z(\P1[329] ) );
  AND U749 ( .A(B[1]), .B(A[327]), .Z(\P1[328] ) );
  AND U750 ( .A(B[1]), .B(A[326]), .Z(\P1[327] ) );
  AND U751 ( .A(B[1]), .B(A[325]), .Z(\P1[326] ) );
  AND U752 ( .A(B[1]), .B(A[324]), .Z(\P1[325] ) );
  AND U753 ( .A(B[1]), .B(A[323]), .Z(\P1[324] ) );
  AND U754 ( .A(B[1]), .B(A[322]), .Z(\P1[323] ) );
  AND U755 ( .A(B[1]), .B(A[321]), .Z(\P1[322] ) );
  AND U756 ( .A(B[1]), .B(A[320]), .Z(\P1[321] ) );
  AND U757 ( .A(B[1]), .B(A[319]), .Z(\P1[320] ) );
  AND U758 ( .A(B[1]), .B(A[30]), .Z(\P1[31] ) );
  AND U759 ( .A(B[1]), .B(A[318]), .Z(\P1[319] ) );
  AND U760 ( .A(B[1]), .B(A[317]), .Z(\P1[318] ) );
  AND U761 ( .A(B[1]), .B(A[316]), .Z(\P1[317] ) );
  AND U762 ( .A(B[1]), .B(A[315]), .Z(\P1[316] ) );
  AND U763 ( .A(B[1]), .B(A[314]), .Z(\P1[315] ) );
  AND U764 ( .A(B[1]), .B(A[313]), .Z(\P1[314] ) );
  AND U765 ( .A(B[1]), .B(A[312]), .Z(\P1[313] ) );
  AND U766 ( .A(B[1]), .B(A[311]), .Z(\P1[312] ) );
  AND U767 ( .A(B[1]), .B(A[310]), .Z(\P1[311] ) );
  AND U768 ( .A(B[1]), .B(A[309]), .Z(\P1[310] ) );
  AND U769 ( .A(B[1]), .B(A[29]), .Z(\P1[30] ) );
  AND U770 ( .A(B[1]), .B(A[308]), .Z(\P1[309] ) );
  AND U771 ( .A(B[1]), .B(A[307]), .Z(\P1[308] ) );
  AND U772 ( .A(B[1]), .B(A[306]), .Z(\P1[307] ) );
  AND U773 ( .A(B[1]), .B(A[305]), .Z(\P1[306] ) );
  AND U774 ( .A(B[1]), .B(A[304]), .Z(\P1[305] ) );
  AND U775 ( .A(B[1]), .B(A[303]), .Z(\P1[304] ) );
  AND U776 ( .A(B[1]), .B(A[302]), .Z(\P1[303] ) );
  AND U777 ( .A(B[1]), .B(A[301]), .Z(\P1[302] ) );
  AND U778 ( .A(B[1]), .B(A[300]), .Z(\P1[301] ) );
  AND U779 ( .A(B[1]), .B(A[299]), .Z(\P1[300] ) );
  AND U780 ( .A(B[1]), .B(A[1]), .Z(\P1[2] ) );
  AND U781 ( .A(B[1]), .B(A[28]), .Z(\P1[29] ) );
  AND U782 ( .A(B[1]), .B(A[298]), .Z(\P1[299] ) );
  AND U783 ( .A(B[1]), .B(A[297]), .Z(\P1[298] ) );
  AND U784 ( .A(B[1]), .B(A[296]), .Z(\P1[297] ) );
  AND U785 ( .A(B[1]), .B(A[295]), .Z(\P1[296] ) );
  AND U786 ( .A(B[1]), .B(A[294]), .Z(\P1[295] ) );
  AND U787 ( .A(B[1]), .B(A[293]), .Z(\P1[294] ) );
  AND U788 ( .A(B[1]), .B(A[292]), .Z(\P1[293] ) );
  AND U789 ( .A(B[1]), .B(A[291]), .Z(\P1[292] ) );
  AND U790 ( .A(B[1]), .B(A[290]), .Z(\P1[291] ) );
  AND U791 ( .A(B[1]), .B(A[289]), .Z(\P1[290] ) );
  AND U792 ( .A(B[1]), .B(A[27]), .Z(\P1[28] ) );
  AND U793 ( .A(B[1]), .B(A[288]), .Z(\P1[289] ) );
  AND U794 ( .A(B[1]), .B(A[287]), .Z(\P1[288] ) );
  AND U795 ( .A(B[1]), .B(A[286]), .Z(\P1[287] ) );
  AND U796 ( .A(B[1]), .B(A[285]), .Z(\P1[286] ) );
  AND U797 ( .A(B[1]), .B(A[284]), .Z(\P1[285] ) );
  AND U798 ( .A(B[1]), .B(A[283]), .Z(\P1[284] ) );
  AND U799 ( .A(B[1]), .B(A[282]), .Z(\P1[283] ) );
  AND U800 ( .A(B[1]), .B(A[281]), .Z(\P1[282] ) );
  AND U801 ( .A(B[1]), .B(A[280]), .Z(\P1[281] ) );
  AND U802 ( .A(B[1]), .B(A[279]), .Z(\P1[280] ) );
  AND U803 ( .A(B[1]), .B(A[26]), .Z(\P1[27] ) );
  AND U804 ( .A(B[1]), .B(A[278]), .Z(\P1[279] ) );
  AND U805 ( .A(B[1]), .B(A[277]), .Z(\P1[278] ) );
  AND U806 ( .A(B[1]), .B(A[276]), .Z(\P1[277] ) );
  AND U807 ( .A(B[1]), .B(A[275]), .Z(\P1[276] ) );
  AND U808 ( .A(B[1]), .B(A[274]), .Z(\P1[275] ) );
  AND U809 ( .A(B[1]), .B(A[273]), .Z(\P1[274] ) );
  AND U810 ( .A(B[1]), .B(A[272]), .Z(\P1[273] ) );
  AND U811 ( .A(B[1]), .B(A[271]), .Z(\P1[272] ) );
  AND U812 ( .A(B[1]), .B(A[270]), .Z(\P1[271] ) );
  AND U813 ( .A(B[1]), .B(A[269]), .Z(\P1[270] ) );
  AND U814 ( .A(B[1]), .B(A[25]), .Z(\P1[26] ) );
  AND U815 ( .A(B[1]), .B(A[268]), .Z(\P1[269] ) );
  AND U816 ( .A(B[1]), .B(A[267]), .Z(\P1[268] ) );
  AND U817 ( .A(B[1]), .B(A[266]), .Z(\P1[267] ) );
  AND U818 ( .A(B[1]), .B(A[265]), .Z(\P1[266] ) );
  AND U819 ( .A(B[1]), .B(A[264]), .Z(\P1[265] ) );
  AND U820 ( .A(B[1]), .B(A[263]), .Z(\P1[264] ) );
  AND U821 ( .A(B[1]), .B(A[262]), .Z(\P1[263] ) );
  AND U822 ( .A(B[1]), .B(A[261]), .Z(\P1[262] ) );
  AND U823 ( .A(B[1]), .B(A[260]), .Z(\P1[261] ) );
  AND U824 ( .A(B[1]), .B(A[259]), .Z(\P1[260] ) );
  AND U825 ( .A(B[1]), .B(A[24]), .Z(\P1[25] ) );
  AND U826 ( .A(B[1]), .B(A[258]), .Z(\P1[259] ) );
  AND U827 ( .A(B[1]), .B(A[257]), .Z(\P1[258] ) );
  AND U828 ( .A(B[1]), .B(A[256]), .Z(\P1[257] ) );
  AND U829 ( .A(B[1]), .B(A[255]), .Z(\P1[256] ) );
  AND U830 ( .A(B[1]), .B(A[254]), .Z(\P1[255] ) );
  AND U831 ( .A(B[1]), .B(A[253]), .Z(\P1[254] ) );
  AND U832 ( .A(B[1]), .B(A[252]), .Z(\P1[253] ) );
  AND U833 ( .A(B[1]), .B(A[251]), .Z(\P1[252] ) );
  AND U834 ( .A(B[1]), .B(A[250]), .Z(\P1[251] ) );
  AND U835 ( .A(B[1]), .B(A[249]), .Z(\P1[250] ) );
  AND U836 ( .A(B[1]), .B(A[23]), .Z(\P1[24] ) );
  AND U837 ( .A(B[1]), .B(A[248]), .Z(\P1[249] ) );
  AND U838 ( .A(B[1]), .B(A[247]), .Z(\P1[248] ) );
  AND U839 ( .A(B[1]), .B(A[246]), .Z(\P1[247] ) );
  AND U840 ( .A(B[1]), .B(A[245]), .Z(\P1[246] ) );
  AND U841 ( .A(B[1]), .B(A[244]), .Z(\P1[245] ) );
  AND U842 ( .A(B[1]), .B(A[243]), .Z(\P1[244] ) );
  AND U843 ( .A(B[1]), .B(A[242]), .Z(\P1[243] ) );
  AND U844 ( .A(B[1]), .B(A[241]), .Z(\P1[242] ) );
  AND U845 ( .A(B[1]), .B(A[240]), .Z(\P1[241] ) );
  AND U846 ( .A(B[1]), .B(A[239]), .Z(\P1[240] ) );
  AND U847 ( .A(B[1]), .B(A[22]), .Z(\P1[23] ) );
  AND U848 ( .A(B[1]), .B(A[238]), .Z(\P1[239] ) );
  AND U849 ( .A(B[1]), .B(A[237]), .Z(\P1[238] ) );
  AND U850 ( .A(B[1]), .B(A[236]), .Z(\P1[237] ) );
  AND U851 ( .A(B[1]), .B(A[235]), .Z(\P1[236] ) );
  AND U852 ( .A(B[1]), .B(A[234]), .Z(\P1[235] ) );
  AND U853 ( .A(B[1]), .B(A[233]), .Z(\P1[234] ) );
  AND U854 ( .A(B[1]), .B(A[232]), .Z(\P1[233] ) );
  AND U855 ( .A(B[1]), .B(A[231]), .Z(\P1[232] ) );
  AND U856 ( .A(B[1]), .B(A[230]), .Z(\P1[231] ) );
  AND U857 ( .A(B[1]), .B(A[229]), .Z(\P1[230] ) );
  AND U858 ( .A(B[1]), .B(A[21]), .Z(\P1[22] ) );
  AND U859 ( .A(B[1]), .B(A[228]), .Z(\P1[229] ) );
  AND U860 ( .A(B[1]), .B(A[227]), .Z(\P1[228] ) );
  AND U861 ( .A(B[1]), .B(A[226]), .Z(\P1[227] ) );
  AND U862 ( .A(B[1]), .B(A[225]), .Z(\P1[226] ) );
  AND U863 ( .A(B[1]), .B(A[224]), .Z(\P1[225] ) );
  AND U864 ( .A(B[1]), .B(A[223]), .Z(\P1[224] ) );
  AND U865 ( .A(B[1]), .B(A[222]), .Z(\P1[223] ) );
  AND U866 ( .A(B[1]), .B(A[221]), .Z(\P1[222] ) );
  AND U867 ( .A(B[1]), .B(A[220]), .Z(\P1[221] ) );
  AND U868 ( .A(B[1]), .B(A[219]), .Z(\P1[220] ) );
  AND U869 ( .A(B[1]), .B(A[20]), .Z(\P1[21] ) );
  AND U870 ( .A(B[1]), .B(A[218]), .Z(\P1[219] ) );
  AND U871 ( .A(B[1]), .B(A[217]), .Z(\P1[218] ) );
  AND U872 ( .A(B[1]), .B(A[216]), .Z(\P1[217] ) );
  AND U873 ( .A(B[1]), .B(A[215]), .Z(\P1[216] ) );
  AND U874 ( .A(B[1]), .B(A[214]), .Z(\P1[215] ) );
  AND U875 ( .A(B[1]), .B(A[213]), .Z(\P1[214] ) );
  AND U876 ( .A(B[1]), .B(A[212]), .Z(\P1[213] ) );
  AND U877 ( .A(B[1]), .B(A[211]), .Z(\P1[212] ) );
  AND U878 ( .A(B[1]), .B(A[210]), .Z(\P1[211] ) );
  AND U879 ( .A(B[1]), .B(A[209]), .Z(\P1[210] ) );
  AND U880 ( .A(B[1]), .B(A[19]), .Z(\P1[20] ) );
  AND U881 ( .A(B[1]), .B(A[208]), .Z(\P1[209] ) );
  AND U882 ( .A(B[1]), .B(A[207]), .Z(\P1[208] ) );
  AND U883 ( .A(B[1]), .B(A[206]), .Z(\P1[207] ) );
  AND U884 ( .A(B[1]), .B(A[205]), .Z(\P1[206] ) );
  AND U885 ( .A(B[1]), .B(A[204]), .Z(\P1[205] ) );
  AND U886 ( .A(B[1]), .B(A[203]), .Z(\P1[204] ) );
  AND U887 ( .A(B[1]), .B(A[202]), .Z(\P1[203] ) );
  AND U888 ( .A(B[1]), .B(A[201]), .Z(\P1[202] ) );
  AND U889 ( .A(B[1]), .B(A[200]), .Z(\P1[201] ) );
  AND U890 ( .A(B[1]), .B(A[199]), .Z(\P1[200] ) );
  AND U891 ( .A(A[0]), .B(B[1]), .Z(\P1[1] ) );
  AND U892 ( .A(B[1]), .B(A[18]), .Z(\P1[19] ) );
  AND U893 ( .A(B[1]), .B(A[198]), .Z(\P1[199] ) );
  AND U894 ( .A(B[1]), .B(A[197]), .Z(\P1[198] ) );
  AND U895 ( .A(B[1]), .B(A[196]), .Z(\P1[197] ) );
  AND U896 ( .A(B[1]), .B(A[195]), .Z(\P1[196] ) );
  AND U897 ( .A(B[1]), .B(A[194]), .Z(\P1[195] ) );
  AND U898 ( .A(B[1]), .B(A[193]), .Z(\P1[194] ) );
  AND U899 ( .A(B[1]), .B(A[192]), .Z(\P1[193] ) );
  AND U900 ( .A(B[1]), .B(A[191]), .Z(\P1[192] ) );
  AND U901 ( .A(B[1]), .B(A[190]), .Z(\P1[191] ) );
  AND U902 ( .A(B[1]), .B(A[189]), .Z(\P1[190] ) );
  AND U903 ( .A(B[1]), .B(A[17]), .Z(\P1[18] ) );
  AND U904 ( .A(B[1]), .B(A[188]), .Z(\P1[189] ) );
  AND U905 ( .A(B[1]), .B(A[187]), .Z(\P1[188] ) );
  AND U906 ( .A(B[1]), .B(A[186]), .Z(\P1[187] ) );
  AND U907 ( .A(B[1]), .B(A[185]), .Z(\P1[186] ) );
  AND U908 ( .A(B[1]), .B(A[184]), .Z(\P1[185] ) );
  AND U909 ( .A(B[1]), .B(A[183]), .Z(\P1[184] ) );
  AND U910 ( .A(B[1]), .B(A[182]), .Z(\P1[183] ) );
  AND U911 ( .A(B[1]), .B(A[181]), .Z(\P1[182] ) );
  AND U912 ( .A(B[1]), .B(A[180]), .Z(\P1[181] ) );
  AND U913 ( .A(B[1]), .B(A[179]), .Z(\P1[180] ) );
  AND U914 ( .A(B[1]), .B(A[16]), .Z(\P1[17] ) );
  AND U915 ( .A(B[1]), .B(A[178]), .Z(\P1[179] ) );
  AND U916 ( .A(B[1]), .B(A[177]), .Z(\P1[178] ) );
  AND U917 ( .A(B[1]), .B(A[176]), .Z(\P1[177] ) );
  AND U918 ( .A(B[1]), .B(A[175]), .Z(\P1[176] ) );
  AND U919 ( .A(B[1]), .B(A[174]), .Z(\P1[175] ) );
  AND U920 ( .A(B[1]), .B(A[173]), .Z(\P1[174] ) );
  AND U921 ( .A(B[1]), .B(A[172]), .Z(\P1[173] ) );
  AND U922 ( .A(B[1]), .B(A[171]), .Z(\P1[172] ) );
  AND U923 ( .A(B[1]), .B(A[170]), .Z(\P1[171] ) );
  AND U924 ( .A(B[1]), .B(A[169]), .Z(\P1[170] ) );
  AND U925 ( .A(B[1]), .B(A[15]), .Z(\P1[16] ) );
  AND U926 ( .A(B[1]), .B(A[168]), .Z(\P1[169] ) );
  AND U927 ( .A(B[1]), .B(A[167]), .Z(\P1[168] ) );
  AND U928 ( .A(B[1]), .B(A[166]), .Z(\P1[167] ) );
  AND U929 ( .A(B[1]), .B(A[165]), .Z(\P1[166] ) );
  AND U930 ( .A(B[1]), .B(A[164]), .Z(\P1[165] ) );
  AND U931 ( .A(B[1]), .B(A[163]), .Z(\P1[164] ) );
  AND U932 ( .A(B[1]), .B(A[162]), .Z(\P1[163] ) );
  AND U933 ( .A(B[1]), .B(A[161]), .Z(\P1[162] ) );
  AND U934 ( .A(B[1]), .B(A[160]), .Z(\P1[161] ) );
  AND U935 ( .A(B[1]), .B(A[159]), .Z(\P1[160] ) );
  AND U936 ( .A(B[1]), .B(A[14]), .Z(\P1[15] ) );
  AND U937 ( .A(B[1]), .B(A[158]), .Z(\P1[159] ) );
  AND U938 ( .A(B[1]), .B(A[157]), .Z(\P1[158] ) );
  AND U939 ( .A(B[1]), .B(A[156]), .Z(\P1[157] ) );
  AND U940 ( .A(B[1]), .B(A[155]), .Z(\P1[156] ) );
  AND U941 ( .A(B[1]), .B(A[154]), .Z(\P1[155] ) );
  AND U942 ( .A(B[1]), .B(A[153]), .Z(\P1[154] ) );
  AND U943 ( .A(B[1]), .B(A[152]), .Z(\P1[153] ) );
  AND U944 ( .A(B[1]), .B(A[151]), .Z(\P1[152] ) );
  AND U945 ( .A(B[1]), .B(A[150]), .Z(\P1[151] ) );
  AND U946 ( .A(B[1]), .B(A[149]), .Z(\P1[150] ) );
  AND U947 ( .A(B[1]), .B(A[13]), .Z(\P1[14] ) );
  AND U948 ( .A(B[1]), .B(A[148]), .Z(\P1[149] ) );
  AND U949 ( .A(B[1]), .B(A[147]), .Z(\P1[148] ) );
  AND U950 ( .A(B[1]), .B(A[146]), .Z(\P1[147] ) );
  AND U951 ( .A(B[1]), .B(A[145]), .Z(\P1[146] ) );
  AND U952 ( .A(B[1]), .B(A[144]), .Z(\P1[145] ) );
  AND U953 ( .A(B[1]), .B(A[143]), .Z(\P1[144] ) );
  AND U954 ( .A(B[1]), .B(A[142]), .Z(\P1[143] ) );
  AND U955 ( .A(B[1]), .B(A[141]), .Z(\P1[142] ) );
  AND U956 ( .A(B[1]), .B(A[140]), .Z(\P1[141] ) );
  AND U957 ( .A(B[1]), .B(A[139]), .Z(\P1[140] ) );
  AND U958 ( .A(B[1]), .B(A[12]), .Z(\P1[13] ) );
  AND U959 ( .A(B[1]), .B(A[138]), .Z(\P1[139] ) );
  AND U960 ( .A(B[1]), .B(A[137]), .Z(\P1[138] ) );
  AND U961 ( .A(B[1]), .B(A[136]), .Z(\P1[137] ) );
  AND U962 ( .A(B[1]), .B(A[135]), .Z(\P1[136] ) );
  AND U963 ( .A(B[1]), .B(A[134]), .Z(\P1[135] ) );
  AND U964 ( .A(B[1]), .B(A[133]), .Z(\P1[134] ) );
  AND U965 ( .A(B[1]), .B(A[132]), .Z(\P1[133] ) );
  AND U966 ( .A(B[1]), .B(A[131]), .Z(\P1[132] ) );
  AND U967 ( .A(B[1]), .B(A[130]), .Z(\P1[131] ) );
  AND U968 ( .A(B[1]), .B(A[129]), .Z(\P1[130] ) );
  AND U969 ( .A(B[1]), .B(A[11]), .Z(\P1[12] ) );
  AND U970 ( .A(B[1]), .B(A[128]), .Z(\P1[129] ) );
  AND U971 ( .A(B[1]), .B(A[127]), .Z(\P1[128] ) );
  AND U972 ( .A(B[1]), .B(A[126]), .Z(\P1[127] ) );
  AND U973 ( .A(B[1]), .B(A[125]), .Z(\P1[126] ) );
  AND U974 ( .A(B[1]), .B(A[124]), .Z(\P1[125] ) );
  AND U975 ( .A(B[1]), .B(A[123]), .Z(\P1[124] ) );
  AND U976 ( .A(B[1]), .B(A[122]), .Z(\P1[123] ) );
  AND U977 ( .A(B[1]), .B(A[121]), .Z(\P1[122] ) );
  AND U978 ( .A(B[1]), .B(A[120]), .Z(\P1[121] ) );
  AND U979 ( .A(B[1]), .B(A[119]), .Z(\P1[120] ) );
  AND U980 ( .A(B[1]), .B(A[10]), .Z(\P1[11] ) );
  AND U981 ( .A(B[1]), .B(A[118]), .Z(\P1[119] ) );
  AND U982 ( .A(B[1]), .B(A[117]), .Z(\P1[118] ) );
  AND U983 ( .A(B[1]), .B(A[116]), .Z(\P1[117] ) );
  AND U984 ( .A(B[1]), .B(A[115]), .Z(\P1[116] ) );
  AND U985 ( .A(B[1]), .B(A[114]), .Z(\P1[115] ) );
  AND U986 ( .A(B[1]), .B(A[113]), .Z(\P1[114] ) );
  AND U987 ( .A(B[1]), .B(A[112]), .Z(\P1[113] ) );
  AND U988 ( .A(B[1]), .B(A[111]), .Z(\P1[112] ) );
  AND U989 ( .A(B[1]), .B(A[110]), .Z(\P1[111] ) );
  AND U990 ( .A(B[1]), .B(A[109]), .Z(\P1[110] ) );
  AND U991 ( .A(B[1]), .B(A[9]), .Z(\P1[10] ) );
  AND U992 ( .A(B[1]), .B(A[108]), .Z(\P1[109] ) );
  AND U993 ( .A(B[1]), .B(A[107]), .Z(\P1[108] ) );
  AND U994 ( .A(B[1]), .B(A[106]), .Z(\P1[107] ) );
  AND U995 ( .A(B[1]), .B(A[105]), .Z(\P1[106] ) );
  AND U996 ( .A(B[1]), .B(A[104]), .Z(\P1[105] ) );
  AND U997 ( .A(B[1]), .B(A[103]), .Z(\P1[104] ) );
  AND U998 ( .A(B[1]), .B(A[102]), .Z(\P1[103] ) );
  AND U999 ( .A(B[1]), .B(A[101]), .Z(\P1[102] ) );
  AND U1000 ( .A(B[1]), .B(A[1023]), .Z(\P1[1024] ) );
  AND U1001 ( .A(B[1]), .B(A[1022]), .Z(\P1[1023] ) );
  AND U1002 ( .A(B[1]), .B(A[1021]), .Z(\P1[1022] ) );
  AND U1003 ( .A(B[1]), .B(A[1020]), .Z(\P1[1021] ) );
  AND U1004 ( .A(B[1]), .B(A[1019]), .Z(\P1[1020] ) );
  AND U1005 ( .A(B[1]), .B(A[100]), .Z(\P1[101] ) );
  AND U1006 ( .A(B[1]), .B(A[1018]), .Z(\P1[1019] ) );
  AND U1007 ( .A(B[1]), .B(A[1017]), .Z(\P1[1018] ) );
  AND U1008 ( .A(B[1]), .B(A[1016]), .Z(\P1[1017] ) );
  AND U1009 ( .A(B[1]), .B(A[1015]), .Z(\P1[1016] ) );
  AND U1010 ( .A(B[1]), .B(A[1014]), .Z(\P1[1015] ) );
  AND U1011 ( .A(B[1]), .B(A[1013]), .Z(\P1[1014] ) );
  AND U1012 ( .A(B[1]), .B(A[1012]), .Z(\P1[1013] ) );
  AND U1013 ( .A(B[1]), .B(A[1011]), .Z(\P1[1012] ) );
  AND U1014 ( .A(B[1]), .B(A[1010]), .Z(\P1[1011] ) );
  AND U1015 ( .A(B[1]), .B(A[1009]), .Z(\P1[1010] ) );
  AND U1016 ( .A(B[1]), .B(A[99]), .Z(\P1[100] ) );
  AND U1017 ( .A(B[1]), .B(A[1008]), .Z(\P1[1009] ) );
  AND U1018 ( .A(B[1]), .B(A[1007]), .Z(\P1[1008] ) );
  AND U1019 ( .A(B[1]), .B(A[1006]), .Z(\P1[1007] ) );
  AND U1020 ( .A(B[1]), .B(A[1005]), .Z(\P1[1006] ) );
  AND U1021 ( .A(B[1]), .B(A[1004]), .Z(\P1[1005] ) );
  AND U1022 ( .A(B[1]), .B(A[1003]), .Z(\P1[1004] ) );
  AND U1023 ( .A(B[1]), .B(A[1002]), .Z(\P1[1003] ) );
  AND U1024 ( .A(B[1]), .B(A[1001]), .Z(\P1[1002] ) );
  AND U1025 ( .A(B[1]), .B(A[1000]), .Z(\P1[1001] ) );
  AND U1026 ( .A(B[1]), .B(A[999]), .Z(\P1[1000] ) );
  AND U1027 ( .A(A[9]), .B(B[0]), .Z(\P0[9] ) );
  AND U1028 ( .A(A[99]), .B(B[0]), .Z(\P0[99] ) );
  AND U1029 ( .A(A[999]), .B(B[0]), .Z(\P0[999] ) );
  AND U1030 ( .A(A[998]), .B(B[0]), .Z(\P0[998] ) );
  AND U1031 ( .A(A[997]), .B(B[0]), .Z(\P0[997] ) );
  AND U1032 ( .A(A[996]), .B(B[0]), .Z(\P0[996] ) );
  AND U1033 ( .A(A[995]), .B(B[0]), .Z(\P0[995] ) );
  AND U1034 ( .A(A[994]), .B(B[0]), .Z(\P0[994] ) );
  AND U1035 ( .A(A[993]), .B(B[0]), .Z(\P0[993] ) );
  AND U1036 ( .A(A[992]), .B(B[0]), .Z(\P0[992] ) );
  AND U1037 ( .A(A[991]), .B(B[0]), .Z(\P0[991] ) );
  AND U1038 ( .A(A[990]), .B(B[0]), .Z(\P0[990] ) );
  AND U1039 ( .A(A[98]), .B(B[0]), .Z(\P0[98] ) );
  AND U1040 ( .A(A[989]), .B(B[0]), .Z(\P0[989] ) );
  AND U1041 ( .A(A[988]), .B(B[0]), .Z(\P0[988] ) );
  AND U1042 ( .A(A[987]), .B(B[0]), .Z(\P0[987] ) );
  AND U1043 ( .A(A[986]), .B(B[0]), .Z(\P0[986] ) );
  AND U1044 ( .A(A[985]), .B(B[0]), .Z(\P0[985] ) );
  AND U1045 ( .A(A[984]), .B(B[0]), .Z(\P0[984] ) );
  AND U1046 ( .A(A[983]), .B(B[0]), .Z(\P0[983] ) );
  AND U1047 ( .A(A[982]), .B(B[0]), .Z(\P0[982] ) );
  AND U1048 ( .A(A[981]), .B(B[0]), .Z(\P0[981] ) );
  AND U1049 ( .A(A[980]), .B(B[0]), .Z(\P0[980] ) );
  AND U1050 ( .A(A[97]), .B(B[0]), .Z(\P0[97] ) );
  AND U1051 ( .A(A[979]), .B(B[0]), .Z(\P0[979] ) );
  AND U1052 ( .A(A[978]), .B(B[0]), .Z(\P0[978] ) );
  AND U1053 ( .A(A[977]), .B(B[0]), .Z(\P0[977] ) );
  AND U1054 ( .A(A[976]), .B(B[0]), .Z(\P0[976] ) );
  AND U1055 ( .A(A[975]), .B(B[0]), .Z(\P0[975] ) );
  AND U1056 ( .A(A[974]), .B(B[0]), .Z(\P0[974] ) );
  AND U1057 ( .A(A[973]), .B(B[0]), .Z(\P0[973] ) );
  AND U1058 ( .A(A[972]), .B(B[0]), .Z(\P0[972] ) );
  AND U1059 ( .A(A[971]), .B(B[0]), .Z(\P0[971] ) );
  AND U1060 ( .A(A[970]), .B(B[0]), .Z(\P0[970] ) );
  AND U1061 ( .A(A[96]), .B(B[0]), .Z(\P0[96] ) );
  AND U1062 ( .A(A[969]), .B(B[0]), .Z(\P0[969] ) );
  AND U1063 ( .A(A[968]), .B(B[0]), .Z(\P0[968] ) );
  AND U1064 ( .A(A[967]), .B(B[0]), .Z(\P0[967] ) );
  AND U1065 ( .A(A[966]), .B(B[0]), .Z(\P0[966] ) );
  AND U1066 ( .A(A[965]), .B(B[0]), .Z(\P0[965] ) );
  AND U1067 ( .A(A[964]), .B(B[0]), .Z(\P0[964] ) );
  AND U1068 ( .A(A[963]), .B(B[0]), .Z(\P0[963] ) );
  AND U1069 ( .A(A[962]), .B(B[0]), .Z(\P0[962] ) );
  AND U1070 ( .A(A[961]), .B(B[0]), .Z(\P0[961] ) );
  AND U1071 ( .A(A[960]), .B(B[0]), .Z(\P0[960] ) );
  AND U1072 ( .A(A[95]), .B(B[0]), .Z(\P0[95] ) );
  AND U1073 ( .A(A[959]), .B(B[0]), .Z(\P0[959] ) );
  AND U1074 ( .A(A[958]), .B(B[0]), .Z(\P0[958] ) );
  AND U1075 ( .A(A[957]), .B(B[0]), .Z(\P0[957] ) );
  AND U1076 ( .A(A[956]), .B(B[0]), .Z(\P0[956] ) );
  AND U1077 ( .A(A[955]), .B(B[0]), .Z(\P0[955] ) );
  AND U1078 ( .A(A[954]), .B(B[0]), .Z(\P0[954] ) );
  AND U1079 ( .A(A[953]), .B(B[0]), .Z(\P0[953] ) );
  AND U1080 ( .A(A[952]), .B(B[0]), .Z(\P0[952] ) );
  AND U1081 ( .A(A[951]), .B(B[0]), .Z(\P0[951] ) );
  AND U1082 ( .A(A[950]), .B(B[0]), .Z(\P0[950] ) );
  AND U1083 ( .A(A[94]), .B(B[0]), .Z(\P0[94] ) );
  AND U1084 ( .A(A[949]), .B(B[0]), .Z(\P0[949] ) );
  AND U1085 ( .A(A[948]), .B(B[0]), .Z(\P0[948] ) );
  AND U1086 ( .A(A[947]), .B(B[0]), .Z(\P0[947] ) );
  AND U1087 ( .A(A[946]), .B(B[0]), .Z(\P0[946] ) );
  AND U1088 ( .A(A[945]), .B(B[0]), .Z(\P0[945] ) );
  AND U1089 ( .A(A[944]), .B(B[0]), .Z(\P0[944] ) );
  AND U1090 ( .A(A[943]), .B(B[0]), .Z(\P0[943] ) );
  AND U1091 ( .A(A[942]), .B(B[0]), .Z(\P0[942] ) );
  AND U1092 ( .A(A[941]), .B(B[0]), .Z(\P0[941] ) );
  AND U1093 ( .A(A[940]), .B(B[0]), .Z(\P0[940] ) );
  AND U1094 ( .A(A[93]), .B(B[0]), .Z(\P0[93] ) );
  AND U1095 ( .A(A[939]), .B(B[0]), .Z(\P0[939] ) );
  AND U1096 ( .A(A[938]), .B(B[0]), .Z(\P0[938] ) );
  AND U1097 ( .A(A[937]), .B(B[0]), .Z(\P0[937] ) );
  AND U1098 ( .A(A[936]), .B(B[0]), .Z(\P0[936] ) );
  AND U1099 ( .A(A[935]), .B(B[0]), .Z(\P0[935] ) );
  AND U1100 ( .A(A[934]), .B(B[0]), .Z(\P0[934] ) );
  AND U1101 ( .A(A[933]), .B(B[0]), .Z(\P0[933] ) );
  AND U1102 ( .A(A[932]), .B(B[0]), .Z(\P0[932] ) );
  AND U1103 ( .A(A[931]), .B(B[0]), .Z(\P0[931] ) );
  AND U1104 ( .A(A[930]), .B(B[0]), .Z(\P0[930] ) );
  AND U1105 ( .A(A[92]), .B(B[0]), .Z(\P0[92] ) );
  AND U1106 ( .A(A[929]), .B(B[0]), .Z(\P0[929] ) );
  AND U1107 ( .A(A[928]), .B(B[0]), .Z(\P0[928] ) );
  AND U1108 ( .A(A[927]), .B(B[0]), .Z(\P0[927] ) );
  AND U1109 ( .A(A[926]), .B(B[0]), .Z(\P0[926] ) );
  AND U1110 ( .A(A[925]), .B(B[0]), .Z(\P0[925] ) );
  AND U1111 ( .A(A[924]), .B(B[0]), .Z(\P0[924] ) );
  AND U1112 ( .A(A[923]), .B(B[0]), .Z(\P0[923] ) );
  AND U1113 ( .A(A[922]), .B(B[0]), .Z(\P0[922] ) );
  AND U1114 ( .A(A[921]), .B(B[0]), .Z(\P0[921] ) );
  AND U1115 ( .A(A[920]), .B(B[0]), .Z(\P0[920] ) );
  AND U1116 ( .A(A[91]), .B(B[0]), .Z(\P0[91] ) );
  AND U1117 ( .A(A[919]), .B(B[0]), .Z(\P0[919] ) );
  AND U1118 ( .A(A[918]), .B(B[0]), .Z(\P0[918] ) );
  AND U1119 ( .A(A[917]), .B(B[0]), .Z(\P0[917] ) );
  AND U1120 ( .A(A[916]), .B(B[0]), .Z(\P0[916] ) );
  AND U1121 ( .A(A[915]), .B(B[0]), .Z(\P0[915] ) );
  AND U1122 ( .A(A[914]), .B(B[0]), .Z(\P0[914] ) );
  AND U1123 ( .A(A[913]), .B(B[0]), .Z(\P0[913] ) );
  AND U1124 ( .A(A[912]), .B(B[0]), .Z(\P0[912] ) );
  AND U1125 ( .A(A[911]), .B(B[0]), .Z(\P0[911] ) );
  AND U1126 ( .A(A[910]), .B(B[0]), .Z(\P0[910] ) );
  AND U1127 ( .A(A[90]), .B(B[0]), .Z(\P0[90] ) );
  AND U1128 ( .A(A[909]), .B(B[0]), .Z(\P0[909] ) );
  AND U1129 ( .A(A[908]), .B(B[0]), .Z(\P0[908] ) );
  AND U1130 ( .A(A[907]), .B(B[0]), .Z(\P0[907] ) );
  AND U1131 ( .A(A[906]), .B(B[0]), .Z(\P0[906] ) );
  AND U1132 ( .A(A[905]), .B(B[0]), .Z(\P0[905] ) );
  AND U1133 ( .A(A[904]), .B(B[0]), .Z(\P0[904] ) );
  AND U1134 ( .A(A[903]), .B(B[0]), .Z(\P0[903] ) );
  AND U1135 ( .A(A[902]), .B(B[0]), .Z(\P0[902] ) );
  AND U1136 ( .A(A[901]), .B(B[0]), .Z(\P0[901] ) );
  AND U1137 ( .A(A[900]), .B(B[0]), .Z(\P0[900] ) );
  AND U1138 ( .A(B[0]), .B(A[8]), .Z(\P0[8] ) );
  AND U1139 ( .A(A[89]), .B(B[0]), .Z(\P0[89] ) );
  AND U1140 ( .A(A[899]), .B(B[0]), .Z(\P0[899] ) );
  AND U1141 ( .A(A[898]), .B(B[0]), .Z(\P0[898] ) );
  AND U1142 ( .A(A[897]), .B(B[0]), .Z(\P0[897] ) );
  AND U1143 ( .A(A[896]), .B(B[0]), .Z(\P0[896] ) );
  AND U1144 ( .A(A[895]), .B(B[0]), .Z(\P0[895] ) );
  AND U1145 ( .A(A[894]), .B(B[0]), .Z(\P0[894] ) );
  AND U1146 ( .A(A[893]), .B(B[0]), .Z(\P0[893] ) );
  AND U1147 ( .A(A[892]), .B(B[0]), .Z(\P0[892] ) );
  AND U1148 ( .A(A[891]), .B(B[0]), .Z(\P0[891] ) );
  AND U1149 ( .A(A[890]), .B(B[0]), .Z(\P0[890] ) );
  AND U1150 ( .A(A[88]), .B(B[0]), .Z(\P0[88] ) );
  AND U1151 ( .A(A[889]), .B(B[0]), .Z(\P0[889] ) );
  AND U1152 ( .A(A[888]), .B(B[0]), .Z(\P0[888] ) );
  AND U1153 ( .A(A[887]), .B(B[0]), .Z(\P0[887] ) );
  AND U1154 ( .A(A[886]), .B(B[0]), .Z(\P0[886] ) );
  AND U1155 ( .A(A[885]), .B(B[0]), .Z(\P0[885] ) );
  AND U1156 ( .A(A[884]), .B(B[0]), .Z(\P0[884] ) );
  AND U1157 ( .A(A[883]), .B(B[0]), .Z(\P0[883] ) );
  AND U1158 ( .A(A[882]), .B(B[0]), .Z(\P0[882] ) );
  AND U1159 ( .A(A[881]), .B(B[0]), .Z(\P0[881] ) );
  AND U1160 ( .A(A[880]), .B(B[0]), .Z(\P0[880] ) );
  AND U1161 ( .A(A[87]), .B(B[0]), .Z(\P0[87] ) );
  AND U1162 ( .A(A[879]), .B(B[0]), .Z(\P0[879] ) );
  AND U1163 ( .A(A[878]), .B(B[0]), .Z(\P0[878] ) );
  AND U1164 ( .A(A[877]), .B(B[0]), .Z(\P0[877] ) );
  AND U1165 ( .A(A[876]), .B(B[0]), .Z(\P0[876] ) );
  AND U1166 ( .A(A[875]), .B(B[0]), .Z(\P0[875] ) );
  AND U1167 ( .A(A[874]), .B(B[0]), .Z(\P0[874] ) );
  AND U1168 ( .A(A[873]), .B(B[0]), .Z(\P0[873] ) );
  AND U1169 ( .A(A[872]), .B(B[0]), .Z(\P0[872] ) );
  AND U1170 ( .A(A[871]), .B(B[0]), .Z(\P0[871] ) );
  AND U1171 ( .A(A[870]), .B(B[0]), .Z(\P0[870] ) );
  AND U1172 ( .A(A[86]), .B(B[0]), .Z(\P0[86] ) );
  AND U1173 ( .A(A[869]), .B(B[0]), .Z(\P0[869] ) );
  AND U1174 ( .A(A[868]), .B(B[0]), .Z(\P0[868] ) );
  AND U1175 ( .A(A[867]), .B(B[0]), .Z(\P0[867] ) );
  AND U1176 ( .A(A[866]), .B(B[0]), .Z(\P0[866] ) );
  AND U1177 ( .A(A[865]), .B(B[0]), .Z(\P0[865] ) );
  AND U1178 ( .A(A[864]), .B(B[0]), .Z(\P0[864] ) );
  AND U1179 ( .A(A[863]), .B(B[0]), .Z(\P0[863] ) );
  AND U1180 ( .A(A[862]), .B(B[0]), .Z(\P0[862] ) );
  AND U1181 ( .A(A[861]), .B(B[0]), .Z(\P0[861] ) );
  AND U1182 ( .A(A[860]), .B(B[0]), .Z(\P0[860] ) );
  AND U1183 ( .A(A[85]), .B(B[0]), .Z(\P0[85] ) );
  AND U1184 ( .A(A[859]), .B(B[0]), .Z(\P0[859] ) );
  AND U1185 ( .A(A[858]), .B(B[0]), .Z(\P0[858] ) );
  AND U1186 ( .A(A[857]), .B(B[0]), .Z(\P0[857] ) );
  AND U1187 ( .A(A[856]), .B(B[0]), .Z(\P0[856] ) );
  AND U1188 ( .A(A[855]), .B(B[0]), .Z(\P0[855] ) );
  AND U1189 ( .A(A[854]), .B(B[0]), .Z(\P0[854] ) );
  AND U1190 ( .A(A[853]), .B(B[0]), .Z(\P0[853] ) );
  AND U1191 ( .A(A[852]), .B(B[0]), .Z(\P0[852] ) );
  AND U1192 ( .A(A[851]), .B(B[0]), .Z(\P0[851] ) );
  AND U1193 ( .A(A[850]), .B(B[0]), .Z(\P0[850] ) );
  AND U1194 ( .A(A[84]), .B(B[0]), .Z(\P0[84] ) );
  AND U1195 ( .A(A[849]), .B(B[0]), .Z(\P0[849] ) );
  AND U1196 ( .A(A[848]), .B(B[0]), .Z(\P0[848] ) );
  AND U1197 ( .A(A[847]), .B(B[0]), .Z(\P0[847] ) );
  AND U1198 ( .A(A[846]), .B(B[0]), .Z(\P0[846] ) );
  AND U1199 ( .A(A[845]), .B(B[0]), .Z(\P0[845] ) );
  AND U1200 ( .A(A[844]), .B(B[0]), .Z(\P0[844] ) );
  AND U1201 ( .A(A[843]), .B(B[0]), .Z(\P0[843] ) );
  AND U1202 ( .A(A[842]), .B(B[0]), .Z(\P0[842] ) );
  AND U1203 ( .A(A[841]), .B(B[0]), .Z(\P0[841] ) );
  AND U1204 ( .A(A[840]), .B(B[0]), .Z(\P0[840] ) );
  AND U1205 ( .A(A[83]), .B(B[0]), .Z(\P0[83] ) );
  AND U1206 ( .A(A[839]), .B(B[0]), .Z(\P0[839] ) );
  AND U1207 ( .A(A[838]), .B(B[0]), .Z(\P0[838] ) );
  AND U1208 ( .A(A[837]), .B(B[0]), .Z(\P0[837] ) );
  AND U1209 ( .A(A[836]), .B(B[0]), .Z(\P0[836] ) );
  AND U1210 ( .A(A[835]), .B(B[0]), .Z(\P0[835] ) );
  AND U1211 ( .A(A[834]), .B(B[0]), .Z(\P0[834] ) );
  AND U1212 ( .A(A[833]), .B(B[0]), .Z(\P0[833] ) );
  AND U1213 ( .A(A[832]), .B(B[0]), .Z(\P0[832] ) );
  AND U1214 ( .A(A[831]), .B(B[0]), .Z(\P0[831] ) );
  AND U1215 ( .A(A[830]), .B(B[0]), .Z(\P0[830] ) );
  AND U1216 ( .A(A[82]), .B(B[0]), .Z(\P0[82] ) );
  AND U1217 ( .A(A[829]), .B(B[0]), .Z(\P0[829] ) );
  AND U1218 ( .A(A[828]), .B(B[0]), .Z(\P0[828] ) );
  AND U1219 ( .A(A[827]), .B(B[0]), .Z(\P0[827] ) );
  AND U1220 ( .A(A[826]), .B(B[0]), .Z(\P0[826] ) );
  AND U1221 ( .A(A[825]), .B(B[0]), .Z(\P0[825] ) );
  AND U1222 ( .A(A[824]), .B(B[0]), .Z(\P0[824] ) );
  AND U1223 ( .A(A[823]), .B(B[0]), .Z(\P0[823] ) );
  AND U1224 ( .A(A[822]), .B(B[0]), .Z(\P0[822] ) );
  AND U1225 ( .A(A[821]), .B(B[0]), .Z(\P0[821] ) );
  AND U1226 ( .A(A[820]), .B(B[0]), .Z(\P0[820] ) );
  AND U1227 ( .A(A[81]), .B(B[0]), .Z(\P0[81] ) );
  AND U1228 ( .A(A[819]), .B(B[0]), .Z(\P0[819] ) );
  AND U1229 ( .A(A[818]), .B(B[0]), .Z(\P0[818] ) );
  AND U1230 ( .A(A[817]), .B(B[0]), .Z(\P0[817] ) );
  AND U1231 ( .A(A[816]), .B(B[0]), .Z(\P0[816] ) );
  AND U1232 ( .A(A[815]), .B(B[0]), .Z(\P0[815] ) );
  AND U1233 ( .A(A[814]), .B(B[0]), .Z(\P0[814] ) );
  AND U1234 ( .A(A[813]), .B(B[0]), .Z(\P0[813] ) );
  AND U1235 ( .A(A[812]), .B(B[0]), .Z(\P0[812] ) );
  AND U1236 ( .A(A[811]), .B(B[0]), .Z(\P0[811] ) );
  AND U1237 ( .A(A[810]), .B(B[0]), .Z(\P0[810] ) );
  AND U1238 ( .A(A[80]), .B(B[0]), .Z(\P0[80] ) );
  AND U1239 ( .A(A[809]), .B(B[0]), .Z(\P0[809] ) );
  AND U1240 ( .A(A[808]), .B(B[0]), .Z(\P0[808] ) );
  AND U1241 ( .A(A[807]), .B(B[0]), .Z(\P0[807] ) );
  AND U1242 ( .A(A[806]), .B(B[0]), .Z(\P0[806] ) );
  AND U1243 ( .A(A[805]), .B(B[0]), .Z(\P0[805] ) );
  AND U1244 ( .A(A[804]), .B(B[0]), .Z(\P0[804] ) );
  AND U1245 ( .A(A[803]), .B(B[0]), .Z(\P0[803] ) );
  AND U1246 ( .A(A[802]), .B(B[0]), .Z(\P0[802] ) );
  AND U1247 ( .A(A[801]), .B(B[0]), .Z(\P0[801] ) );
  AND U1248 ( .A(A[800]), .B(B[0]), .Z(\P0[800] ) );
  AND U1249 ( .A(A[7]), .B(B[0]), .Z(\P0[7] ) );
  AND U1250 ( .A(A[79]), .B(B[0]), .Z(\P0[79] ) );
  AND U1251 ( .A(A[799]), .B(B[0]), .Z(\P0[799] ) );
  AND U1252 ( .A(A[798]), .B(B[0]), .Z(\P0[798] ) );
  AND U1253 ( .A(A[797]), .B(B[0]), .Z(\P0[797] ) );
  AND U1254 ( .A(A[796]), .B(B[0]), .Z(\P0[796] ) );
  AND U1255 ( .A(A[795]), .B(B[0]), .Z(\P0[795] ) );
  AND U1256 ( .A(A[794]), .B(B[0]), .Z(\P0[794] ) );
  AND U1257 ( .A(A[793]), .B(B[0]), .Z(\P0[793] ) );
  AND U1258 ( .A(A[792]), .B(B[0]), .Z(\P0[792] ) );
  AND U1259 ( .A(A[791]), .B(B[0]), .Z(\P0[791] ) );
  AND U1260 ( .A(A[790]), .B(B[0]), .Z(\P0[790] ) );
  AND U1261 ( .A(A[78]), .B(B[0]), .Z(\P0[78] ) );
  AND U1262 ( .A(A[789]), .B(B[0]), .Z(\P0[789] ) );
  AND U1263 ( .A(A[788]), .B(B[0]), .Z(\P0[788] ) );
  AND U1264 ( .A(A[787]), .B(B[0]), .Z(\P0[787] ) );
  AND U1265 ( .A(A[786]), .B(B[0]), .Z(\P0[786] ) );
  AND U1266 ( .A(A[785]), .B(B[0]), .Z(\P0[785] ) );
  AND U1267 ( .A(A[784]), .B(B[0]), .Z(\P0[784] ) );
  AND U1268 ( .A(A[783]), .B(B[0]), .Z(\P0[783] ) );
  AND U1269 ( .A(A[782]), .B(B[0]), .Z(\P0[782] ) );
  AND U1270 ( .A(A[781]), .B(B[0]), .Z(\P0[781] ) );
  AND U1271 ( .A(A[780]), .B(B[0]), .Z(\P0[780] ) );
  AND U1272 ( .A(A[77]), .B(B[0]), .Z(\P0[77] ) );
  AND U1273 ( .A(A[779]), .B(B[0]), .Z(\P0[779] ) );
  AND U1274 ( .A(A[778]), .B(B[0]), .Z(\P0[778] ) );
  AND U1275 ( .A(A[777]), .B(B[0]), .Z(\P0[777] ) );
  AND U1276 ( .A(A[776]), .B(B[0]), .Z(\P0[776] ) );
  AND U1277 ( .A(A[775]), .B(B[0]), .Z(\P0[775] ) );
  AND U1278 ( .A(A[774]), .B(B[0]), .Z(\P0[774] ) );
  AND U1279 ( .A(A[773]), .B(B[0]), .Z(\P0[773] ) );
  AND U1280 ( .A(A[772]), .B(B[0]), .Z(\P0[772] ) );
  AND U1281 ( .A(A[771]), .B(B[0]), .Z(\P0[771] ) );
  AND U1282 ( .A(A[770]), .B(B[0]), .Z(\P0[770] ) );
  AND U1283 ( .A(A[76]), .B(B[0]), .Z(\P0[76] ) );
  AND U1284 ( .A(A[769]), .B(B[0]), .Z(\P0[769] ) );
  AND U1285 ( .A(A[768]), .B(B[0]), .Z(\P0[768] ) );
  AND U1286 ( .A(A[767]), .B(B[0]), .Z(\P0[767] ) );
  AND U1287 ( .A(A[766]), .B(B[0]), .Z(\P0[766] ) );
  AND U1288 ( .A(A[765]), .B(B[0]), .Z(\P0[765] ) );
  AND U1289 ( .A(A[764]), .B(B[0]), .Z(\P0[764] ) );
  AND U1290 ( .A(A[763]), .B(B[0]), .Z(\P0[763] ) );
  AND U1291 ( .A(A[762]), .B(B[0]), .Z(\P0[762] ) );
  AND U1292 ( .A(A[761]), .B(B[0]), .Z(\P0[761] ) );
  AND U1293 ( .A(A[760]), .B(B[0]), .Z(\P0[760] ) );
  AND U1294 ( .A(A[75]), .B(B[0]), .Z(\P0[75] ) );
  AND U1295 ( .A(A[759]), .B(B[0]), .Z(\P0[759] ) );
  AND U1296 ( .A(A[758]), .B(B[0]), .Z(\P0[758] ) );
  AND U1297 ( .A(A[757]), .B(B[0]), .Z(\P0[757] ) );
  AND U1298 ( .A(A[756]), .B(B[0]), .Z(\P0[756] ) );
  AND U1299 ( .A(A[755]), .B(B[0]), .Z(\P0[755] ) );
  AND U1300 ( .A(A[754]), .B(B[0]), .Z(\P0[754] ) );
  AND U1301 ( .A(A[753]), .B(B[0]), .Z(\P0[753] ) );
  AND U1302 ( .A(A[752]), .B(B[0]), .Z(\P0[752] ) );
  AND U1303 ( .A(A[751]), .B(B[0]), .Z(\P0[751] ) );
  AND U1304 ( .A(A[750]), .B(B[0]), .Z(\P0[750] ) );
  AND U1305 ( .A(A[74]), .B(B[0]), .Z(\P0[74] ) );
  AND U1306 ( .A(A[749]), .B(B[0]), .Z(\P0[749] ) );
  AND U1307 ( .A(A[748]), .B(B[0]), .Z(\P0[748] ) );
  AND U1308 ( .A(A[747]), .B(B[0]), .Z(\P0[747] ) );
  AND U1309 ( .A(A[746]), .B(B[0]), .Z(\P0[746] ) );
  AND U1310 ( .A(A[745]), .B(B[0]), .Z(\P0[745] ) );
  AND U1311 ( .A(A[744]), .B(B[0]), .Z(\P0[744] ) );
  AND U1312 ( .A(A[743]), .B(B[0]), .Z(\P0[743] ) );
  AND U1313 ( .A(A[742]), .B(B[0]), .Z(\P0[742] ) );
  AND U1314 ( .A(A[741]), .B(B[0]), .Z(\P0[741] ) );
  AND U1315 ( .A(A[740]), .B(B[0]), .Z(\P0[740] ) );
  AND U1316 ( .A(A[73]), .B(B[0]), .Z(\P0[73] ) );
  AND U1317 ( .A(A[739]), .B(B[0]), .Z(\P0[739] ) );
  AND U1318 ( .A(A[738]), .B(B[0]), .Z(\P0[738] ) );
  AND U1319 ( .A(A[737]), .B(B[0]), .Z(\P0[737] ) );
  AND U1320 ( .A(A[736]), .B(B[0]), .Z(\P0[736] ) );
  AND U1321 ( .A(A[735]), .B(B[0]), .Z(\P0[735] ) );
  AND U1322 ( .A(A[734]), .B(B[0]), .Z(\P0[734] ) );
  AND U1323 ( .A(A[733]), .B(B[0]), .Z(\P0[733] ) );
  AND U1324 ( .A(A[732]), .B(B[0]), .Z(\P0[732] ) );
  AND U1325 ( .A(A[731]), .B(B[0]), .Z(\P0[731] ) );
  AND U1326 ( .A(A[730]), .B(B[0]), .Z(\P0[730] ) );
  AND U1327 ( .A(A[72]), .B(B[0]), .Z(\P0[72] ) );
  AND U1328 ( .A(A[729]), .B(B[0]), .Z(\P0[729] ) );
  AND U1329 ( .A(A[728]), .B(B[0]), .Z(\P0[728] ) );
  AND U1330 ( .A(A[727]), .B(B[0]), .Z(\P0[727] ) );
  AND U1331 ( .A(A[726]), .B(B[0]), .Z(\P0[726] ) );
  AND U1332 ( .A(A[725]), .B(B[0]), .Z(\P0[725] ) );
  AND U1333 ( .A(A[724]), .B(B[0]), .Z(\P0[724] ) );
  AND U1334 ( .A(A[723]), .B(B[0]), .Z(\P0[723] ) );
  AND U1335 ( .A(A[722]), .B(B[0]), .Z(\P0[722] ) );
  AND U1336 ( .A(A[721]), .B(B[0]), .Z(\P0[721] ) );
  AND U1337 ( .A(A[720]), .B(B[0]), .Z(\P0[720] ) );
  AND U1338 ( .A(A[71]), .B(B[0]), .Z(\P0[71] ) );
  AND U1339 ( .A(A[719]), .B(B[0]), .Z(\P0[719] ) );
  AND U1340 ( .A(A[718]), .B(B[0]), .Z(\P0[718] ) );
  AND U1341 ( .A(A[717]), .B(B[0]), .Z(\P0[717] ) );
  AND U1342 ( .A(A[716]), .B(B[0]), .Z(\P0[716] ) );
  AND U1343 ( .A(A[715]), .B(B[0]), .Z(\P0[715] ) );
  AND U1344 ( .A(A[714]), .B(B[0]), .Z(\P0[714] ) );
  AND U1345 ( .A(A[713]), .B(B[0]), .Z(\P0[713] ) );
  AND U1346 ( .A(A[712]), .B(B[0]), .Z(\P0[712] ) );
  AND U1347 ( .A(A[711]), .B(B[0]), .Z(\P0[711] ) );
  AND U1348 ( .A(A[710]), .B(B[0]), .Z(\P0[710] ) );
  AND U1349 ( .A(A[70]), .B(B[0]), .Z(\P0[70] ) );
  AND U1350 ( .A(A[709]), .B(B[0]), .Z(\P0[709] ) );
  AND U1351 ( .A(A[708]), .B(B[0]), .Z(\P0[708] ) );
  AND U1352 ( .A(A[707]), .B(B[0]), .Z(\P0[707] ) );
  AND U1353 ( .A(A[706]), .B(B[0]), .Z(\P0[706] ) );
  AND U1354 ( .A(A[705]), .B(B[0]), .Z(\P0[705] ) );
  AND U1355 ( .A(A[704]), .B(B[0]), .Z(\P0[704] ) );
  AND U1356 ( .A(A[703]), .B(B[0]), .Z(\P0[703] ) );
  AND U1357 ( .A(A[702]), .B(B[0]), .Z(\P0[702] ) );
  AND U1358 ( .A(A[701]), .B(B[0]), .Z(\P0[701] ) );
  AND U1359 ( .A(A[700]), .B(B[0]), .Z(\P0[700] ) );
  AND U1360 ( .A(A[6]), .B(B[0]), .Z(\P0[6] ) );
  AND U1361 ( .A(A[69]), .B(B[0]), .Z(\P0[69] ) );
  AND U1362 ( .A(A[699]), .B(B[0]), .Z(\P0[699] ) );
  AND U1363 ( .A(A[698]), .B(B[0]), .Z(\P0[698] ) );
  AND U1364 ( .A(A[697]), .B(B[0]), .Z(\P0[697] ) );
  AND U1365 ( .A(A[696]), .B(B[0]), .Z(\P0[696] ) );
  AND U1366 ( .A(A[695]), .B(B[0]), .Z(\P0[695] ) );
  AND U1367 ( .A(A[694]), .B(B[0]), .Z(\P0[694] ) );
  AND U1368 ( .A(A[693]), .B(B[0]), .Z(\P0[693] ) );
  AND U1369 ( .A(A[692]), .B(B[0]), .Z(\P0[692] ) );
  AND U1370 ( .A(A[691]), .B(B[0]), .Z(\P0[691] ) );
  AND U1371 ( .A(A[690]), .B(B[0]), .Z(\P0[690] ) );
  AND U1372 ( .A(A[68]), .B(B[0]), .Z(\P0[68] ) );
  AND U1373 ( .A(A[689]), .B(B[0]), .Z(\P0[689] ) );
  AND U1374 ( .A(A[688]), .B(B[0]), .Z(\P0[688] ) );
  AND U1375 ( .A(A[687]), .B(B[0]), .Z(\P0[687] ) );
  AND U1376 ( .A(A[686]), .B(B[0]), .Z(\P0[686] ) );
  AND U1377 ( .A(A[685]), .B(B[0]), .Z(\P0[685] ) );
  AND U1378 ( .A(A[684]), .B(B[0]), .Z(\P0[684] ) );
  AND U1379 ( .A(A[683]), .B(B[0]), .Z(\P0[683] ) );
  AND U1380 ( .A(A[682]), .B(B[0]), .Z(\P0[682] ) );
  AND U1381 ( .A(A[681]), .B(B[0]), .Z(\P0[681] ) );
  AND U1382 ( .A(A[680]), .B(B[0]), .Z(\P0[680] ) );
  AND U1383 ( .A(A[67]), .B(B[0]), .Z(\P0[67] ) );
  AND U1384 ( .A(A[679]), .B(B[0]), .Z(\P0[679] ) );
  AND U1385 ( .A(A[678]), .B(B[0]), .Z(\P0[678] ) );
  AND U1386 ( .A(A[677]), .B(B[0]), .Z(\P0[677] ) );
  AND U1387 ( .A(A[676]), .B(B[0]), .Z(\P0[676] ) );
  AND U1388 ( .A(A[675]), .B(B[0]), .Z(\P0[675] ) );
  AND U1389 ( .A(A[674]), .B(B[0]), .Z(\P0[674] ) );
  AND U1390 ( .A(A[673]), .B(B[0]), .Z(\P0[673] ) );
  AND U1391 ( .A(A[672]), .B(B[0]), .Z(\P0[672] ) );
  AND U1392 ( .A(A[671]), .B(B[0]), .Z(\P0[671] ) );
  AND U1393 ( .A(A[670]), .B(B[0]), .Z(\P0[670] ) );
  AND U1394 ( .A(A[66]), .B(B[0]), .Z(\P0[66] ) );
  AND U1395 ( .A(A[669]), .B(B[0]), .Z(\P0[669] ) );
  AND U1396 ( .A(A[668]), .B(B[0]), .Z(\P0[668] ) );
  AND U1397 ( .A(A[667]), .B(B[0]), .Z(\P0[667] ) );
  AND U1398 ( .A(A[666]), .B(B[0]), .Z(\P0[666] ) );
  AND U1399 ( .A(A[665]), .B(B[0]), .Z(\P0[665] ) );
  AND U1400 ( .A(A[664]), .B(B[0]), .Z(\P0[664] ) );
  AND U1401 ( .A(A[663]), .B(B[0]), .Z(\P0[663] ) );
  AND U1402 ( .A(A[662]), .B(B[0]), .Z(\P0[662] ) );
  AND U1403 ( .A(A[661]), .B(B[0]), .Z(\P0[661] ) );
  AND U1404 ( .A(A[660]), .B(B[0]), .Z(\P0[660] ) );
  AND U1405 ( .A(A[65]), .B(B[0]), .Z(\P0[65] ) );
  AND U1406 ( .A(A[659]), .B(B[0]), .Z(\P0[659] ) );
  AND U1407 ( .A(A[658]), .B(B[0]), .Z(\P0[658] ) );
  AND U1408 ( .A(A[657]), .B(B[0]), .Z(\P0[657] ) );
  AND U1409 ( .A(A[656]), .B(B[0]), .Z(\P0[656] ) );
  AND U1410 ( .A(A[655]), .B(B[0]), .Z(\P0[655] ) );
  AND U1411 ( .A(A[654]), .B(B[0]), .Z(\P0[654] ) );
  AND U1412 ( .A(A[653]), .B(B[0]), .Z(\P0[653] ) );
  AND U1413 ( .A(A[652]), .B(B[0]), .Z(\P0[652] ) );
  AND U1414 ( .A(A[651]), .B(B[0]), .Z(\P0[651] ) );
  AND U1415 ( .A(A[650]), .B(B[0]), .Z(\P0[650] ) );
  AND U1416 ( .A(A[64]), .B(B[0]), .Z(\P0[64] ) );
  AND U1417 ( .A(A[649]), .B(B[0]), .Z(\P0[649] ) );
  AND U1418 ( .A(A[648]), .B(B[0]), .Z(\P0[648] ) );
  AND U1419 ( .A(A[647]), .B(B[0]), .Z(\P0[647] ) );
  AND U1420 ( .A(A[646]), .B(B[0]), .Z(\P0[646] ) );
  AND U1421 ( .A(A[645]), .B(B[0]), .Z(\P0[645] ) );
  AND U1422 ( .A(A[644]), .B(B[0]), .Z(\P0[644] ) );
  AND U1423 ( .A(A[643]), .B(B[0]), .Z(\P0[643] ) );
  AND U1424 ( .A(A[642]), .B(B[0]), .Z(\P0[642] ) );
  AND U1425 ( .A(A[641]), .B(B[0]), .Z(\P0[641] ) );
  AND U1426 ( .A(A[640]), .B(B[0]), .Z(\P0[640] ) );
  AND U1427 ( .A(A[63]), .B(B[0]), .Z(\P0[63] ) );
  AND U1428 ( .A(A[639]), .B(B[0]), .Z(\P0[639] ) );
  AND U1429 ( .A(A[638]), .B(B[0]), .Z(\P0[638] ) );
  AND U1430 ( .A(A[637]), .B(B[0]), .Z(\P0[637] ) );
  AND U1431 ( .A(A[636]), .B(B[0]), .Z(\P0[636] ) );
  AND U1432 ( .A(A[635]), .B(B[0]), .Z(\P0[635] ) );
  AND U1433 ( .A(A[634]), .B(B[0]), .Z(\P0[634] ) );
  AND U1434 ( .A(A[633]), .B(B[0]), .Z(\P0[633] ) );
  AND U1435 ( .A(A[632]), .B(B[0]), .Z(\P0[632] ) );
  AND U1436 ( .A(A[631]), .B(B[0]), .Z(\P0[631] ) );
  AND U1437 ( .A(A[630]), .B(B[0]), .Z(\P0[630] ) );
  AND U1438 ( .A(A[62]), .B(B[0]), .Z(\P0[62] ) );
  AND U1439 ( .A(A[629]), .B(B[0]), .Z(\P0[629] ) );
  AND U1440 ( .A(A[628]), .B(B[0]), .Z(\P0[628] ) );
  AND U1441 ( .A(A[627]), .B(B[0]), .Z(\P0[627] ) );
  AND U1442 ( .A(A[626]), .B(B[0]), .Z(\P0[626] ) );
  AND U1443 ( .A(A[625]), .B(B[0]), .Z(\P0[625] ) );
  AND U1444 ( .A(A[624]), .B(B[0]), .Z(\P0[624] ) );
  AND U1445 ( .A(A[623]), .B(B[0]), .Z(\P0[623] ) );
  AND U1446 ( .A(A[622]), .B(B[0]), .Z(\P0[622] ) );
  AND U1447 ( .A(A[621]), .B(B[0]), .Z(\P0[621] ) );
  AND U1448 ( .A(A[620]), .B(B[0]), .Z(\P0[620] ) );
  AND U1449 ( .A(A[61]), .B(B[0]), .Z(\P0[61] ) );
  AND U1450 ( .A(A[619]), .B(B[0]), .Z(\P0[619] ) );
  AND U1451 ( .A(A[618]), .B(B[0]), .Z(\P0[618] ) );
  AND U1452 ( .A(A[617]), .B(B[0]), .Z(\P0[617] ) );
  AND U1453 ( .A(A[616]), .B(B[0]), .Z(\P0[616] ) );
  AND U1454 ( .A(A[615]), .B(B[0]), .Z(\P0[615] ) );
  AND U1455 ( .A(A[614]), .B(B[0]), .Z(\P0[614] ) );
  AND U1456 ( .A(A[613]), .B(B[0]), .Z(\P0[613] ) );
  AND U1457 ( .A(A[612]), .B(B[0]), .Z(\P0[612] ) );
  AND U1458 ( .A(A[611]), .B(B[0]), .Z(\P0[611] ) );
  AND U1459 ( .A(A[610]), .B(B[0]), .Z(\P0[610] ) );
  AND U1460 ( .A(A[60]), .B(B[0]), .Z(\P0[60] ) );
  AND U1461 ( .A(A[609]), .B(B[0]), .Z(\P0[609] ) );
  AND U1462 ( .A(A[608]), .B(B[0]), .Z(\P0[608] ) );
  AND U1463 ( .A(A[607]), .B(B[0]), .Z(\P0[607] ) );
  AND U1464 ( .A(A[606]), .B(B[0]), .Z(\P0[606] ) );
  AND U1465 ( .A(A[605]), .B(B[0]), .Z(\P0[605] ) );
  AND U1466 ( .A(A[604]), .B(B[0]), .Z(\P0[604] ) );
  AND U1467 ( .A(A[603]), .B(B[0]), .Z(\P0[603] ) );
  AND U1468 ( .A(A[602]), .B(B[0]), .Z(\P0[602] ) );
  AND U1469 ( .A(A[601]), .B(B[0]), .Z(\P0[601] ) );
  AND U1470 ( .A(A[600]), .B(B[0]), .Z(\P0[600] ) );
  AND U1471 ( .A(A[5]), .B(B[0]), .Z(\P0[5] ) );
  AND U1472 ( .A(A[59]), .B(B[0]), .Z(\P0[59] ) );
  AND U1473 ( .A(A[599]), .B(B[0]), .Z(\P0[599] ) );
  AND U1474 ( .A(A[598]), .B(B[0]), .Z(\P0[598] ) );
  AND U1475 ( .A(A[597]), .B(B[0]), .Z(\P0[597] ) );
  AND U1476 ( .A(A[596]), .B(B[0]), .Z(\P0[596] ) );
  AND U1477 ( .A(A[595]), .B(B[0]), .Z(\P0[595] ) );
  AND U1478 ( .A(A[594]), .B(B[0]), .Z(\P0[594] ) );
  AND U1479 ( .A(A[593]), .B(B[0]), .Z(\P0[593] ) );
  AND U1480 ( .A(A[592]), .B(B[0]), .Z(\P0[592] ) );
  AND U1481 ( .A(A[591]), .B(B[0]), .Z(\P0[591] ) );
  AND U1482 ( .A(A[590]), .B(B[0]), .Z(\P0[590] ) );
  AND U1483 ( .A(A[58]), .B(B[0]), .Z(\P0[58] ) );
  AND U1484 ( .A(A[589]), .B(B[0]), .Z(\P0[589] ) );
  AND U1485 ( .A(A[588]), .B(B[0]), .Z(\P0[588] ) );
  AND U1486 ( .A(A[587]), .B(B[0]), .Z(\P0[587] ) );
  AND U1487 ( .A(A[586]), .B(B[0]), .Z(\P0[586] ) );
  AND U1488 ( .A(A[585]), .B(B[0]), .Z(\P0[585] ) );
  AND U1489 ( .A(A[584]), .B(B[0]), .Z(\P0[584] ) );
  AND U1490 ( .A(A[583]), .B(B[0]), .Z(\P0[583] ) );
  AND U1491 ( .A(A[582]), .B(B[0]), .Z(\P0[582] ) );
  AND U1492 ( .A(A[581]), .B(B[0]), .Z(\P0[581] ) );
  AND U1493 ( .A(A[580]), .B(B[0]), .Z(\P0[580] ) );
  AND U1494 ( .A(A[57]), .B(B[0]), .Z(\P0[57] ) );
  AND U1495 ( .A(A[579]), .B(B[0]), .Z(\P0[579] ) );
  AND U1496 ( .A(A[578]), .B(B[0]), .Z(\P0[578] ) );
  AND U1497 ( .A(A[577]), .B(B[0]), .Z(\P0[577] ) );
  AND U1498 ( .A(A[576]), .B(B[0]), .Z(\P0[576] ) );
  AND U1499 ( .A(A[575]), .B(B[0]), .Z(\P0[575] ) );
  AND U1500 ( .A(A[574]), .B(B[0]), .Z(\P0[574] ) );
  AND U1501 ( .A(A[573]), .B(B[0]), .Z(\P0[573] ) );
  AND U1502 ( .A(A[572]), .B(B[0]), .Z(\P0[572] ) );
  AND U1503 ( .A(A[571]), .B(B[0]), .Z(\P0[571] ) );
  AND U1504 ( .A(A[570]), .B(B[0]), .Z(\P0[570] ) );
  AND U1505 ( .A(A[56]), .B(B[0]), .Z(\P0[56] ) );
  AND U1506 ( .A(A[569]), .B(B[0]), .Z(\P0[569] ) );
  AND U1507 ( .A(A[568]), .B(B[0]), .Z(\P0[568] ) );
  AND U1508 ( .A(A[567]), .B(B[0]), .Z(\P0[567] ) );
  AND U1509 ( .A(A[566]), .B(B[0]), .Z(\P0[566] ) );
  AND U1510 ( .A(A[565]), .B(B[0]), .Z(\P0[565] ) );
  AND U1511 ( .A(A[564]), .B(B[0]), .Z(\P0[564] ) );
  AND U1512 ( .A(A[563]), .B(B[0]), .Z(\P0[563] ) );
  AND U1513 ( .A(A[562]), .B(B[0]), .Z(\P0[562] ) );
  AND U1514 ( .A(A[561]), .B(B[0]), .Z(\P0[561] ) );
  AND U1515 ( .A(A[560]), .B(B[0]), .Z(\P0[560] ) );
  AND U1516 ( .A(A[55]), .B(B[0]), .Z(\P0[55] ) );
  AND U1517 ( .A(A[559]), .B(B[0]), .Z(\P0[559] ) );
  AND U1518 ( .A(A[558]), .B(B[0]), .Z(\P0[558] ) );
  AND U1519 ( .A(A[557]), .B(B[0]), .Z(\P0[557] ) );
  AND U1520 ( .A(A[556]), .B(B[0]), .Z(\P0[556] ) );
  AND U1521 ( .A(A[555]), .B(B[0]), .Z(\P0[555] ) );
  AND U1522 ( .A(A[554]), .B(B[0]), .Z(\P0[554] ) );
  AND U1523 ( .A(A[553]), .B(B[0]), .Z(\P0[553] ) );
  AND U1524 ( .A(A[552]), .B(B[0]), .Z(\P0[552] ) );
  AND U1525 ( .A(A[551]), .B(B[0]), .Z(\P0[551] ) );
  AND U1526 ( .A(A[550]), .B(B[0]), .Z(\P0[550] ) );
  AND U1527 ( .A(A[54]), .B(B[0]), .Z(\P0[54] ) );
  AND U1528 ( .A(A[549]), .B(B[0]), .Z(\P0[549] ) );
  AND U1529 ( .A(A[548]), .B(B[0]), .Z(\P0[548] ) );
  AND U1530 ( .A(A[547]), .B(B[0]), .Z(\P0[547] ) );
  AND U1531 ( .A(A[546]), .B(B[0]), .Z(\P0[546] ) );
  AND U1532 ( .A(A[545]), .B(B[0]), .Z(\P0[545] ) );
  AND U1533 ( .A(A[544]), .B(B[0]), .Z(\P0[544] ) );
  AND U1534 ( .A(A[543]), .B(B[0]), .Z(\P0[543] ) );
  AND U1535 ( .A(A[542]), .B(B[0]), .Z(\P0[542] ) );
  AND U1536 ( .A(A[541]), .B(B[0]), .Z(\P0[541] ) );
  AND U1537 ( .A(A[540]), .B(B[0]), .Z(\P0[540] ) );
  AND U1538 ( .A(A[53]), .B(B[0]), .Z(\P0[53] ) );
  AND U1539 ( .A(A[539]), .B(B[0]), .Z(\P0[539] ) );
  AND U1540 ( .A(A[538]), .B(B[0]), .Z(\P0[538] ) );
  AND U1541 ( .A(A[537]), .B(B[0]), .Z(\P0[537] ) );
  AND U1542 ( .A(A[536]), .B(B[0]), .Z(\P0[536] ) );
  AND U1543 ( .A(A[535]), .B(B[0]), .Z(\P0[535] ) );
  AND U1544 ( .A(A[534]), .B(B[0]), .Z(\P0[534] ) );
  AND U1545 ( .A(A[533]), .B(B[0]), .Z(\P0[533] ) );
  AND U1546 ( .A(A[532]), .B(B[0]), .Z(\P0[532] ) );
  AND U1547 ( .A(A[531]), .B(B[0]), .Z(\P0[531] ) );
  AND U1548 ( .A(A[530]), .B(B[0]), .Z(\P0[530] ) );
  AND U1549 ( .A(A[52]), .B(B[0]), .Z(\P0[52] ) );
  AND U1550 ( .A(A[529]), .B(B[0]), .Z(\P0[529] ) );
  AND U1551 ( .A(A[528]), .B(B[0]), .Z(\P0[528] ) );
  AND U1552 ( .A(A[527]), .B(B[0]), .Z(\P0[527] ) );
  AND U1553 ( .A(A[526]), .B(B[0]), .Z(\P0[526] ) );
  AND U1554 ( .A(A[525]), .B(B[0]), .Z(\P0[525] ) );
  AND U1555 ( .A(A[524]), .B(B[0]), .Z(\P0[524] ) );
  AND U1556 ( .A(A[523]), .B(B[0]), .Z(\P0[523] ) );
  AND U1557 ( .A(A[522]), .B(B[0]), .Z(\P0[522] ) );
  AND U1558 ( .A(A[521]), .B(B[0]), .Z(\P0[521] ) );
  AND U1559 ( .A(A[520]), .B(B[0]), .Z(\P0[520] ) );
  AND U1560 ( .A(A[51]), .B(B[0]), .Z(\P0[51] ) );
  AND U1561 ( .A(A[519]), .B(B[0]), .Z(\P0[519] ) );
  AND U1562 ( .A(A[518]), .B(B[0]), .Z(\P0[518] ) );
  AND U1563 ( .A(A[517]), .B(B[0]), .Z(\P0[517] ) );
  AND U1564 ( .A(A[516]), .B(B[0]), .Z(\P0[516] ) );
  AND U1565 ( .A(A[515]), .B(B[0]), .Z(\P0[515] ) );
  AND U1566 ( .A(A[514]), .B(B[0]), .Z(\P0[514] ) );
  AND U1567 ( .A(A[513]), .B(B[0]), .Z(\P0[513] ) );
  AND U1568 ( .A(A[512]), .B(B[0]), .Z(\P0[512] ) );
  AND U1569 ( .A(A[511]), .B(B[0]), .Z(\P0[511] ) );
  AND U1570 ( .A(A[510]), .B(B[0]), .Z(\P0[510] ) );
  AND U1571 ( .A(A[50]), .B(B[0]), .Z(\P0[50] ) );
  AND U1572 ( .A(A[509]), .B(B[0]), .Z(\P0[509] ) );
  AND U1573 ( .A(A[508]), .B(B[0]), .Z(\P0[508] ) );
  AND U1574 ( .A(A[507]), .B(B[0]), .Z(\P0[507] ) );
  AND U1575 ( .A(A[506]), .B(B[0]), .Z(\P0[506] ) );
  AND U1576 ( .A(A[505]), .B(B[0]), .Z(\P0[505] ) );
  AND U1577 ( .A(A[504]), .B(B[0]), .Z(\P0[504] ) );
  AND U1578 ( .A(A[503]), .B(B[0]), .Z(\P0[503] ) );
  AND U1579 ( .A(A[502]), .B(B[0]), .Z(\P0[502] ) );
  AND U1580 ( .A(A[501]), .B(B[0]), .Z(\P0[501] ) );
  AND U1581 ( .A(A[500]), .B(B[0]), .Z(\P0[500] ) );
  AND U1582 ( .A(A[4]), .B(B[0]), .Z(\P0[4] ) );
  AND U1583 ( .A(A[49]), .B(B[0]), .Z(\P0[49] ) );
  AND U1584 ( .A(A[499]), .B(B[0]), .Z(\P0[499] ) );
  AND U1585 ( .A(A[498]), .B(B[0]), .Z(\P0[498] ) );
  AND U1586 ( .A(A[497]), .B(B[0]), .Z(\P0[497] ) );
  AND U1587 ( .A(A[496]), .B(B[0]), .Z(\P0[496] ) );
  AND U1588 ( .A(A[495]), .B(B[0]), .Z(\P0[495] ) );
  AND U1589 ( .A(A[494]), .B(B[0]), .Z(\P0[494] ) );
  AND U1590 ( .A(A[493]), .B(B[0]), .Z(\P0[493] ) );
  AND U1591 ( .A(A[492]), .B(B[0]), .Z(\P0[492] ) );
  AND U1592 ( .A(A[491]), .B(B[0]), .Z(\P0[491] ) );
  AND U1593 ( .A(A[490]), .B(B[0]), .Z(\P0[490] ) );
  AND U1594 ( .A(A[48]), .B(B[0]), .Z(\P0[48] ) );
  AND U1595 ( .A(A[489]), .B(B[0]), .Z(\P0[489] ) );
  AND U1596 ( .A(A[488]), .B(B[0]), .Z(\P0[488] ) );
  AND U1597 ( .A(A[487]), .B(B[0]), .Z(\P0[487] ) );
  AND U1598 ( .A(A[486]), .B(B[0]), .Z(\P0[486] ) );
  AND U1599 ( .A(A[485]), .B(B[0]), .Z(\P0[485] ) );
  AND U1600 ( .A(A[484]), .B(B[0]), .Z(\P0[484] ) );
  AND U1601 ( .A(A[483]), .B(B[0]), .Z(\P0[483] ) );
  AND U1602 ( .A(A[482]), .B(B[0]), .Z(\P0[482] ) );
  AND U1603 ( .A(A[481]), .B(B[0]), .Z(\P0[481] ) );
  AND U1604 ( .A(A[480]), .B(B[0]), .Z(\P0[480] ) );
  AND U1605 ( .A(A[47]), .B(B[0]), .Z(\P0[47] ) );
  AND U1606 ( .A(A[479]), .B(B[0]), .Z(\P0[479] ) );
  AND U1607 ( .A(A[478]), .B(B[0]), .Z(\P0[478] ) );
  AND U1608 ( .A(A[477]), .B(B[0]), .Z(\P0[477] ) );
  AND U1609 ( .A(A[476]), .B(B[0]), .Z(\P0[476] ) );
  AND U1610 ( .A(A[475]), .B(B[0]), .Z(\P0[475] ) );
  AND U1611 ( .A(A[474]), .B(B[0]), .Z(\P0[474] ) );
  AND U1612 ( .A(A[473]), .B(B[0]), .Z(\P0[473] ) );
  AND U1613 ( .A(A[472]), .B(B[0]), .Z(\P0[472] ) );
  AND U1614 ( .A(A[471]), .B(B[0]), .Z(\P0[471] ) );
  AND U1615 ( .A(A[470]), .B(B[0]), .Z(\P0[470] ) );
  AND U1616 ( .A(A[46]), .B(B[0]), .Z(\P0[46] ) );
  AND U1617 ( .A(A[469]), .B(B[0]), .Z(\P0[469] ) );
  AND U1618 ( .A(A[468]), .B(B[0]), .Z(\P0[468] ) );
  AND U1619 ( .A(A[467]), .B(B[0]), .Z(\P0[467] ) );
  AND U1620 ( .A(A[466]), .B(B[0]), .Z(\P0[466] ) );
  AND U1621 ( .A(A[465]), .B(B[0]), .Z(\P0[465] ) );
  AND U1622 ( .A(A[464]), .B(B[0]), .Z(\P0[464] ) );
  AND U1623 ( .A(A[463]), .B(B[0]), .Z(\P0[463] ) );
  AND U1624 ( .A(A[462]), .B(B[0]), .Z(\P0[462] ) );
  AND U1625 ( .A(A[461]), .B(B[0]), .Z(\P0[461] ) );
  AND U1626 ( .A(A[460]), .B(B[0]), .Z(\P0[460] ) );
  AND U1627 ( .A(A[45]), .B(B[0]), .Z(\P0[45] ) );
  AND U1628 ( .A(A[459]), .B(B[0]), .Z(\P0[459] ) );
  AND U1629 ( .A(A[458]), .B(B[0]), .Z(\P0[458] ) );
  AND U1630 ( .A(A[457]), .B(B[0]), .Z(\P0[457] ) );
  AND U1631 ( .A(A[456]), .B(B[0]), .Z(\P0[456] ) );
  AND U1632 ( .A(A[455]), .B(B[0]), .Z(\P0[455] ) );
  AND U1633 ( .A(A[454]), .B(B[0]), .Z(\P0[454] ) );
  AND U1634 ( .A(A[453]), .B(B[0]), .Z(\P0[453] ) );
  AND U1635 ( .A(A[452]), .B(B[0]), .Z(\P0[452] ) );
  AND U1636 ( .A(A[451]), .B(B[0]), .Z(\P0[451] ) );
  AND U1637 ( .A(A[450]), .B(B[0]), .Z(\P0[450] ) );
  AND U1638 ( .A(A[44]), .B(B[0]), .Z(\P0[44] ) );
  AND U1639 ( .A(A[449]), .B(B[0]), .Z(\P0[449] ) );
  AND U1640 ( .A(A[448]), .B(B[0]), .Z(\P0[448] ) );
  AND U1641 ( .A(A[447]), .B(B[0]), .Z(\P0[447] ) );
  AND U1642 ( .A(A[446]), .B(B[0]), .Z(\P0[446] ) );
  AND U1643 ( .A(A[445]), .B(B[0]), .Z(\P0[445] ) );
  AND U1644 ( .A(A[444]), .B(B[0]), .Z(\P0[444] ) );
  AND U1645 ( .A(A[443]), .B(B[0]), .Z(\P0[443] ) );
  AND U1646 ( .A(A[442]), .B(B[0]), .Z(\P0[442] ) );
  AND U1647 ( .A(A[441]), .B(B[0]), .Z(\P0[441] ) );
  AND U1648 ( .A(A[440]), .B(B[0]), .Z(\P0[440] ) );
  AND U1649 ( .A(A[43]), .B(B[0]), .Z(\P0[43] ) );
  AND U1650 ( .A(A[439]), .B(B[0]), .Z(\P0[439] ) );
  AND U1651 ( .A(A[438]), .B(B[0]), .Z(\P0[438] ) );
  AND U1652 ( .A(A[437]), .B(B[0]), .Z(\P0[437] ) );
  AND U1653 ( .A(A[436]), .B(B[0]), .Z(\P0[436] ) );
  AND U1654 ( .A(A[435]), .B(B[0]), .Z(\P0[435] ) );
  AND U1655 ( .A(A[434]), .B(B[0]), .Z(\P0[434] ) );
  AND U1656 ( .A(A[433]), .B(B[0]), .Z(\P0[433] ) );
  AND U1657 ( .A(A[432]), .B(B[0]), .Z(\P0[432] ) );
  AND U1658 ( .A(A[431]), .B(B[0]), .Z(\P0[431] ) );
  AND U1659 ( .A(A[430]), .B(B[0]), .Z(\P0[430] ) );
  AND U1660 ( .A(A[42]), .B(B[0]), .Z(\P0[42] ) );
  AND U1661 ( .A(A[429]), .B(B[0]), .Z(\P0[429] ) );
  AND U1662 ( .A(A[428]), .B(B[0]), .Z(\P0[428] ) );
  AND U1663 ( .A(A[427]), .B(B[0]), .Z(\P0[427] ) );
  AND U1664 ( .A(A[426]), .B(B[0]), .Z(\P0[426] ) );
  AND U1665 ( .A(A[425]), .B(B[0]), .Z(\P0[425] ) );
  AND U1666 ( .A(A[424]), .B(B[0]), .Z(\P0[424] ) );
  AND U1667 ( .A(A[423]), .B(B[0]), .Z(\P0[423] ) );
  AND U1668 ( .A(A[422]), .B(B[0]), .Z(\P0[422] ) );
  AND U1669 ( .A(A[421]), .B(B[0]), .Z(\P0[421] ) );
  AND U1670 ( .A(A[420]), .B(B[0]), .Z(\P0[420] ) );
  AND U1671 ( .A(A[41]), .B(B[0]), .Z(\P0[41] ) );
  AND U1672 ( .A(A[419]), .B(B[0]), .Z(\P0[419] ) );
  AND U1673 ( .A(A[418]), .B(B[0]), .Z(\P0[418] ) );
  AND U1674 ( .A(A[417]), .B(B[0]), .Z(\P0[417] ) );
  AND U1675 ( .A(A[416]), .B(B[0]), .Z(\P0[416] ) );
  AND U1676 ( .A(A[415]), .B(B[0]), .Z(\P0[415] ) );
  AND U1677 ( .A(A[414]), .B(B[0]), .Z(\P0[414] ) );
  AND U1678 ( .A(A[413]), .B(B[0]), .Z(\P0[413] ) );
  AND U1679 ( .A(A[412]), .B(B[0]), .Z(\P0[412] ) );
  AND U1680 ( .A(A[411]), .B(B[0]), .Z(\P0[411] ) );
  AND U1681 ( .A(A[410]), .B(B[0]), .Z(\P0[410] ) );
  AND U1682 ( .A(A[40]), .B(B[0]), .Z(\P0[40] ) );
  AND U1683 ( .A(A[409]), .B(B[0]), .Z(\P0[409] ) );
  AND U1684 ( .A(A[408]), .B(B[0]), .Z(\P0[408] ) );
  AND U1685 ( .A(A[407]), .B(B[0]), .Z(\P0[407] ) );
  AND U1686 ( .A(A[406]), .B(B[0]), .Z(\P0[406] ) );
  AND U1687 ( .A(A[405]), .B(B[0]), .Z(\P0[405] ) );
  AND U1688 ( .A(A[404]), .B(B[0]), .Z(\P0[404] ) );
  AND U1689 ( .A(A[403]), .B(B[0]), .Z(\P0[403] ) );
  AND U1690 ( .A(A[402]), .B(B[0]), .Z(\P0[402] ) );
  AND U1691 ( .A(A[401]), .B(B[0]), .Z(\P0[401] ) );
  AND U1692 ( .A(A[400]), .B(B[0]), .Z(\P0[400] ) );
  AND U1693 ( .A(A[3]), .B(B[0]), .Z(\P0[3] ) );
  AND U1694 ( .A(A[39]), .B(B[0]), .Z(\P0[39] ) );
  AND U1695 ( .A(A[399]), .B(B[0]), .Z(\P0[399] ) );
  AND U1696 ( .A(A[398]), .B(B[0]), .Z(\P0[398] ) );
  AND U1697 ( .A(A[397]), .B(B[0]), .Z(\P0[397] ) );
  AND U1698 ( .A(A[396]), .B(B[0]), .Z(\P0[396] ) );
  AND U1699 ( .A(A[395]), .B(B[0]), .Z(\P0[395] ) );
  AND U1700 ( .A(A[394]), .B(B[0]), .Z(\P0[394] ) );
  AND U1701 ( .A(A[393]), .B(B[0]), .Z(\P0[393] ) );
  AND U1702 ( .A(A[392]), .B(B[0]), .Z(\P0[392] ) );
  AND U1703 ( .A(A[391]), .B(B[0]), .Z(\P0[391] ) );
  AND U1704 ( .A(A[390]), .B(B[0]), .Z(\P0[390] ) );
  AND U1705 ( .A(A[38]), .B(B[0]), .Z(\P0[38] ) );
  AND U1706 ( .A(A[389]), .B(B[0]), .Z(\P0[389] ) );
  AND U1707 ( .A(A[388]), .B(B[0]), .Z(\P0[388] ) );
  AND U1708 ( .A(A[387]), .B(B[0]), .Z(\P0[387] ) );
  AND U1709 ( .A(A[386]), .B(B[0]), .Z(\P0[386] ) );
  AND U1710 ( .A(A[385]), .B(B[0]), .Z(\P0[385] ) );
  AND U1711 ( .A(A[384]), .B(B[0]), .Z(\P0[384] ) );
  AND U1712 ( .A(A[383]), .B(B[0]), .Z(\P0[383] ) );
  AND U1713 ( .A(A[382]), .B(B[0]), .Z(\P0[382] ) );
  AND U1714 ( .A(A[381]), .B(B[0]), .Z(\P0[381] ) );
  AND U1715 ( .A(A[380]), .B(B[0]), .Z(\P0[380] ) );
  AND U1716 ( .A(A[37]), .B(B[0]), .Z(\P0[37] ) );
  AND U1717 ( .A(A[379]), .B(B[0]), .Z(\P0[379] ) );
  AND U1718 ( .A(A[378]), .B(B[0]), .Z(\P0[378] ) );
  AND U1719 ( .A(A[377]), .B(B[0]), .Z(\P0[377] ) );
  AND U1720 ( .A(A[376]), .B(B[0]), .Z(\P0[376] ) );
  AND U1721 ( .A(A[375]), .B(B[0]), .Z(\P0[375] ) );
  AND U1722 ( .A(A[374]), .B(B[0]), .Z(\P0[374] ) );
  AND U1723 ( .A(A[373]), .B(B[0]), .Z(\P0[373] ) );
  AND U1724 ( .A(A[372]), .B(B[0]), .Z(\P0[372] ) );
  AND U1725 ( .A(A[371]), .B(B[0]), .Z(\P0[371] ) );
  AND U1726 ( .A(A[370]), .B(B[0]), .Z(\P0[370] ) );
  AND U1727 ( .A(A[36]), .B(B[0]), .Z(\P0[36] ) );
  AND U1728 ( .A(A[369]), .B(B[0]), .Z(\P0[369] ) );
  AND U1729 ( .A(A[368]), .B(B[0]), .Z(\P0[368] ) );
  AND U1730 ( .A(A[367]), .B(B[0]), .Z(\P0[367] ) );
  AND U1731 ( .A(A[366]), .B(B[0]), .Z(\P0[366] ) );
  AND U1732 ( .A(A[365]), .B(B[0]), .Z(\P0[365] ) );
  AND U1733 ( .A(A[364]), .B(B[0]), .Z(\P0[364] ) );
  AND U1734 ( .A(A[363]), .B(B[0]), .Z(\P0[363] ) );
  AND U1735 ( .A(A[362]), .B(B[0]), .Z(\P0[362] ) );
  AND U1736 ( .A(A[361]), .B(B[0]), .Z(\P0[361] ) );
  AND U1737 ( .A(A[360]), .B(B[0]), .Z(\P0[360] ) );
  AND U1738 ( .A(A[35]), .B(B[0]), .Z(\P0[35] ) );
  AND U1739 ( .A(A[359]), .B(B[0]), .Z(\P0[359] ) );
  AND U1740 ( .A(A[358]), .B(B[0]), .Z(\P0[358] ) );
  AND U1741 ( .A(A[357]), .B(B[0]), .Z(\P0[357] ) );
  AND U1742 ( .A(A[356]), .B(B[0]), .Z(\P0[356] ) );
  AND U1743 ( .A(A[355]), .B(B[0]), .Z(\P0[355] ) );
  AND U1744 ( .A(A[354]), .B(B[0]), .Z(\P0[354] ) );
  AND U1745 ( .A(A[353]), .B(B[0]), .Z(\P0[353] ) );
  AND U1746 ( .A(A[352]), .B(B[0]), .Z(\P0[352] ) );
  AND U1747 ( .A(A[351]), .B(B[0]), .Z(\P0[351] ) );
  AND U1748 ( .A(A[350]), .B(B[0]), .Z(\P0[350] ) );
  AND U1749 ( .A(A[34]), .B(B[0]), .Z(\P0[34] ) );
  AND U1750 ( .A(A[349]), .B(B[0]), .Z(\P0[349] ) );
  AND U1751 ( .A(A[348]), .B(B[0]), .Z(\P0[348] ) );
  AND U1752 ( .A(A[347]), .B(B[0]), .Z(\P0[347] ) );
  AND U1753 ( .A(A[346]), .B(B[0]), .Z(\P0[346] ) );
  AND U1754 ( .A(A[345]), .B(B[0]), .Z(\P0[345] ) );
  AND U1755 ( .A(A[344]), .B(B[0]), .Z(\P0[344] ) );
  AND U1756 ( .A(A[343]), .B(B[0]), .Z(\P0[343] ) );
  AND U1757 ( .A(A[342]), .B(B[0]), .Z(\P0[342] ) );
  AND U1758 ( .A(A[341]), .B(B[0]), .Z(\P0[341] ) );
  AND U1759 ( .A(A[340]), .B(B[0]), .Z(\P0[340] ) );
  AND U1760 ( .A(A[33]), .B(B[0]), .Z(\P0[33] ) );
  AND U1761 ( .A(A[339]), .B(B[0]), .Z(\P0[339] ) );
  AND U1762 ( .A(A[338]), .B(B[0]), .Z(\P0[338] ) );
  AND U1763 ( .A(A[337]), .B(B[0]), .Z(\P0[337] ) );
  AND U1764 ( .A(A[336]), .B(B[0]), .Z(\P0[336] ) );
  AND U1765 ( .A(A[335]), .B(B[0]), .Z(\P0[335] ) );
  AND U1766 ( .A(A[334]), .B(B[0]), .Z(\P0[334] ) );
  AND U1767 ( .A(A[333]), .B(B[0]), .Z(\P0[333] ) );
  AND U1768 ( .A(A[332]), .B(B[0]), .Z(\P0[332] ) );
  AND U1769 ( .A(A[331]), .B(B[0]), .Z(\P0[331] ) );
  AND U1770 ( .A(A[330]), .B(B[0]), .Z(\P0[330] ) );
  AND U1771 ( .A(A[32]), .B(B[0]), .Z(\P0[32] ) );
  AND U1772 ( .A(A[329]), .B(B[0]), .Z(\P0[329] ) );
  AND U1773 ( .A(A[328]), .B(B[0]), .Z(\P0[328] ) );
  AND U1774 ( .A(A[327]), .B(B[0]), .Z(\P0[327] ) );
  AND U1775 ( .A(A[326]), .B(B[0]), .Z(\P0[326] ) );
  AND U1776 ( .A(A[325]), .B(B[0]), .Z(\P0[325] ) );
  AND U1777 ( .A(A[324]), .B(B[0]), .Z(\P0[324] ) );
  AND U1778 ( .A(A[323]), .B(B[0]), .Z(\P0[323] ) );
  AND U1779 ( .A(A[322]), .B(B[0]), .Z(\P0[322] ) );
  AND U1780 ( .A(A[321]), .B(B[0]), .Z(\P0[321] ) );
  AND U1781 ( .A(A[320]), .B(B[0]), .Z(\P0[320] ) );
  AND U1782 ( .A(A[31]), .B(B[0]), .Z(\P0[31] ) );
  AND U1783 ( .A(A[319]), .B(B[0]), .Z(\P0[319] ) );
  AND U1784 ( .A(A[318]), .B(B[0]), .Z(\P0[318] ) );
  AND U1785 ( .A(A[317]), .B(B[0]), .Z(\P0[317] ) );
  AND U1786 ( .A(A[316]), .B(B[0]), .Z(\P0[316] ) );
  AND U1787 ( .A(A[315]), .B(B[0]), .Z(\P0[315] ) );
  AND U1788 ( .A(A[314]), .B(B[0]), .Z(\P0[314] ) );
  AND U1789 ( .A(A[313]), .B(B[0]), .Z(\P0[313] ) );
  AND U1790 ( .A(A[312]), .B(B[0]), .Z(\P0[312] ) );
  AND U1791 ( .A(A[311]), .B(B[0]), .Z(\P0[311] ) );
  AND U1792 ( .A(A[310]), .B(B[0]), .Z(\P0[310] ) );
  AND U1793 ( .A(A[30]), .B(B[0]), .Z(\P0[30] ) );
  AND U1794 ( .A(A[309]), .B(B[0]), .Z(\P0[309] ) );
  AND U1795 ( .A(A[308]), .B(B[0]), .Z(\P0[308] ) );
  AND U1796 ( .A(A[307]), .B(B[0]), .Z(\P0[307] ) );
  AND U1797 ( .A(A[306]), .B(B[0]), .Z(\P0[306] ) );
  AND U1798 ( .A(A[305]), .B(B[0]), .Z(\P0[305] ) );
  AND U1799 ( .A(A[304]), .B(B[0]), .Z(\P0[304] ) );
  AND U1800 ( .A(A[303]), .B(B[0]), .Z(\P0[303] ) );
  AND U1801 ( .A(A[302]), .B(B[0]), .Z(\P0[302] ) );
  AND U1802 ( .A(A[301]), .B(B[0]), .Z(\P0[301] ) );
  AND U1803 ( .A(A[300]), .B(B[0]), .Z(\P0[300] ) );
  AND U1804 ( .A(A[2]), .B(B[0]), .Z(\P0[2] ) );
  AND U1805 ( .A(A[29]), .B(B[0]), .Z(\P0[29] ) );
  AND U1806 ( .A(A[299]), .B(B[0]), .Z(\P0[299] ) );
  AND U1807 ( .A(A[298]), .B(B[0]), .Z(\P0[298] ) );
  AND U1808 ( .A(A[297]), .B(B[0]), .Z(\P0[297] ) );
  AND U1809 ( .A(A[296]), .B(B[0]), .Z(\P0[296] ) );
  AND U1810 ( .A(A[295]), .B(B[0]), .Z(\P0[295] ) );
  AND U1811 ( .A(A[294]), .B(B[0]), .Z(\P0[294] ) );
  AND U1812 ( .A(A[293]), .B(B[0]), .Z(\P0[293] ) );
  AND U1813 ( .A(A[292]), .B(B[0]), .Z(\P0[292] ) );
  AND U1814 ( .A(A[291]), .B(B[0]), .Z(\P0[291] ) );
  AND U1815 ( .A(A[290]), .B(B[0]), .Z(\P0[290] ) );
  AND U1816 ( .A(A[28]), .B(B[0]), .Z(\P0[28] ) );
  AND U1817 ( .A(A[289]), .B(B[0]), .Z(\P0[289] ) );
  AND U1818 ( .A(A[288]), .B(B[0]), .Z(\P0[288] ) );
  AND U1819 ( .A(A[287]), .B(B[0]), .Z(\P0[287] ) );
  AND U1820 ( .A(A[286]), .B(B[0]), .Z(\P0[286] ) );
  AND U1821 ( .A(A[285]), .B(B[0]), .Z(\P0[285] ) );
  AND U1822 ( .A(A[284]), .B(B[0]), .Z(\P0[284] ) );
  AND U1823 ( .A(A[283]), .B(B[0]), .Z(\P0[283] ) );
  AND U1824 ( .A(A[282]), .B(B[0]), .Z(\P0[282] ) );
  AND U1825 ( .A(A[281]), .B(B[0]), .Z(\P0[281] ) );
  AND U1826 ( .A(A[280]), .B(B[0]), .Z(\P0[280] ) );
  AND U1827 ( .A(A[27]), .B(B[0]), .Z(\P0[27] ) );
  AND U1828 ( .A(A[279]), .B(B[0]), .Z(\P0[279] ) );
  AND U1829 ( .A(A[278]), .B(B[0]), .Z(\P0[278] ) );
  AND U1830 ( .A(A[277]), .B(B[0]), .Z(\P0[277] ) );
  AND U1831 ( .A(A[276]), .B(B[0]), .Z(\P0[276] ) );
  AND U1832 ( .A(A[275]), .B(B[0]), .Z(\P0[275] ) );
  AND U1833 ( .A(A[274]), .B(B[0]), .Z(\P0[274] ) );
  AND U1834 ( .A(A[273]), .B(B[0]), .Z(\P0[273] ) );
  AND U1835 ( .A(A[272]), .B(B[0]), .Z(\P0[272] ) );
  AND U1836 ( .A(A[271]), .B(B[0]), .Z(\P0[271] ) );
  AND U1837 ( .A(A[270]), .B(B[0]), .Z(\P0[270] ) );
  AND U1838 ( .A(A[26]), .B(B[0]), .Z(\P0[26] ) );
  AND U1839 ( .A(A[269]), .B(B[0]), .Z(\P0[269] ) );
  AND U1840 ( .A(A[268]), .B(B[0]), .Z(\P0[268] ) );
  AND U1841 ( .A(A[267]), .B(B[0]), .Z(\P0[267] ) );
  AND U1842 ( .A(A[266]), .B(B[0]), .Z(\P0[266] ) );
  AND U1843 ( .A(A[265]), .B(B[0]), .Z(\P0[265] ) );
  AND U1844 ( .A(A[264]), .B(B[0]), .Z(\P0[264] ) );
  AND U1845 ( .A(A[263]), .B(B[0]), .Z(\P0[263] ) );
  AND U1846 ( .A(A[262]), .B(B[0]), .Z(\P0[262] ) );
  AND U1847 ( .A(A[261]), .B(B[0]), .Z(\P0[261] ) );
  AND U1848 ( .A(A[260]), .B(B[0]), .Z(\P0[260] ) );
  AND U1849 ( .A(A[25]), .B(B[0]), .Z(\P0[25] ) );
  AND U1850 ( .A(A[259]), .B(B[0]), .Z(\P0[259] ) );
  AND U1851 ( .A(A[258]), .B(B[0]), .Z(\P0[258] ) );
  AND U1852 ( .A(A[257]), .B(B[0]), .Z(\P0[257] ) );
  AND U1853 ( .A(A[256]), .B(B[0]), .Z(\P0[256] ) );
  AND U1854 ( .A(A[255]), .B(B[0]), .Z(\P0[255] ) );
  AND U1855 ( .A(A[254]), .B(B[0]), .Z(\P0[254] ) );
  AND U1856 ( .A(A[253]), .B(B[0]), .Z(\P0[253] ) );
  AND U1857 ( .A(A[252]), .B(B[0]), .Z(\P0[252] ) );
  AND U1858 ( .A(A[251]), .B(B[0]), .Z(\P0[251] ) );
  AND U1859 ( .A(A[250]), .B(B[0]), .Z(\P0[250] ) );
  AND U1860 ( .A(A[24]), .B(B[0]), .Z(\P0[24] ) );
  AND U1861 ( .A(A[249]), .B(B[0]), .Z(\P0[249] ) );
  AND U1862 ( .A(A[248]), .B(B[0]), .Z(\P0[248] ) );
  AND U1863 ( .A(A[247]), .B(B[0]), .Z(\P0[247] ) );
  AND U1864 ( .A(A[246]), .B(B[0]), .Z(\P0[246] ) );
  AND U1865 ( .A(A[245]), .B(B[0]), .Z(\P0[245] ) );
  AND U1866 ( .A(A[244]), .B(B[0]), .Z(\P0[244] ) );
  AND U1867 ( .A(A[243]), .B(B[0]), .Z(\P0[243] ) );
  AND U1868 ( .A(A[242]), .B(B[0]), .Z(\P0[242] ) );
  AND U1869 ( .A(A[241]), .B(B[0]), .Z(\P0[241] ) );
  AND U1870 ( .A(A[240]), .B(B[0]), .Z(\P0[240] ) );
  AND U1871 ( .A(A[23]), .B(B[0]), .Z(\P0[23] ) );
  AND U1872 ( .A(A[239]), .B(B[0]), .Z(\P0[239] ) );
  AND U1873 ( .A(A[238]), .B(B[0]), .Z(\P0[238] ) );
  AND U1874 ( .A(A[237]), .B(B[0]), .Z(\P0[237] ) );
  AND U1875 ( .A(A[236]), .B(B[0]), .Z(\P0[236] ) );
  AND U1876 ( .A(A[235]), .B(B[0]), .Z(\P0[235] ) );
  AND U1877 ( .A(A[234]), .B(B[0]), .Z(\P0[234] ) );
  AND U1878 ( .A(A[233]), .B(B[0]), .Z(\P0[233] ) );
  AND U1879 ( .A(A[232]), .B(B[0]), .Z(\P0[232] ) );
  AND U1880 ( .A(A[231]), .B(B[0]), .Z(\P0[231] ) );
  AND U1881 ( .A(A[230]), .B(B[0]), .Z(\P0[230] ) );
  AND U1882 ( .A(A[22]), .B(B[0]), .Z(\P0[22] ) );
  AND U1883 ( .A(A[229]), .B(B[0]), .Z(\P0[229] ) );
  AND U1884 ( .A(A[228]), .B(B[0]), .Z(\P0[228] ) );
  AND U1885 ( .A(A[227]), .B(B[0]), .Z(\P0[227] ) );
  AND U1886 ( .A(A[226]), .B(B[0]), .Z(\P0[226] ) );
  AND U1887 ( .A(A[225]), .B(B[0]), .Z(\P0[225] ) );
  AND U1888 ( .A(A[224]), .B(B[0]), .Z(\P0[224] ) );
  AND U1889 ( .A(A[223]), .B(B[0]), .Z(\P0[223] ) );
  AND U1890 ( .A(A[222]), .B(B[0]), .Z(\P0[222] ) );
  AND U1891 ( .A(A[221]), .B(B[0]), .Z(\P0[221] ) );
  AND U1892 ( .A(A[220]), .B(B[0]), .Z(\P0[220] ) );
  AND U1893 ( .A(A[21]), .B(B[0]), .Z(\P0[21] ) );
  AND U1894 ( .A(A[219]), .B(B[0]), .Z(\P0[219] ) );
  AND U1895 ( .A(A[218]), .B(B[0]), .Z(\P0[218] ) );
  AND U1896 ( .A(A[217]), .B(B[0]), .Z(\P0[217] ) );
  AND U1897 ( .A(A[216]), .B(B[0]), .Z(\P0[216] ) );
  AND U1898 ( .A(A[215]), .B(B[0]), .Z(\P0[215] ) );
  AND U1899 ( .A(A[214]), .B(B[0]), .Z(\P0[214] ) );
  AND U1900 ( .A(A[213]), .B(B[0]), .Z(\P0[213] ) );
  AND U1901 ( .A(A[212]), .B(B[0]), .Z(\P0[212] ) );
  AND U1902 ( .A(A[211]), .B(B[0]), .Z(\P0[211] ) );
  AND U1903 ( .A(A[210]), .B(B[0]), .Z(\P0[210] ) );
  AND U1904 ( .A(A[20]), .B(B[0]), .Z(\P0[20] ) );
  AND U1905 ( .A(A[209]), .B(B[0]), .Z(\P0[209] ) );
  AND U1906 ( .A(A[208]), .B(B[0]), .Z(\P0[208] ) );
  AND U1907 ( .A(A[207]), .B(B[0]), .Z(\P0[207] ) );
  AND U1908 ( .A(A[206]), .B(B[0]), .Z(\P0[206] ) );
  AND U1909 ( .A(A[205]), .B(B[0]), .Z(\P0[205] ) );
  AND U1910 ( .A(A[204]), .B(B[0]), .Z(\P0[204] ) );
  AND U1911 ( .A(A[203]), .B(B[0]), .Z(\P0[203] ) );
  AND U1912 ( .A(A[202]), .B(B[0]), .Z(\P0[202] ) );
  AND U1913 ( .A(A[201]), .B(B[0]), .Z(\P0[201] ) );
  AND U1914 ( .A(A[200]), .B(B[0]), .Z(\P0[200] ) );
  AND U1915 ( .A(A[1]), .B(B[0]), .Z(\P0[1] ) );
  AND U1916 ( .A(A[19]), .B(B[0]), .Z(\P0[19] ) );
  AND U1917 ( .A(A[199]), .B(B[0]), .Z(\P0[199] ) );
  AND U1918 ( .A(A[198]), .B(B[0]), .Z(\P0[198] ) );
  AND U1919 ( .A(A[197]), .B(B[0]), .Z(\P0[197] ) );
  AND U1920 ( .A(A[196]), .B(B[0]), .Z(\P0[196] ) );
  AND U1921 ( .A(A[195]), .B(B[0]), .Z(\P0[195] ) );
  AND U1922 ( .A(A[194]), .B(B[0]), .Z(\P0[194] ) );
  AND U1923 ( .A(A[193]), .B(B[0]), .Z(\P0[193] ) );
  AND U1924 ( .A(A[192]), .B(B[0]), .Z(\P0[192] ) );
  AND U1925 ( .A(A[191]), .B(B[0]), .Z(\P0[191] ) );
  AND U1926 ( .A(A[190]), .B(B[0]), .Z(\P0[190] ) );
  AND U1927 ( .A(A[18]), .B(B[0]), .Z(\P0[18] ) );
  AND U1928 ( .A(A[189]), .B(B[0]), .Z(\P0[189] ) );
  AND U1929 ( .A(A[188]), .B(B[0]), .Z(\P0[188] ) );
  AND U1930 ( .A(A[187]), .B(B[0]), .Z(\P0[187] ) );
  AND U1931 ( .A(A[186]), .B(B[0]), .Z(\P0[186] ) );
  AND U1932 ( .A(A[185]), .B(B[0]), .Z(\P0[185] ) );
  AND U1933 ( .A(A[184]), .B(B[0]), .Z(\P0[184] ) );
  AND U1934 ( .A(A[183]), .B(B[0]), .Z(\P0[183] ) );
  AND U1935 ( .A(A[182]), .B(B[0]), .Z(\P0[182] ) );
  AND U1936 ( .A(A[181]), .B(B[0]), .Z(\P0[181] ) );
  AND U1937 ( .A(A[180]), .B(B[0]), .Z(\P0[180] ) );
  AND U1938 ( .A(A[17]), .B(B[0]), .Z(\P0[17] ) );
  AND U1939 ( .A(A[179]), .B(B[0]), .Z(\P0[179] ) );
  AND U1940 ( .A(A[178]), .B(B[0]), .Z(\P0[178] ) );
  AND U1941 ( .A(A[177]), .B(B[0]), .Z(\P0[177] ) );
  AND U1942 ( .A(A[176]), .B(B[0]), .Z(\P0[176] ) );
  AND U1943 ( .A(A[175]), .B(B[0]), .Z(\P0[175] ) );
  AND U1944 ( .A(A[174]), .B(B[0]), .Z(\P0[174] ) );
  AND U1945 ( .A(A[173]), .B(B[0]), .Z(\P0[173] ) );
  AND U1946 ( .A(A[172]), .B(B[0]), .Z(\P0[172] ) );
  AND U1947 ( .A(A[171]), .B(B[0]), .Z(\P0[171] ) );
  AND U1948 ( .A(A[170]), .B(B[0]), .Z(\P0[170] ) );
  AND U1949 ( .A(A[16]), .B(B[0]), .Z(\P0[16] ) );
  AND U1950 ( .A(A[169]), .B(B[0]), .Z(\P0[169] ) );
  AND U1951 ( .A(A[168]), .B(B[0]), .Z(\P0[168] ) );
  AND U1952 ( .A(A[167]), .B(B[0]), .Z(\P0[167] ) );
  AND U1953 ( .A(A[166]), .B(B[0]), .Z(\P0[166] ) );
  AND U1954 ( .A(A[165]), .B(B[0]), .Z(\P0[165] ) );
  AND U1955 ( .A(A[164]), .B(B[0]), .Z(\P0[164] ) );
  AND U1956 ( .A(A[163]), .B(B[0]), .Z(\P0[163] ) );
  AND U1957 ( .A(A[162]), .B(B[0]), .Z(\P0[162] ) );
  AND U1958 ( .A(A[161]), .B(B[0]), .Z(\P0[161] ) );
  AND U1959 ( .A(A[160]), .B(B[0]), .Z(\P0[160] ) );
  AND U1960 ( .A(A[15]), .B(B[0]), .Z(\P0[15] ) );
  AND U1961 ( .A(A[159]), .B(B[0]), .Z(\P0[159] ) );
  AND U1962 ( .A(A[158]), .B(B[0]), .Z(\P0[158] ) );
  AND U1963 ( .A(A[157]), .B(B[0]), .Z(\P0[157] ) );
  AND U1964 ( .A(A[156]), .B(B[0]), .Z(\P0[156] ) );
  AND U1965 ( .A(A[155]), .B(B[0]), .Z(\P0[155] ) );
  AND U1966 ( .A(A[154]), .B(B[0]), .Z(\P0[154] ) );
  AND U1967 ( .A(A[153]), .B(B[0]), .Z(\P0[153] ) );
  AND U1968 ( .A(A[152]), .B(B[0]), .Z(\P0[152] ) );
  AND U1969 ( .A(A[151]), .B(B[0]), .Z(\P0[151] ) );
  AND U1970 ( .A(A[150]), .B(B[0]), .Z(\P0[150] ) );
  AND U1971 ( .A(A[14]), .B(B[0]), .Z(\P0[14] ) );
  AND U1972 ( .A(A[149]), .B(B[0]), .Z(\P0[149] ) );
  AND U1973 ( .A(A[148]), .B(B[0]), .Z(\P0[148] ) );
  AND U1974 ( .A(A[147]), .B(B[0]), .Z(\P0[147] ) );
  AND U1975 ( .A(A[146]), .B(B[0]), .Z(\P0[146] ) );
  AND U1976 ( .A(A[145]), .B(B[0]), .Z(\P0[145] ) );
  AND U1977 ( .A(A[144]), .B(B[0]), .Z(\P0[144] ) );
  AND U1978 ( .A(A[143]), .B(B[0]), .Z(\P0[143] ) );
  AND U1979 ( .A(A[142]), .B(B[0]), .Z(\P0[142] ) );
  AND U1980 ( .A(A[141]), .B(B[0]), .Z(\P0[141] ) );
  AND U1981 ( .A(A[140]), .B(B[0]), .Z(\P0[140] ) );
  AND U1982 ( .A(A[13]), .B(B[0]), .Z(\P0[13] ) );
  AND U1983 ( .A(A[139]), .B(B[0]), .Z(\P0[139] ) );
  AND U1984 ( .A(A[138]), .B(B[0]), .Z(\P0[138] ) );
  AND U1985 ( .A(A[137]), .B(B[0]), .Z(\P0[137] ) );
  AND U1986 ( .A(A[136]), .B(B[0]), .Z(\P0[136] ) );
  AND U1987 ( .A(A[135]), .B(B[0]), .Z(\P0[135] ) );
  AND U1988 ( .A(A[134]), .B(B[0]), .Z(\P0[134] ) );
  AND U1989 ( .A(A[133]), .B(B[0]), .Z(\P0[133] ) );
  AND U1990 ( .A(A[132]), .B(B[0]), .Z(\P0[132] ) );
  AND U1991 ( .A(A[131]), .B(B[0]), .Z(\P0[131] ) );
  AND U1992 ( .A(A[130]), .B(B[0]), .Z(\P0[130] ) );
  AND U1993 ( .A(A[12]), .B(B[0]), .Z(\P0[12] ) );
  AND U1994 ( .A(A[129]), .B(B[0]), .Z(\P0[129] ) );
  AND U1995 ( .A(A[128]), .B(B[0]), .Z(\P0[128] ) );
  AND U1996 ( .A(A[127]), .B(B[0]), .Z(\P0[127] ) );
  AND U1997 ( .A(A[126]), .B(B[0]), .Z(\P0[126] ) );
  AND U1998 ( .A(A[125]), .B(B[0]), .Z(\P0[125] ) );
  AND U1999 ( .A(A[124]), .B(B[0]), .Z(\P0[124] ) );
  AND U2000 ( .A(A[123]), .B(B[0]), .Z(\P0[123] ) );
  AND U2001 ( .A(A[122]), .B(B[0]), .Z(\P0[122] ) );
  AND U2002 ( .A(A[121]), .B(B[0]), .Z(\P0[121] ) );
  AND U2003 ( .A(A[120]), .B(B[0]), .Z(\P0[120] ) );
  AND U2004 ( .A(A[11]), .B(B[0]), .Z(\P0[11] ) );
  AND U2005 ( .A(A[119]), .B(B[0]), .Z(\P0[119] ) );
  AND U2006 ( .A(A[118]), .B(B[0]), .Z(\P0[118] ) );
  AND U2007 ( .A(A[117]), .B(B[0]), .Z(\P0[117] ) );
  AND U2008 ( .A(A[116]), .B(B[0]), .Z(\P0[116] ) );
  AND U2009 ( .A(A[115]), .B(B[0]), .Z(\P0[115] ) );
  AND U2010 ( .A(A[114]), .B(B[0]), .Z(\P0[114] ) );
  AND U2011 ( .A(A[113]), .B(B[0]), .Z(\P0[113] ) );
  AND U2012 ( .A(A[112]), .B(B[0]), .Z(\P0[112] ) );
  AND U2013 ( .A(A[111]), .B(B[0]), .Z(\P0[111] ) );
  AND U2014 ( .A(A[110]), .B(B[0]), .Z(\P0[110] ) );
  AND U2015 ( .A(A[10]), .B(B[0]), .Z(\P0[10] ) );
  AND U2016 ( .A(A[109]), .B(B[0]), .Z(\P0[109] ) );
  AND U2017 ( .A(A[108]), .B(B[0]), .Z(\P0[108] ) );
  AND U2018 ( .A(A[107]), .B(B[0]), .Z(\P0[107] ) );
  AND U2019 ( .A(A[106]), .B(B[0]), .Z(\P0[106] ) );
  AND U2020 ( .A(A[105]), .B(B[0]), .Z(\P0[105] ) );
  AND U2021 ( .A(A[104]), .B(B[0]), .Z(\P0[104] ) );
  AND U2022 ( .A(A[103]), .B(B[0]), .Z(\P0[103] ) );
  AND U2023 ( .A(A[102]), .B(B[0]), .Z(\P0[102] ) );
  AND U2024 ( .A(A[1023]), .B(B[0]), .Z(\P0[1023] ) );
  AND U2025 ( .A(A[1022]), .B(B[0]), .Z(\P0[1022] ) );
  AND U2026 ( .A(A[1021]), .B(B[0]), .Z(\P0[1021] ) );
  AND U2027 ( .A(A[1020]), .B(B[0]), .Z(\P0[1020] ) );
  AND U2028 ( .A(A[101]), .B(B[0]), .Z(\P0[101] ) );
  AND U2029 ( .A(A[1019]), .B(B[0]), .Z(\P0[1019] ) );
  AND U2030 ( .A(A[1018]), .B(B[0]), .Z(\P0[1018] ) );
  AND U2031 ( .A(A[1017]), .B(B[0]), .Z(\P0[1017] ) );
  AND U2032 ( .A(A[1016]), .B(B[0]), .Z(\P0[1016] ) );
  AND U2033 ( .A(A[1015]), .B(B[0]), .Z(\P0[1015] ) );
  AND U2034 ( .A(A[1014]), .B(B[0]), .Z(\P0[1014] ) );
  AND U2035 ( .A(A[1013]), .B(B[0]), .Z(\P0[1013] ) );
  AND U2036 ( .A(A[1012]), .B(B[0]), .Z(\P0[1012] ) );
  AND U2037 ( .A(A[1011]), .B(B[0]), .Z(\P0[1011] ) );
  AND U2038 ( .A(A[1010]), .B(B[0]), .Z(\P0[1010] ) );
  AND U2039 ( .A(A[100]), .B(B[0]), .Z(\P0[100] ) );
  AND U2040 ( .A(A[1009]), .B(B[0]), .Z(\P0[1009] ) );
  AND U2041 ( .A(A[1008]), .B(B[0]), .Z(\P0[1008] ) );
  AND U2042 ( .A(A[1007]), .B(B[0]), .Z(\P0[1007] ) );
  AND U2043 ( .A(A[1006]), .B(B[0]), .Z(\P0[1006] ) );
  AND U2044 ( .A(A[1005]), .B(B[0]), .Z(\P0[1005] ) );
  AND U2045 ( .A(A[1004]), .B(B[0]), .Z(\P0[1004] ) );
  AND U2046 ( .A(A[1003]), .B(B[0]), .Z(\P0[1003] ) );
  AND U2047 ( .A(A[1002]), .B(B[0]), .Z(\P0[1002] ) );
  AND U2048 ( .A(A[1001]), .B(B[0]), .Z(\P0[1001] ) );
  AND U2049 ( .A(A[1000]), .B(B[0]), .Z(\P0[1000] ) );
endmodule


module mult_N1024_CC512 ( clk, rst, a, b, c );
  input [1023:0] a;
  input [1:0] b;
  output [1023:0] c;
  input clk, rst;

  wire   [1023:2] swire;
  wire   [1023:0] clocal;
  wire   [2047:1024] sreg;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;

  DFF \sreg_reg[1024]  ( .D(swire[2]), .CLK(clk), .RST(rst), .Q(sreg[1024]) );
  DFF \sreg_reg[1025]  ( .D(swire[3]), .CLK(clk), .RST(rst), .Q(sreg[1025]) );
  DFF \sreg_reg[1026]  ( .D(swire[4]), .CLK(clk), .RST(rst), .Q(sreg[1026]) );
  DFF \sreg_reg[1027]  ( .D(swire[5]), .CLK(clk), .RST(rst), .Q(sreg[1027]) );
  DFF \sreg_reg[1028]  ( .D(swire[6]), .CLK(clk), .RST(rst), .Q(sreg[1028]) );
  DFF \sreg_reg[1029]  ( .D(swire[7]), .CLK(clk), .RST(rst), .Q(sreg[1029]) );
  DFF \sreg_reg[1030]  ( .D(swire[8]), .CLK(clk), .RST(rst), .Q(sreg[1030]) );
  DFF \sreg_reg[1031]  ( .D(swire[9]), .CLK(clk), .RST(rst), .Q(sreg[1031]) );
  DFF \sreg_reg[1032]  ( .D(swire[10]), .CLK(clk), .RST(rst), .Q(sreg[1032])
         );
  DFF \sreg_reg[1033]  ( .D(swire[11]), .CLK(clk), .RST(rst), .Q(sreg[1033])
         );
  DFF \sreg_reg[1034]  ( .D(swire[12]), .CLK(clk), .RST(rst), .Q(sreg[1034])
         );
  DFF \sreg_reg[1035]  ( .D(swire[13]), .CLK(clk), .RST(rst), .Q(sreg[1035])
         );
  DFF \sreg_reg[1036]  ( .D(swire[14]), .CLK(clk), .RST(rst), .Q(sreg[1036])
         );
  DFF \sreg_reg[1037]  ( .D(swire[15]), .CLK(clk), .RST(rst), .Q(sreg[1037])
         );
  DFF \sreg_reg[1038]  ( .D(swire[16]), .CLK(clk), .RST(rst), .Q(sreg[1038])
         );
  DFF \sreg_reg[1039]  ( .D(swire[17]), .CLK(clk), .RST(rst), .Q(sreg[1039])
         );
  DFF \sreg_reg[1040]  ( .D(swire[18]), .CLK(clk), .RST(rst), .Q(sreg[1040])
         );
  DFF \sreg_reg[1041]  ( .D(swire[19]), .CLK(clk), .RST(rst), .Q(sreg[1041])
         );
  DFF \sreg_reg[1042]  ( .D(swire[20]), .CLK(clk), .RST(rst), .Q(sreg[1042])
         );
  DFF \sreg_reg[1043]  ( .D(swire[21]), .CLK(clk), .RST(rst), .Q(sreg[1043])
         );
  DFF \sreg_reg[1044]  ( .D(swire[22]), .CLK(clk), .RST(rst), .Q(sreg[1044])
         );
  DFF \sreg_reg[1045]  ( .D(swire[23]), .CLK(clk), .RST(rst), .Q(sreg[1045])
         );
  DFF \sreg_reg[1046]  ( .D(swire[24]), .CLK(clk), .RST(rst), .Q(sreg[1046])
         );
  DFF \sreg_reg[1047]  ( .D(swire[25]), .CLK(clk), .RST(rst), .Q(sreg[1047])
         );
  DFF \sreg_reg[1048]  ( .D(swire[26]), .CLK(clk), .RST(rst), .Q(sreg[1048])
         );
  DFF \sreg_reg[1049]  ( .D(swire[27]), .CLK(clk), .RST(rst), .Q(sreg[1049])
         );
  DFF \sreg_reg[1050]  ( .D(swire[28]), .CLK(clk), .RST(rst), .Q(sreg[1050])
         );
  DFF \sreg_reg[1051]  ( .D(swire[29]), .CLK(clk), .RST(rst), .Q(sreg[1051])
         );
  DFF \sreg_reg[1052]  ( .D(swire[30]), .CLK(clk), .RST(rst), .Q(sreg[1052])
         );
  DFF \sreg_reg[1053]  ( .D(swire[31]), .CLK(clk), .RST(rst), .Q(sreg[1053])
         );
  DFF \sreg_reg[1054]  ( .D(swire[32]), .CLK(clk), .RST(rst), .Q(sreg[1054])
         );
  DFF \sreg_reg[1055]  ( .D(swire[33]), .CLK(clk), .RST(rst), .Q(sreg[1055])
         );
  DFF \sreg_reg[1056]  ( .D(swire[34]), .CLK(clk), .RST(rst), .Q(sreg[1056])
         );
  DFF \sreg_reg[1057]  ( .D(swire[35]), .CLK(clk), .RST(rst), .Q(sreg[1057])
         );
  DFF \sreg_reg[1058]  ( .D(swire[36]), .CLK(clk), .RST(rst), .Q(sreg[1058])
         );
  DFF \sreg_reg[1059]  ( .D(swire[37]), .CLK(clk), .RST(rst), .Q(sreg[1059])
         );
  DFF \sreg_reg[1060]  ( .D(swire[38]), .CLK(clk), .RST(rst), .Q(sreg[1060])
         );
  DFF \sreg_reg[1061]  ( .D(swire[39]), .CLK(clk), .RST(rst), .Q(sreg[1061])
         );
  DFF \sreg_reg[1062]  ( .D(swire[40]), .CLK(clk), .RST(rst), .Q(sreg[1062])
         );
  DFF \sreg_reg[1063]  ( .D(swire[41]), .CLK(clk), .RST(rst), .Q(sreg[1063])
         );
  DFF \sreg_reg[1064]  ( .D(swire[42]), .CLK(clk), .RST(rst), .Q(sreg[1064])
         );
  DFF \sreg_reg[1065]  ( .D(swire[43]), .CLK(clk), .RST(rst), .Q(sreg[1065])
         );
  DFF \sreg_reg[1066]  ( .D(swire[44]), .CLK(clk), .RST(rst), .Q(sreg[1066])
         );
  DFF \sreg_reg[1067]  ( .D(swire[45]), .CLK(clk), .RST(rst), .Q(sreg[1067])
         );
  DFF \sreg_reg[1068]  ( .D(swire[46]), .CLK(clk), .RST(rst), .Q(sreg[1068])
         );
  DFF \sreg_reg[1069]  ( .D(swire[47]), .CLK(clk), .RST(rst), .Q(sreg[1069])
         );
  DFF \sreg_reg[1070]  ( .D(swire[48]), .CLK(clk), .RST(rst), .Q(sreg[1070])
         );
  DFF \sreg_reg[1071]  ( .D(swire[49]), .CLK(clk), .RST(rst), .Q(sreg[1071])
         );
  DFF \sreg_reg[1072]  ( .D(swire[50]), .CLK(clk), .RST(rst), .Q(sreg[1072])
         );
  DFF \sreg_reg[1073]  ( .D(swire[51]), .CLK(clk), .RST(rst), .Q(sreg[1073])
         );
  DFF \sreg_reg[1074]  ( .D(swire[52]), .CLK(clk), .RST(rst), .Q(sreg[1074])
         );
  DFF \sreg_reg[1075]  ( .D(swire[53]), .CLK(clk), .RST(rst), .Q(sreg[1075])
         );
  DFF \sreg_reg[1076]  ( .D(swire[54]), .CLK(clk), .RST(rst), .Q(sreg[1076])
         );
  DFF \sreg_reg[1077]  ( .D(swire[55]), .CLK(clk), .RST(rst), .Q(sreg[1077])
         );
  DFF \sreg_reg[1078]  ( .D(swire[56]), .CLK(clk), .RST(rst), .Q(sreg[1078])
         );
  DFF \sreg_reg[1079]  ( .D(swire[57]), .CLK(clk), .RST(rst), .Q(sreg[1079])
         );
  DFF \sreg_reg[1080]  ( .D(swire[58]), .CLK(clk), .RST(rst), .Q(sreg[1080])
         );
  DFF \sreg_reg[1081]  ( .D(swire[59]), .CLK(clk), .RST(rst), .Q(sreg[1081])
         );
  DFF \sreg_reg[1082]  ( .D(swire[60]), .CLK(clk), .RST(rst), .Q(sreg[1082])
         );
  DFF \sreg_reg[1083]  ( .D(swire[61]), .CLK(clk), .RST(rst), .Q(sreg[1083])
         );
  DFF \sreg_reg[1084]  ( .D(swire[62]), .CLK(clk), .RST(rst), .Q(sreg[1084])
         );
  DFF \sreg_reg[1085]  ( .D(swire[63]), .CLK(clk), .RST(rst), .Q(sreg[1085])
         );
  DFF \sreg_reg[1086]  ( .D(swire[64]), .CLK(clk), .RST(rst), .Q(sreg[1086])
         );
  DFF \sreg_reg[1087]  ( .D(swire[65]), .CLK(clk), .RST(rst), .Q(sreg[1087])
         );
  DFF \sreg_reg[1088]  ( .D(swire[66]), .CLK(clk), .RST(rst), .Q(sreg[1088])
         );
  DFF \sreg_reg[1089]  ( .D(swire[67]), .CLK(clk), .RST(rst), .Q(sreg[1089])
         );
  DFF \sreg_reg[1090]  ( .D(swire[68]), .CLK(clk), .RST(rst), .Q(sreg[1090])
         );
  DFF \sreg_reg[1091]  ( .D(swire[69]), .CLK(clk), .RST(rst), .Q(sreg[1091])
         );
  DFF \sreg_reg[1092]  ( .D(swire[70]), .CLK(clk), .RST(rst), .Q(sreg[1092])
         );
  DFF \sreg_reg[1093]  ( .D(swire[71]), .CLK(clk), .RST(rst), .Q(sreg[1093])
         );
  DFF \sreg_reg[1094]  ( .D(swire[72]), .CLK(clk), .RST(rst), .Q(sreg[1094])
         );
  DFF \sreg_reg[1095]  ( .D(swire[73]), .CLK(clk), .RST(rst), .Q(sreg[1095])
         );
  DFF \sreg_reg[1096]  ( .D(swire[74]), .CLK(clk), .RST(rst), .Q(sreg[1096])
         );
  DFF \sreg_reg[1097]  ( .D(swire[75]), .CLK(clk), .RST(rst), .Q(sreg[1097])
         );
  DFF \sreg_reg[1098]  ( .D(swire[76]), .CLK(clk), .RST(rst), .Q(sreg[1098])
         );
  DFF \sreg_reg[1099]  ( .D(swire[77]), .CLK(clk), .RST(rst), .Q(sreg[1099])
         );
  DFF \sreg_reg[1100]  ( .D(swire[78]), .CLK(clk), .RST(rst), .Q(sreg[1100])
         );
  DFF \sreg_reg[1101]  ( .D(swire[79]), .CLK(clk), .RST(rst), .Q(sreg[1101])
         );
  DFF \sreg_reg[1102]  ( .D(swire[80]), .CLK(clk), .RST(rst), .Q(sreg[1102])
         );
  DFF \sreg_reg[1103]  ( .D(swire[81]), .CLK(clk), .RST(rst), .Q(sreg[1103])
         );
  DFF \sreg_reg[1104]  ( .D(swire[82]), .CLK(clk), .RST(rst), .Q(sreg[1104])
         );
  DFF \sreg_reg[1105]  ( .D(swire[83]), .CLK(clk), .RST(rst), .Q(sreg[1105])
         );
  DFF \sreg_reg[1106]  ( .D(swire[84]), .CLK(clk), .RST(rst), .Q(sreg[1106])
         );
  DFF \sreg_reg[1107]  ( .D(swire[85]), .CLK(clk), .RST(rst), .Q(sreg[1107])
         );
  DFF \sreg_reg[1108]  ( .D(swire[86]), .CLK(clk), .RST(rst), .Q(sreg[1108])
         );
  DFF \sreg_reg[1109]  ( .D(swire[87]), .CLK(clk), .RST(rst), .Q(sreg[1109])
         );
  DFF \sreg_reg[1110]  ( .D(swire[88]), .CLK(clk), .RST(rst), .Q(sreg[1110])
         );
  DFF \sreg_reg[1111]  ( .D(swire[89]), .CLK(clk), .RST(rst), .Q(sreg[1111])
         );
  DFF \sreg_reg[1112]  ( .D(swire[90]), .CLK(clk), .RST(rst), .Q(sreg[1112])
         );
  DFF \sreg_reg[1113]  ( .D(swire[91]), .CLK(clk), .RST(rst), .Q(sreg[1113])
         );
  DFF \sreg_reg[1114]  ( .D(swire[92]), .CLK(clk), .RST(rst), .Q(sreg[1114])
         );
  DFF \sreg_reg[1115]  ( .D(swire[93]), .CLK(clk), .RST(rst), .Q(sreg[1115])
         );
  DFF \sreg_reg[1116]  ( .D(swire[94]), .CLK(clk), .RST(rst), .Q(sreg[1116])
         );
  DFF \sreg_reg[1117]  ( .D(swire[95]), .CLK(clk), .RST(rst), .Q(sreg[1117])
         );
  DFF \sreg_reg[1118]  ( .D(swire[96]), .CLK(clk), .RST(rst), .Q(sreg[1118])
         );
  DFF \sreg_reg[1119]  ( .D(swire[97]), .CLK(clk), .RST(rst), .Q(sreg[1119])
         );
  DFF \sreg_reg[1120]  ( .D(swire[98]), .CLK(clk), .RST(rst), .Q(sreg[1120])
         );
  DFF \sreg_reg[1121]  ( .D(swire[99]), .CLK(clk), .RST(rst), .Q(sreg[1121])
         );
  DFF \sreg_reg[1122]  ( .D(swire[100]), .CLK(clk), .RST(rst), .Q(sreg[1122])
         );
  DFF \sreg_reg[1123]  ( .D(swire[101]), .CLK(clk), .RST(rst), .Q(sreg[1123])
         );
  DFF \sreg_reg[1124]  ( .D(swire[102]), .CLK(clk), .RST(rst), .Q(sreg[1124])
         );
  DFF \sreg_reg[1125]  ( .D(swire[103]), .CLK(clk), .RST(rst), .Q(sreg[1125])
         );
  DFF \sreg_reg[1126]  ( .D(swire[104]), .CLK(clk), .RST(rst), .Q(sreg[1126])
         );
  DFF \sreg_reg[1127]  ( .D(swire[105]), .CLK(clk), .RST(rst), .Q(sreg[1127])
         );
  DFF \sreg_reg[1128]  ( .D(swire[106]), .CLK(clk), .RST(rst), .Q(sreg[1128])
         );
  DFF \sreg_reg[1129]  ( .D(swire[107]), .CLK(clk), .RST(rst), .Q(sreg[1129])
         );
  DFF \sreg_reg[1130]  ( .D(swire[108]), .CLK(clk), .RST(rst), .Q(sreg[1130])
         );
  DFF \sreg_reg[1131]  ( .D(swire[109]), .CLK(clk), .RST(rst), .Q(sreg[1131])
         );
  DFF \sreg_reg[1132]  ( .D(swire[110]), .CLK(clk), .RST(rst), .Q(sreg[1132])
         );
  DFF \sreg_reg[1133]  ( .D(swire[111]), .CLK(clk), .RST(rst), .Q(sreg[1133])
         );
  DFF \sreg_reg[1134]  ( .D(swire[112]), .CLK(clk), .RST(rst), .Q(sreg[1134])
         );
  DFF \sreg_reg[1135]  ( .D(swire[113]), .CLK(clk), .RST(rst), .Q(sreg[1135])
         );
  DFF \sreg_reg[1136]  ( .D(swire[114]), .CLK(clk), .RST(rst), .Q(sreg[1136])
         );
  DFF \sreg_reg[1137]  ( .D(swire[115]), .CLK(clk), .RST(rst), .Q(sreg[1137])
         );
  DFF \sreg_reg[1138]  ( .D(swire[116]), .CLK(clk), .RST(rst), .Q(sreg[1138])
         );
  DFF \sreg_reg[1139]  ( .D(swire[117]), .CLK(clk), .RST(rst), .Q(sreg[1139])
         );
  DFF \sreg_reg[1140]  ( .D(swire[118]), .CLK(clk), .RST(rst), .Q(sreg[1140])
         );
  DFF \sreg_reg[1141]  ( .D(swire[119]), .CLK(clk), .RST(rst), .Q(sreg[1141])
         );
  DFF \sreg_reg[1142]  ( .D(swire[120]), .CLK(clk), .RST(rst), .Q(sreg[1142])
         );
  DFF \sreg_reg[1143]  ( .D(swire[121]), .CLK(clk), .RST(rst), .Q(sreg[1143])
         );
  DFF \sreg_reg[1144]  ( .D(swire[122]), .CLK(clk), .RST(rst), .Q(sreg[1144])
         );
  DFF \sreg_reg[1145]  ( .D(swire[123]), .CLK(clk), .RST(rst), .Q(sreg[1145])
         );
  DFF \sreg_reg[1146]  ( .D(swire[124]), .CLK(clk), .RST(rst), .Q(sreg[1146])
         );
  DFF \sreg_reg[1147]  ( .D(swire[125]), .CLK(clk), .RST(rst), .Q(sreg[1147])
         );
  DFF \sreg_reg[1148]  ( .D(swire[126]), .CLK(clk), .RST(rst), .Q(sreg[1148])
         );
  DFF \sreg_reg[1149]  ( .D(swire[127]), .CLK(clk), .RST(rst), .Q(sreg[1149])
         );
  DFF \sreg_reg[1150]  ( .D(swire[128]), .CLK(clk), .RST(rst), .Q(sreg[1150])
         );
  DFF \sreg_reg[1151]  ( .D(swire[129]), .CLK(clk), .RST(rst), .Q(sreg[1151])
         );
  DFF \sreg_reg[1152]  ( .D(swire[130]), .CLK(clk), .RST(rst), .Q(sreg[1152])
         );
  DFF \sreg_reg[1153]  ( .D(swire[131]), .CLK(clk), .RST(rst), .Q(sreg[1153])
         );
  DFF \sreg_reg[1154]  ( .D(swire[132]), .CLK(clk), .RST(rst), .Q(sreg[1154])
         );
  DFF \sreg_reg[1155]  ( .D(swire[133]), .CLK(clk), .RST(rst), .Q(sreg[1155])
         );
  DFF \sreg_reg[1156]  ( .D(swire[134]), .CLK(clk), .RST(rst), .Q(sreg[1156])
         );
  DFF \sreg_reg[1157]  ( .D(swire[135]), .CLK(clk), .RST(rst), .Q(sreg[1157])
         );
  DFF \sreg_reg[1158]  ( .D(swire[136]), .CLK(clk), .RST(rst), .Q(sreg[1158])
         );
  DFF \sreg_reg[1159]  ( .D(swire[137]), .CLK(clk), .RST(rst), .Q(sreg[1159])
         );
  DFF \sreg_reg[1160]  ( .D(swire[138]), .CLK(clk), .RST(rst), .Q(sreg[1160])
         );
  DFF \sreg_reg[1161]  ( .D(swire[139]), .CLK(clk), .RST(rst), .Q(sreg[1161])
         );
  DFF \sreg_reg[1162]  ( .D(swire[140]), .CLK(clk), .RST(rst), .Q(sreg[1162])
         );
  DFF \sreg_reg[1163]  ( .D(swire[141]), .CLK(clk), .RST(rst), .Q(sreg[1163])
         );
  DFF \sreg_reg[1164]  ( .D(swire[142]), .CLK(clk), .RST(rst), .Q(sreg[1164])
         );
  DFF \sreg_reg[1165]  ( .D(swire[143]), .CLK(clk), .RST(rst), .Q(sreg[1165])
         );
  DFF \sreg_reg[1166]  ( .D(swire[144]), .CLK(clk), .RST(rst), .Q(sreg[1166])
         );
  DFF \sreg_reg[1167]  ( .D(swire[145]), .CLK(clk), .RST(rst), .Q(sreg[1167])
         );
  DFF \sreg_reg[1168]  ( .D(swire[146]), .CLK(clk), .RST(rst), .Q(sreg[1168])
         );
  DFF \sreg_reg[1169]  ( .D(swire[147]), .CLK(clk), .RST(rst), .Q(sreg[1169])
         );
  DFF \sreg_reg[1170]  ( .D(swire[148]), .CLK(clk), .RST(rst), .Q(sreg[1170])
         );
  DFF \sreg_reg[1171]  ( .D(swire[149]), .CLK(clk), .RST(rst), .Q(sreg[1171])
         );
  DFF \sreg_reg[1172]  ( .D(swire[150]), .CLK(clk), .RST(rst), .Q(sreg[1172])
         );
  DFF \sreg_reg[1173]  ( .D(swire[151]), .CLK(clk), .RST(rst), .Q(sreg[1173])
         );
  DFF \sreg_reg[1174]  ( .D(swire[152]), .CLK(clk), .RST(rst), .Q(sreg[1174])
         );
  DFF \sreg_reg[1175]  ( .D(swire[153]), .CLK(clk), .RST(rst), .Q(sreg[1175])
         );
  DFF \sreg_reg[1176]  ( .D(swire[154]), .CLK(clk), .RST(rst), .Q(sreg[1176])
         );
  DFF \sreg_reg[1177]  ( .D(swire[155]), .CLK(clk), .RST(rst), .Q(sreg[1177])
         );
  DFF \sreg_reg[1178]  ( .D(swire[156]), .CLK(clk), .RST(rst), .Q(sreg[1178])
         );
  DFF \sreg_reg[1179]  ( .D(swire[157]), .CLK(clk), .RST(rst), .Q(sreg[1179])
         );
  DFF \sreg_reg[1180]  ( .D(swire[158]), .CLK(clk), .RST(rst), .Q(sreg[1180])
         );
  DFF \sreg_reg[1181]  ( .D(swire[159]), .CLK(clk), .RST(rst), .Q(sreg[1181])
         );
  DFF \sreg_reg[1182]  ( .D(swire[160]), .CLK(clk), .RST(rst), .Q(sreg[1182])
         );
  DFF \sreg_reg[1183]  ( .D(swire[161]), .CLK(clk), .RST(rst), .Q(sreg[1183])
         );
  DFF \sreg_reg[1184]  ( .D(swire[162]), .CLK(clk), .RST(rst), .Q(sreg[1184])
         );
  DFF \sreg_reg[1185]  ( .D(swire[163]), .CLK(clk), .RST(rst), .Q(sreg[1185])
         );
  DFF \sreg_reg[1186]  ( .D(swire[164]), .CLK(clk), .RST(rst), .Q(sreg[1186])
         );
  DFF \sreg_reg[1187]  ( .D(swire[165]), .CLK(clk), .RST(rst), .Q(sreg[1187])
         );
  DFF \sreg_reg[1188]  ( .D(swire[166]), .CLK(clk), .RST(rst), .Q(sreg[1188])
         );
  DFF \sreg_reg[1189]  ( .D(swire[167]), .CLK(clk), .RST(rst), .Q(sreg[1189])
         );
  DFF \sreg_reg[1190]  ( .D(swire[168]), .CLK(clk), .RST(rst), .Q(sreg[1190])
         );
  DFF \sreg_reg[1191]  ( .D(swire[169]), .CLK(clk), .RST(rst), .Q(sreg[1191])
         );
  DFF \sreg_reg[1192]  ( .D(swire[170]), .CLK(clk), .RST(rst), .Q(sreg[1192])
         );
  DFF \sreg_reg[1193]  ( .D(swire[171]), .CLK(clk), .RST(rst), .Q(sreg[1193])
         );
  DFF \sreg_reg[1194]  ( .D(swire[172]), .CLK(clk), .RST(rst), .Q(sreg[1194])
         );
  DFF \sreg_reg[1195]  ( .D(swire[173]), .CLK(clk), .RST(rst), .Q(sreg[1195])
         );
  DFF \sreg_reg[1196]  ( .D(swire[174]), .CLK(clk), .RST(rst), .Q(sreg[1196])
         );
  DFF \sreg_reg[1197]  ( .D(swire[175]), .CLK(clk), .RST(rst), .Q(sreg[1197])
         );
  DFF \sreg_reg[1198]  ( .D(swire[176]), .CLK(clk), .RST(rst), .Q(sreg[1198])
         );
  DFF \sreg_reg[1199]  ( .D(swire[177]), .CLK(clk), .RST(rst), .Q(sreg[1199])
         );
  DFF \sreg_reg[1200]  ( .D(swire[178]), .CLK(clk), .RST(rst), .Q(sreg[1200])
         );
  DFF \sreg_reg[1201]  ( .D(swire[179]), .CLK(clk), .RST(rst), .Q(sreg[1201])
         );
  DFF \sreg_reg[1202]  ( .D(swire[180]), .CLK(clk), .RST(rst), .Q(sreg[1202])
         );
  DFF \sreg_reg[1203]  ( .D(swire[181]), .CLK(clk), .RST(rst), .Q(sreg[1203])
         );
  DFF \sreg_reg[1204]  ( .D(swire[182]), .CLK(clk), .RST(rst), .Q(sreg[1204])
         );
  DFF \sreg_reg[1205]  ( .D(swire[183]), .CLK(clk), .RST(rst), .Q(sreg[1205])
         );
  DFF \sreg_reg[1206]  ( .D(swire[184]), .CLK(clk), .RST(rst), .Q(sreg[1206])
         );
  DFF \sreg_reg[1207]  ( .D(swire[185]), .CLK(clk), .RST(rst), .Q(sreg[1207])
         );
  DFF \sreg_reg[1208]  ( .D(swire[186]), .CLK(clk), .RST(rst), .Q(sreg[1208])
         );
  DFF \sreg_reg[1209]  ( .D(swire[187]), .CLK(clk), .RST(rst), .Q(sreg[1209])
         );
  DFF \sreg_reg[1210]  ( .D(swire[188]), .CLK(clk), .RST(rst), .Q(sreg[1210])
         );
  DFF \sreg_reg[1211]  ( .D(swire[189]), .CLK(clk), .RST(rst), .Q(sreg[1211])
         );
  DFF \sreg_reg[1212]  ( .D(swire[190]), .CLK(clk), .RST(rst), .Q(sreg[1212])
         );
  DFF \sreg_reg[1213]  ( .D(swire[191]), .CLK(clk), .RST(rst), .Q(sreg[1213])
         );
  DFF \sreg_reg[1214]  ( .D(swire[192]), .CLK(clk), .RST(rst), .Q(sreg[1214])
         );
  DFF \sreg_reg[1215]  ( .D(swire[193]), .CLK(clk), .RST(rst), .Q(sreg[1215])
         );
  DFF \sreg_reg[1216]  ( .D(swire[194]), .CLK(clk), .RST(rst), .Q(sreg[1216])
         );
  DFF \sreg_reg[1217]  ( .D(swire[195]), .CLK(clk), .RST(rst), .Q(sreg[1217])
         );
  DFF \sreg_reg[1218]  ( .D(swire[196]), .CLK(clk), .RST(rst), .Q(sreg[1218])
         );
  DFF \sreg_reg[1219]  ( .D(swire[197]), .CLK(clk), .RST(rst), .Q(sreg[1219])
         );
  DFF \sreg_reg[1220]  ( .D(swire[198]), .CLK(clk), .RST(rst), .Q(sreg[1220])
         );
  DFF \sreg_reg[1221]  ( .D(swire[199]), .CLK(clk), .RST(rst), .Q(sreg[1221])
         );
  DFF \sreg_reg[1222]  ( .D(swire[200]), .CLK(clk), .RST(rst), .Q(sreg[1222])
         );
  DFF \sreg_reg[1223]  ( .D(swire[201]), .CLK(clk), .RST(rst), .Q(sreg[1223])
         );
  DFF \sreg_reg[1224]  ( .D(swire[202]), .CLK(clk), .RST(rst), .Q(sreg[1224])
         );
  DFF \sreg_reg[1225]  ( .D(swire[203]), .CLK(clk), .RST(rst), .Q(sreg[1225])
         );
  DFF \sreg_reg[1226]  ( .D(swire[204]), .CLK(clk), .RST(rst), .Q(sreg[1226])
         );
  DFF \sreg_reg[1227]  ( .D(swire[205]), .CLK(clk), .RST(rst), .Q(sreg[1227])
         );
  DFF \sreg_reg[1228]  ( .D(swire[206]), .CLK(clk), .RST(rst), .Q(sreg[1228])
         );
  DFF \sreg_reg[1229]  ( .D(swire[207]), .CLK(clk), .RST(rst), .Q(sreg[1229])
         );
  DFF \sreg_reg[1230]  ( .D(swire[208]), .CLK(clk), .RST(rst), .Q(sreg[1230])
         );
  DFF \sreg_reg[1231]  ( .D(swire[209]), .CLK(clk), .RST(rst), .Q(sreg[1231])
         );
  DFF \sreg_reg[1232]  ( .D(swire[210]), .CLK(clk), .RST(rst), .Q(sreg[1232])
         );
  DFF \sreg_reg[1233]  ( .D(swire[211]), .CLK(clk), .RST(rst), .Q(sreg[1233])
         );
  DFF \sreg_reg[1234]  ( .D(swire[212]), .CLK(clk), .RST(rst), .Q(sreg[1234])
         );
  DFF \sreg_reg[1235]  ( .D(swire[213]), .CLK(clk), .RST(rst), .Q(sreg[1235])
         );
  DFF \sreg_reg[1236]  ( .D(swire[214]), .CLK(clk), .RST(rst), .Q(sreg[1236])
         );
  DFF \sreg_reg[1237]  ( .D(swire[215]), .CLK(clk), .RST(rst), .Q(sreg[1237])
         );
  DFF \sreg_reg[1238]  ( .D(swire[216]), .CLK(clk), .RST(rst), .Q(sreg[1238])
         );
  DFF \sreg_reg[1239]  ( .D(swire[217]), .CLK(clk), .RST(rst), .Q(sreg[1239])
         );
  DFF \sreg_reg[1240]  ( .D(swire[218]), .CLK(clk), .RST(rst), .Q(sreg[1240])
         );
  DFF \sreg_reg[1241]  ( .D(swire[219]), .CLK(clk), .RST(rst), .Q(sreg[1241])
         );
  DFF \sreg_reg[1242]  ( .D(swire[220]), .CLK(clk), .RST(rst), .Q(sreg[1242])
         );
  DFF \sreg_reg[1243]  ( .D(swire[221]), .CLK(clk), .RST(rst), .Q(sreg[1243])
         );
  DFF \sreg_reg[1244]  ( .D(swire[222]), .CLK(clk), .RST(rst), .Q(sreg[1244])
         );
  DFF \sreg_reg[1245]  ( .D(swire[223]), .CLK(clk), .RST(rst), .Q(sreg[1245])
         );
  DFF \sreg_reg[1246]  ( .D(swire[224]), .CLK(clk), .RST(rst), .Q(sreg[1246])
         );
  DFF \sreg_reg[1247]  ( .D(swire[225]), .CLK(clk), .RST(rst), .Q(sreg[1247])
         );
  DFF \sreg_reg[1248]  ( .D(swire[226]), .CLK(clk), .RST(rst), .Q(sreg[1248])
         );
  DFF \sreg_reg[1249]  ( .D(swire[227]), .CLK(clk), .RST(rst), .Q(sreg[1249])
         );
  DFF \sreg_reg[1250]  ( .D(swire[228]), .CLK(clk), .RST(rst), .Q(sreg[1250])
         );
  DFF \sreg_reg[1251]  ( .D(swire[229]), .CLK(clk), .RST(rst), .Q(sreg[1251])
         );
  DFF \sreg_reg[1252]  ( .D(swire[230]), .CLK(clk), .RST(rst), .Q(sreg[1252])
         );
  DFF \sreg_reg[1253]  ( .D(swire[231]), .CLK(clk), .RST(rst), .Q(sreg[1253])
         );
  DFF \sreg_reg[1254]  ( .D(swire[232]), .CLK(clk), .RST(rst), .Q(sreg[1254])
         );
  DFF \sreg_reg[1255]  ( .D(swire[233]), .CLK(clk), .RST(rst), .Q(sreg[1255])
         );
  DFF \sreg_reg[1256]  ( .D(swire[234]), .CLK(clk), .RST(rst), .Q(sreg[1256])
         );
  DFF \sreg_reg[1257]  ( .D(swire[235]), .CLK(clk), .RST(rst), .Q(sreg[1257])
         );
  DFF \sreg_reg[1258]  ( .D(swire[236]), .CLK(clk), .RST(rst), .Q(sreg[1258])
         );
  DFF \sreg_reg[1259]  ( .D(swire[237]), .CLK(clk), .RST(rst), .Q(sreg[1259])
         );
  DFF \sreg_reg[1260]  ( .D(swire[238]), .CLK(clk), .RST(rst), .Q(sreg[1260])
         );
  DFF \sreg_reg[1261]  ( .D(swire[239]), .CLK(clk), .RST(rst), .Q(sreg[1261])
         );
  DFF \sreg_reg[1262]  ( .D(swire[240]), .CLK(clk), .RST(rst), .Q(sreg[1262])
         );
  DFF \sreg_reg[1263]  ( .D(swire[241]), .CLK(clk), .RST(rst), .Q(sreg[1263])
         );
  DFF \sreg_reg[1264]  ( .D(swire[242]), .CLK(clk), .RST(rst), .Q(sreg[1264])
         );
  DFF \sreg_reg[1265]  ( .D(swire[243]), .CLK(clk), .RST(rst), .Q(sreg[1265])
         );
  DFF \sreg_reg[1266]  ( .D(swire[244]), .CLK(clk), .RST(rst), .Q(sreg[1266])
         );
  DFF \sreg_reg[1267]  ( .D(swire[245]), .CLK(clk), .RST(rst), .Q(sreg[1267])
         );
  DFF \sreg_reg[1268]  ( .D(swire[246]), .CLK(clk), .RST(rst), .Q(sreg[1268])
         );
  DFF \sreg_reg[1269]  ( .D(swire[247]), .CLK(clk), .RST(rst), .Q(sreg[1269])
         );
  DFF \sreg_reg[1270]  ( .D(swire[248]), .CLK(clk), .RST(rst), .Q(sreg[1270])
         );
  DFF \sreg_reg[1271]  ( .D(swire[249]), .CLK(clk), .RST(rst), .Q(sreg[1271])
         );
  DFF \sreg_reg[1272]  ( .D(swire[250]), .CLK(clk), .RST(rst), .Q(sreg[1272])
         );
  DFF \sreg_reg[1273]  ( .D(swire[251]), .CLK(clk), .RST(rst), .Q(sreg[1273])
         );
  DFF \sreg_reg[1274]  ( .D(swire[252]), .CLK(clk), .RST(rst), .Q(sreg[1274])
         );
  DFF \sreg_reg[1275]  ( .D(swire[253]), .CLK(clk), .RST(rst), .Q(sreg[1275])
         );
  DFF \sreg_reg[1276]  ( .D(swire[254]), .CLK(clk), .RST(rst), .Q(sreg[1276])
         );
  DFF \sreg_reg[1277]  ( .D(swire[255]), .CLK(clk), .RST(rst), .Q(sreg[1277])
         );
  DFF \sreg_reg[1278]  ( .D(swire[256]), .CLK(clk), .RST(rst), .Q(sreg[1278])
         );
  DFF \sreg_reg[1279]  ( .D(swire[257]), .CLK(clk), .RST(rst), .Q(sreg[1279])
         );
  DFF \sreg_reg[1280]  ( .D(swire[258]), .CLK(clk), .RST(rst), .Q(sreg[1280])
         );
  DFF \sreg_reg[1281]  ( .D(swire[259]), .CLK(clk), .RST(rst), .Q(sreg[1281])
         );
  DFF \sreg_reg[1282]  ( .D(swire[260]), .CLK(clk), .RST(rst), .Q(sreg[1282])
         );
  DFF \sreg_reg[1283]  ( .D(swire[261]), .CLK(clk), .RST(rst), .Q(sreg[1283])
         );
  DFF \sreg_reg[1284]  ( .D(swire[262]), .CLK(clk), .RST(rst), .Q(sreg[1284])
         );
  DFF \sreg_reg[1285]  ( .D(swire[263]), .CLK(clk), .RST(rst), .Q(sreg[1285])
         );
  DFF \sreg_reg[1286]  ( .D(swire[264]), .CLK(clk), .RST(rst), .Q(sreg[1286])
         );
  DFF \sreg_reg[1287]  ( .D(swire[265]), .CLK(clk), .RST(rst), .Q(sreg[1287])
         );
  DFF \sreg_reg[1288]  ( .D(swire[266]), .CLK(clk), .RST(rst), .Q(sreg[1288])
         );
  DFF \sreg_reg[1289]  ( .D(swire[267]), .CLK(clk), .RST(rst), .Q(sreg[1289])
         );
  DFF \sreg_reg[1290]  ( .D(swire[268]), .CLK(clk), .RST(rst), .Q(sreg[1290])
         );
  DFF \sreg_reg[1291]  ( .D(swire[269]), .CLK(clk), .RST(rst), .Q(sreg[1291])
         );
  DFF \sreg_reg[1292]  ( .D(swire[270]), .CLK(clk), .RST(rst), .Q(sreg[1292])
         );
  DFF \sreg_reg[1293]  ( .D(swire[271]), .CLK(clk), .RST(rst), .Q(sreg[1293])
         );
  DFF \sreg_reg[1294]  ( .D(swire[272]), .CLK(clk), .RST(rst), .Q(sreg[1294])
         );
  DFF \sreg_reg[1295]  ( .D(swire[273]), .CLK(clk), .RST(rst), .Q(sreg[1295])
         );
  DFF \sreg_reg[1296]  ( .D(swire[274]), .CLK(clk), .RST(rst), .Q(sreg[1296])
         );
  DFF \sreg_reg[1297]  ( .D(swire[275]), .CLK(clk), .RST(rst), .Q(sreg[1297])
         );
  DFF \sreg_reg[1298]  ( .D(swire[276]), .CLK(clk), .RST(rst), .Q(sreg[1298])
         );
  DFF \sreg_reg[1299]  ( .D(swire[277]), .CLK(clk), .RST(rst), .Q(sreg[1299])
         );
  DFF \sreg_reg[1300]  ( .D(swire[278]), .CLK(clk), .RST(rst), .Q(sreg[1300])
         );
  DFF \sreg_reg[1301]  ( .D(swire[279]), .CLK(clk), .RST(rst), .Q(sreg[1301])
         );
  DFF \sreg_reg[1302]  ( .D(swire[280]), .CLK(clk), .RST(rst), .Q(sreg[1302])
         );
  DFF \sreg_reg[1303]  ( .D(swire[281]), .CLK(clk), .RST(rst), .Q(sreg[1303])
         );
  DFF \sreg_reg[1304]  ( .D(swire[282]), .CLK(clk), .RST(rst), .Q(sreg[1304])
         );
  DFF \sreg_reg[1305]  ( .D(swire[283]), .CLK(clk), .RST(rst), .Q(sreg[1305])
         );
  DFF \sreg_reg[1306]  ( .D(swire[284]), .CLK(clk), .RST(rst), .Q(sreg[1306])
         );
  DFF \sreg_reg[1307]  ( .D(swire[285]), .CLK(clk), .RST(rst), .Q(sreg[1307])
         );
  DFF \sreg_reg[1308]  ( .D(swire[286]), .CLK(clk), .RST(rst), .Q(sreg[1308])
         );
  DFF \sreg_reg[1309]  ( .D(swire[287]), .CLK(clk), .RST(rst), .Q(sreg[1309])
         );
  DFF \sreg_reg[1310]  ( .D(swire[288]), .CLK(clk), .RST(rst), .Q(sreg[1310])
         );
  DFF \sreg_reg[1311]  ( .D(swire[289]), .CLK(clk), .RST(rst), .Q(sreg[1311])
         );
  DFF \sreg_reg[1312]  ( .D(swire[290]), .CLK(clk), .RST(rst), .Q(sreg[1312])
         );
  DFF \sreg_reg[1313]  ( .D(swire[291]), .CLK(clk), .RST(rst), .Q(sreg[1313])
         );
  DFF \sreg_reg[1314]  ( .D(swire[292]), .CLK(clk), .RST(rst), .Q(sreg[1314])
         );
  DFF \sreg_reg[1315]  ( .D(swire[293]), .CLK(clk), .RST(rst), .Q(sreg[1315])
         );
  DFF \sreg_reg[1316]  ( .D(swire[294]), .CLK(clk), .RST(rst), .Q(sreg[1316])
         );
  DFF \sreg_reg[1317]  ( .D(swire[295]), .CLK(clk), .RST(rst), .Q(sreg[1317])
         );
  DFF \sreg_reg[1318]  ( .D(swire[296]), .CLK(clk), .RST(rst), .Q(sreg[1318])
         );
  DFF \sreg_reg[1319]  ( .D(swire[297]), .CLK(clk), .RST(rst), .Q(sreg[1319])
         );
  DFF \sreg_reg[1320]  ( .D(swire[298]), .CLK(clk), .RST(rst), .Q(sreg[1320])
         );
  DFF \sreg_reg[1321]  ( .D(swire[299]), .CLK(clk), .RST(rst), .Q(sreg[1321])
         );
  DFF \sreg_reg[1322]  ( .D(swire[300]), .CLK(clk), .RST(rst), .Q(sreg[1322])
         );
  DFF \sreg_reg[1323]  ( .D(swire[301]), .CLK(clk), .RST(rst), .Q(sreg[1323])
         );
  DFF \sreg_reg[1324]  ( .D(swire[302]), .CLK(clk), .RST(rst), .Q(sreg[1324])
         );
  DFF \sreg_reg[1325]  ( .D(swire[303]), .CLK(clk), .RST(rst), .Q(sreg[1325])
         );
  DFF \sreg_reg[1326]  ( .D(swire[304]), .CLK(clk), .RST(rst), .Q(sreg[1326])
         );
  DFF \sreg_reg[1327]  ( .D(swire[305]), .CLK(clk), .RST(rst), .Q(sreg[1327])
         );
  DFF \sreg_reg[1328]  ( .D(swire[306]), .CLK(clk), .RST(rst), .Q(sreg[1328])
         );
  DFF \sreg_reg[1329]  ( .D(swire[307]), .CLK(clk), .RST(rst), .Q(sreg[1329])
         );
  DFF \sreg_reg[1330]  ( .D(swire[308]), .CLK(clk), .RST(rst), .Q(sreg[1330])
         );
  DFF \sreg_reg[1331]  ( .D(swire[309]), .CLK(clk), .RST(rst), .Q(sreg[1331])
         );
  DFF \sreg_reg[1332]  ( .D(swire[310]), .CLK(clk), .RST(rst), .Q(sreg[1332])
         );
  DFF \sreg_reg[1333]  ( .D(swire[311]), .CLK(clk), .RST(rst), .Q(sreg[1333])
         );
  DFF \sreg_reg[1334]  ( .D(swire[312]), .CLK(clk), .RST(rst), .Q(sreg[1334])
         );
  DFF \sreg_reg[1335]  ( .D(swire[313]), .CLK(clk), .RST(rst), .Q(sreg[1335])
         );
  DFF \sreg_reg[1336]  ( .D(swire[314]), .CLK(clk), .RST(rst), .Q(sreg[1336])
         );
  DFF \sreg_reg[1337]  ( .D(swire[315]), .CLK(clk), .RST(rst), .Q(sreg[1337])
         );
  DFF \sreg_reg[1338]  ( .D(swire[316]), .CLK(clk), .RST(rst), .Q(sreg[1338])
         );
  DFF \sreg_reg[1339]  ( .D(swire[317]), .CLK(clk), .RST(rst), .Q(sreg[1339])
         );
  DFF \sreg_reg[1340]  ( .D(swire[318]), .CLK(clk), .RST(rst), .Q(sreg[1340])
         );
  DFF \sreg_reg[1341]  ( .D(swire[319]), .CLK(clk), .RST(rst), .Q(sreg[1341])
         );
  DFF \sreg_reg[1342]  ( .D(swire[320]), .CLK(clk), .RST(rst), .Q(sreg[1342])
         );
  DFF \sreg_reg[1343]  ( .D(swire[321]), .CLK(clk), .RST(rst), .Q(sreg[1343])
         );
  DFF \sreg_reg[1344]  ( .D(swire[322]), .CLK(clk), .RST(rst), .Q(sreg[1344])
         );
  DFF \sreg_reg[1345]  ( .D(swire[323]), .CLK(clk), .RST(rst), .Q(sreg[1345])
         );
  DFF \sreg_reg[1346]  ( .D(swire[324]), .CLK(clk), .RST(rst), .Q(sreg[1346])
         );
  DFF \sreg_reg[1347]  ( .D(swire[325]), .CLK(clk), .RST(rst), .Q(sreg[1347])
         );
  DFF \sreg_reg[1348]  ( .D(swire[326]), .CLK(clk), .RST(rst), .Q(sreg[1348])
         );
  DFF \sreg_reg[1349]  ( .D(swire[327]), .CLK(clk), .RST(rst), .Q(sreg[1349])
         );
  DFF \sreg_reg[1350]  ( .D(swire[328]), .CLK(clk), .RST(rst), .Q(sreg[1350])
         );
  DFF \sreg_reg[1351]  ( .D(swire[329]), .CLK(clk), .RST(rst), .Q(sreg[1351])
         );
  DFF \sreg_reg[1352]  ( .D(swire[330]), .CLK(clk), .RST(rst), .Q(sreg[1352])
         );
  DFF \sreg_reg[1353]  ( .D(swire[331]), .CLK(clk), .RST(rst), .Q(sreg[1353])
         );
  DFF \sreg_reg[1354]  ( .D(swire[332]), .CLK(clk), .RST(rst), .Q(sreg[1354])
         );
  DFF \sreg_reg[1355]  ( .D(swire[333]), .CLK(clk), .RST(rst), .Q(sreg[1355])
         );
  DFF \sreg_reg[1356]  ( .D(swire[334]), .CLK(clk), .RST(rst), .Q(sreg[1356])
         );
  DFF \sreg_reg[1357]  ( .D(swire[335]), .CLK(clk), .RST(rst), .Q(sreg[1357])
         );
  DFF \sreg_reg[1358]  ( .D(swire[336]), .CLK(clk), .RST(rst), .Q(sreg[1358])
         );
  DFF \sreg_reg[1359]  ( .D(swire[337]), .CLK(clk), .RST(rst), .Q(sreg[1359])
         );
  DFF \sreg_reg[1360]  ( .D(swire[338]), .CLK(clk), .RST(rst), .Q(sreg[1360])
         );
  DFF \sreg_reg[1361]  ( .D(swire[339]), .CLK(clk), .RST(rst), .Q(sreg[1361])
         );
  DFF \sreg_reg[1362]  ( .D(swire[340]), .CLK(clk), .RST(rst), .Q(sreg[1362])
         );
  DFF \sreg_reg[1363]  ( .D(swire[341]), .CLK(clk), .RST(rst), .Q(sreg[1363])
         );
  DFF \sreg_reg[1364]  ( .D(swire[342]), .CLK(clk), .RST(rst), .Q(sreg[1364])
         );
  DFF \sreg_reg[1365]  ( .D(swire[343]), .CLK(clk), .RST(rst), .Q(sreg[1365])
         );
  DFF \sreg_reg[1366]  ( .D(swire[344]), .CLK(clk), .RST(rst), .Q(sreg[1366])
         );
  DFF \sreg_reg[1367]  ( .D(swire[345]), .CLK(clk), .RST(rst), .Q(sreg[1367])
         );
  DFF \sreg_reg[1368]  ( .D(swire[346]), .CLK(clk), .RST(rst), .Q(sreg[1368])
         );
  DFF \sreg_reg[1369]  ( .D(swire[347]), .CLK(clk), .RST(rst), .Q(sreg[1369])
         );
  DFF \sreg_reg[1370]  ( .D(swire[348]), .CLK(clk), .RST(rst), .Q(sreg[1370])
         );
  DFF \sreg_reg[1371]  ( .D(swire[349]), .CLK(clk), .RST(rst), .Q(sreg[1371])
         );
  DFF \sreg_reg[1372]  ( .D(swire[350]), .CLK(clk), .RST(rst), .Q(sreg[1372])
         );
  DFF \sreg_reg[1373]  ( .D(swire[351]), .CLK(clk), .RST(rst), .Q(sreg[1373])
         );
  DFF \sreg_reg[1374]  ( .D(swire[352]), .CLK(clk), .RST(rst), .Q(sreg[1374])
         );
  DFF \sreg_reg[1375]  ( .D(swire[353]), .CLK(clk), .RST(rst), .Q(sreg[1375])
         );
  DFF \sreg_reg[1376]  ( .D(swire[354]), .CLK(clk), .RST(rst), .Q(sreg[1376])
         );
  DFF \sreg_reg[1377]  ( .D(swire[355]), .CLK(clk), .RST(rst), .Q(sreg[1377])
         );
  DFF \sreg_reg[1378]  ( .D(swire[356]), .CLK(clk), .RST(rst), .Q(sreg[1378])
         );
  DFF \sreg_reg[1379]  ( .D(swire[357]), .CLK(clk), .RST(rst), .Q(sreg[1379])
         );
  DFF \sreg_reg[1380]  ( .D(swire[358]), .CLK(clk), .RST(rst), .Q(sreg[1380])
         );
  DFF \sreg_reg[1381]  ( .D(swire[359]), .CLK(clk), .RST(rst), .Q(sreg[1381])
         );
  DFF \sreg_reg[1382]  ( .D(swire[360]), .CLK(clk), .RST(rst), .Q(sreg[1382])
         );
  DFF \sreg_reg[1383]  ( .D(swire[361]), .CLK(clk), .RST(rst), .Q(sreg[1383])
         );
  DFF \sreg_reg[1384]  ( .D(swire[362]), .CLK(clk), .RST(rst), .Q(sreg[1384])
         );
  DFF \sreg_reg[1385]  ( .D(swire[363]), .CLK(clk), .RST(rst), .Q(sreg[1385])
         );
  DFF \sreg_reg[1386]  ( .D(swire[364]), .CLK(clk), .RST(rst), .Q(sreg[1386])
         );
  DFF \sreg_reg[1387]  ( .D(swire[365]), .CLK(clk), .RST(rst), .Q(sreg[1387])
         );
  DFF \sreg_reg[1388]  ( .D(swire[366]), .CLK(clk), .RST(rst), .Q(sreg[1388])
         );
  DFF \sreg_reg[1389]  ( .D(swire[367]), .CLK(clk), .RST(rst), .Q(sreg[1389])
         );
  DFF \sreg_reg[1390]  ( .D(swire[368]), .CLK(clk), .RST(rst), .Q(sreg[1390])
         );
  DFF \sreg_reg[1391]  ( .D(swire[369]), .CLK(clk), .RST(rst), .Q(sreg[1391])
         );
  DFF \sreg_reg[1392]  ( .D(swire[370]), .CLK(clk), .RST(rst), .Q(sreg[1392])
         );
  DFF \sreg_reg[1393]  ( .D(swire[371]), .CLK(clk), .RST(rst), .Q(sreg[1393])
         );
  DFF \sreg_reg[1394]  ( .D(swire[372]), .CLK(clk), .RST(rst), .Q(sreg[1394])
         );
  DFF \sreg_reg[1395]  ( .D(swire[373]), .CLK(clk), .RST(rst), .Q(sreg[1395])
         );
  DFF \sreg_reg[1396]  ( .D(swire[374]), .CLK(clk), .RST(rst), .Q(sreg[1396])
         );
  DFF \sreg_reg[1397]  ( .D(swire[375]), .CLK(clk), .RST(rst), .Q(sreg[1397])
         );
  DFF \sreg_reg[1398]  ( .D(swire[376]), .CLK(clk), .RST(rst), .Q(sreg[1398])
         );
  DFF \sreg_reg[1399]  ( .D(swire[377]), .CLK(clk), .RST(rst), .Q(sreg[1399])
         );
  DFF \sreg_reg[1400]  ( .D(swire[378]), .CLK(clk), .RST(rst), .Q(sreg[1400])
         );
  DFF \sreg_reg[1401]  ( .D(swire[379]), .CLK(clk), .RST(rst), .Q(sreg[1401])
         );
  DFF \sreg_reg[1402]  ( .D(swire[380]), .CLK(clk), .RST(rst), .Q(sreg[1402])
         );
  DFF \sreg_reg[1403]  ( .D(swire[381]), .CLK(clk), .RST(rst), .Q(sreg[1403])
         );
  DFF \sreg_reg[1404]  ( .D(swire[382]), .CLK(clk), .RST(rst), .Q(sreg[1404])
         );
  DFF \sreg_reg[1405]  ( .D(swire[383]), .CLK(clk), .RST(rst), .Q(sreg[1405])
         );
  DFF \sreg_reg[1406]  ( .D(swire[384]), .CLK(clk), .RST(rst), .Q(sreg[1406])
         );
  DFF \sreg_reg[1407]  ( .D(swire[385]), .CLK(clk), .RST(rst), .Q(sreg[1407])
         );
  DFF \sreg_reg[1408]  ( .D(swire[386]), .CLK(clk), .RST(rst), .Q(sreg[1408])
         );
  DFF \sreg_reg[1409]  ( .D(swire[387]), .CLK(clk), .RST(rst), .Q(sreg[1409])
         );
  DFF \sreg_reg[1410]  ( .D(swire[388]), .CLK(clk), .RST(rst), .Q(sreg[1410])
         );
  DFF \sreg_reg[1411]  ( .D(swire[389]), .CLK(clk), .RST(rst), .Q(sreg[1411])
         );
  DFF \sreg_reg[1412]  ( .D(swire[390]), .CLK(clk), .RST(rst), .Q(sreg[1412])
         );
  DFF \sreg_reg[1413]  ( .D(swire[391]), .CLK(clk), .RST(rst), .Q(sreg[1413])
         );
  DFF \sreg_reg[1414]  ( .D(swire[392]), .CLK(clk), .RST(rst), .Q(sreg[1414])
         );
  DFF \sreg_reg[1415]  ( .D(swire[393]), .CLK(clk), .RST(rst), .Q(sreg[1415])
         );
  DFF \sreg_reg[1416]  ( .D(swire[394]), .CLK(clk), .RST(rst), .Q(sreg[1416])
         );
  DFF \sreg_reg[1417]  ( .D(swire[395]), .CLK(clk), .RST(rst), .Q(sreg[1417])
         );
  DFF \sreg_reg[1418]  ( .D(swire[396]), .CLK(clk), .RST(rst), .Q(sreg[1418])
         );
  DFF \sreg_reg[1419]  ( .D(swire[397]), .CLK(clk), .RST(rst), .Q(sreg[1419])
         );
  DFF \sreg_reg[1420]  ( .D(swire[398]), .CLK(clk), .RST(rst), .Q(sreg[1420])
         );
  DFF \sreg_reg[1421]  ( .D(swire[399]), .CLK(clk), .RST(rst), .Q(sreg[1421])
         );
  DFF \sreg_reg[1422]  ( .D(swire[400]), .CLK(clk), .RST(rst), .Q(sreg[1422])
         );
  DFF \sreg_reg[1423]  ( .D(swire[401]), .CLK(clk), .RST(rst), .Q(sreg[1423])
         );
  DFF \sreg_reg[1424]  ( .D(swire[402]), .CLK(clk), .RST(rst), .Q(sreg[1424])
         );
  DFF \sreg_reg[1425]  ( .D(swire[403]), .CLK(clk), .RST(rst), .Q(sreg[1425])
         );
  DFF \sreg_reg[1426]  ( .D(swire[404]), .CLK(clk), .RST(rst), .Q(sreg[1426])
         );
  DFF \sreg_reg[1427]  ( .D(swire[405]), .CLK(clk), .RST(rst), .Q(sreg[1427])
         );
  DFF \sreg_reg[1428]  ( .D(swire[406]), .CLK(clk), .RST(rst), .Q(sreg[1428])
         );
  DFF \sreg_reg[1429]  ( .D(swire[407]), .CLK(clk), .RST(rst), .Q(sreg[1429])
         );
  DFF \sreg_reg[1430]  ( .D(swire[408]), .CLK(clk), .RST(rst), .Q(sreg[1430])
         );
  DFF \sreg_reg[1431]  ( .D(swire[409]), .CLK(clk), .RST(rst), .Q(sreg[1431])
         );
  DFF \sreg_reg[1432]  ( .D(swire[410]), .CLK(clk), .RST(rst), .Q(sreg[1432])
         );
  DFF \sreg_reg[1433]  ( .D(swire[411]), .CLK(clk), .RST(rst), .Q(sreg[1433])
         );
  DFF \sreg_reg[1434]  ( .D(swire[412]), .CLK(clk), .RST(rst), .Q(sreg[1434])
         );
  DFF \sreg_reg[1435]  ( .D(swire[413]), .CLK(clk), .RST(rst), .Q(sreg[1435])
         );
  DFF \sreg_reg[1436]  ( .D(swire[414]), .CLK(clk), .RST(rst), .Q(sreg[1436])
         );
  DFF \sreg_reg[1437]  ( .D(swire[415]), .CLK(clk), .RST(rst), .Q(sreg[1437])
         );
  DFF \sreg_reg[1438]  ( .D(swire[416]), .CLK(clk), .RST(rst), .Q(sreg[1438])
         );
  DFF \sreg_reg[1439]  ( .D(swire[417]), .CLK(clk), .RST(rst), .Q(sreg[1439])
         );
  DFF \sreg_reg[1440]  ( .D(swire[418]), .CLK(clk), .RST(rst), .Q(sreg[1440])
         );
  DFF \sreg_reg[1441]  ( .D(swire[419]), .CLK(clk), .RST(rst), .Q(sreg[1441])
         );
  DFF \sreg_reg[1442]  ( .D(swire[420]), .CLK(clk), .RST(rst), .Q(sreg[1442])
         );
  DFF \sreg_reg[1443]  ( .D(swire[421]), .CLK(clk), .RST(rst), .Q(sreg[1443])
         );
  DFF \sreg_reg[1444]  ( .D(swire[422]), .CLK(clk), .RST(rst), .Q(sreg[1444])
         );
  DFF \sreg_reg[1445]  ( .D(swire[423]), .CLK(clk), .RST(rst), .Q(sreg[1445])
         );
  DFF \sreg_reg[1446]  ( .D(swire[424]), .CLK(clk), .RST(rst), .Q(sreg[1446])
         );
  DFF \sreg_reg[1447]  ( .D(swire[425]), .CLK(clk), .RST(rst), .Q(sreg[1447])
         );
  DFF \sreg_reg[1448]  ( .D(swire[426]), .CLK(clk), .RST(rst), .Q(sreg[1448])
         );
  DFF \sreg_reg[1449]  ( .D(swire[427]), .CLK(clk), .RST(rst), .Q(sreg[1449])
         );
  DFF \sreg_reg[1450]  ( .D(swire[428]), .CLK(clk), .RST(rst), .Q(sreg[1450])
         );
  DFF \sreg_reg[1451]  ( .D(swire[429]), .CLK(clk), .RST(rst), .Q(sreg[1451])
         );
  DFF \sreg_reg[1452]  ( .D(swire[430]), .CLK(clk), .RST(rst), .Q(sreg[1452])
         );
  DFF \sreg_reg[1453]  ( .D(swire[431]), .CLK(clk), .RST(rst), .Q(sreg[1453])
         );
  DFF \sreg_reg[1454]  ( .D(swire[432]), .CLK(clk), .RST(rst), .Q(sreg[1454])
         );
  DFF \sreg_reg[1455]  ( .D(swire[433]), .CLK(clk), .RST(rst), .Q(sreg[1455])
         );
  DFF \sreg_reg[1456]  ( .D(swire[434]), .CLK(clk), .RST(rst), .Q(sreg[1456])
         );
  DFF \sreg_reg[1457]  ( .D(swire[435]), .CLK(clk), .RST(rst), .Q(sreg[1457])
         );
  DFF \sreg_reg[1458]  ( .D(swire[436]), .CLK(clk), .RST(rst), .Q(sreg[1458])
         );
  DFF \sreg_reg[1459]  ( .D(swire[437]), .CLK(clk), .RST(rst), .Q(sreg[1459])
         );
  DFF \sreg_reg[1460]  ( .D(swire[438]), .CLK(clk), .RST(rst), .Q(sreg[1460])
         );
  DFF \sreg_reg[1461]  ( .D(swire[439]), .CLK(clk), .RST(rst), .Q(sreg[1461])
         );
  DFF \sreg_reg[1462]  ( .D(swire[440]), .CLK(clk), .RST(rst), .Q(sreg[1462])
         );
  DFF \sreg_reg[1463]  ( .D(swire[441]), .CLK(clk), .RST(rst), .Q(sreg[1463])
         );
  DFF \sreg_reg[1464]  ( .D(swire[442]), .CLK(clk), .RST(rst), .Q(sreg[1464])
         );
  DFF \sreg_reg[1465]  ( .D(swire[443]), .CLK(clk), .RST(rst), .Q(sreg[1465])
         );
  DFF \sreg_reg[1466]  ( .D(swire[444]), .CLK(clk), .RST(rst), .Q(sreg[1466])
         );
  DFF \sreg_reg[1467]  ( .D(swire[445]), .CLK(clk), .RST(rst), .Q(sreg[1467])
         );
  DFF \sreg_reg[1468]  ( .D(swire[446]), .CLK(clk), .RST(rst), .Q(sreg[1468])
         );
  DFF \sreg_reg[1469]  ( .D(swire[447]), .CLK(clk), .RST(rst), .Q(sreg[1469])
         );
  DFF \sreg_reg[1470]  ( .D(swire[448]), .CLK(clk), .RST(rst), .Q(sreg[1470])
         );
  DFF \sreg_reg[1471]  ( .D(swire[449]), .CLK(clk), .RST(rst), .Q(sreg[1471])
         );
  DFF \sreg_reg[1472]  ( .D(swire[450]), .CLK(clk), .RST(rst), .Q(sreg[1472])
         );
  DFF \sreg_reg[1473]  ( .D(swire[451]), .CLK(clk), .RST(rst), .Q(sreg[1473])
         );
  DFF \sreg_reg[1474]  ( .D(swire[452]), .CLK(clk), .RST(rst), .Q(sreg[1474])
         );
  DFF \sreg_reg[1475]  ( .D(swire[453]), .CLK(clk), .RST(rst), .Q(sreg[1475])
         );
  DFF \sreg_reg[1476]  ( .D(swire[454]), .CLK(clk), .RST(rst), .Q(sreg[1476])
         );
  DFF \sreg_reg[1477]  ( .D(swire[455]), .CLK(clk), .RST(rst), .Q(sreg[1477])
         );
  DFF \sreg_reg[1478]  ( .D(swire[456]), .CLK(clk), .RST(rst), .Q(sreg[1478])
         );
  DFF \sreg_reg[1479]  ( .D(swire[457]), .CLK(clk), .RST(rst), .Q(sreg[1479])
         );
  DFF \sreg_reg[1480]  ( .D(swire[458]), .CLK(clk), .RST(rst), .Q(sreg[1480])
         );
  DFF \sreg_reg[1481]  ( .D(swire[459]), .CLK(clk), .RST(rst), .Q(sreg[1481])
         );
  DFF \sreg_reg[1482]  ( .D(swire[460]), .CLK(clk), .RST(rst), .Q(sreg[1482])
         );
  DFF \sreg_reg[1483]  ( .D(swire[461]), .CLK(clk), .RST(rst), .Q(sreg[1483])
         );
  DFF \sreg_reg[1484]  ( .D(swire[462]), .CLK(clk), .RST(rst), .Q(sreg[1484])
         );
  DFF \sreg_reg[1485]  ( .D(swire[463]), .CLK(clk), .RST(rst), .Q(sreg[1485])
         );
  DFF \sreg_reg[1486]  ( .D(swire[464]), .CLK(clk), .RST(rst), .Q(sreg[1486])
         );
  DFF \sreg_reg[1487]  ( .D(swire[465]), .CLK(clk), .RST(rst), .Q(sreg[1487])
         );
  DFF \sreg_reg[1488]  ( .D(swire[466]), .CLK(clk), .RST(rst), .Q(sreg[1488])
         );
  DFF \sreg_reg[1489]  ( .D(swire[467]), .CLK(clk), .RST(rst), .Q(sreg[1489])
         );
  DFF \sreg_reg[1490]  ( .D(swire[468]), .CLK(clk), .RST(rst), .Q(sreg[1490])
         );
  DFF \sreg_reg[1491]  ( .D(swire[469]), .CLK(clk), .RST(rst), .Q(sreg[1491])
         );
  DFF \sreg_reg[1492]  ( .D(swire[470]), .CLK(clk), .RST(rst), .Q(sreg[1492])
         );
  DFF \sreg_reg[1493]  ( .D(swire[471]), .CLK(clk), .RST(rst), .Q(sreg[1493])
         );
  DFF \sreg_reg[1494]  ( .D(swire[472]), .CLK(clk), .RST(rst), .Q(sreg[1494])
         );
  DFF \sreg_reg[1495]  ( .D(swire[473]), .CLK(clk), .RST(rst), .Q(sreg[1495])
         );
  DFF \sreg_reg[1496]  ( .D(swire[474]), .CLK(clk), .RST(rst), .Q(sreg[1496])
         );
  DFF \sreg_reg[1497]  ( .D(swire[475]), .CLK(clk), .RST(rst), .Q(sreg[1497])
         );
  DFF \sreg_reg[1498]  ( .D(swire[476]), .CLK(clk), .RST(rst), .Q(sreg[1498])
         );
  DFF \sreg_reg[1499]  ( .D(swire[477]), .CLK(clk), .RST(rst), .Q(sreg[1499])
         );
  DFF \sreg_reg[1500]  ( .D(swire[478]), .CLK(clk), .RST(rst), .Q(sreg[1500])
         );
  DFF \sreg_reg[1501]  ( .D(swire[479]), .CLK(clk), .RST(rst), .Q(sreg[1501])
         );
  DFF \sreg_reg[1502]  ( .D(swire[480]), .CLK(clk), .RST(rst), .Q(sreg[1502])
         );
  DFF \sreg_reg[1503]  ( .D(swire[481]), .CLK(clk), .RST(rst), .Q(sreg[1503])
         );
  DFF \sreg_reg[1504]  ( .D(swire[482]), .CLK(clk), .RST(rst), .Q(sreg[1504])
         );
  DFF \sreg_reg[1505]  ( .D(swire[483]), .CLK(clk), .RST(rst), .Q(sreg[1505])
         );
  DFF \sreg_reg[1506]  ( .D(swire[484]), .CLK(clk), .RST(rst), .Q(sreg[1506])
         );
  DFF \sreg_reg[1507]  ( .D(swire[485]), .CLK(clk), .RST(rst), .Q(sreg[1507])
         );
  DFF \sreg_reg[1508]  ( .D(swire[486]), .CLK(clk), .RST(rst), .Q(sreg[1508])
         );
  DFF \sreg_reg[1509]  ( .D(swire[487]), .CLK(clk), .RST(rst), .Q(sreg[1509])
         );
  DFF \sreg_reg[1510]  ( .D(swire[488]), .CLK(clk), .RST(rst), .Q(sreg[1510])
         );
  DFF \sreg_reg[1511]  ( .D(swire[489]), .CLK(clk), .RST(rst), .Q(sreg[1511])
         );
  DFF \sreg_reg[1512]  ( .D(swire[490]), .CLK(clk), .RST(rst), .Q(sreg[1512])
         );
  DFF \sreg_reg[1513]  ( .D(swire[491]), .CLK(clk), .RST(rst), .Q(sreg[1513])
         );
  DFF \sreg_reg[1514]  ( .D(swire[492]), .CLK(clk), .RST(rst), .Q(sreg[1514])
         );
  DFF \sreg_reg[1515]  ( .D(swire[493]), .CLK(clk), .RST(rst), .Q(sreg[1515])
         );
  DFF \sreg_reg[1516]  ( .D(swire[494]), .CLK(clk), .RST(rst), .Q(sreg[1516])
         );
  DFF \sreg_reg[1517]  ( .D(swire[495]), .CLK(clk), .RST(rst), .Q(sreg[1517])
         );
  DFF \sreg_reg[1518]  ( .D(swire[496]), .CLK(clk), .RST(rst), .Q(sreg[1518])
         );
  DFF \sreg_reg[1519]  ( .D(swire[497]), .CLK(clk), .RST(rst), .Q(sreg[1519])
         );
  DFF \sreg_reg[1520]  ( .D(swire[498]), .CLK(clk), .RST(rst), .Q(sreg[1520])
         );
  DFF \sreg_reg[1521]  ( .D(swire[499]), .CLK(clk), .RST(rst), .Q(sreg[1521])
         );
  DFF \sreg_reg[1522]  ( .D(swire[500]), .CLK(clk), .RST(rst), .Q(sreg[1522])
         );
  DFF \sreg_reg[1523]  ( .D(swire[501]), .CLK(clk), .RST(rst), .Q(sreg[1523])
         );
  DFF \sreg_reg[1524]  ( .D(swire[502]), .CLK(clk), .RST(rst), .Q(sreg[1524])
         );
  DFF \sreg_reg[1525]  ( .D(swire[503]), .CLK(clk), .RST(rst), .Q(sreg[1525])
         );
  DFF \sreg_reg[1526]  ( .D(swire[504]), .CLK(clk), .RST(rst), .Q(sreg[1526])
         );
  DFF \sreg_reg[1527]  ( .D(swire[505]), .CLK(clk), .RST(rst), .Q(sreg[1527])
         );
  DFF \sreg_reg[1528]  ( .D(swire[506]), .CLK(clk), .RST(rst), .Q(sreg[1528])
         );
  DFF \sreg_reg[1529]  ( .D(swire[507]), .CLK(clk), .RST(rst), .Q(sreg[1529])
         );
  DFF \sreg_reg[1530]  ( .D(swire[508]), .CLK(clk), .RST(rst), .Q(sreg[1530])
         );
  DFF \sreg_reg[1531]  ( .D(swire[509]), .CLK(clk), .RST(rst), .Q(sreg[1531])
         );
  DFF \sreg_reg[1532]  ( .D(swire[510]), .CLK(clk), .RST(rst), .Q(sreg[1532])
         );
  DFF \sreg_reg[1533]  ( .D(swire[511]), .CLK(clk), .RST(rst), .Q(sreg[1533])
         );
  DFF \sreg_reg[1534]  ( .D(swire[512]), .CLK(clk), .RST(rst), .Q(sreg[1534])
         );
  DFF \sreg_reg[1535]  ( .D(swire[513]), .CLK(clk), .RST(rst), .Q(sreg[1535])
         );
  DFF \sreg_reg[1536]  ( .D(swire[514]), .CLK(clk), .RST(rst), .Q(sreg[1536])
         );
  DFF \sreg_reg[1537]  ( .D(swire[515]), .CLK(clk), .RST(rst), .Q(sreg[1537])
         );
  DFF \sreg_reg[1538]  ( .D(swire[516]), .CLK(clk), .RST(rst), .Q(sreg[1538])
         );
  DFF \sreg_reg[1539]  ( .D(swire[517]), .CLK(clk), .RST(rst), .Q(sreg[1539])
         );
  DFF \sreg_reg[1540]  ( .D(swire[518]), .CLK(clk), .RST(rst), .Q(sreg[1540])
         );
  DFF \sreg_reg[1541]  ( .D(swire[519]), .CLK(clk), .RST(rst), .Q(sreg[1541])
         );
  DFF \sreg_reg[1542]  ( .D(swire[520]), .CLK(clk), .RST(rst), .Q(sreg[1542])
         );
  DFF \sreg_reg[1543]  ( .D(swire[521]), .CLK(clk), .RST(rst), .Q(sreg[1543])
         );
  DFF \sreg_reg[1544]  ( .D(swire[522]), .CLK(clk), .RST(rst), .Q(sreg[1544])
         );
  DFF \sreg_reg[1545]  ( .D(swire[523]), .CLK(clk), .RST(rst), .Q(sreg[1545])
         );
  DFF \sreg_reg[1546]  ( .D(swire[524]), .CLK(clk), .RST(rst), .Q(sreg[1546])
         );
  DFF \sreg_reg[1547]  ( .D(swire[525]), .CLK(clk), .RST(rst), .Q(sreg[1547])
         );
  DFF \sreg_reg[1548]  ( .D(swire[526]), .CLK(clk), .RST(rst), .Q(sreg[1548])
         );
  DFF \sreg_reg[1549]  ( .D(swire[527]), .CLK(clk), .RST(rst), .Q(sreg[1549])
         );
  DFF \sreg_reg[1550]  ( .D(swire[528]), .CLK(clk), .RST(rst), .Q(sreg[1550])
         );
  DFF \sreg_reg[1551]  ( .D(swire[529]), .CLK(clk), .RST(rst), .Q(sreg[1551])
         );
  DFF \sreg_reg[1552]  ( .D(swire[530]), .CLK(clk), .RST(rst), .Q(sreg[1552])
         );
  DFF \sreg_reg[1553]  ( .D(swire[531]), .CLK(clk), .RST(rst), .Q(sreg[1553])
         );
  DFF \sreg_reg[1554]  ( .D(swire[532]), .CLK(clk), .RST(rst), .Q(sreg[1554])
         );
  DFF \sreg_reg[1555]  ( .D(swire[533]), .CLK(clk), .RST(rst), .Q(sreg[1555])
         );
  DFF \sreg_reg[1556]  ( .D(swire[534]), .CLK(clk), .RST(rst), .Q(sreg[1556])
         );
  DFF \sreg_reg[1557]  ( .D(swire[535]), .CLK(clk), .RST(rst), .Q(sreg[1557])
         );
  DFF \sreg_reg[1558]  ( .D(swire[536]), .CLK(clk), .RST(rst), .Q(sreg[1558])
         );
  DFF \sreg_reg[1559]  ( .D(swire[537]), .CLK(clk), .RST(rst), .Q(sreg[1559])
         );
  DFF \sreg_reg[1560]  ( .D(swire[538]), .CLK(clk), .RST(rst), .Q(sreg[1560])
         );
  DFF \sreg_reg[1561]  ( .D(swire[539]), .CLK(clk), .RST(rst), .Q(sreg[1561])
         );
  DFF \sreg_reg[1562]  ( .D(swire[540]), .CLK(clk), .RST(rst), .Q(sreg[1562])
         );
  DFF \sreg_reg[1563]  ( .D(swire[541]), .CLK(clk), .RST(rst), .Q(sreg[1563])
         );
  DFF \sreg_reg[1564]  ( .D(swire[542]), .CLK(clk), .RST(rst), .Q(sreg[1564])
         );
  DFF \sreg_reg[1565]  ( .D(swire[543]), .CLK(clk), .RST(rst), .Q(sreg[1565])
         );
  DFF \sreg_reg[1566]  ( .D(swire[544]), .CLK(clk), .RST(rst), .Q(sreg[1566])
         );
  DFF \sreg_reg[1567]  ( .D(swire[545]), .CLK(clk), .RST(rst), .Q(sreg[1567])
         );
  DFF \sreg_reg[1568]  ( .D(swire[546]), .CLK(clk), .RST(rst), .Q(sreg[1568])
         );
  DFF \sreg_reg[1569]  ( .D(swire[547]), .CLK(clk), .RST(rst), .Q(sreg[1569])
         );
  DFF \sreg_reg[1570]  ( .D(swire[548]), .CLK(clk), .RST(rst), .Q(sreg[1570])
         );
  DFF \sreg_reg[1571]  ( .D(swire[549]), .CLK(clk), .RST(rst), .Q(sreg[1571])
         );
  DFF \sreg_reg[1572]  ( .D(swire[550]), .CLK(clk), .RST(rst), .Q(sreg[1572])
         );
  DFF \sreg_reg[1573]  ( .D(swire[551]), .CLK(clk), .RST(rst), .Q(sreg[1573])
         );
  DFF \sreg_reg[1574]  ( .D(swire[552]), .CLK(clk), .RST(rst), .Q(sreg[1574])
         );
  DFF \sreg_reg[1575]  ( .D(swire[553]), .CLK(clk), .RST(rst), .Q(sreg[1575])
         );
  DFF \sreg_reg[1576]  ( .D(swire[554]), .CLK(clk), .RST(rst), .Q(sreg[1576])
         );
  DFF \sreg_reg[1577]  ( .D(swire[555]), .CLK(clk), .RST(rst), .Q(sreg[1577])
         );
  DFF \sreg_reg[1578]  ( .D(swire[556]), .CLK(clk), .RST(rst), .Q(sreg[1578])
         );
  DFF \sreg_reg[1579]  ( .D(swire[557]), .CLK(clk), .RST(rst), .Q(sreg[1579])
         );
  DFF \sreg_reg[1580]  ( .D(swire[558]), .CLK(clk), .RST(rst), .Q(sreg[1580])
         );
  DFF \sreg_reg[1581]  ( .D(swire[559]), .CLK(clk), .RST(rst), .Q(sreg[1581])
         );
  DFF \sreg_reg[1582]  ( .D(swire[560]), .CLK(clk), .RST(rst), .Q(sreg[1582])
         );
  DFF \sreg_reg[1583]  ( .D(swire[561]), .CLK(clk), .RST(rst), .Q(sreg[1583])
         );
  DFF \sreg_reg[1584]  ( .D(swire[562]), .CLK(clk), .RST(rst), .Q(sreg[1584])
         );
  DFF \sreg_reg[1585]  ( .D(swire[563]), .CLK(clk), .RST(rst), .Q(sreg[1585])
         );
  DFF \sreg_reg[1586]  ( .D(swire[564]), .CLK(clk), .RST(rst), .Q(sreg[1586])
         );
  DFF \sreg_reg[1587]  ( .D(swire[565]), .CLK(clk), .RST(rst), .Q(sreg[1587])
         );
  DFF \sreg_reg[1588]  ( .D(swire[566]), .CLK(clk), .RST(rst), .Q(sreg[1588])
         );
  DFF \sreg_reg[1589]  ( .D(swire[567]), .CLK(clk), .RST(rst), .Q(sreg[1589])
         );
  DFF \sreg_reg[1590]  ( .D(swire[568]), .CLK(clk), .RST(rst), .Q(sreg[1590])
         );
  DFF \sreg_reg[1591]  ( .D(swire[569]), .CLK(clk), .RST(rst), .Q(sreg[1591])
         );
  DFF \sreg_reg[1592]  ( .D(swire[570]), .CLK(clk), .RST(rst), .Q(sreg[1592])
         );
  DFF \sreg_reg[1593]  ( .D(swire[571]), .CLK(clk), .RST(rst), .Q(sreg[1593])
         );
  DFF \sreg_reg[1594]  ( .D(swire[572]), .CLK(clk), .RST(rst), .Q(sreg[1594])
         );
  DFF \sreg_reg[1595]  ( .D(swire[573]), .CLK(clk), .RST(rst), .Q(sreg[1595])
         );
  DFF \sreg_reg[1596]  ( .D(swire[574]), .CLK(clk), .RST(rst), .Q(sreg[1596])
         );
  DFF \sreg_reg[1597]  ( .D(swire[575]), .CLK(clk), .RST(rst), .Q(sreg[1597])
         );
  DFF \sreg_reg[1598]  ( .D(swire[576]), .CLK(clk), .RST(rst), .Q(sreg[1598])
         );
  DFF \sreg_reg[1599]  ( .D(swire[577]), .CLK(clk), .RST(rst), .Q(sreg[1599])
         );
  DFF \sreg_reg[1600]  ( .D(swire[578]), .CLK(clk), .RST(rst), .Q(sreg[1600])
         );
  DFF \sreg_reg[1601]  ( .D(swire[579]), .CLK(clk), .RST(rst), .Q(sreg[1601])
         );
  DFF \sreg_reg[1602]  ( .D(swire[580]), .CLK(clk), .RST(rst), .Q(sreg[1602])
         );
  DFF \sreg_reg[1603]  ( .D(swire[581]), .CLK(clk), .RST(rst), .Q(sreg[1603])
         );
  DFF \sreg_reg[1604]  ( .D(swire[582]), .CLK(clk), .RST(rst), .Q(sreg[1604])
         );
  DFF \sreg_reg[1605]  ( .D(swire[583]), .CLK(clk), .RST(rst), .Q(sreg[1605])
         );
  DFF \sreg_reg[1606]  ( .D(swire[584]), .CLK(clk), .RST(rst), .Q(sreg[1606])
         );
  DFF \sreg_reg[1607]  ( .D(swire[585]), .CLK(clk), .RST(rst), .Q(sreg[1607])
         );
  DFF \sreg_reg[1608]  ( .D(swire[586]), .CLK(clk), .RST(rst), .Q(sreg[1608])
         );
  DFF \sreg_reg[1609]  ( .D(swire[587]), .CLK(clk), .RST(rst), .Q(sreg[1609])
         );
  DFF \sreg_reg[1610]  ( .D(swire[588]), .CLK(clk), .RST(rst), .Q(sreg[1610])
         );
  DFF \sreg_reg[1611]  ( .D(swire[589]), .CLK(clk), .RST(rst), .Q(sreg[1611])
         );
  DFF \sreg_reg[1612]  ( .D(swire[590]), .CLK(clk), .RST(rst), .Q(sreg[1612])
         );
  DFF \sreg_reg[1613]  ( .D(swire[591]), .CLK(clk), .RST(rst), .Q(sreg[1613])
         );
  DFF \sreg_reg[1614]  ( .D(swire[592]), .CLK(clk), .RST(rst), .Q(sreg[1614])
         );
  DFF \sreg_reg[1615]  ( .D(swire[593]), .CLK(clk), .RST(rst), .Q(sreg[1615])
         );
  DFF \sreg_reg[1616]  ( .D(swire[594]), .CLK(clk), .RST(rst), .Q(sreg[1616])
         );
  DFF \sreg_reg[1617]  ( .D(swire[595]), .CLK(clk), .RST(rst), .Q(sreg[1617])
         );
  DFF \sreg_reg[1618]  ( .D(swire[596]), .CLK(clk), .RST(rst), .Q(sreg[1618])
         );
  DFF \sreg_reg[1619]  ( .D(swire[597]), .CLK(clk), .RST(rst), .Q(sreg[1619])
         );
  DFF \sreg_reg[1620]  ( .D(swire[598]), .CLK(clk), .RST(rst), .Q(sreg[1620])
         );
  DFF \sreg_reg[1621]  ( .D(swire[599]), .CLK(clk), .RST(rst), .Q(sreg[1621])
         );
  DFF \sreg_reg[1622]  ( .D(swire[600]), .CLK(clk), .RST(rst), .Q(sreg[1622])
         );
  DFF \sreg_reg[1623]  ( .D(swire[601]), .CLK(clk), .RST(rst), .Q(sreg[1623])
         );
  DFF \sreg_reg[1624]  ( .D(swire[602]), .CLK(clk), .RST(rst), .Q(sreg[1624])
         );
  DFF \sreg_reg[1625]  ( .D(swire[603]), .CLK(clk), .RST(rst), .Q(sreg[1625])
         );
  DFF \sreg_reg[1626]  ( .D(swire[604]), .CLK(clk), .RST(rst), .Q(sreg[1626])
         );
  DFF \sreg_reg[1627]  ( .D(swire[605]), .CLK(clk), .RST(rst), .Q(sreg[1627])
         );
  DFF \sreg_reg[1628]  ( .D(swire[606]), .CLK(clk), .RST(rst), .Q(sreg[1628])
         );
  DFF \sreg_reg[1629]  ( .D(swire[607]), .CLK(clk), .RST(rst), .Q(sreg[1629])
         );
  DFF \sreg_reg[1630]  ( .D(swire[608]), .CLK(clk), .RST(rst), .Q(sreg[1630])
         );
  DFF \sreg_reg[1631]  ( .D(swire[609]), .CLK(clk), .RST(rst), .Q(sreg[1631])
         );
  DFF \sreg_reg[1632]  ( .D(swire[610]), .CLK(clk), .RST(rst), .Q(sreg[1632])
         );
  DFF \sreg_reg[1633]  ( .D(swire[611]), .CLK(clk), .RST(rst), .Q(sreg[1633])
         );
  DFF \sreg_reg[1634]  ( .D(swire[612]), .CLK(clk), .RST(rst), .Q(sreg[1634])
         );
  DFF \sreg_reg[1635]  ( .D(swire[613]), .CLK(clk), .RST(rst), .Q(sreg[1635])
         );
  DFF \sreg_reg[1636]  ( .D(swire[614]), .CLK(clk), .RST(rst), .Q(sreg[1636])
         );
  DFF \sreg_reg[1637]  ( .D(swire[615]), .CLK(clk), .RST(rst), .Q(sreg[1637])
         );
  DFF \sreg_reg[1638]  ( .D(swire[616]), .CLK(clk), .RST(rst), .Q(sreg[1638])
         );
  DFF \sreg_reg[1639]  ( .D(swire[617]), .CLK(clk), .RST(rst), .Q(sreg[1639])
         );
  DFF \sreg_reg[1640]  ( .D(swire[618]), .CLK(clk), .RST(rst), .Q(sreg[1640])
         );
  DFF \sreg_reg[1641]  ( .D(swire[619]), .CLK(clk), .RST(rst), .Q(sreg[1641])
         );
  DFF \sreg_reg[1642]  ( .D(swire[620]), .CLK(clk), .RST(rst), .Q(sreg[1642])
         );
  DFF \sreg_reg[1643]  ( .D(swire[621]), .CLK(clk), .RST(rst), .Q(sreg[1643])
         );
  DFF \sreg_reg[1644]  ( .D(swire[622]), .CLK(clk), .RST(rst), .Q(sreg[1644])
         );
  DFF \sreg_reg[1645]  ( .D(swire[623]), .CLK(clk), .RST(rst), .Q(sreg[1645])
         );
  DFF \sreg_reg[1646]  ( .D(swire[624]), .CLK(clk), .RST(rst), .Q(sreg[1646])
         );
  DFF \sreg_reg[1647]  ( .D(swire[625]), .CLK(clk), .RST(rst), .Q(sreg[1647])
         );
  DFF \sreg_reg[1648]  ( .D(swire[626]), .CLK(clk), .RST(rst), .Q(sreg[1648])
         );
  DFF \sreg_reg[1649]  ( .D(swire[627]), .CLK(clk), .RST(rst), .Q(sreg[1649])
         );
  DFF \sreg_reg[1650]  ( .D(swire[628]), .CLK(clk), .RST(rst), .Q(sreg[1650])
         );
  DFF \sreg_reg[1651]  ( .D(swire[629]), .CLK(clk), .RST(rst), .Q(sreg[1651])
         );
  DFF \sreg_reg[1652]  ( .D(swire[630]), .CLK(clk), .RST(rst), .Q(sreg[1652])
         );
  DFF \sreg_reg[1653]  ( .D(swire[631]), .CLK(clk), .RST(rst), .Q(sreg[1653])
         );
  DFF \sreg_reg[1654]  ( .D(swire[632]), .CLK(clk), .RST(rst), .Q(sreg[1654])
         );
  DFF \sreg_reg[1655]  ( .D(swire[633]), .CLK(clk), .RST(rst), .Q(sreg[1655])
         );
  DFF \sreg_reg[1656]  ( .D(swire[634]), .CLK(clk), .RST(rst), .Q(sreg[1656])
         );
  DFF \sreg_reg[1657]  ( .D(swire[635]), .CLK(clk), .RST(rst), .Q(sreg[1657])
         );
  DFF \sreg_reg[1658]  ( .D(swire[636]), .CLK(clk), .RST(rst), .Q(sreg[1658])
         );
  DFF \sreg_reg[1659]  ( .D(swire[637]), .CLK(clk), .RST(rst), .Q(sreg[1659])
         );
  DFF \sreg_reg[1660]  ( .D(swire[638]), .CLK(clk), .RST(rst), .Q(sreg[1660])
         );
  DFF \sreg_reg[1661]  ( .D(swire[639]), .CLK(clk), .RST(rst), .Q(sreg[1661])
         );
  DFF \sreg_reg[1662]  ( .D(swire[640]), .CLK(clk), .RST(rst), .Q(sreg[1662])
         );
  DFF \sreg_reg[1663]  ( .D(swire[641]), .CLK(clk), .RST(rst), .Q(sreg[1663])
         );
  DFF \sreg_reg[1664]  ( .D(swire[642]), .CLK(clk), .RST(rst), .Q(sreg[1664])
         );
  DFF \sreg_reg[1665]  ( .D(swire[643]), .CLK(clk), .RST(rst), .Q(sreg[1665])
         );
  DFF \sreg_reg[1666]  ( .D(swire[644]), .CLK(clk), .RST(rst), .Q(sreg[1666])
         );
  DFF \sreg_reg[1667]  ( .D(swire[645]), .CLK(clk), .RST(rst), .Q(sreg[1667])
         );
  DFF \sreg_reg[1668]  ( .D(swire[646]), .CLK(clk), .RST(rst), .Q(sreg[1668])
         );
  DFF \sreg_reg[1669]  ( .D(swire[647]), .CLK(clk), .RST(rst), .Q(sreg[1669])
         );
  DFF \sreg_reg[1670]  ( .D(swire[648]), .CLK(clk), .RST(rst), .Q(sreg[1670])
         );
  DFF \sreg_reg[1671]  ( .D(swire[649]), .CLK(clk), .RST(rst), .Q(sreg[1671])
         );
  DFF \sreg_reg[1672]  ( .D(swire[650]), .CLK(clk), .RST(rst), .Q(sreg[1672])
         );
  DFF \sreg_reg[1673]  ( .D(swire[651]), .CLK(clk), .RST(rst), .Q(sreg[1673])
         );
  DFF \sreg_reg[1674]  ( .D(swire[652]), .CLK(clk), .RST(rst), .Q(sreg[1674])
         );
  DFF \sreg_reg[1675]  ( .D(swire[653]), .CLK(clk), .RST(rst), .Q(sreg[1675])
         );
  DFF \sreg_reg[1676]  ( .D(swire[654]), .CLK(clk), .RST(rst), .Q(sreg[1676])
         );
  DFF \sreg_reg[1677]  ( .D(swire[655]), .CLK(clk), .RST(rst), .Q(sreg[1677])
         );
  DFF \sreg_reg[1678]  ( .D(swire[656]), .CLK(clk), .RST(rst), .Q(sreg[1678])
         );
  DFF \sreg_reg[1679]  ( .D(swire[657]), .CLK(clk), .RST(rst), .Q(sreg[1679])
         );
  DFF \sreg_reg[1680]  ( .D(swire[658]), .CLK(clk), .RST(rst), .Q(sreg[1680])
         );
  DFF \sreg_reg[1681]  ( .D(swire[659]), .CLK(clk), .RST(rst), .Q(sreg[1681])
         );
  DFF \sreg_reg[1682]  ( .D(swire[660]), .CLK(clk), .RST(rst), .Q(sreg[1682])
         );
  DFF \sreg_reg[1683]  ( .D(swire[661]), .CLK(clk), .RST(rst), .Q(sreg[1683])
         );
  DFF \sreg_reg[1684]  ( .D(swire[662]), .CLK(clk), .RST(rst), .Q(sreg[1684])
         );
  DFF \sreg_reg[1685]  ( .D(swire[663]), .CLK(clk), .RST(rst), .Q(sreg[1685])
         );
  DFF \sreg_reg[1686]  ( .D(swire[664]), .CLK(clk), .RST(rst), .Q(sreg[1686])
         );
  DFF \sreg_reg[1687]  ( .D(swire[665]), .CLK(clk), .RST(rst), .Q(sreg[1687])
         );
  DFF \sreg_reg[1688]  ( .D(swire[666]), .CLK(clk), .RST(rst), .Q(sreg[1688])
         );
  DFF \sreg_reg[1689]  ( .D(swire[667]), .CLK(clk), .RST(rst), .Q(sreg[1689])
         );
  DFF \sreg_reg[1690]  ( .D(swire[668]), .CLK(clk), .RST(rst), .Q(sreg[1690])
         );
  DFF \sreg_reg[1691]  ( .D(swire[669]), .CLK(clk), .RST(rst), .Q(sreg[1691])
         );
  DFF \sreg_reg[1692]  ( .D(swire[670]), .CLK(clk), .RST(rst), .Q(sreg[1692])
         );
  DFF \sreg_reg[1693]  ( .D(swire[671]), .CLK(clk), .RST(rst), .Q(sreg[1693])
         );
  DFF \sreg_reg[1694]  ( .D(swire[672]), .CLK(clk), .RST(rst), .Q(sreg[1694])
         );
  DFF \sreg_reg[1695]  ( .D(swire[673]), .CLK(clk), .RST(rst), .Q(sreg[1695])
         );
  DFF \sreg_reg[1696]  ( .D(swire[674]), .CLK(clk), .RST(rst), .Q(sreg[1696])
         );
  DFF \sreg_reg[1697]  ( .D(swire[675]), .CLK(clk), .RST(rst), .Q(sreg[1697])
         );
  DFF \sreg_reg[1698]  ( .D(swire[676]), .CLK(clk), .RST(rst), .Q(sreg[1698])
         );
  DFF \sreg_reg[1699]  ( .D(swire[677]), .CLK(clk), .RST(rst), .Q(sreg[1699])
         );
  DFF \sreg_reg[1700]  ( .D(swire[678]), .CLK(clk), .RST(rst), .Q(sreg[1700])
         );
  DFF \sreg_reg[1701]  ( .D(swire[679]), .CLK(clk), .RST(rst), .Q(sreg[1701])
         );
  DFF \sreg_reg[1702]  ( .D(swire[680]), .CLK(clk), .RST(rst), .Q(sreg[1702])
         );
  DFF \sreg_reg[1703]  ( .D(swire[681]), .CLK(clk), .RST(rst), .Q(sreg[1703])
         );
  DFF \sreg_reg[1704]  ( .D(swire[682]), .CLK(clk), .RST(rst), .Q(sreg[1704])
         );
  DFF \sreg_reg[1705]  ( .D(swire[683]), .CLK(clk), .RST(rst), .Q(sreg[1705])
         );
  DFF \sreg_reg[1706]  ( .D(swire[684]), .CLK(clk), .RST(rst), .Q(sreg[1706])
         );
  DFF \sreg_reg[1707]  ( .D(swire[685]), .CLK(clk), .RST(rst), .Q(sreg[1707])
         );
  DFF \sreg_reg[1708]  ( .D(swire[686]), .CLK(clk), .RST(rst), .Q(sreg[1708])
         );
  DFF \sreg_reg[1709]  ( .D(swire[687]), .CLK(clk), .RST(rst), .Q(sreg[1709])
         );
  DFF \sreg_reg[1710]  ( .D(swire[688]), .CLK(clk), .RST(rst), .Q(sreg[1710])
         );
  DFF \sreg_reg[1711]  ( .D(swire[689]), .CLK(clk), .RST(rst), .Q(sreg[1711])
         );
  DFF \sreg_reg[1712]  ( .D(swire[690]), .CLK(clk), .RST(rst), .Q(sreg[1712])
         );
  DFF \sreg_reg[1713]  ( .D(swire[691]), .CLK(clk), .RST(rst), .Q(sreg[1713])
         );
  DFF \sreg_reg[1714]  ( .D(swire[692]), .CLK(clk), .RST(rst), .Q(sreg[1714])
         );
  DFF \sreg_reg[1715]  ( .D(swire[693]), .CLK(clk), .RST(rst), .Q(sreg[1715])
         );
  DFF \sreg_reg[1716]  ( .D(swire[694]), .CLK(clk), .RST(rst), .Q(sreg[1716])
         );
  DFF \sreg_reg[1717]  ( .D(swire[695]), .CLK(clk), .RST(rst), .Q(sreg[1717])
         );
  DFF \sreg_reg[1718]  ( .D(swire[696]), .CLK(clk), .RST(rst), .Q(sreg[1718])
         );
  DFF \sreg_reg[1719]  ( .D(swire[697]), .CLK(clk), .RST(rst), .Q(sreg[1719])
         );
  DFF \sreg_reg[1720]  ( .D(swire[698]), .CLK(clk), .RST(rst), .Q(sreg[1720])
         );
  DFF \sreg_reg[1721]  ( .D(swire[699]), .CLK(clk), .RST(rst), .Q(sreg[1721])
         );
  DFF \sreg_reg[1722]  ( .D(swire[700]), .CLK(clk), .RST(rst), .Q(sreg[1722])
         );
  DFF \sreg_reg[1723]  ( .D(swire[701]), .CLK(clk), .RST(rst), .Q(sreg[1723])
         );
  DFF \sreg_reg[1724]  ( .D(swire[702]), .CLK(clk), .RST(rst), .Q(sreg[1724])
         );
  DFF \sreg_reg[1725]  ( .D(swire[703]), .CLK(clk), .RST(rst), .Q(sreg[1725])
         );
  DFF \sreg_reg[1726]  ( .D(swire[704]), .CLK(clk), .RST(rst), .Q(sreg[1726])
         );
  DFF \sreg_reg[1727]  ( .D(swire[705]), .CLK(clk), .RST(rst), .Q(sreg[1727])
         );
  DFF \sreg_reg[1728]  ( .D(swire[706]), .CLK(clk), .RST(rst), .Q(sreg[1728])
         );
  DFF \sreg_reg[1729]  ( .D(swire[707]), .CLK(clk), .RST(rst), .Q(sreg[1729])
         );
  DFF \sreg_reg[1730]  ( .D(swire[708]), .CLK(clk), .RST(rst), .Q(sreg[1730])
         );
  DFF \sreg_reg[1731]  ( .D(swire[709]), .CLK(clk), .RST(rst), .Q(sreg[1731])
         );
  DFF \sreg_reg[1732]  ( .D(swire[710]), .CLK(clk), .RST(rst), .Q(sreg[1732])
         );
  DFF \sreg_reg[1733]  ( .D(swire[711]), .CLK(clk), .RST(rst), .Q(sreg[1733])
         );
  DFF \sreg_reg[1734]  ( .D(swire[712]), .CLK(clk), .RST(rst), .Q(sreg[1734])
         );
  DFF \sreg_reg[1735]  ( .D(swire[713]), .CLK(clk), .RST(rst), .Q(sreg[1735])
         );
  DFF \sreg_reg[1736]  ( .D(swire[714]), .CLK(clk), .RST(rst), .Q(sreg[1736])
         );
  DFF \sreg_reg[1737]  ( .D(swire[715]), .CLK(clk), .RST(rst), .Q(sreg[1737])
         );
  DFF \sreg_reg[1738]  ( .D(swire[716]), .CLK(clk), .RST(rst), .Q(sreg[1738])
         );
  DFF \sreg_reg[1739]  ( .D(swire[717]), .CLK(clk), .RST(rst), .Q(sreg[1739])
         );
  DFF \sreg_reg[1740]  ( .D(swire[718]), .CLK(clk), .RST(rst), .Q(sreg[1740])
         );
  DFF \sreg_reg[1741]  ( .D(swire[719]), .CLK(clk), .RST(rst), .Q(sreg[1741])
         );
  DFF \sreg_reg[1742]  ( .D(swire[720]), .CLK(clk), .RST(rst), .Q(sreg[1742])
         );
  DFF \sreg_reg[1743]  ( .D(swire[721]), .CLK(clk), .RST(rst), .Q(sreg[1743])
         );
  DFF \sreg_reg[1744]  ( .D(swire[722]), .CLK(clk), .RST(rst), .Q(sreg[1744])
         );
  DFF \sreg_reg[1745]  ( .D(swire[723]), .CLK(clk), .RST(rst), .Q(sreg[1745])
         );
  DFF \sreg_reg[1746]  ( .D(swire[724]), .CLK(clk), .RST(rst), .Q(sreg[1746])
         );
  DFF \sreg_reg[1747]  ( .D(swire[725]), .CLK(clk), .RST(rst), .Q(sreg[1747])
         );
  DFF \sreg_reg[1748]  ( .D(swire[726]), .CLK(clk), .RST(rst), .Q(sreg[1748])
         );
  DFF \sreg_reg[1749]  ( .D(swire[727]), .CLK(clk), .RST(rst), .Q(sreg[1749])
         );
  DFF \sreg_reg[1750]  ( .D(swire[728]), .CLK(clk), .RST(rst), .Q(sreg[1750])
         );
  DFF \sreg_reg[1751]  ( .D(swire[729]), .CLK(clk), .RST(rst), .Q(sreg[1751])
         );
  DFF \sreg_reg[1752]  ( .D(swire[730]), .CLK(clk), .RST(rst), .Q(sreg[1752])
         );
  DFF \sreg_reg[1753]  ( .D(swire[731]), .CLK(clk), .RST(rst), .Q(sreg[1753])
         );
  DFF \sreg_reg[1754]  ( .D(swire[732]), .CLK(clk), .RST(rst), .Q(sreg[1754])
         );
  DFF \sreg_reg[1755]  ( .D(swire[733]), .CLK(clk), .RST(rst), .Q(sreg[1755])
         );
  DFF \sreg_reg[1756]  ( .D(swire[734]), .CLK(clk), .RST(rst), .Q(sreg[1756])
         );
  DFF \sreg_reg[1757]  ( .D(swire[735]), .CLK(clk), .RST(rst), .Q(sreg[1757])
         );
  DFF \sreg_reg[1758]  ( .D(swire[736]), .CLK(clk), .RST(rst), .Q(sreg[1758])
         );
  DFF \sreg_reg[1759]  ( .D(swire[737]), .CLK(clk), .RST(rst), .Q(sreg[1759])
         );
  DFF \sreg_reg[1760]  ( .D(swire[738]), .CLK(clk), .RST(rst), .Q(sreg[1760])
         );
  DFF \sreg_reg[1761]  ( .D(swire[739]), .CLK(clk), .RST(rst), .Q(sreg[1761])
         );
  DFF \sreg_reg[1762]  ( .D(swire[740]), .CLK(clk), .RST(rst), .Q(sreg[1762])
         );
  DFF \sreg_reg[1763]  ( .D(swire[741]), .CLK(clk), .RST(rst), .Q(sreg[1763])
         );
  DFF \sreg_reg[1764]  ( .D(swire[742]), .CLK(clk), .RST(rst), .Q(sreg[1764])
         );
  DFF \sreg_reg[1765]  ( .D(swire[743]), .CLK(clk), .RST(rst), .Q(sreg[1765])
         );
  DFF \sreg_reg[1766]  ( .D(swire[744]), .CLK(clk), .RST(rst), .Q(sreg[1766])
         );
  DFF \sreg_reg[1767]  ( .D(swire[745]), .CLK(clk), .RST(rst), .Q(sreg[1767])
         );
  DFF \sreg_reg[1768]  ( .D(swire[746]), .CLK(clk), .RST(rst), .Q(sreg[1768])
         );
  DFF \sreg_reg[1769]  ( .D(swire[747]), .CLK(clk), .RST(rst), .Q(sreg[1769])
         );
  DFF \sreg_reg[1770]  ( .D(swire[748]), .CLK(clk), .RST(rst), .Q(sreg[1770])
         );
  DFF \sreg_reg[1771]  ( .D(swire[749]), .CLK(clk), .RST(rst), .Q(sreg[1771])
         );
  DFF \sreg_reg[1772]  ( .D(swire[750]), .CLK(clk), .RST(rst), .Q(sreg[1772])
         );
  DFF \sreg_reg[1773]  ( .D(swire[751]), .CLK(clk), .RST(rst), .Q(sreg[1773])
         );
  DFF \sreg_reg[1774]  ( .D(swire[752]), .CLK(clk), .RST(rst), .Q(sreg[1774])
         );
  DFF \sreg_reg[1775]  ( .D(swire[753]), .CLK(clk), .RST(rst), .Q(sreg[1775])
         );
  DFF \sreg_reg[1776]  ( .D(swire[754]), .CLK(clk), .RST(rst), .Q(sreg[1776])
         );
  DFF \sreg_reg[1777]  ( .D(swire[755]), .CLK(clk), .RST(rst), .Q(sreg[1777])
         );
  DFF \sreg_reg[1778]  ( .D(swire[756]), .CLK(clk), .RST(rst), .Q(sreg[1778])
         );
  DFF \sreg_reg[1779]  ( .D(swire[757]), .CLK(clk), .RST(rst), .Q(sreg[1779])
         );
  DFF \sreg_reg[1780]  ( .D(swire[758]), .CLK(clk), .RST(rst), .Q(sreg[1780])
         );
  DFF \sreg_reg[1781]  ( .D(swire[759]), .CLK(clk), .RST(rst), .Q(sreg[1781])
         );
  DFF \sreg_reg[1782]  ( .D(swire[760]), .CLK(clk), .RST(rst), .Q(sreg[1782])
         );
  DFF \sreg_reg[1783]  ( .D(swire[761]), .CLK(clk), .RST(rst), .Q(sreg[1783])
         );
  DFF \sreg_reg[1784]  ( .D(swire[762]), .CLK(clk), .RST(rst), .Q(sreg[1784])
         );
  DFF \sreg_reg[1785]  ( .D(swire[763]), .CLK(clk), .RST(rst), .Q(sreg[1785])
         );
  DFF \sreg_reg[1786]  ( .D(swire[764]), .CLK(clk), .RST(rst), .Q(sreg[1786])
         );
  DFF \sreg_reg[1787]  ( .D(swire[765]), .CLK(clk), .RST(rst), .Q(sreg[1787])
         );
  DFF \sreg_reg[1788]  ( .D(swire[766]), .CLK(clk), .RST(rst), .Q(sreg[1788])
         );
  DFF \sreg_reg[1789]  ( .D(swire[767]), .CLK(clk), .RST(rst), .Q(sreg[1789])
         );
  DFF \sreg_reg[1790]  ( .D(swire[768]), .CLK(clk), .RST(rst), .Q(sreg[1790])
         );
  DFF \sreg_reg[1791]  ( .D(swire[769]), .CLK(clk), .RST(rst), .Q(sreg[1791])
         );
  DFF \sreg_reg[1792]  ( .D(swire[770]), .CLK(clk), .RST(rst), .Q(sreg[1792])
         );
  DFF \sreg_reg[1793]  ( .D(swire[771]), .CLK(clk), .RST(rst), .Q(sreg[1793])
         );
  DFF \sreg_reg[1794]  ( .D(swire[772]), .CLK(clk), .RST(rst), .Q(sreg[1794])
         );
  DFF \sreg_reg[1795]  ( .D(swire[773]), .CLK(clk), .RST(rst), .Q(sreg[1795])
         );
  DFF \sreg_reg[1796]  ( .D(swire[774]), .CLK(clk), .RST(rst), .Q(sreg[1796])
         );
  DFF \sreg_reg[1797]  ( .D(swire[775]), .CLK(clk), .RST(rst), .Q(sreg[1797])
         );
  DFF \sreg_reg[1798]  ( .D(swire[776]), .CLK(clk), .RST(rst), .Q(sreg[1798])
         );
  DFF \sreg_reg[1799]  ( .D(swire[777]), .CLK(clk), .RST(rst), .Q(sreg[1799])
         );
  DFF \sreg_reg[1800]  ( .D(swire[778]), .CLK(clk), .RST(rst), .Q(sreg[1800])
         );
  DFF \sreg_reg[1801]  ( .D(swire[779]), .CLK(clk), .RST(rst), .Q(sreg[1801])
         );
  DFF \sreg_reg[1802]  ( .D(swire[780]), .CLK(clk), .RST(rst), .Q(sreg[1802])
         );
  DFF \sreg_reg[1803]  ( .D(swire[781]), .CLK(clk), .RST(rst), .Q(sreg[1803])
         );
  DFF \sreg_reg[1804]  ( .D(swire[782]), .CLK(clk), .RST(rst), .Q(sreg[1804])
         );
  DFF \sreg_reg[1805]  ( .D(swire[783]), .CLK(clk), .RST(rst), .Q(sreg[1805])
         );
  DFF \sreg_reg[1806]  ( .D(swire[784]), .CLK(clk), .RST(rst), .Q(sreg[1806])
         );
  DFF \sreg_reg[1807]  ( .D(swire[785]), .CLK(clk), .RST(rst), .Q(sreg[1807])
         );
  DFF \sreg_reg[1808]  ( .D(swire[786]), .CLK(clk), .RST(rst), .Q(sreg[1808])
         );
  DFF \sreg_reg[1809]  ( .D(swire[787]), .CLK(clk), .RST(rst), .Q(sreg[1809])
         );
  DFF \sreg_reg[1810]  ( .D(swire[788]), .CLK(clk), .RST(rst), .Q(sreg[1810])
         );
  DFF \sreg_reg[1811]  ( .D(swire[789]), .CLK(clk), .RST(rst), .Q(sreg[1811])
         );
  DFF \sreg_reg[1812]  ( .D(swire[790]), .CLK(clk), .RST(rst), .Q(sreg[1812])
         );
  DFF \sreg_reg[1813]  ( .D(swire[791]), .CLK(clk), .RST(rst), .Q(sreg[1813])
         );
  DFF \sreg_reg[1814]  ( .D(swire[792]), .CLK(clk), .RST(rst), .Q(sreg[1814])
         );
  DFF \sreg_reg[1815]  ( .D(swire[793]), .CLK(clk), .RST(rst), .Q(sreg[1815])
         );
  DFF \sreg_reg[1816]  ( .D(swire[794]), .CLK(clk), .RST(rst), .Q(sreg[1816])
         );
  DFF \sreg_reg[1817]  ( .D(swire[795]), .CLK(clk), .RST(rst), .Q(sreg[1817])
         );
  DFF \sreg_reg[1818]  ( .D(swire[796]), .CLK(clk), .RST(rst), .Q(sreg[1818])
         );
  DFF \sreg_reg[1819]  ( .D(swire[797]), .CLK(clk), .RST(rst), .Q(sreg[1819])
         );
  DFF \sreg_reg[1820]  ( .D(swire[798]), .CLK(clk), .RST(rst), .Q(sreg[1820])
         );
  DFF \sreg_reg[1821]  ( .D(swire[799]), .CLK(clk), .RST(rst), .Q(sreg[1821])
         );
  DFF \sreg_reg[1822]  ( .D(swire[800]), .CLK(clk), .RST(rst), .Q(sreg[1822])
         );
  DFF \sreg_reg[1823]  ( .D(swire[801]), .CLK(clk), .RST(rst), .Q(sreg[1823])
         );
  DFF \sreg_reg[1824]  ( .D(swire[802]), .CLK(clk), .RST(rst), .Q(sreg[1824])
         );
  DFF \sreg_reg[1825]  ( .D(swire[803]), .CLK(clk), .RST(rst), .Q(sreg[1825])
         );
  DFF \sreg_reg[1826]  ( .D(swire[804]), .CLK(clk), .RST(rst), .Q(sreg[1826])
         );
  DFF \sreg_reg[1827]  ( .D(swire[805]), .CLK(clk), .RST(rst), .Q(sreg[1827])
         );
  DFF \sreg_reg[1828]  ( .D(swire[806]), .CLK(clk), .RST(rst), .Q(sreg[1828])
         );
  DFF \sreg_reg[1829]  ( .D(swire[807]), .CLK(clk), .RST(rst), .Q(sreg[1829])
         );
  DFF \sreg_reg[1830]  ( .D(swire[808]), .CLK(clk), .RST(rst), .Q(sreg[1830])
         );
  DFF \sreg_reg[1831]  ( .D(swire[809]), .CLK(clk), .RST(rst), .Q(sreg[1831])
         );
  DFF \sreg_reg[1832]  ( .D(swire[810]), .CLK(clk), .RST(rst), .Q(sreg[1832])
         );
  DFF \sreg_reg[1833]  ( .D(swire[811]), .CLK(clk), .RST(rst), .Q(sreg[1833])
         );
  DFF \sreg_reg[1834]  ( .D(swire[812]), .CLK(clk), .RST(rst), .Q(sreg[1834])
         );
  DFF \sreg_reg[1835]  ( .D(swire[813]), .CLK(clk), .RST(rst), .Q(sreg[1835])
         );
  DFF \sreg_reg[1836]  ( .D(swire[814]), .CLK(clk), .RST(rst), .Q(sreg[1836])
         );
  DFF \sreg_reg[1837]  ( .D(swire[815]), .CLK(clk), .RST(rst), .Q(sreg[1837])
         );
  DFF \sreg_reg[1838]  ( .D(swire[816]), .CLK(clk), .RST(rst), .Q(sreg[1838])
         );
  DFF \sreg_reg[1839]  ( .D(swire[817]), .CLK(clk), .RST(rst), .Q(sreg[1839])
         );
  DFF \sreg_reg[1840]  ( .D(swire[818]), .CLK(clk), .RST(rst), .Q(sreg[1840])
         );
  DFF \sreg_reg[1841]  ( .D(swire[819]), .CLK(clk), .RST(rst), .Q(sreg[1841])
         );
  DFF \sreg_reg[1842]  ( .D(swire[820]), .CLK(clk), .RST(rst), .Q(sreg[1842])
         );
  DFF \sreg_reg[1843]  ( .D(swire[821]), .CLK(clk), .RST(rst), .Q(sreg[1843])
         );
  DFF \sreg_reg[1844]  ( .D(swire[822]), .CLK(clk), .RST(rst), .Q(sreg[1844])
         );
  DFF \sreg_reg[1845]  ( .D(swire[823]), .CLK(clk), .RST(rst), .Q(sreg[1845])
         );
  DFF \sreg_reg[1846]  ( .D(swire[824]), .CLK(clk), .RST(rst), .Q(sreg[1846])
         );
  DFF \sreg_reg[1847]  ( .D(swire[825]), .CLK(clk), .RST(rst), .Q(sreg[1847])
         );
  DFF \sreg_reg[1848]  ( .D(swire[826]), .CLK(clk), .RST(rst), .Q(sreg[1848])
         );
  DFF \sreg_reg[1849]  ( .D(swire[827]), .CLK(clk), .RST(rst), .Q(sreg[1849])
         );
  DFF \sreg_reg[1850]  ( .D(swire[828]), .CLK(clk), .RST(rst), .Q(sreg[1850])
         );
  DFF \sreg_reg[1851]  ( .D(swire[829]), .CLK(clk), .RST(rst), .Q(sreg[1851])
         );
  DFF \sreg_reg[1852]  ( .D(swire[830]), .CLK(clk), .RST(rst), .Q(sreg[1852])
         );
  DFF \sreg_reg[1853]  ( .D(swire[831]), .CLK(clk), .RST(rst), .Q(sreg[1853])
         );
  DFF \sreg_reg[1854]  ( .D(swire[832]), .CLK(clk), .RST(rst), .Q(sreg[1854])
         );
  DFF \sreg_reg[1855]  ( .D(swire[833]), .CLK(clk), .RST(rst), .Q(sreg[1855])
         );
  DFF \sreg_reg[1856]  ( .D(swire[834]), .CLK(clk), .RST(rst), .Q(sreg[1856])
         );
  DFF \sreg_reg[1857]  ( .D(swire[835]), .CLK(clk), .RST(rst), .Q(sreg[1857])
         );
  DFF \sreg_reg[1858]  ( .D(swire[836]), .CLK(clk), .RST(rst), .Q(sreg[1858])
         );
  DFF \sreg_reg[1859]  ( .D(swire[837]), .CLK(clk), .RST(rst), .Q(sreg[1859])
         );
  DFF \sreg_reg[1860]  ( .D(swire[838]), .CLK(clk), .RST(rst), .Q(sreg[1860])
         );
  DFF \sreg_reg[1861]  ( .D(swire[839]), .CLK(clk), .RST(rst), .Q(sreg[1861])
         );
  DFF \sreg_reg[1862]  ( .D(swire[840]), .CLK(clk), .RST(rst), .Q(sreg[1862])
         );
  DFF \sreg_reg[1863]  ( .D(swire[841]), .CLK(clk), .RST(rst), .Q(sreg[1863])
         );
  DFF \sreg_reg[1864]  ( .D(swire[842]), .CLK(clk), .RST(rst), .Q(sreg[1864])
         );
  DFF \sreg_reg[1865]  ( .D(swire[843]), .CLK(clk), .RST(rst), .Q(sreg[1865])
         );
  DFF \sreg_reg[1866]  ( .D(swire[844]), .CLK(clk), .RST(rst), .Q(sreg[1866])
         );
  DFF \sreg_reg[1867]  ( .D(swire[845]), .CLK(clk), .RST(rst), .Q(sreg[1867])
         );
  DFF \sreg_reg[1868]  ( .D(swire[846]), .CLK(clk), .RST(rst), .Q(sreg[1868])
         );
  DFF \sreg_reg[1869]  ( .D(swire[847]), .CLK(clk), .RST(rst), .Q(sreg[1869])
         );
  DFF \sreg_reg[1870]  ( .D(swire[848]), .CLK(clk), .RST(rst), .Q(sreg[1870])
         );
  DFF \sreg_reg[1871]  ( .D(swire[849]), .CLK(clk), .RST(rst), .Q(sreg[1871])
         );
  DFF \sreg_reg[1872]  ( .D(swire[850]), .CLK(clk), .RST(rst), .Q(sreg[1872])
         );
  DFF \sreg_reg[1873]  ( .D(swire[851]), .CLK(clk), .RST(rst), .Q(sreg[1873])
         );
  DFF \sreg_reg[1874]  ( .D(swire[852]), .CLK(clk), .RST(rst), .Q(sreg[1874])
         );
  DFF \sreg_reg[1875]  ( .D(swire[853]), .CLK(clk), .RST(rst), .Q(sreg[1875])
         );
  DFF \sreg_reg[1876]  ( .D(swire[854]), .CLK(clk), .RST(rst), .Q(sreg[1876])
         );
  DFF \sreg_reg[1877]  ( .D(swire[855]), .CLK(clk), .RST(rst), .Q(sreg[1877])
         );
  DFF \sreg_reg[1878]  ( .D(swire[856]), .CLK(clk), .RST(rst), .Q(sreg[1878])
         );
  DFF \sreg_reg[1879]  ( .D(swire[857]), .CLK(clk), .RST(rst), .Q(sreg[1879])
         );
  DFF \sreg_reg[1880]  ( .D(swire[858]), .CLK(clk), .RST(rst), .Q(sreg[1880])
         );
  DFF \sreg_reg[1881]  ( .D(swire[859]), .CLK(clk), .RST(rst), .Q(sreg[1881])
         );
  DFF \sreg_reg[1882]  ( .D(swire[860]), .CLK(clk), .RST(rst), .Q(sreg[1882])
         );
  DFF \sreg_reg[1883]  ( .D(swire[861]), .CLK(clk), .RST(rst), .Q(sreg[1883])
         );
  DFF \sreg_reg[1884]  ( .D(swire[862]), .CLK(clk), .RST(rst), .Q(sreg[1884])
         );
  DFF \sreg_reg[1885]  ( .D(swire[863]), .CLK(clk), .RST(rst), .Q(sreg[1885])
         );
  DFF \sreg_reg[1886]  ( .D(swire[864]), .CLK(clk), .RST(rst), .Q(sreg[1886])
         );
  DFF \sreg_reg[1887]  ( .D(swire[865]), .CLK(clk), .RST(rst), .Q(sreg[1887])
         );
  DFF \sreg_reg[1888]  ( .D(swire[866]), .CLK(clk), .RST(rst), .Q(sreg[1888])
         );
  DFF \sreg_reg[1889]  ( .D(swire[867]), .CLK(clk), .RST(rst), .Q(sreg[1889])
         );
  DFF \sreg_reg[1890]  ( .D(swire[868]), .CLK(clk), .RST(rst), .Q(sreg[1890])
         );
  DFF \sreg_reg[1891]  ( .D(swire[869]), .CLK(clk), .RST(rst), .Q(sreg[1891])
         );
  DFF \sreg_reg[1892]  ( .D(swire[870]), .CLK(clk), .RST(rst), .Q(sreg[1892])
         );
  DFF \sreg_reg[1893]  ( .D(swire[871]), .CLK(clk), .RST(rst), .Q(sreg[1893])
         );
  DFF \sreg_reg[1894]  ( .D(swire[872]), .CLK(clk), .RST(rst), .Q(sreg[1894])
         );
  DFF \sreg_reg[1895]  ( .D(swire[873]), .CLK(clk), .RST(rst), .Q(sreg[1895])
         );
  DFF \sreg_reg[1896]  ( .D(swire[874]), .CLK(clk), .RST(rst), .Q(sreg[1896])
         );
  DFF \sreg_reg[1897]  ( .D(swire[875]), .CLK(clk), .RST(rst), .Q(sreg[1897])
         );
  DFF \sreg_reg[1898]  ( .D(swire[876]), .CLK(clk), .RST(rst), .Q(sreg[1898])
         );
  DFF \sreg_reg[1899]  ( .D(swire[877]), .CLK(clk), .RST(rst), .Q(sreg[1899])
         );
  DFF \sreg_reg[1900]  ( .D(swire[878]), .CLK(clk), .RST(rst), .Q(sreg[1900])
         );
  DFF \sreg_reg[1901]  ( .D(swire[879]), .CLK(clk), .RST(rst), .Q(sreg[1901])
         );
  DFF \sreg_reg[1902]  ( .D(swire[880]), .CLK(clk), .RST(rst), .Q(sreg[1902])
         );
  DFF \sreg_reg[1903]  ( .D(swire[881]), .CLK(clk), .RST(rst), .Q(sreg[1903])
         );
  DFF \sreg_reg[1904]  ( .D(swire[882]), .CLK(clk), .RST(rst), .Q(sreg[1904])
         );
  DFF \sreg_reg[1905]  ( .D(swire[883]), .CLK(clk), .RST(rst), .Q(sreg[1905])
         );
  DFF \sreg_reg[1906]  ( .D(swire[884]), .CLK(clk), .RST(rst), .Q(sreg[1906])
         );
  DFF \sreg_reg[1907]  ( .D(swire[885]), .CLK(clk), .RST(rst), .Q(sreg[1907])
         );
  DFF \sreg_reg[1908]  ( .D(swire[886]), .CLK(clk), .RST(rst), .Q(sreg[1908])
         );
  DFF \sreg_reg[1909]  ( .D(swire[887]), .CLK(clk), .RST(rst), .Q(sreg[1909])
         );
  DFF \sreg_reg[1910]  ( .D(swire[888]), .CLK(clk), .RST(rst), .Q(sreg[1910])
         );
  DFF \sreg_reg[1911]  ( .D(swire[889]), .CLK(clk), .RST(rst), .Q(sreg[1911])
         );
  DFF \sreg_reg[1912]  ( .D(swire[890]), .CLK(clk), .RST(rst), .Q(sreg[1912])
         );
  DFF \sreg_reg[1913]  ( .D(swire[891]), .CLK(clk), .RST(rst), .Q(sreg[1913])
         );
  DFF \sreg_reg[1914]  ( .D(swire[892]), .CLK(clk), .RST(rst), .Q(sreg[1914])
         );
  DFF \sreg_reg[1915]  ( .D(swire[893]), .CLK(clk), .RST(rst), .Q(sreg[1915])
         );
  DFF \sreg_reg[1916]  ( .D(swire[894]), .CLK(clk), .RST(rst), .Q(sreg[1916])
         );
  DFF \sreg_reg[1917]  ( .D(swire[895]), .CLK(clk), .RST(rst), .Q(sreg[1917])
         );
  DFF \sreg_reg[1918]  ( .D(swire[896]), .CLK(clk), .RST(rst), .Q(sreg[1918])
         );
  DFF \sreg_reg[1919]  ( .D(swire[897]), .CLK(clk), .RST(rst), .Q(sreg[1919])
         );
  DFF \sreg_reg[1920]  ( .D(swire[898]), .CLK(clk), .RST(rst), .Q(sreg[1920])
         );
  DFF \sreg_reg[1921]  ( .D(swire[899]), .CLK(clk), .RST(rst), .Q(sreg[1921])
         );
  DFF \sreg_reg[1922]  ( .D(swire[900]), .CLK(clk), .RST(rst), .Q(sreg[1922])
         );
  DFF \sreg_reg[1923]  ( .D(swire[901]), .CLK(clk), .RST(rst), .Q(sreg[1923])
         );
  DFF \sreg_reg[1924]  ( .D(swire[902]), .CLK(clk), .RST(rst), .Q(sreg[1924])
         );
  DFF \sreg_reg[1925]  ( .D(swire[903]), .CLK(clk), .RST(rst), .Q(sreg[1925])
         );
  DFF \sreg_reg[1926]  ( .D(swire[904]), .CLK(clk), .RST(rst), .Q(sreg[1926])
         );
  DFF \sreg_reg[1927]  ( .D(swire[905]), .CLK(clk), .RST(rst), .Q(sreg[1927])
         );
  DFF \sreg_reg[1928]  ( .D(swire[906]), .CLK(clk), .RST(rst), .Q(sreg[1928])
         );
  DFF \sreg_reg[1929]  ( .D(swire[907]), .CLK(clk), .RST(rst), .Q(sreg[1929])
         );
  DFF \sreg_reg[1930]  ( .D(swire[908]), .CLK(clk), .RST(rst), .Q(sreg[1930])
         );
  DFF \sreg_reg[1931]  ( .D(swire[909]), .CLK(clk), .RST(rst), .Q(sreg[1931])
         );
  DFF \sreg_reg[1932]  ( .D(swire[910]), .CLK(clk), .RST(rst), .Q(sreg[1932])
         );
  DFF \sreg_reg[1933]  ( .D(swire[911]), .CLK(clk), .RST(rst), .Q(sreg[1933])
         );
  DFF \sreg_reg[1934]  ( .D(swire[912]), .CLK(clk), .RST(rst), .Q(sreg[1934])
         );
  DFF \sreg_reg[1935]  ( .D(swire[913]), .CLK(clk), .RST(rst), .Q(sreg[1935])
         );
  DFF \sreg_reg[1936]  ( .D(swire[914]), .CLK(clk), .RST(rst), .Q(sreg[1936])
         );
  DFF \sreg_reg[1937]  ( .D(swire[915]), .CLK(clk), .RST(rst), .Q(sreg[1937])
         );
  DFF \sreg_reg[1938]  ( .D(swire[916]), .CLK(clk), .RST(rst), .Q(sreg[1938])
         );
  DFF \sreg_reg[1939]  ( .D(swire[917]), .CLK(clk), .RST(rst), .Q(sreg[1939])
         );
  DFF \sreg_reg[1940]  ( .D(swire[918]), .CLK(clk), .RST(rst), .Q(sreg[1940])
         );
  DFF \sreg_reg[1941]  ( .D(swire[919]), .CLK(clk), .RST(rst), .Q(sreg[1941])
         );
  DFF \sreg_reg[1942]  ( .D(swire[920]), .CLK(clk), .RST(rst), .Q(sreg[1942])
         );
  DFF \sreg_reg[1943]  ( .D(swire[921]), .CLK(clk), .RST(rst), .Q(sreg[1943])
         );
  DFF \sreg_reg[1944]  ( .D(swire[922]), .CLK(clk), .RST(rst), .Q(sreg[1944])
         );
  DFF \sreg_reg[1945]  ( .D(swire[923]), .CLK(clk), .RST(rst), .Q(sreg[1945])
         );
  DFF \sreg_reg[1946]  ( .D(swire[924]), .CLK(clk), .RST(rst), .Q(sreg[1946])
         );
  DFF \sreg_reg[1947]  ( .D(swire[925]), .CLK(clk), .RST(rst), .Q(sreg[1947])
         );
  DFF \sreg_reg[1948]  ( .D(swire[926]), .CLK(clk), .RST(rst), .Q(sreg[1948])
         );
  DFF \sreg_reg[1949]  ( .D(swire[927]), .CLK(clk), .RST(rst), .Q(sreg[1949])
         );
  DFF \sreg_reg[1950]  ( .D(swire[928]), .CLK(clk), .RST(rst), .Q(sreg[1950])
         );
  DFF \sreg_reg[1951]  ( .D(swire[929]), .CLK(clk), .RST(rst), .Q(sreg[1951])
         );
  DFF \sreg_reg[1952]  ( .D(swire[930]), .CLK(clk), .RST(rst), .Q(sreg[1952])
         );
  DFF \sreg_reg[1953]  ( .D(swire[931]), .CLK(clk), .RST(rst), .Q(sreg[1953])
         );
  DFF \sreg_reg[1954]  ( .D(swire[932]), .CLK(clk), .RST(rst), .Q(sreg[1954])
         );
  DFF \sreg_reg[1955]  ( .D(swire[933]), .CLK(clk), .RST(rst), .Q(sreg[1955])
         );
  DFF \sreg_reg[1956]  ( .D(swire[934]), .CLK(clk), .RST(rst), .Q(sreg[1956])
         );
  DFF \sreg_reg[1957]  ( .D(swire[935]), .CLK(clk), .RST(rst), .Q(sreg[1957])
         );
  DFF \sreg_reg[1958]  ( .D(swire[936]), .CLK(clk), .RST(rst), .Q(sreg[1958])
         );
  DFF \sreg_reg[1959]  ( .D(swire[937]), .CLK(clk), .RST(rst), .Q(sreg[1959])
         );
  DFF \sreg_reg[1960]  ( .D(swire[938]), .CLK(clk), .RST(rst), .Q(sreg[1960])
         );
  DFF \sreg_reg[1961]  ( .D(swire[939]), .CLK(clk), .RST(rst), .Q(sreg[1961])
         );
  DFF \sreg_reg[1962]  ( .D(swire[940]), .CLK(clk), .RST(rst), .Q(sreg[1962])
         );
  DFF \sreg_reg[1963]  ( .D(swire[941]), .CLK(clk), .RST(rst), .Q(sreg[1963])
         );
  DFF \sreg_reg[1964]  ( .D(swire[942]), .CLK(clk), .RST(rst), .Q(sreg[1964])
         );
  DFF \sreg_reg[1965]  ( .D(swire[943]), .CLK(clk), .RST(rst), .Q(sreg[1965])
         );
  DFF \sreg_reg[1966]  ( .D(swire[944]), .CLK(clk), .RST(rst), .Q(sreg[1966])
         );
  DFF \sreg_reg[1967]  ( .D(swire[945]), .CLK(clk), .RST(rst), .Q(sreg[1967])
         );
  DFF \sreg_reg[1968]  ( .D(swire[946]), .CLK(clk), .RST(rst), .Q(sreg[1968])
         );
  DFF \sreg_reg[1969]  ( .D(swire[947]), .CLK(clk), .RST(rst), .Q(sreg[1969])
         );
  DFF \sreg_reg[1970]  ( .D(swire[948]), .CLK(clk), .RST(rst), .Q(sreg[1970])
         );
  DFF \sreg_reg[1971]  ( .D(swire[949]), .CLK(clk), .RST(rst), .Q(sreg[1971])
         );
  DFF \sreg_reg[1972]  ( .D(swire[950]), .CLK(clk), .RST(rst), .Q(sreg[1972])
         );
  DFF \sreg_reg[1973]  ( .D(swire[951]), .CLK(clk), .RST(rst), .Q(sreg[1973])
         );
  DFF \sreg_reg[1974]  ( .D(swire[952]), .CLK(clk), .RST(rst), .Q(sreg[1974])
         );
  DFF \sreg_reg[1975]  ( .D(swire[953]), .CLK(clk), .RST(rst), .Q(sreg[1975])
         );
  DFF \sreg_reg[1976]  ( .D(swire[954]), .CLK(clk), .RST(rst), .Q(sreg[1976])
         );
  DFF \sreg_reg[1977]  ( .D(swire[955]), .CLK(clk), .RST(rst), .Q(sreg[1977])
         );
  DFF \sreg_reg[1978]  ( .D(swire[956]), .CLK(clk), .RST(rst), .Q(sreg[1978])
         );
  DFF \sreg_reg[1979]  ( .D(swire[957]), .CLK(clk), .RST(rst), .Q(sreg[1979])
         );
  DFF \sreg_reg[1980]  ( .D(swire[958]), .CLK(clk), .RST(rst), .Q(sreg[1980])
         );
  DFF \sreg_reg[1981]  ( .D(swire[959]), .CLK(clk), .RST(rst), .Q(sreg[1981])
         );
  DFF \sreg_reg[1982]  ( .D(swire[960]), .CLK(clk), .RST(rst), .Q(sreg[1982])
         );
  DFF \sreg_reg[1983]  ( .D(swire[961]), .CLK(clk), .RST(rst), .Q(sreg[1983])
         );
  DFF \sreg_reg[1984]  ( .D(swire[962]), .CLK(clk), .RST(rst), .Q(sreg[1984])
         );
  DFF \sreg_reg[1985]  ( .D(swire[963]), .CLK(clk), .RST(rst), .Q(sreg[1985])
         );
  DFF \sreg_reg[1986]  ( .D(swire[964]), .CLK(clk), .RST(rst), .Q(sreg[1986])
         );
  DFF \sreg_reg[1987]  ( .D(swire[965]), .CLK(clk), .RST(rst), .Q(sreg[1987])
         );
  DFF \sreg_reg[1988]  ( .D(swire[966]), .CLK(clk), .RST(rst), .Q(sreg[1988])
         );
  DFF \sreg_reg[1989]  ( .D(swire[967]), .CLK(clk), .RST(rst), .Q(sreg[1989])
         );
  DFF \sreg_reg[1990]  ( .D(swire[968]), .CLK(clk), .RST(rst), .Q(sreg[1990])
         );
  DFF \sreg_reg[1991]  ( .D(swire[969]), .CLK(clk), .RST(rst), .Q(sreg[1991])
         );
  DFF \sreg_reg[1992]  ( .D(swire[970]), .CLK(clk), .RST(rst), .Q(sreg[1992])
         );
  DFF \sreg_reg[1993]  ( .D(swire[971]), .CLK(clk), .RST(rst), .Q(sreg[1993])
         );
  DFF \sreg_reg[1994]  ( .D(swire[972]), .CLK(clk), .RST(rst), .Q(sreg[1994])
         );
  DFF \sreg_reg[1995]  ( .D(swire[973]), .CLK(clk), .RST(rst), .Q(sreg[1995])
         );
  DFF \sreg_reg[1996]  ( .D(swire[974]), .CLK(clk), .RST(rst), .Q(sreg[1996])
         );
  DFF \sreg_reg[1997]  ( .D(swire[975]), .CLK(clk), .RST(rst), .Q(sreg[1997])
         );
  DFF \sreg_reg[1998]  ( .D(swire[976]), .CLK(clk), .RST(rst), .Q(sreg[1998])
         );
  DFF \sreg_reg[1999]  ( .D(swire[977]), .CLK(clk), .RST(rst), .Q(sreg[1999])
         );
  DFF \sreg_reg[2000]  ( .D(swire[978]), .CLK(clk), .RST(rst), .Q(sreg[2000])
         );
  DFF \sreg_reg[2001]  ( .D(swire[979]), .CLK(clk), .RST(rst), .Q(sreg[2001])
         );
  DFF \sreg_reg[2002]  ( .D(swire[980]), .CLK(clk), .RST(rst), .Q(sreg[2002])
         );
  DFF \sreg_reg[2003]  ( .D(swire[981]), .CLK(clk), .RST(rst), .Q(sreg[2003])
         );
  DFF \sreg_reg[2004]  ( .D(swire[982]), .CLK(clk), .RST(rst), .Q(sreg[2004])
         );
  DFF \sreg_reg[2005]  ( .D(swire[983]), .CLK(clk), .RST(rst), .Q(sreg[2005])
         );
  DFF \sreg_reg[2006]  ( .D(swire[984]), .CLK(clk), .RST(rst), .Q(sreg[2006])
         );
  DFF \sreg_reg[2007]  ( .D(swire[985]), .CLK(clk), .RST(rst), .Q(sreg[2007])
         );
  DFF \sreg_reg[2008]  ( .D(swire[986]), .CLK(clk), .RST(rst), .Q(sreg[2008])
         );
  DFF \sreg_reg[2009]  ( .D(swire[987]), .CLK(clk), .RST(rst), .Q(sreg[2009])
         );
  DFF \sreg_reg[2010]  ( .D(swire[988]), .CLK(clk), .RST(rst), .Q(sreg[2010])
         );
  DFF \sreg_reg[2011]  ( .D(swire[989]), .CLK(clk), .RST(rst), .Q(sreg[2011])
         );
  DFF \sreg_reg[2012]  ( .D(swire[990]), .CLK(clk), .RST(rst), .Q(sreg[2012])
         );
  DFF \sreg_reg[2013]  ( .D(swire[991]), .CLK(clk), .RST(rst), .Q(sreg[2013])
         );
  DFF \sreg_reg[2014]  ( .D(swire[992]), .CLK(clk), .RST(rst), .Q(sreg[2014])
         );
  DFF \sreg_reg[2015]  ( .D(swire[993]), .CLK(clk), .RST(rst), .Q(sreg[2015])
         );
  DFF \sreg_reg[2016]  ( .D(swire[994]), .CLK(clk), .RST(rst), .Q(sreg[2016])
         );
  DFF \sreg_reg[2017]  ( .D(swire[995]), .CLK(clk), .RST(rst), .Q(sreg[2017])
         );
  DFF \sreg_reg[2018]  ( .D(swire[996]), .CLK(clk), .RST(rst), .Q(sreg[2018])
         );
  DFF \sreg_reg[2019]  ( .D(swire[997]), .CLK(clk), .RST(rst), .Q(sreg[2019])
         );
  DFF \sreg_reg[2020]  ( .D(swire[998]), .CLK(clk), .RST(rst), .Q(sreg[2020])
         );
  DFF \sreg_reg[2021]  ( .D(swire[999]), .CLK(clk), .RST(rst), .Q(sreg[2021])
         );
  DFF \sreg_reg[2022]  ( .D(swire[1000]), .CLK(clk), .RST(rst), .Q(sreg[2022])
         );
  DFF \sreg_reg[2023]  ( .D(swire[1001]), .CLK(clk), .RST(rst), .Q(sreg[2023])
         );
  DFF \sreg_reg[2024]  ( .D(swire[1002]), .CLK(clk), .RST(rst), .Q(sreg[2024])
         );
  DFF \sreg_reg[2025]  ( .D(swire[1003]), .CLK(clk), .RST(rst), .Q(sreg[2025])
         );
  DFF \sreg_reg[2026]  ( .D(swire[1004]), .CLK(clk), .RST(rst), .Q(sreg[2026])
         );
  DFF \sreg_reg[2027]  ( .D(swire[1005]), .CLK(clk), .RST(rst), .Q(sreg[2027])
         );
  DFF \sreg_reg[2028]  ( .D(swire[1006]), .CLK(clk), .RST(rst), .Q(sreg[2028])
         );
  DFF \sreg_reg[2029]  ( .D(swire[1007]), .CLK(clk), .RST(rst), .Q(sreg[2029])
         );
  DFF \sreg_reg[2030]  ( .D(swire[1008]), .CLK(clk), .RST(rst), .Q(sreg[2030])
         );
  DFF \sreg_reg[2031]  ( .D(swire[1009]), .CLK(clk), .RST(rst), .Q(sreg[2031])
         );
  DFF \sreg_reg[2032]  ( .D(swire[1010]), .CLK(clk), .RST(rst), .Q(sreg[2032])
         );
  DFF \sreg_reg[2033]  ( .D(swire[1011]), .CLK(clk), .RST(rst), .Q(sreg[2033])
         );
  DFF \sreg_reg[2034]  ( .D(swire[1012]), .CLK(clk), .RST(rst), .Q(sreg[2034])
         );
  DFF \sreg_reg[2035]  ( .D(swire[1013]), .CLK(clk), .RST(rst), .Q(sreg[2035])
         );
  DFF \sreg_reg[2036]  ( .D(swire[1014]), .CLK(clk), .RST(rst), .Q(sreg[2036])
         );
  DFF \sreg_reg[2037]  ( .D(swire[1015]), .CLK(clk), .RST(rst), .Q(sreg[2037])
         );
  DFF \sreg_reg[2038]  ( .D(swire[1016]), .CLK(clk), .RST(rst), .Q(sreg[2038])
         );
  DFF \sreg_reg[2039]  ( .D(swire[1017]), .CLK(clk), .RST(rst), .Q(sreg[2039])
         );
  DFF \sreg_reg[2040]  ( .D(swire[1018]), .CLK(clk), .RST(rst), .Q(sreg[2040])
         );
  DFF \sreg_reg[2041]  ( .D(swire[1019]), .CLK(clk), .RST(rst), .Q(sreg[2041])
         );
  DFF \sreg_reg[2042]  ( .D(swire[1020]), .CLK(clk), .RST(rst), .Q(sreg[2042])
         );
  DFF \sreg_reg[2043]  ( .D(swire[1021]), .CLK(clk), .RST(rst), .Q(sreg[2043])
         );
  DFF \sreg_reg[2044]  ( .D(swire[1022]), .CLK(clk), .RST(rst), .Q(sreg[2044])
         );
  DFF \sreg_reg[2045]  ( .D(swire[1023]), .CLK(clk), .RST(rst), .Q(sreg[2045])
         );
  DFF \sreg_reg[1023]  ( .D(c[1023]), .CLK(clk), .RST(rst), .Q(c[1021]) );
  DFF \sreg_reg[1022]  ( .D(c[1022]), .CLK(clk), .RST(rst), .Q(c[1020]) );
  DFF \sreg_reg[1021]  ( .D(c[1021]), .CLK(clk), .RST(rst), .Q(c[1019]) );
  DFF \sreg_reg[1020]  ( .D(c[1020]), .CLK(clk), .RST(rst), .Q(c[1018]) );
  DFF \sreg_reg[1019]  ( .D(c[1019]), .CLK(clk), .RST(rst), .Q(c[1017]) );
  DFF \sreg_reg[1018]  ( .D(c[1018]), .CLK(clk), .RST(rst), .Q(c[1016]) );
  DFF \sreg_reg[1017]  ( .D(c[1017]), .CLK(clk), .RST(rst), .Q(c[1015]) );
  DFF \sreg_reg[1016]  ( .D(c[1016]), .CLK(clk), .RST(rst), .Q(c[1014]) );
  DFF \sreg_reg[1015]  ( .D(c[1015]), .CLK(clk), .RST(rst), .Q(c[1013]) );
  DFF \sreg_reg[1014]  ( .D(c[1014]), .CLK(clk), .RST(rst), .Q(c[1012]) );
  DFF \sreg_reg[1013]  ( .D(c[1013]), .CLK(clk), .RST(rst), .Q(c[1011]) );
  DFF \sreg_reg[1012]  ( .D(c[1012]), .CLK(clk), .RST(rst), .Q(c[1010]) );
  DFF \sreg_reg[1011]  ( .D(c[1011]), .CLK(clk), .RST(rst), .Q(c[1009]) );
  DFF \sreg_reg[1010]  ( .D(c[1010]), .CLK(clk), .RST(rst), .Q(c[1008]) );
  DFF \sreg_reg[1009]  ( .D(c[1009]), .CLK(clk), .RST(rst), .Q(c[1007]) );
  DFF \sreg_reg[1008]  ( .D(c[1008]), .CLK(clk), .RST(rst), .Q(c[1006]) );
  DFF \sreg_reg[1007]  ( .D(c[1007]), .CLK(clk), .RST(rst), .Q(c[1005]) );
  DFF \sreg_reg[1006]  ( .D(c[1006]), .CLK(clk), .RST(rst), .Q(c[1004]) );
  DFF \sreg_reg[1005]  ( .D(c[1005]), .CLK(clk), .RST(rst), .Q(c[1003]) );
  DFF \sreg_reg[1004]  ( .D(c[1004]), .CLK(clk), .RST(rst), .Q(c[1002]) );
  DFF \sreg_reg[1003]  ( .D(c[1003]), .CLK(clk), .RST(rst), .Q(c[1001]) );
  DFF \sreg_reg[1002]  ( .D(c[1002]), .CLK(clk), .RST(rst), .Q(c[1000]) );
  DFF \sreg_reg[1001]  ( .D(c[1001]), .CLK(clk), .RST(rst), .Q(c[999]) );
  DFF \sreg_reg[1000]  ( .D(c[1000]), .CLK(clk), .RST(rst), .Q(c[998]) );
  DFF \sreg_reg[999]  ( .D(c[999]), .CLK(clk), .RST(rst), .Q(c[997]) );
  DFF \sreg_reg[998]  ( .D(c[998]), .CLK(clk), .RST(rst), .Q(c[996]) );
  DFF \sreg_reg[997]  ( .D(c[997]), .CLK(clk), .RST(rst), .Q(c[995]) );
  DFF \sreg_reg[996]  ( .D(c[996]), .CLK(clk), .RST(rst), .Q(c[994]) );
  DFF \sreg_reg[995]  ( .D(c[995]), .CLK(clk), .RST(rst), .Q(c[993]) );
  DFF \sreg_reg[994]  ( .D(c[994]), .CLK(clk), .RST(rst), .Q(c[992]) );
  DFF \sreg_reg[993]  ( .D(c[993]), .CLK(clk), .RST(rst), .Q(c[991]) );
  DFF \sreg_reg[992]  ( .D(c[992]), .CLK(clk), .RST(rst), .Q(c[990]) );
  DFF \sreg_reg[991]  ( .D(c[991]), .CLK(clk), .RST(rst), .Q(c[989]) );
  DFF \sreg_reg[990]  ( .D(c[990]), .CLK(clk), .RST(rst), .Q(c[988]) );
  DFF \sreg_reg[989]  ( .D(c[989]), .CLK(clk), .RST(rst), .Q(c[987]) );
  DFF \sreg_reg[988]  ( .D(c[988]), .CLK(clk), .RST(rst), .Q(c[986]) );
  DFF \sreg_reg[987]  ( .D(c[987]), .CLK(clk), .RST(rst), .Q(c[985]) );
  DFF \sreg_reg[986]  ( .D(c[986]), .CLK(clk), .RST(rst), .Q(c[984]) );
  DFF \sreg_reg[985]  ( .D(c[985]), .CLK(clk), .RST(rst), .Q(c[983]) );
  DFF \sreg_reg[984]  ( .D(c[984]), .CLK(clk), .RST(rst), .Q(c[982]) );
  DFF \sreg_reg[983]  ( .D(c[983]), .CLK(clk), .RST(rst), .Q(c[981]) );
  DFF \sreg_reg[982]  ( .D(c[982]), .CLK(clk), .RST(rst), .Q(c[980]) );
  DFF \sreg_reg[981]  ( .D(c[981]), .CLK(clk), .RST(rst), .Q(c[979]) );
  DFF \sreg_reg[980]  ( .D(c[980]), .CLK(clk), .RST(rst), .Q(c[978]) );
  DFF \sreg_reg[979]  ( .D(c[979]), .CLK(clk), .RST(rst), .Q(c[977]) );
  DFF \sreg_reg[978]  ( .D(c[978]), .CLK(clk), .RST(rst), .Q(c[976]) );
  DFF \sreg_reg[977]  ( .D(c[977]), .CLK(clk), .RST(rst), .Q(c[975]) );
  DFF \sreg_reg[976]  ( .D(c[976]), .CLK(clk), .RST(rst), .Q(c[974]) );
  DFF \sreg_reg[975]  ( .D(c[975]), .CLK(clk), .RST(rst), .Q(c[973]) );
  DFF \sreg_reg[974]  ( .D(c[974]), .CLK(clk), .RST(rst), .Q(c[972]) );
  DFF \sreg_reg[973]  ( .D(c[973]), .CLK(clk), .RST(rst), .Q(c[971]) );
  DFF \sreg_reg[972]  ( .D(c[972]), .CLK(clk), .RST(rst), .Q(c[970]) );
  DFF \sreg_reg[971]  ( .D(c[971]), .CLK(clk), .RST(rst), .Q(c[969]) );
  DFF \sreg_reg[970]  ( .D(c[970]), .CLK(clk), .RST(rst), .Q(c[968]) );
  DFF \sreg_reg[969]  ( .D(c[969]), .CLK(clk), .RST(rst), .Q(c[967]) );
  DFF \sreg_reg[968]  ( .D(c[968]), .CLK(clk), .RST(rst), .Q(c[966]) );
  DFF \sreg_reg[967]  ( .D(c[967]), .CLK(clk), .RST(rst), .Q(c[965]) );
  DFF \sreg_reg[966]  ( .D(c[966]), .CLK(clk), .RST(rst), .Q(c[964]) );
  DFF \sreg_reg[965]  ( .D(c[965]), .CLK(clk), .RST(rst), .Q(c[963]) );
  DFF \sreg_reg[964]  ( .D(c[964]), .CLK(clk), .RST(rst), .Q(c[962]) );
  DFF \sreg_reg[963]  ( .D(c[963]), .CLK(clk), .RST(rst), .Q(c[961]) );
  DFF \sreg_reg[962]  ( .D(c[962]), .CLK(clk), .RST(rst), .Q(c[960]) );
  DFF \sreg_reg[961]  ( .D(c[961]), .CLK(clk), .RST(rst), .Q(c[959]) );
  DFF \sreg_reg[960]  ( .D(c[960]), .CLK(clk), .RST(rst), .Q(c[958]) );
  DFF \sreg_reg[959]  ( .D(c[959]), .CLK(clk), .RST(rst), .Q(c[957]) );
  DFF \sreg_reg[958]  ( .D(c[958]), .CLK(clk), .RST(rst), .Q(c[956]) );
  DFF \sreg_reg[957]  ( .D(c[957]), .CLK(clk), .RST(rst), .Q(c[955]) );
  DFF \sreg_reg[956]  ( .D(c[956]), .CLK(clk), .RST(rst), .Q(c[954]) );
  DFF \sreg_reg[955]  ( .D(c[955]), .CLK(clk), .RST(rst), .Q(c[953]) );
  DFF \sreg_reg[954]  ( .D(c[954]), .CLK(clk), .RST(rst), .Q(c[952]) );
  DFF \sreg_reg[953]  ( .D(c[953]), .CLK(clk), .RST(rst), .Q(c[951]) );
  DFF \sreg_reg[952]  ( .D(c[952]), .CLK(clk), .RST(rst), .Q(c[950]) );
  DFF \sreg_reg[951]  ( .D(c[951]), .CLK(clk), .RST(rst), .Q(c[949]) );
  DFF \sreg_reg[950]  ( .D(c[950]), .CLK(clk), .RST(rst), .Q(c[948]) );
  DFF \sreg_reg[949]  ( .D(c[949]), .CLK(clk), .RST(rst), .Q(c[947]) );
  DFF \sreg_reg[948]  ( .D(c[948]), .CLK(clk), .RST(rst), .Q(c[946]) );
  DFF \sreg_reg[947]  ( .D(c[947]), .CLK(clk), .RST(rst), .Q(c[945]) );
  DFF \sreg_reg[946]  ( .D(c[946]), .CLK(clk), .RST(rst), .Q(c[944]) );
  DFF \sreg_reg[945]  ( .D(c[945]), .CLK(clk), .RST(rst), .Q(c[943]) );
  DFF \sreg_reg[944]  ( .D(c[944]), .CLK(clk), .RST(rst), .Q(c[942]) );
  DFF \sreg_reg[943]  ( .D(c[943]), .CLK(clk), .RST(rst), .Q(c[941]) );
  DFF \sreg_reg[942]  ( .D(c[942]), .CLK(clk), .RST(rst), .Q(c[940]) );
  DFF \sreg_reg[941]  ( .D(c[941]), .CLK(clk), .RST(rst), .Q(c[939]) );
  DFF \sreg_reg[940]  ( .D(c[940]), .CLK(clk), .RST(rst), .Q(c[938]) );
  DFF \sreg_reg[939]  ( .D(c[939]), .CLK(clk), .RST(rst), .Q(c[937]) );
  DFF \sreg_reg[938]  ( .D(c[938]), .CLK(clk), .RST(rst), .Q(c[936]) );
  DFF \sreg_reg[937]  ( .D(c[937]), .CLK(clk), .RST(rst), .Q(c[935]) );
  DFF \sreg_reg[936]  ( .D(c[936]), .CLK(clk), .RST(rst), .Q(c[934]) );
  DFF \sreg_reg[935]  ( .D(c[935]), .CLK(clk), .RST(rst), .Q(c[933]) );
  DFF \sreg_reg[934]  ( .D(c[934]), .CLK(clk), .RST(rst), .Q(c[932]) );
  DFF \sreg_reg[933]  ( .D(c[933]), .CLK(clk), .RST(rst), .Q(c[931]) );
  DFF \sreg_reg[932]  ( .D(c[932]), .CLK(clk), .RST(rst), .Q(c[930]) );
  DFF \sreg_reg[931]  ( .D(c[931]), .CLK(clk), .RST(rst), .Q(c[929]) );
  DFF \sreg_reg[930]  ( .D(c[930]), .CLK(clk), .RST(rst), .Q(c[928]) );
  DFF \sreg_reg[929]  ( .D(c[929]), .CLK(clk), .RST(rst), .Q(c[927]) );
  DFF \sreg_reg[928]  ( .D(c[928]), .CLK(clk), .RST(rst), .Q(c[926]) );
  DFF \sreg_reg[927]  ( .D(c[927]), .CLK(clk), .RST(rst), .Q(c[925]) );
  DFF \sreg_reg[926]  ( .D(c[926]), .CLK(clk), .RST(rst), .Q(c[924]) );
  DFF \sreg_reg[925]  ( .D(c[925]), .CLK(clk), .RST(rst), .Q(c[923]) );
  DFF \sreg_reg[924]  ( .D(c[924]), .CLK(clk), .RST(rst), .Q(c[922]) );
  DFF \sreg_reg[923]  ( .D(c[923]), .CLK(clk), .RST(rst), .Q(c[921]) );
  DFF \sreg_reg[922]  ( .D(c[922]), .CLK(clk), .RST(rst), .Q(c[920]) );
  DFF \sreg_reg[921]  ( .D(c[921]), .CLK(clk), .RST(rst), .Q(c[919]) );
  DFF \sreg_reg[920]  ( .D(c[920]), .CLK(clk), .RST(rst), .Q(c[918]) );
  DFF \sreg_reg[919]  ( .D(c[919]), .CLK(clk), .RST(rst), .Q(c[917]) );
  DFF \sreg_reg[918]  ( .D(c[918]), .CLK(clk), .RST(rst), .Q(c[916]) );
  DFF \sreg_reg[917]  ( .D(c[917]), .CLK(clk), .RST(rst), .Q(c[915]) );
  DFF \sreg_reg[916]  ( .D(c[916]), .CLK(clk), .RST(rst), .Q(c[914]) );
  DFF \sreg_reg[915]  ( .D(c[915]), .CLK(clk), .RST(rst), .Q(c[913]) );
  DFF \sreg_reg[914]  ( .D(c[914]), .CLK(clk), .RST(rst), .Q(c[912]) );
  DFF \sreg_reg[913]  ( .D(c[913]), .CLK(clk), .RST(rst), .Q(c[911]) );
  DFF \sreg_reg[912]  ( .D(c[912]), .CLK(clk), .RST(rst), .Q(c[910]) );
  DFF \sreg_reg[911]  ( .D(c[911]), .CLK(clk), .RST(rst), .Q(c[909]) );
  DFF \sreg_reg[910]  ( .D(c[910]), .CLK(clk), .RST(rst), .Q(c[908]) );
  DFF \sreg_reg[909]  ( .D(c[909]), .CLK(clk), .RST(rst), .Q(c[907]) );
  DFF \sreg_reg[908]  ( .D(c[908]), .CLK(clk), .RST(rst), .Q(c[906]) );
  DFF \sreg_reg[907]  ( .D(c[907]), .CLK(clk), .RST(rst), .Q(c[905]) );
  DFF \sreg_reg[906]  ( .D(c[906]), .CLK(clk), .RST(rst), .Q(c[904]) );
  DFF \sreg_reg[905]  ( .D(c[905]), .CLK(clk), .RST(rst), .Q(c[903]) );
  DFF \sreg_reg[904]  ( .D(c[904]), .CLK(clk), .RST(rst), .Q(c[902]) );
  DFF \sreg_reg[903]  ( .D(c[903]), .CLK(clk), .RST(rst), .Q(c[901]) );
  DFF \sreg_reg[902]  ( .D(c[902]), .CLK(clk), .RST(rst), .Q(c[900]) );
  DFF \sreg_reg[901]  ( .D(c[901]), .CLK(clk), .RST(rst), .Q(c[899]) );
  DFF \sreg_reg[900]  ( .D(c[900]), .CLK(clk), .RST(rst), .Q(c[898]) );
  DFF \sreg_reg[899]  ( .D(c[899]), .CLK(clk), .RST(rst), .Q(c[897]) );
  DFF \sreg_reg[898]  ( .D(c[898]), .CLK(clk), .RST(rst), .Q(c[896]) );
  DFF \sreg_reg[897]  ( .D(c[897]), .CLK(clk), .RST(rst), .Q(c[895]) );
  DFF \sreg_reg[896]  ( .D(c[896]), .CLK(clk), .RST(rst), .Q(c[894]) );
  DFF \sreg_reg[895]  ( .D(c[895]), .CLK(clk), .RST(rst), .Q(c[893]) );
  DFF \sreg_reg[894]  ( .D(c[894]), .CLK(clk), .RST(rst), .Q(c[892]) );
  DFF \sreg_reg[893]  ( .D(c[893]), .CLK(clk), .RST(rst), .Q(c[891]) );
  DFF \sreg_reg[892]  ( .D(c[892]), .CLK(clk), .RST(rst), .Q(c[890]) );
  DFF \sreg_reg[891]  ( .D(c[891]), .CLK(clk), .RST(rst), .Q(c[889]) );
  DFF \sreg_reg[890]  ( .D(c[890]), .CLK(clk), .RST(rst), .Q(c[888]) );
  DFF \sreg_reg[889]  ( .D(c[889]), .CLK(clk), .RST(rst), .Q(c[887]) );
  DFF \sreg_reg[888]  ( .D(c[888]), .CLK(clk), .RST(rst), .Q(c[886]) );
  DFF \sreg_reg[887]  ( .D(c[887]), .CLK(clk), .RST(rst), .Q(c[885]) );
  DFF \sreg_reg[886]  ( .D(c[886]), .CLK(clk), .RST(rst), .Q(c[884]) );
  DFF \sreg_reg[885]  ( .D(c[885]), .CLK(clk), .RST(rst), .Q(c[883]) );
  DFF \sreg_reg[884]  ( .D(c[884]), .CLK(clk), .RST(rst), .Q(c[882]) );
  DFF \sreg_reg[883]  ( .D(c[883]), .CLK(clk), .RST(rst), .Q(c[881]) );
  DFF \sreg_reg[882]  ( .D(c[882]), .CLK(clk), .RST(rst), .Q(c[880]) );
  DFF \sreg_reg[881]  ( .D(c[881]), .CLK(clk), .RST(rst), .Q(c[879]) );
  DFF \sreg_reg[880]  ( .D(c[880]), .CLK(clk), .RST(rst), .Q(c[878]) );
  DFF \sreg_reg[879]  ( .D(c[879]), .CLK(clk), .RST(rst), .Q(c[877]) );
  DFF \sreg_reg[878]  ( .D(c[878]), .CLK(clk), .RST(rst), .Q(c[876]) );
  DFF \sreg_reg[877]  ( .D(c[877]), .CLK(clk), .RST(rst), .Q(c[875]) );
  DFF \sreg_reg[876]  ( .D(c[876]), .CLK(clk), .RST(rst), .Q(c[874]) );
  DFF \sreg_reg[875]  ( .D(c[875]), .CLK(clk), .RST(rst), .Q(c[873]) );
  DFF \sreg_reg[874]  ( .D(c[874]), .CLK(clk), .RST(rst), .Q(c[872]) );
  DFF \sreg_reg[873]  ( .D(c[873]), .CLK(clk), .RST(rst), .Q(c[871]) );
  DFF \sreg_reg[872]  ( .D(c[872]), .CLK(clk), .RST(rst), .Q(c[870]) );
  DFF \sreg_reg[871]  ( .D(c[871]), .CLK(clk), .RST(rst), .Q(c[869]) );
  DFF \sreg_reg[870]  ( .D(c[870]), .CLK(clk), .RST(rst), .Q(c[868]) );
  DFF \sreg_reg[869]  ( .D(c[869]), .CLK(clk), .RST(rst), .Q(c[867]) );
  DFF \sreg_reg[868]  ( .D(c[868]), .CLK(clk), .RST(rst), .Q(c[866]) );
  DFF \sreg_reg[867]  ( .D(c[867]), .CLK(clk), .RST(rst), .Q(c[865]) );
  DFF \sreg_reg[866]  ( .D(c[866]), .CLK(clk), .RST(rst), .Q(c[864]) );
  DFF \sreg_reg[865]  ( .D(c[865]), .CLK(clk), .RST(rst), .Q(c[863]) );
  DFF \sreg_reg[864]  ( .D(c[864]), .CLK(clk), .RST(rst), .Q(c[862]) );
  DFF \sreg_reg[863]  ( .D(c[863]), .CLK(clk), .RST(rst), .Q(c[861]) );
  DFF \sreg_reg[862]  ( .D(c[862]), .CLK(clk), .RST(rst), .Q(c[860]) );
  DFF \sreg_reg[861]  ( .D(c[861]), .CLK(clk), .RST(rst), .Q(c[859]) );
  DFF \sreg_reg[860]  ( .D(c[860]), .CLK(clk), .RST(rst), .Q(c[858]) );
  DFF \sreg_reg[859]  ( .D(c[859]), .CLK(clk), .RST(rst), .Q(c[857]) );
  DFF \sreg_reg[858]  ( .D(c[858]), .CLK(clk), .RST(rst), .Q(c[856]) );
  DFF \sreg_reg[857]  ( .D(c[857]), .CLK(clk), .RST(rst), .Q(c[855]) );
  DFF \sreg_reg[856]  ( .D(c[856]), .CLK(clk), .RST(rst), .Q(c[854]) );
  DFF \sreg_reg[855]  ( .D(c[855]), .CLK(clk), .RST(rst), .Q(c[853]) );
  DFF \sreg_reg[854]  ( .D(c[854]), .CLK(clk), .RST(rst), .Q(c[852]) );
  DFF \sreg_reg[853]  ( .D(c[853]), .CLK(clk), .RST(rst), .Q(c[851]) );
  DFF \sreg_reg[852]  ( .D(c[852]), .CLK(clk), .RST(rst), .Q(c[850]) );
  DFF \sreg_reg[851]  ( .D(c[851]), .CLK(clk), .RST(rst), .Q(c[849]) );
  DFF \sreg_reg[850]  ( .D(c[850]), .CLK(clk), .RST(rst), .Q(c[848]) );
  DFF \sreg_reg[849]  ( .D(c[849]), .CLK(clk), .RST(rst), .Q(c[847]) );
  DFF \sreg_reg[848]  ( .D(c[848]), .CLK(clk), .RST(rst), .Q(c[846]) );
  DFF \sreg_reg[847]  ( .D(c[847]), .CLK(clk), .RST(rst), .Q(c[845]) );
  DFF \sreg_reg[846]  ( .D(c[846]), .CLK(clk), .RST(rst), .Q(c[844]) );
  DFF \sreg_reg[845]  ( .D(c[845]), .CLK(clk), .RST(rst), .Q(c[843]) );
  DFF \sreg_reg[844]  ( .D(c[844]), .CLK(clk), .RST(rst), .Q(c[842]) );
  DFF \sreg_reg[843]  ( .D(c[843]), .CLK(clk), .RST(rst), .Q(c[841]) );
  DFF \sreg_reg[842]  ( .D(c[842]), .CLK(clk), .RST(rst), .Q(c[840]) );
  DFF \sreg_reg[841]  ( .D(c[841]), .CLK(clk), .RST(rst), .Q(c[839]) );
  DFF \sreg_reg[840]  ( .D(c[840]), .CLK(clk), .RST(rst), .Q(c[838]) );
  DFF \sreg_reg[839]  ( .D(c[839]), .CLK(clk), .RST(rst), .Q(c[837]) );
  DFF \sreg_reg[838]  ( .D(c[838]), .CLK(clk), .RST(rst), .Q(c[836]) );
  DFF \sreg_reg[837]  ( .D(c[837]), .CLK(clk), .RST(rst), .Q(c[835]) );
  DFF \sreg_reg[836]  ( .D(c[836]), .CLK(clk), .RST(rst), .Q(c[834]) );
  DFF \sreg_reg[835]  ( .D(c[835]), .CLK(clk), .RST(rst), .Q(c[833]) );
  DFF \sreg_reg[834]  ( .D(c[834]), .CLK(clk), .RST(rst), .Q(c[832]) );
  DFF \sreg_reg[833]  ( .D(c[833]), .CLK(clk), .RST(rst), .Q(c[831]) );
  DFF \sreg_reg[832]  ( .D(c[832]), .CLK(clk), .RST(rst), .Q(c[830]) );
  DFF \sreg_reg[831]  ( .D(c[831]), .CLK(clk), .RST(rst), .Q(c[829]) );
  DFF \sreg_reg[830]  ( .D(c[830]), .CLK(clk), .RST(rst), .Q(c[828]) );
  DFF \sreg_reg[829]  ( .D(c[829]), .CLK(clk), .RST(rst), .Q(c[827]) );
  DFF \sreg_reg[828]  ( .D(c[828]), .CLK(clk), .RST(rst), .Q(c[826]) );
  DFF \sreg_reg[827]  ( .D(c[827]), .CLK(clk), .RST(rst), .Q(c[825]) );
  DFF \sreg_reg[826]  ( .D(c[826]), .CLK(clk), .RST(rst), .Q(c[824]) );
  DFF \sreg_reg[825]  ( .D(c[825]), .CLK(clk), .RST(rst), .Q(c[823]) );
  DFF \sreg_reg[824]  ( .D(c[824]), .CLK(clk), .RST(rst), .Q(c[822]) );
  DFF \sreg_reg[823]  ( .D(c[823]), .CLK(clk), .RST(rst), .Q(c[821]) );
  DFF \sreg_reg[822]  ( .D(c[822]), .CLK(clk), .RST(rst), .Q(c[820]) );
  DFF \sreg_reg[821]  ( .D(c[821]), .CLK(clk), .RST(rst), .Q(c[819]) );
  DFF \sreg_reg[820]  ( .D(c[820]), .CLK(clk), .RST(rst), .Q(c[818]) );
  DFF \sreg_reg[819]  ( .D(c[819]), .CLK(clk), .RST(rst), .Q(c[817]) );
  DFF \sreg_reg[818]  ( .D(c[818]), .CLK(clk), .RST(rst), .Q(c[816]) );
  DFF \sreg_reg[817]  ( .D(c[817]), .CLK(clk), .RST(rst), .Q(c[815]) );
  DFF \sreg_reg[816]  ( .D(c[816]), .CLK(clk), .RST(rst), .Q(c[814]) );
  DFF \sreg_reg[815]  ( .D(c[815]), .CLK(clk), .RST(rst), .Q(c[813]) );
  DFF \sreg_reg[814]  ( .D(c[814]), .CLK(clk), .RST(rst), .Q(c[812]) );
  DFF \sreg_reg[813]  ( .D(c[813]), .CLK(clk), .RST(rst), .Q(c[811]) );
  DFF \sreg_reg[812]  ( .D(c[812]), .CLK(clk), .RST(rst), .Q(c[810]) );
  DFF \sreg_reg[811]  ( .D(c[811]), .CLK(clk), .RST(rst), .Q(c[809]) );
  DFF \sreg_reg[810]  ( .D(c[810]), .CLK(clk), .RST(rst), .Q(c[808]) );
  DFF \sreg_reg[809]  ( .D(c[809]), .CLK(clk), .RST(rst), .Q(c[807]) );
  DFF \sreg_reg[808]  ( .D(c[808]), .CLK(clk), .RST(rst), .Q(c[806]) );
  DFF \sreg_reg[807]  ( .D(c[807]), .CLK(clk), .RST(rst), .Q(c[805]) );
  DFF \sreg_reg[806]  ( .D(c[806]), .CLK(clk), .RST(rst), .Q(c[804]) );
  DFF \sreg_reg[805]  ( .D(c[805]), .CLK(clk), .RST(rst), .Q(c[803]) );
  DFF \sreg_reg[804]  ( .D(c[804]), .CLK(clk), .RST(rst), .Q(c[802]) );
  DFF \sreg_reg[803]  ( .D(c[803]), .CLK(clk), .RST(rst), .Q(c[801]) );
  DFF \sreg_reg[802]  ( .D(c[802]), .CLK(clk), .RST(rst), .Q(c[800]) );
  DFF \sreg_reg[801]  ( .D(c[801]), .CLK(clk), .RST(rst), .Q(c[799]) );
  DFF \sreg_reg[800]  ( .D(c[800]), .CLK(clk), .RST(rst), .Q(c[798]) );
  DFF \sreg_reg[799]  ( .D(c[799]), .CLK(clk), .RST(rst), .Q(c[797]) );
  DFF \sreg_reg[798]  ( .D(c[798]), .CLK(clk), .RST(rst), .Q(c[796]) );
  DFF \sreg_reg[797]  ( .D(c[797]), .CLK(clk), .RST(rst), .Q(c[795]) );
  DFF \sreg_reg[796]  ( .D(c[796]), .CLK(clk), .RST(rst), .Q(c[794]) );
  DFF \sreg_reg[795]  ( .D(c[795]), .CLK(clk), .RST(rst), .Q(c[793]) );
  DFF \sreg_reg[794]  ( .D(c[794]), .CLK(clk), .RST(rst), .Q(c[792]) );
  DFF \sreg_reg[793]  ( .D(c[793]), .CLK(clk), .RST(rst), .Q(c[791]) );
  DFF \sreg_reg[792]  ( .D(c[792]), .CLK(clk), .RST(rst), .Q(c[790]) );
  DFF \sreg_reg[791]  ( .D(c[791]), .CLK(clk), .RST(rst), .Q(c[789]) );
  DFF \sreg_reg[790]  ( .D(c[790]), .CLK(clk), .RST(rst), .Q(c[788]) );
  DFF \sreg_reg[789]  ( .D(c[789]), .CLK(clk), .RST(rst), .Q(c[787]) );
  DFF \sreg_reg[788]  ( .D(c[788]), .CLK(clk), .RST(rst), .Q(c[786]) );
  DFF \sreg_reg[787]  ( .D(c[787]), .CLK(clk), .RST(rst), .Q(c[785]) );
  DFF \sreg_reg[786]  ( .D(c[786]), .CLK(clk), .RST(rst), .Q(c[784]) );
  DFF \sreg_reg[785]  ( .D(c[785]), .CLK(clk), .RST(rst), .Q(c[783]) );
  DFF \sreg_reg[784]  ( .D(c[784]), .CLK(clk), .RST(rst), .Q(c[782]) );
  DFF \sreg_reg[783]  ( .D(c[783]), .CLK(clk), .RST(rst), .Q(c[781]) );
  DFF \sreg_reg[782]  ( .D(c[782]), .CLK(clk), .RST(rst), .Q(c[780]) );
  DFF \sreg_reg[781]  ( .D(c[781]), .CLK(clk), .RST(rst), .Q(c[779]) );
  DFF \sreg_reg[780]  ( .D(c[780]), .CLK(clk), .RST(rst), .Q(c[778]) );
  DFF \sreg_reg[779]  ( .D(c[779]), .CLK(clk), .RST(rst), .Q(c[777]) );
  DFF \sreg_reg[778]  ( .D(c[778]), .CLK(clk), .RST(rst), .Q(c[776]) );
  DFF \sreg_reg[777]  ( .D(c[777]), .CLK(clk), .RST(rst), .Q(c[775]) );
  DFF \sreg_reg[776]  ( .D(c[776]), .CLK(clk), .RST(rst), .Q(c[774]) );
  DFF \sreg_reg[775]  ( .D(c[775]), .CLK(clk), .RST(rst), .Q(c[773]) );
  DFF \sreg_reg[774]  ( .D(c[774]), .CLK(clk), .RST(rst), .Q(c[772]) );
  DFF \sreg_reg[773]  ( .D(c[773]), .CLK(clk), .RST(rst), .Q(c[771]) );
  DFF \sreg_reg[772]  ( .D(c[772]), .CLK(clk), .RST(rst), .Q(c[770]) );
  DFF \sreg_reg[771]  ( .D(c[771]), .CLK(clk), .RST(rst), .Q(c[769]) );
  DFF \sreg_reg[770]  ( .D(c[770]), .CLK(clk), .RST(rst), .Q(c[768]) );
  DFF \sreg_reg[769]  ( .D(c[769]), .CLK(clk), .RST(rst), .Q(c[767]) );
  DFF \sreg_reg[768]  ( .D(c[768]), .CLK(clk), .RST(rst), .Q(c[766]) );
  DFF \sreg_reg[767]  ( .D(c[767]), .CLK(clk), .RST(rst), .Q(c[765]) );
  DFF \sreg_reg[766]  ( .D(c[766]), .CLK(clk), .RST(rst), .Q(c[764]) );
  DFF \sreg_reg[765]  ( .D(c[765]), .CLK(clk), .RST(rst), .Q(c[763]) );
  DFF \sreg_reg[764]  ( .D(c[764]), .CLK(clk), .RST(rst), .Q(c[762]) );
  DFF \sreg_reg[763]  ( .D(c[763]), .CLK(clk), .RST(rst), .Q(c[761]) );
  DFF \sreg_reg[762]  ( .D(c[762]), .CLK(clk), .RST(rst), .Q(c[760]) );
  DFF \sreg_reg[761]  ( .D(c[761]), .CLK(clk), .RST(rst), .Q(c[759]) );
  DFF \sreg_reg[760]  ( .D(c[760]), .CLK(clk), .RST(rst), .Q(c[758]) );
  DFF \sreg_reg[759]  ( .D(c[759]), .CLK(clk), .RST(rst), .Q(c[757]) );
  DFF \sreg_reg[758]  ( .D(c[758]), .CLK(clk), .RST(rst), .Q(c[756]) );
  DFF \sreg_reg[757]  ( .D(c[757]), .CLK(clk), .RST(rst), .Q(c[755]) );
  DFF \sreg_reg[756]  ( .D(c[756]), .CLK(clk), .RST(rst), .Q(c[754]) );
  DFF \sreg_reg[755]  ( .D(c[755]), .CLK(clk), .RST(rst), .Q(c[753]) );
  DFF \sreg_reg[754]  ( .D(c[754]), .CLK(clk), .RST(rst), .Q(c[752]) );
  DFF \sreg_reg[753]  ( .D(c[753]), .CLK(clk), .RST(rst), .Q(c[751]) );
  DFF \sreg_reg[752]  ( .D(c[752]), .CLK(clk), .RST(rst), .Q(c[750]) );
  DFF \sreg_reg[751]  ( .D(c[751]), .CLK(clk), .RST(rst), .Q(c[749]) );
  DFF \sreg_reg[750]  ( .D(c[750]), .CLK(clk), .RST(rst), .Q(c[748]) );
  DFF \sreg_reg[749]  ( .D(c[749]), .CLK(clk), .RST(rst), .Q(c[747]) );
  DFF \sreg_reg[748]  ( .D(c[748]), .CLK(clk), .RST(rst), .Q(c[746]) );
  DFF \sreg_reg[747]  ( .D(c[747]), .CLK(clk), .RST(rst), .Q(c[745]) );
  DFF \sreg_reg[746]  ( .D(c[746]), .CLK(clk), .RST(rst), .Q(c[744]) );
  DFF \sreg_reg[745]  ( .D(c[745]), .CLK(clk), .RST(rst), .Q(c[743]) );
  DFF \sreg_reg[744]  ( .D(c[744]), .CLK(clk), .RST(rst), .Q(c[742]) );
  DFF \sreg_reg[743]  ( .D(c[743]), .CLK(clk), .RST(rst), .Q(c[741]) );
  DFF \sreg_reg[742]  ( .D(c[742]), .CLK(clk), .RST(rst), .Q(c[740]) );
  DFF \sreg_reg[741]  ( .D(c[741]), .CLK(clk), .RST(rst), .Q(c[739]) );
  DFF \sreg_reg[740]  ( .D(c[740]), .CLK(clk), .RST(rst), .Q(c[738]) );
  DFF \sreg_reg[739]  ( .D(c[739]), .CLK(clk), .RST(rst), .Q(c[737]) );
  DFF \sreg_reg[738]  ( .D(c[738]), .CLK(clk), .RST(rst), .Q(c[736]) );
  DFF \sreg_reg[737]  ( .D(c[737]), .CLK(clk), .RST(rst), .Q(c[735]) );
  DFF \sreg_reg[736]  ( .D(c[736]), .CLK(clk), .RST(rst), .Q(c[734]) );
  DFF \sreg_reg[735]  ( .D(c[735]), .CLK(clk), .RST(rst), .Q(c[733]) );
  DFF \sreg_reg[734]  ( .D(c[734]), .CLK(clk), .RST(rst), .Q(c[732]) );
  DFF \sreg_reg[733]  ( .D(c[733]), .CLK(clk), .RST(rst), .Q(c[731]) );
  DFF \sreg_reg[732]  ( .D(c[732]), .CLK(clk), .RST(rst), .Q(c[730]) );
  DFF \sreg_reg[731]  ( .D(c[731]), .CLK(clk), .RST(rst), .Q(c[729]) );
  DFF \sreg_reg[730]  ( .D(c[730]), .CLK(clk), .RST(rst), .Q(c[728]) );
  DFF \sreg_reg[729]  ( .D(c[729]), .CLK(clk), .RST(rst), .Q(c[727]) );
  DFF \sreg_reg[728]  ( .D(c[728]), .CLK(clk), .RST(rst), .Q(c[726]) );
  DFF \sreg_reg[727]  ( .D(c[727]), .CLK(clk), .RST(rst), .Q(c[725]) );
  DFF \sreg_reg[726]  ( .D(c[726]), .CLK(clk), .RST(rst), .Q(c[724]) );
  DFF \sreg_reg[725]  ( .D(c[725]), .CLK(clk), .RST(rst), .Q(c[723]) );
  DFF \sreg_reg[724]  ( .D(c[724]), .CLK(clk), .RST(rst), .Q(c[722]) );
  DFF \sreg_reg[723]  ( .D(c[723]), .CLK(clk), .RST(rst), .Q(c[721]) );
  DFF \sreg_reg[722]  ( .D(c[722]), .CLK(clk), .RST(rst), .Q(c[720]) );
  DFF \sreg_reg[721]  ( .D(c[721]), .CLK(clk), .RST(rst), .Q(c[719]) );
  DFF \sreg_reg[720]  ( .D(c[720]), .CLK(clk), .RST(rst), .Q(c[718]) );
  DFF \sreg_reg[719]  ( .D(c[719]), .CLK(clk), .RST(rst), .Q(c[717]) );
  DFF \sreg_reg[718]  ( .D(c[718]), .CLK(clk), .RST(rst), .Q(c[716]) );
  DFF \sreg_reg[717]  ( .D(c[717]), .CLK(clk), .RST(rst), .Q(c[715]) );
  DFF \sreg_reg[716]  ( .D(c[716]), .CLK(clk), .RST(rst), .Q(c[714]) );
  DFF \sreg_reg[715]  ( .D(c[715]), .CLK(clk), .RST(rst), .Q(c[713]) );
  DFF \sreg_reg[714]  ( .D(c[714]), .CLK(clk), .RST(rst), .Q(c[712]) );
  DFF \sreg_reg[713]  ( .D(c[713]), .CLK(clk), .RST(rst), .Q(c[711]) );
  DFF \sreg_reg[712]  ( .D(c[712]), .CLK(clk), .RST(rst), .Q(c[710]) );
  DFF \sreg_reg[711]  ( .D(c[711]), .CLK(clk), .RST(rst), .Q(c[709]) );
  DFF \sreg_reg[710]  ( .D(c[710]), .CLK(clk), .RST(rst), .Q(c[708]) );
  DFF \sreg_reg[709]  ( .D(c[709]), .CLK(clk), .RST(rst), .Q(c[707]) );
  DFF \sreg_reg[708]  ( .D(c[708]), .CLK(clk), .RST(rst), .Q(c[706]) );
  DFF \sreg_reg[707]  ( .D(c[707]), .CLK(clk), .RST(rst), .Q(c[705]) );
  DFF \sreg_reg[706]  ( .D(c[706]), .CLK(clk), .RST(rst), .Q(c[704]) );
  DFF \sreg_reg[705]  ( .D(c[705]), .CLK(clk), .RST(rst), .Q(c[703]) );
  DFF \sreg_reg[704]  ( .D(c[704]), .CLK(clk), .RST(rst), .Q(c[702]) );
  DFF \sreg_reg[703]  ( .D(c[703]), .CLK(clk), .RST(rst), .Q(c[701]) );
  DFF \sreg_reg[702]  ( .D(c[702]), .CLK(clk), .RST(rst), .Q(c[700]) );
  DFF \sreg_reg[701]  ( .D(c[701]), .CLK(clk), .RST(rst), .Q(c[699]) );
  DFF \sreg_reg[700]  ( .D(c[700]), .CLK(clk), .RST(rst), .Q(c[698]) );
  DFF \sreg_reg[699]  ( .D(c[699]), .CLK(clk), .RST(rst), .Q(c[697]) );
  DFF \sreg_reg[698]  ( .D(c[698]), .CLK(clk), .RST(rst), .Q(c[696]) );
  DFF \sreg_reg[697]  ( .D(c[697]), .CLK(clk), .RST(rst), .Q(c[695]) );
  DFF \sreg_reg[696]  ( .D(c[696]), .CLK(clk), .RST(rst), .Q(c[694]) );
  DFF \sreg_reg[695]  ( .D(c[695]), .CLK(clk), .RST(rst), .Q(c[693]) );
  DFF \sreg_reg[694]  ( .D(c[694]), .CLK(clk), .RST(rst), .Q(c[692]) );
  DFF \sreg_reg[693]  ( .D(c[693]), .CLK(clk), .RST(rst), .Q(c[691]) );
  DFF \sreg_reg[692]  ( .D(c[692]), .CLK(clk), .RST(rst), .Q(c[690]) );
  DFF \sreg_reg[691]  ( .D(c[691]), .CLK(clk), .RST(rst), .Q(c[689]) );
  DFF \sreg_reg[690]  ( .D(c[690]), .CLK(clk), .RST(rst), .Q(c[688]) );
  DFF \sreg_reg[689]  ( .D(c[689]), .CLK(clk), .RST(rst), .Q(c[687]) );
  DFF \sreg_reg[688]  ( .D(c[688]), .CLK(clk), .RST(rst), .Q(c[686]) );
  DFF \sreg_reg[687]  ( .D(c[687]), .CLK(clk), .RST(rst), .Q(c[685]) );
  DFF \sreg_reg[686]  ( .D(c[686]), .CLK(clk), .RST(rst), .Q(c[684]) );
  DFF \sreg_reg[685]  ( .D(c[685]), .CLK(clk), .RST(rst), .Q(c[683]) );
  DFF \sreg_reg[684]  ( .D(c[684]), .CLK(clk), .RST(rst), .Q(c[682]) );
  DFF \sreg_reg[683]  ( .D(c[683]), .CLK(clk), .RST(rst), .Q(c[681]) );
  DFF \sreg_reg[682]  ( .D(c[682]), .CLK(clk), .RST(rst), .Q(c[680]) );
  DFF \sreg_reg[681]  ( .D(c[681]), .CLK(clk), .RST(rst), .Q(c[679]) );
  DFF \sreg_reg[680]  ( .D(c[680]), .CLK(clk), .RST(rst), .Q(c[678]) );
  DFF \sreg_reg[679]  ( .D(c[679]), .CLK(clk), .RST(rst), .Q(c[677]) );
  DFF \sreg_reg[678]  ( .D(c[678]), .CLK(clk), .RST(rst), .Q(c[676]) );
  DFF \sreg_reg[677]  ( .D(c[677]), .CLK(clk), .RST(rst), .Q(c[675]) );
  DFF \sreg_reg[676]  ( .D(c[676]), .CLK(clk), .RST(rst), .Q(c[674]) );
  DFF \sreg_reg[675]  ( .D(c[675]), .CLK(clk), .RST(rst), .Q(c[673]) );
  DFF \sreg_reg[674]  ( .D(c[674]), .CLK(clk), .RST(rst), .Q(c[672]) );
  DFF \sreg_reg[673]  ( .D(c[673]), .CLK(clk), .RST(rst), .Q(c[671]) );
  DFF \sreg_reg[672]  ( .D(c[672]), .CLK(clk), .RST(rst), .Q(c[670]) );
  DFF \sreg_reg[671]  ( .D(c[671]), .CLK(clk), .RST(rst), .Q(c[669]) );
  DFF \sreg_reg[670]  ( .D(c[670]), .CLK(clk), .RST(rst), .Q(c[668]) );
  DFF \sreg_reg[669]  ( .D(c[669]), .CLK(clk), .RST(rst), .Q(c[667]) );
  DFF \sreg_reg[668]  ( .D(c[668]), .CLK(clk), .RST(rst), .Q(c[666]) );
  DFF \sreg_reg[667]  ( .D(c[667]), .CLK(clk), .RST(rst), .Q(c[665]) );
  DFF \sreg_reg[666]  ( .D(c[666]), .CLK(clk), .RST(rst), .Q(c[664]) );
  DFF \sreg_reg[665]  ( .D(c[665]), .CLK(clk), .RST(rst), .Q(c[663]) );
  DFF \sreg_reg[664]  ( .D(c[664]), .CLK(clk), .RST(rst), .Q(c[662]) );
  DFF \sreg_reg[663]  ( .D(c[663]), .CLK(clk), .RST(rst), .Q(c[661]) );
  DFF \sreg_reg[662]  ( .D(c[662]), .CLK(clk), .RST(rst), .Q(c[660]) );
  DFF \sreg_reg[661]  ( .D(c[661]), .CLK(clk), .RST(rst), .Q(c[659]) );
  DFF \sreg_reg[660]  ( .D(c[660]), .CLK(clk), .RST(rst), .Q(c[658]) );
  DFF \sreg_reg[659]  ( .D(c[659]), .CLK(clk), .RST(rst), .Q(c[657]) );
  DFF \sreg_reg[658]  ( .D(c[658]), .CLK(clk), .RST(rst), .Q(c[656]) );
  DFF \sreg_reg[657]  ( .D(c[657]), .CLK(clk), .RST(rst), .Q(c[655]) );
  DFF \sreg_reg[656]  ( .D(c[656]), .CLK(clk), .RST(rst), .Q(c[654]) );
  DFF \sreg_reg[655]  ( .D(c[655]), .CLK(clk), .RST(rst), .Q(c[653]) );
  DFF \sreg_reg[654]  ( .D(c[654]), .CLK(clk), .RST(rst), .Q(c[652]) );
  DFF \sreg_reg[653]  ( .D(c[653]), .CLK(clk), .RST(rst), .Q(c[651]) );
  DFF \sreg_reg[652]  ( .D(c[652]), .CLK(clk), .RST(rst), .Q(c[650]) );
  DFF \sreg_reg[651]  ( .D(c[651]), .CLK(clk), .RST(rst), .Q(c[649]) );
  DFF \sreg_reg[650]  ( .D(c[650]), .CLK(clk), .RST(rst), .Q(c[648]) );
  DFF \sreg_reg[649]  ( .D(c[649]), .CLK(clk), .RST(rst), .Q(c[647]) );
  DFF \sreg_reg[648]  ( .D(c[648]), .CLK(clk), .RST(rst), .Q(c[646]) );
  DFF \sreg_reg[647]  ( .D(c[647]), .CLK(clk), .RST(rst), .Q(c[645]) );
  DFF \sreg_reg[646]  ( .D(c[646]), .CLK(clk), .RST(rst), .Q(c[644]) );
  DFF \sreg_reg[645]  ( .D(c[645]), .CLK(clk), .RST(rst), .Q(c[643]) );
  DFF \sreg_reg[644]  ( .D(c[644]), .CLK(clk), .RST(rst), .Q(c[642]) );
  DFF \sreg_reg[643]  ( .D(c[643]), .CLK(clk), .RST(rst), .Q(c[641]) );
  DFF \sreg_reg[642]  ( .D(c[642]), .CLK(clk), .RST(rst), .Q(c[640]) );
  DFF \sreg_reg[641]  ( .D(c[641]), .CLK(clk), .RST(rst), .Q(c[639]) );
  DFF \sreg_reg[640]  ( .D(c[640]), .CLK(clk), .RST(rst), .Q(c[638]) );
  DFF \sreg_reg[639]  ( .D(c[639]), .CLK(clk), .RST(rst), .Q(c[637]) );
  DFF \sreg_reg[638]  ( .D(c[638]), .CLK(clk), .RST(rst), .Q(c[636]) );
  DFF \sreg_reg[637]  ( .D(c[637]), .CLK(clk), .RST(rst), .Q(c[635]) );
  DFF \sreg_reg[636]  ( .D(c[636]), .CLK(clk), .RST(rst), .Q(c[634]) );
  DFF \sreg_reg[635]  ( .D(c[635]), .CLK(clk), .RST(rst), .Q(c[633]) );
  DFF \sreg_reg[634]  ( .D(c[634]), .CLK(clk), .RST(rst), .Q(c[632]) );
  DFF \sreg_reg[633]  ( .D(c[633]), .CLK(clk), .RST(rst), .Q(c[631]) );
  DFF \sreg_reg[632]  ( .D(c[632]), .CLK(clk), .RST(rst), .Q(c[630]) );
  DFF \sreg_reg[631]  ( .D(c[631]), .CLK(clk), .RST(rst), .Q(c[629]) );
  DFF \sreg_reg[630]  ( .D(c[630]), .CLK(clk), .RST(rst), .Q(c[628]) );
  DFF \sreg_reg[629]  ( .D(c[629]), .CLK(clk), .RST(rst), .Q(c[627]) );
  DFF \sreg_reg[628]  ( .D(c[628]), .CLK(clk), .RST(rst), .Q(c[626]) );
  DFF \sreg_reg[627]  ( .D(c[627]), .CLK(clk), .RST(rst), .Q(c[625]) );
  DFF \sreg_reg[626]  ( .D(c[626]), .CLK(clk), .RST(rst), .Q(c[624]) );
  DFF \sreg_reg[625]  ( .D(c[625]), .CLK(clk), .RST(rst), .Q(c[623]) );
  DFF \sreg_reg[624]  ( .D(c[624]), .CLK(clk), .RST(rst), .Q(c[622]) );
  DFF \sreg_reg[623]  ( .D(c[623]), .CLK(clk), .RST(rst), .Q(c[621]) );
  DFF \sreg_reg[622]  ( .D(c[622]), .CLK(clk), .RST(rst), .Q(c[620]) );
  DFF \sreg_reg[621]  ( .D(c[621]), .CLK(clk), .RST(rst), .Q(c[619]) );
  DFF \sreg_reg[620]  ( .D(c[620]), .CLK(clk), .RST(rst), .Q(c[618]) );
  DFF \sreg_reg[619]  ( .D(c[619]), .CLK(clk), .RST(rst), .Q(c[617]) );
  DFF \sreg_reg[618]  ( .D(c[618]), .CLK(clk), .RST(rst), .Q(c[616]) );
  DFF \sreg_reg[617]  ( .D(c[617]), .CLK(clk), .RST(rst), .Q(c[615]) );
  DFF \sreg_reg[616]  ( .D(c[616]), .CLK(clk), .RST(rst), .Q(c[614]) );
  DFF \sreg_reg[615]  ( .D(c[615]), .CLK(clk), .RST(rst), .Q(c[613]) );
  DFF \sreg_reg[614]  ( .D(c[614]), .CLK(clk), .RST(rst), .Q(c[612]) );
  DFF \sreg_reg[613]  ( .D(c[613]), .CLK(clk), .RST(rst), .Q(c[611]) );
  DFF \sreg_reg[612]  ( .D(c[612]), .CLK(clk), .RST(rst), .Q(c[610]) );
  DFF \sreg_reg[611]  ( .D(c[611]), .CLK(clk), .RST(rst), .Q(c[609]) );
  DFF \sreg_reg[610]  ( .D(c[610]), .CLK(clk), .RST(rst), .Q(c[608]) );
  DFF \sreg_reg[609]  ( .D(c[609]), .CLK(clk), .RST(rst), .Q(c[607]) );
  DFF \sreg_reg[608]  ( .D(c[608]), .CLK(clk), .RST(rst), .Q(c[606]) );
  DFF \sreg_reg[607]  ( .D(c[607]), .CLK(clk), .RST(rst), .Q(c[605]) );
  DFF \sreg_reg[606]  ( .D(c[606]), .CLK(clk), .RST(rst), .Q(c[604]) );
  DFF \sreg_reg[605]  ( .D(c[605]), .CLK(clk), .RST(rst), .Q(c[603]) );
  DFF \sreg_reg[604]  ( .D(c[604]), .CLK(clk), .RST(rst), .Q(c[602]) );
  DFF \sreg_reg[603]  ( .D(c[603]), .CLK(clk), .RST(rst), .Q(c[601]) );
  DFF \sreg_reg[602]  ( .D(c[602]), .CLK(clk), .RST(rst), .Q(c[600]) );
  DFF \sreg_reg[601]  ( .D(c[601]), .CLK(clk), .RST(rst), .Q(c[599]) );
  DFF \sreg_reg[600]  ( .D(c[600]), .CLK(clk), .RST(rst), .Q(c[598]) );
  DFF \sreg_reg[599]  ( .D(c[599]), .CLK(clk), .RST(rst), .Q(c[597]) );
  DFF \sreg_reg[598]  ( .D(c[598]), .CLK(clk), .RST(rst), .Q(c[596]) );
  DFF \sreg_reg[597]  ( .D(c[597]), .CLK(clk), .RST(rst), .Q(c[595]) );
  DFF \sreg_reg[596]  ( .D(c[596]), .CLK(clk), .RST(rst), .Q(c[594]) );
  DFF \sreg_reg[595]  ( .D(c[595]), .CLK(clk), .RST(rst), .Q(c[593]) );
  DFF \sreg_reg[594]  ( .D(c[594]), .CLK(clk), .RST(rst), .Q(c[592]) );
  DFF \sreg_reg[593]  ( .D(c[593]), .CLK(clk), .RST(rst), .Q(c[591]) );
  DFF \sreg_reg[592]  ( .D(c[592]), .CLK(clk), .RST(rst), .Q(c[590]) );
  DFF \sreg_reg[591]  ( .D(c[591]), .CLK(clk), .RST(rst), .Q(c[589]) );
  DFF \sreg_reg[590]  ( .D(c[590]), .CLK(clk), .RST(rst), .Q(c[588]) );
  DFF \sreg_reg[589]  ( .D(c[589]), .CLK(clk), .RST(rst), .Q(c[587]) );
  DFF \sreg_reg[588]  ( .D(c[588]), .CLK(clk), .RST(rst), .Q(c[586]) );
  DFF \sreg_reg[587]  ( .D(c[587]), .CLK(clk), .RST(rst), .Q(c[585]) );
  DFF \sreg_reg[586]  ( .D(c[586]), .CLK(clk), .RST(rst), .Q(c[584]) );
  DFF \sreg_reg[585]  ( .D(c[585]), .CLK(clk), .RST(rst), .Q(c[583]) );
  DFF \sreg_reg[584]  ( .D(c[584]), .CLK(clk), .RST(rst), .Q(c[582]) );
  DFF \sreg_reg[583]  ( .D(c[583]), .CLK(clk), .RST(rst), .Q(c[581]) );
  DFF \sreg_reg[582]  ( .D(c[582]), .CLK(clk), .RST(rst), .Q(c[580]) );
  DFF \sreg_reg[581]  ( .D(c[581]), .CLK(clk), .RST(rst), .Q(c[579]) );
  DFF \sreg_reg[580]  ( .D(c[580]), .CLK(clk), .RST(rst), .Q(c[578]) );
  DFF \sreg_reg[579]  ( .D(c[579]), .CLK(clk), .RST(rst), .Q(c[577]) );
  DFF \sreg_reg[578]  ( .D(c[578]), .CLK(clk), .RST(rst), .Q(c[576]) );
  DFF \sreg_reg[577]  ( .D(c[577]), .CLK(clk), .RST(rst), .Q(c[575]) );
  DFF \sreg_reg[576]  ( .D(c[576]), .CLK(clk), .RST(rst), .Q(c[574]) );
  DFF \sreg_reg[575]  ( .D(c[575]), .CLK(clk), .RST(rst), .Q(c[573]) );
  DFF \sreg_reg[574]  ( .D(c[574]), .CLK(clk), .RST(rst), .Q(c[572]) );
  DFF \sreg_reg[573]  ( .D(c[573]), .CLK(clk), .RST(rst), .Q(c[571]) );
  DFF \sreg_reg[572]  ( .D(c[572]), .CLK(clk), .RST(rst), .Q(c[570]) );
  DFF \sreg_reg[571]  ( .D(c[571]), .CLK(clk), .RST(rst), .Q(c[569]) );
  DFF \sreg_reg[570]  ( .D(c[570]), .CLK(clk), .RST(rst), .Q(c[568]) );
  DFF \sreg_reg[569]  ( .D(c[569]), .CLK(clk), .RST(rst), .Q(c[567]) );
  DFF \sreg_reg[568]  ( .D(c[568]), .CLK(clk), .RST(rst), .Q(c[566]) );
  DFF \sreg_reg[567]  ( .D(c[567]), .CLK(clk), .RST(rst), .Q(c[565]) );
  DFF \sreg_reg[566]  ( .D(c[566]), .CLK(clk), .RST(rst), .Q(c[564]) );
  DFF \sreg_reg[565]  ( .D(c[565]), .CLK(clk), .RST(rst), .Q(c[563]) );
  DFF \sreg_reg[564]  ( .D(c[564]), .CLK(clk), .RST(rst), .Q(c[562]) );
  DFF \sreg_reg[563]  ( .D(c[563]), .CLK(clk), .RST(rst), .Q(c[561]) );
  DFF \sreg_reg[562]  ( .D(c[562]), .CLK(clk), .RST(rst), .Q(c[560]) );
  DFF \sreg_reg[561]  ( .D(c[561]), .CLK(clk), .RST(rst), .Q(c[559]) );
  DFF \sreg_reg[560]  ( .D(c[560]), .CLK(clk), .RST(rst), .Q(c[558]) );
  DFF \sreg_reg[559]  ( .D(c[559]), .CLK(clk), .RST(rst), .Q(c[557]) );
  DFF \sreg_reg[558]  ( .D(c[558]), .CLK(clk), .RST(rst), .Q(c[556]) );
  DFF \sreg_reg[557]  ( .D(c[557]), .CLK(clk), .RST(rst), .Q(c[555]) );
  DFF \sreg_reg[556]  ( .D(c[556]), .CLK(clk), .RST(rst), .Q(c[554]) );
  DFF \sreg_reg[555]  ( .D(c[555]), .CLK(clk), .RST(rst), .Q(c[553]) );
  DFF \sreg_reg[554]  ( .D(c[554]), .CLK(clk), .RST(rst), .Q(c[552]) );
  DFF \sreg_reg[553]  ( .D(c[553]), .CLK(clk), .RST(rst), .Q(c[551]) );
  DFF \sreg_reg[552]  ( .D(c[552]), .CLK(clk), .RST(rst), .Q(c[550]) );
  DFF \sreg_reg[551]  ( .D(c[551]), .CLK(clk), .RST(rst), .Q(c[549]) );
  DFF \sreg_reg[550]  ( .D(c[550]), .CLK(clk), .RST(rst), .Q(c[548]) );
  DFF \sreg_reg[549]  ( .D(c[549]), .CLK(clk), .RST(rst), .Q(c[547]) );
  DFF \sreg_reg[548]  ( .D(c[548]), .CLK(clk), .RST(rst), .Q(c[546]) );
  DFF \sreg_reg[547]  ( .D(c[547]), .CLK(clk), .RST(rst), .Q(c[545]) );
  DFF \sreg_reg[546]  ( .D(c[546]), .CLK(clk), .RST(rst), .Q(c[544]) );
  DFF \sreg_reg[545]  ( .D(c[545]), .CLK(clk), .RST(rst), .Q(c[543]) );
  DFF \sreg_reg[544]  ( .D(c[544]), .CLK(clk), .RST(rst), .Q(c[542]) );
  DFF \sreg_reg[543]  ( .D(c[543]), .CLK(clk), .RST(rst), .Q(c[541]) );
  DFF \sreg_reg[542]  ( .D(c[542]), .CLK(clk), .RST(rst), .Q(c[540]) );
  DFF \sreg_reg[541]  ( .D(c[541]), .CLK(clk), .RST(rst), .Q(c[539]) );
  DFF \sreg_reg[540]  ( .D(c[540]), .CLK(clk), .RST(rst), .Q(c[538]) );
  DFF \sreg_reg[539]  ( .D(c[539]), .CLK(clk), .RST(rst), .Q(c[537]) );
  DFF \sreg_reg[538]  ( .D(c[538]), .CLK(clk), .RST(rst), .Q(c[536]) );
  DFF \sreg_reg[537]  ( .D(c[537]), .CLK(clk), .RST(rst), .Q(c[535]) );
  DFF \sreg_reg[536]  ( .D(c[536]), .CLK(clk), .RST(rst), .Q(c[534]) );
  DFF \sreg_reg[535]  ( .D(c[535]), .CLK(clk), .RST(rst), .Q(c[533]) );
  DFF \sreg_reg[534]  ( .D(c[534]), .CLK(clk), .RST(rst), .Q(c[532]) );
  DFF \sreg_reg[533]  ( .D(c[533]), .CLK(clk), .RST(rst), .Q(c[531]) );
  DFF \sreg_reg[532]  ( .D(c[532]), .CLK(clk), .RST(rst), .Q(c[530]) );
  DFF \sreg_reg[531]  ( .D(c[531]), .CLK(clk), .RST(rst), .Q(c[529]) );
  DFF \sreg_reg[530]  ( .D(c[530]), .CLK(clk), .RST(rst), .Q(c[528]) );
  DFF \sreg_reg[529]  ( .D(c[529]), .CLK(clk), .RST(rst), .Q(c[527]) );
  DFF \sreg_reg[528]  ( .D(c[528]), .CLK(clk), .RST(rst), .Q(c[526]) );
  DFF \sreg_reg[527]  ( .D(c[527]), .CLK(clk), .RST(rst), .Q(c[525]) );
  DFF \sreg_reg[526]  ( .D(c[526]), .CLK(clk), .RST(rst), .Q(c[524]) );
  DFF \sreg_reg[525]  ( .D(c[525]), .CLK(clk), .RST(rst), .Q(c[523]) );
  DFF \sreg_reg[524]  ( .D(c[524]), .CLK(clk), .RST(rst), .Q(c[522]) );
  DFF \sreg_reg[523]  ( .D(c[523]), .CLK(clk), .RST(rst), .Q(c[521]) );
  DFF \sreg_reg[522]  ( .D(c[522]), .CLK(clk), .RST(rst), .Q(c[520]) );
  DFF \sreg_reg[521]  ( .D(c[521]), .CLK(clk), .RST(rst), .Q(c[519]) );
  DFF \sreg_reg[520]  ( .D(c[520]), .CLK(clk), .RST(rst), .Q(c[518]) );
  DFF \sreg_reg[519]  ( .D(c[519]), .CLK(clk), .RST(rst), .Q(c[517]) );
  DFF \sreg_reg[518]  ( .D(c[518]), .CLK(clk), .RST(rst), .Q(c[516]) );
  DFF \sreg_reg[517]  ( .D(c[517]), .CLK(clk), .RST(rst), .Q(c[515]) );
  DFF \sreg_reg[516]  ( .D(c[516]), .CLK(clk), .RST(rst), .Q(c[514]) );
  DFF \sreg_reg[515]  ( .D(c[515]), .CLK(clk), .RST(rst), .Q(c[513]) );
  DFF \sreg_reg[514]  ( .D(c[514]), .CLK(clk), .RST(rst), .Q(c[512]) );
  DFF \sreg_reg[513]  ( .D(c[513]), .CLK(clk), .RST(rst), .Q(c[511]) );
  DFF \sreg_reg[512]  ( .D(c[512]), .CLK(clk), .RST(rst), .Q(c[510]) );
  DFF \sreg_reg[511]  ( .D(c[511]), .CLK(clk), .RST(rst), .Q(c[509]) );
  DFF \sreg_reg[510]  ( .D(c[510]), .CLK(clk), .RST(rst), .Q(c[508]) );
  DFF \sreg_reg[509]  ( .D(c[509]), .CLK(clk), .RST(rst), .Q(c[507]) );
  DFF \sreg_reg[508]  ( .D(c[508]), .CLK(clk), .RST(rst), .Q(c[506]) );
  DFF \sreg_reg[507]  ( .D(c[507]), .CLK(clk), .RST(rst), .Q(c[505]) );
  DFF \sreg_reg[506]  ( .D(c[506]), .CLK(clk), .RST(rst), .Q(c[504]) );
  DFF \sreg_reg[505]  ( .D(c[505]), .CLK(clk), .RST(rst), .Q(c[503]) );
  DFF \sreg_reg[504]  ( .D(c[504]), .CLK(clk), .RST(rst), .Q(c[502]) );
  DFF \sreg_reg[503]  ( .D(c[503]), .CLK(clk), .RST(rst), .Q(c[501]) );
  DFF \sreg_reg[502]  ( .D(c[502]), .CLK(clk), .RST(rst), .Q(c[500]) );
  DFF \sreg_reg[501]  ( .D(c[501]), .CLK(clk), .RST(rst), .Q(c[499]) );
  DFF \sreg_reg[500]  ( .D(c[500]), .CLK(clk), .RST(rst), .Q(c[498]) );
  DFF \sreg_reg[499]  ( .D(c[499]), .CLK(clk), .RST(rst), .Q(c[497]) );
  DFF \sreg_reg[498]  ( .D(c[498]), .CLK(clk), .RST(rst), .Q(c[496]) );
  DFF \sreg_reg[497]  ( .D(c[497]), .CLK(clk), .RST(rst), .Q(c[495]) );
  DFF \sreg_reg[496]  ( .D(c[496]), .CLK(clk), .RST(rst), .Q(c[494]) );
  DFF \sreg_reg[495]  ( .D(c[495]), .CLK(clk), .RST(rst), .Q(c[493]) );
  DFF \sreg_reg[494]  ( .D(c[494]), .CLK(clk), .RST(rst), .Q(c[492]) );
  DFF \sreg_reg[493]  ( .D(c[493]), .CLK(clk), .RST(rst), .Q(c[491]) );
  DFF \sreg_reg[492]  ( .D(c[492]), .CLK(clk), .RST(rst), .Q(c[490]) );
  DFF \sreg_reg[491]  ( .D(c[491]), .CLK(clk), .RST(rst), .Q(c[489]) );
  DFF \sreg_reg[490]  ( .D(c[490]), .CLK(clk), .RST(rst), .Q(c[488]) );
  DFF \sreg_reg[489]  ( .D(c[489]), .CLK(clk), .RST(rst), .Q(c[487]) );
  DFF \sreg_reg[488]  ( .D(c[488]), .CLK(clk), .RST(rst), .Q(c[486]) );
  DFF \sreg_reg[487]  ( .D(c[487]), .CLK(clk), .RST(rst), .Q(c[485]) );
  DFF \sreg_reg[486]  ( .D(c[486]), .CLK(clk), .RST(rst), .Q(c[484]) );
  DFF \sreg_reg[485]  ( .D(c[485]), .CLK(clk), .RST(rst), .Q(c[483]) );
  DFF \sreg_reg[484]  ( .D(c[484]), .CLK(clk), .RST(rst), .Q(c[482]) );
  DFF \sreg_reg[483]  ( .D(c[483]), .CLK(clk), .RST(rst), .Q(c[481]) );
  DFF \sreg_reg[482]  ( .D(c[482]), .CLK(clk), .RST(rst), .Q(c[480]) );
  DFF \sreg_reg[481]  ( .D(c[481]), .CLK(clk), .RST(rst), .Q(c[479]) );
  DFF \sreg_reg[480]  ( .D(c[480]), .CLK(clk), .RST(rst), .Q(c[478]) );
  DFF \sreg_reg[479]  ( .D(c[479]), .CLK(clk), .RST(rst), .Q(c[477]) );
  DFF \sreg_reg[478]  ( .D(c[478]), .CLK(clk), .RST(rst), .Q(c[476]) );
  DFF \sreg_reg[477]  ( .D(c[477]), .CLK(clk), .RST(rst), .Q(c[475]) );
  DFF \sreg_reg[476]  ( .D(c[476]), .CLK(clk), .RST(rst), .Q(c[474]) );
  DFF \sreg_reg[475]  ( .D(c[475]), .CLK(clk), .RST(rst), .Q(c[473]) );
  DFF \sreg_reg[474]  ( .D(c[474]), .CLK(clk), .RST(rst), .Q(c[472]) );
  DFF \sreg_reg[473]  ( .D(c[473]), .CLK(clk), .RST(rst), .Q(c[471]) );
  DFF \sreg_reg[472]  ( .D(c[472]), .CLK(clk), .RST(rst), .Q(c[470]) );
  DFF \sreg_reg[471]  ( .D(c[471]), .CLK(clk), .RST(rst), .Q(c[469]) );
  DFF \sreg_reg[470]  ( .D(c[470]), .CLK(clk), .RST(rst), .Q(c[468]) );
  DFF \sreg_reg[469]  ( .D(c[469]), .CLK(clk), .RST(rst), .Q(c[467]) );
  DFF \sreg_reg[468]  ( .D(c[468]), .CLK(clk), .RST(rst), .Q(c[466]) );
  DFF \sreg_reg[467]  ( .D(c[467]), .CLK(clk), .RST(rst), .Q(c[465]) );
  DFF \sreg_reg[466]  ( .D(c[466]), .CLK(clk), .RST(rst), .Q(c[464]) );
  DFF \sreg_reg[465]  ( .D(c[465]), .CLK(clk), .RST(rst), .Q(c[463]) );
  DFF \sreg_reg[464]  ( .D(c[464]), .CLK(clk), .RST(rst), .Q(c[462]) );
  DFF \sreg_reg[463]  ( .D(c[463]), .CLK(clk), .RST(rst), .Q(c[461]) );
  DFF \sreg_reg[462]  ( .D(c[462]), .CLK(clk), .RST(rst), .Q(c[460]) );
  DFF \sreg_reg[461]  ( .D(c[461]), .CLK(clk), .RST(rst), .Q(c[459]) );
  DFF \sreg_reg[460]  ( .D(c[460]), .CLK(clk), .RST(rst), .Q(c[458]) );
  DFF \sreg_reg[459]  ( .D(c[459]), .CLK(clk), .RST(rst), .Q(c[457]) );
  DFF \sreg_reg[458]  ( .D(c[458]), .CLK(clk), .RST(rst), .Q(c[456]) );
  DFF \sreg_reg[457]  ( .D(c[457]), .CLK(clk), .RST(rst), .Q(c[455]) );
  DFF \sreg_reg[456]  ( .D(c[456]), .CLK(clk), .RST(rst), .Q(c[454]) );
  DFF \sreg_reg[455]  ( .D(c[455]), .CLK(clk), .RST(rst), .Q(c[453]) );
  DFF \sreg_reg[454]  ( .D(c[454]), .CLK(clk), .RST(rst), .Q(c[452]) );
  DFF \sreg_reg[453]  ( .D(c[453]), .CLK(clk), .RST(rst), .Q(c[451]) );
  DFF \sreg_reg[452]  ( .D(c[452]), .CLK(clk), .RST(rst), .Q(c[450]) );
  DFF \sreg_reg[451]  ( .D(c[451]), .CLK(clk), .RST(rst), .Q(c[449]) );
  DFF \sreg_reg[450]  ( .D(c[450]), .CLK(clk), .RST(rst), .Q(c[448]) );
  DFF \sreg_reg[449]  ( .D(c[449]), .CLK(clk), .RST(rst), .Q(c[447]) );
  DFF \sreg_reg[448]  ( .D(c[448]), .CLK(clk), .RST(rst), .Q(c[446]) );
  DFF \sreg_reg[447]  ( .D(c[447]), .CLK(clk), .RST(rst), .Q(c[445]) );
  DFF \sreg_reg[446]  ( .D(c[446]), .CLK(clk), .RST(rst), .Q(c[444]) );
  DFF \sreg_reg[445]  ( .D(c[445]), .CLK(clk), .RST(rst), .Q(c[443]) );
  DFF \sreg_reg[444]  ( .D(c[444]), .CLK(clk), .RST(rst), .Q(c[442]) );
  DFF \sreg_reg[443]  ( .D(c[443]), .CLK(clk), .RST(rst), .Q(c[441]) );
  DFF \sreg_reg[442]  ( .D(c[442]), .CLK(clk), .RST(rst), .Q(c[440]) );
  DFF \sreg_reg[441]  ( .D(c[441]), .CLK(clk), .RST(rst), .Q(c[439]) );
  DFF \sreg_reg[440]  ( .D(c[440]), .CLK(clk), .RST(rst), .Q(c[438]) );
  DFF \sreg_reg[439]  ( .D(c[439]), .CLK(clk), .RST(rst), .Q(c[437]) );
  DFF \sreg_reg[438]  ( .D(c[438]), .CLK(clk), .RST(rst), .Q(c[436]) );
  DFF \sreg_reg[437]  ( .D(c[437]), .CLK(clk), .RST(rst), .Q(c[435]) );
  DFF \sreg_reg[436]  ( .D(c[436]), .CLK(clk), .RST(rst), .Q(c[434]) );
  DFF \sreg_reg[435]  ( .D(c[435]), .CLK(clk), .RST(rst), .Q(c[433]) );
  DFF \sreg_reg[434]  ( .D(c[434]), .CLK(clk), .RST(rst), .Q(c[432]) );
  DFF \sreg_reg[433]  ( .D(c[433]), .CLK(clk), .RST(rst), .Q(c[431]) );
  DFF \sreg_reg[432]  ( .D(c[432]), .CLK(clk), .RST(rst), .Q(c[430]) );
  DFF \sreg_reg[431]  ( .D(c[431]), .CLK(clk), .RST(rst), .Q(c[429]) );
  DFF \sreg_reg[430]  ( .D(c[430]), .CLK(clk), .RST(rst), .Q(c[428]) );
  DFF \sreg_reg[429]  ( .D(c[429]), .CLK(clk), .RST(rst), .Q(c[427]) );
  DFF \sreg_reg[428]  ( .D(c[428]), .CLK(clk), .RST(rst), .Q(c[426]) );
  DFF \sreg_reg[427]  ( .D(c[427]), .CLK(clk), .RST(rst), .Q(c[425]) );
  DFF \sreg_reg[426]  ( .D(c[426]), .CLK(clk), .RST(rst), .Q(c[424]) );
  DFF \sreg_reg[425]  ( .D(c[425]), .CLK(clk), .RST(rst), .Q(c[423]) );
  DFF \sreg_reg[424]  ( .D(c[424]), .CLK(clk), .RST(rst), .Q(c[422]) );
  DFF \sreg_reg[423]  ( .D(c[423]), .CLK(clk), .RST(rst), .Q(c[421]) );
  DFF \sreg_reg[422]  ( .D(c[422]), .CLK(clk), .RST(rst), .Q(c[420]) );
  DFF \sreg_reg[421]  ( .D(c[421]), .CLK(clk), .RST(rst), .Q(c[419]) );
  DFF \sreg_reg[420]  ( .D(c[420]), .CLK(clk), .RST(rst), .Q(c[418]) );
  DFF \sreg_reg[419]  ( .D(c[419]), .CLK(clk), .RST(rst), .Q(c[417]) );
  DFF \sreg_reg[418]  ( .D(c[418]), .CLK(clk), .RST(rst), .Q(c[416]) );
  DFF \sreg_reg[417]  ( .D(c[417]), .CLK(clk), .RST(rst), .Q(c[415]) );
  DFF \sreg_reg[416]  ( .D(c[416]), .CLK(clk), .RST(rst), .Q(c[414]) );
  DFF \sreg_reg[415]  ( .D(c[415]), .CLK(clk), .RST(rst), .Q(c[413]) );
  DFF \sreg_reg[414]  ( .D(c[414]), .CLK(clk), .RST(rst), .Q(c[412]) );
  DFF \sreg_reg[413]  ( .D(c[413]), .CLK(clk), .RST(rst), .Q(c[411]) );
  DFF \sreg_reg[412]  ( .D(c[412]), .CLK(clk), .RST(rst), .Q(c[410]) );
  DFF \sreg_reg[411]  ( .D(c[411]), .CLK(clk), .RST(rst), .Q(c[409]) );
  DFF \sreg_reg[410]  ( .D(c[410]), .CLK(clk), .RST(rst), .Q(c[408]) );
  DFF \sreg_reg[409]  ( .D(c[409]), .CLK(clk), .RST(rst), .Q(c[407]) );
  DFF \sreg_reg[408]  ( .D(c[408]), .CLK(clk), .RST(rst), .Q(c[406]) );
  DFF \sreg_reg[407]  ( .D(c[407]), .CLK(clk), .RST(rst), .Q(c[405]) );
  DFF \sreg_reg[406]  ( .D(c[406]), .CLK(clk), .RST(rst), .Q(c[404]) );
  DFF \sreg_reg[405]  ( .D(c[405]), .CLK(clk), .RST(rst), .Q(c[403]) );
  DFF \sreg_reg[404]  ( .D(c[404]), .CLK(clk), .RST(rst), .Q(c[402]) );
  DFF \sreg_reg[403]  ( .D(c[403]), .CLK(clk), .RST(rst), .Q(c[401]) );
  DFF \sreg_reg[402]  ( .D(c[402]), .CLK(clk), .RST(rst), .Q(c[400]) );
  DFF \sreg_reg[401]  ( .D(c[401]), .CLK(clk), .RST(rst), .Q(c[399]) );
  DFF \sreg_reg[400]  ( .D(c[400]), .CLK(clk), .RST(rst), .Q(c[398]) );
  DFF \sreg_reg[399]  ( .D(c[399]), .CLK(clk), .RST(rst), .Q(c[397]) );
  DFF \sreg_reg[398]  ( .D(c[398]), .CLK(clk), .RST(rst), .Q(c[396]) );
  DFF \sreg_reg[397]  ( .D(c[397]), .CLK(clk), .RST(rst), .Q(c[395]) );
  DFF \sreg_reg[396]  ( .D(c[396]), .CLK(clk), .RST(rst), .Q(c[394]) );
  DFF \sreg_reg[395]  ( .D(c[395]), .CLK(clk), .RST(rst), .Q(c[393]) );
  DFF \sreg_reg[394]  ( .D(c[394]), .CLK(clk), .RST(rst), .Q(c[392]) );
  DFF \sreg_reg[393]  ( .D(c[393]), .CLK(clk), .RST(rst), .Q(c[391]) );
  DFF \sreg_reg[392]  ( .D(c[392]), .CLK(clk), .RST(rst), .Q(c[390]) );
  DFF \sreg_reg[391]  ( .D(c[391]), .CLK(clk), .RST(rst), .Q(c[389]) );
  DFF \sreg_reg[390]  ( .D(c[390]), .CLK(clk), .RST(rst), .Q(c[388]) );
  DFF \sreg_reg[389]  ( .D(c[389]), .CLK(clk), .RST(rst), .Q(c[387]) );
  DFF \sreg_reg[388]  ( .D(c[388]), .CLK(clk), .RST(rst), .Q(c[386]) );
  DFF \sreg_reg[387]  ( .D(c[387]), .CLK(clk), .RST(rst), .Q(c[385]) );
  DFF \sreg_reg[386]  ( .D(c[386]), .CLK(clk), .RST(rst), .Q(c[384]) );
  DFF \sreg_reg[385]  ( .D(c[385]), .CLK(clk), .RST(rst), .Q(c[383]) );
  DFF \sreg_reg[384]  ( .D(c[384]), .CLK(clk), .RST(rst), .Q(c[382]) );
  DFF \sreg_reg[383]  ( .D(c[383]), .CLK(clk), .RST(rst), .Q(c[381]) );
  DFF \sreg_reg[382]  ( .D(c[382]), .CLK(clk), .RST(rst), .Q(c[380]) );
  DFF \sreg_reg[381]  ( .D(c[381]), .CLK(clk), .RST(rst), .Q(c[379]) );
  DFF \sreg_reg[380]  ( .D(c[380]), .CLK(clk), .RST(rst), .Q(c[378]) );
  DFF \sreg_reg[379]  ( .D(c[379]), .CLK(clk), .RST(rst), .Q(c[377]) );
  DFF \sreg_reg[378]  ( .D(c[378]), .CLK(clk), .RST(rst), .Q(c[376]) );
  DFF \sreg_reg[377]  ( .D(c[377]), .CLK(clk), .RST(rst), .Q(c[375]) );
  DFF \sreg_reg[376]  ( .D(c[376]), .CLK(clk), .RST(rst), .Q(c[374]) );
  DFF \sreg_reg[375]  ( .D(c[375]), .CLK(clk), .RST(rst), .Q(c[373]) );
  DFF \sreg_reg[374]  ( .D(c[374]), .CLK(clk), .RST(rst), .Q(c[372]) );
  DFF \sreg_reg[373]  ( .D(c[373]), .CLK(clk), .RST(rst), .Q(c[371]) );
  DFF \sreg_reg[372]  ( .D(c[372]), .CLK(clk), .RST(rst), .Q(c[370]) );
  DFF \sreg_reg[371]  ( .D(c[371]), .CLK(clk), .RST(rst), .Q(c[369]) );
  DFF \sreg_reg[370]  ( .D(c[370]), .CLK(clk), .RST(rst), .Q(c[368]) );
  DFF \sreg_reg[369]  ( .D(c[369]), .CLK(clk), .RST(rst), .Q(c[367]) );
  DFF \sreg_reg[368]  ( .D(c[368]), .CLK(clk), .RST(rst), .Q(c[366]) );
  DFF \sreg_reg[367]  ( .D(c[367]), .CLK(clk), .RST(rst), .Q(c[365]) );
  DFF \sreg_reg[366]  ( .D(c[366]), .CLK(clk), .RST(rst), .Q(c[364]) );
  DFF \sreg_reg[365]  ( .D(c[365]), .CLK(clk), .RST(rst), .Q(c[363]) );
  DFF \sreg_reg[364]  ( .D(c[364]), .CLK(clk), .RST(rst), .Q(c[362]) );
  DFF \sreg_reg[363]  ( .D(c[363]), .CLK(clk), .RST(rst), .Q(c[361]) );
  DFF \sreg_reg[362]  ( .D(c[362]), .CLK(clk), .RST(rst), .Q(c[360]) );
  DFF \sreg_reg[361]  ( .D(c[361]), .CLK(clk), .RST(rst), .Q(c[359]) );
  DFF \sreg_reg[360]  ( .D(c[360]), .CLK(clk), .RST(rst), .Q(c[358]) );
  DFF \sreg_reg[359]  ( .D(c[359]), .CLK(clk), .RST(rst), .Q(c[357]) );
  DFF \sreg_reg[358]  ( .D(c[358]), .CLK(clk), .RST(rst), .Q(c[356]) );
  DFF \sreg_reg[357]  ( .D(c[357]), .CLK(clk), .RST(rst), .Q(c[355]) );
  DFF \sreg_reg[356]  ( .D(c[356]), .CLK(clk), .RST(rst), .Q(c[354]) );
  DFF \sreg_reg[355]  ( .D(c[355]), .CLK(clk), .RST(rst), .Q(c[353]) );
  DFF \sreg_reg[354]  ( .D(c[354]), .CLK(clk), .RST(rst), .Q(c[352]) );
  DFF \sreg_reg[353]  ( .D(c[353]), .CLK(clk), .RST(rst), .Q(c[351]) );
  DFF \sreg_reg[352]  ( .D(c[352]), .CLK(clk), .RST(rst), .Q(c[350]) );
  DFF \sreg_reg[351]  ( .D(c[351]), .CLK(clk), .RST(rst), .Q(c[349]) );
  DFF \sreg_reg[350]  ( .D(c[350]), .CLK(clk), .RST(rst), .Q(c[348]) );
  DFF \sreg_reg[349]  ( .D(c[349]), .CLK(clk), .RST(rst), .Q(c[347]) );
  DFF \sreg_reg[348]  ( .D(c[348]), .CLK(clk), .RST(rst), .Q(c[346]) );
  DFF \sreg_reg[347]  ( .D(c[347]), .CLK(clk), .RST(rst), .Q(c[345]) );
  DFF \sreg_reg[346]  ( .D(c[346]), .CLK(clk), .RST(rst), .Q(c[344]) );
  DFF \sreg_reg[345]  ( .D(c[345]), .CLK(clk), .RST(rst), .Q(c[343]) );
  DFF \sreg_reg[344]  ( .D(c[344]), .CLK(clk), .RST(rst), .Q(c[342]) );
  DFF \sreg_reg[343]  ( .D(c[343]), .CLK(clk), .RST(rst), .Q(c[341]) );
  DFF \sreg_reg[342]  ( .D(c[342]), .CLK(clk), .RST(rst), .Q(c[340]) );
  DFF \sreg_reg[341]  ( .D(c[341]), .CLK(clk), .RST(rst), .Q(c[339]) );
  DFF \sreg_reg[340]  ( .D(c[340]), .CLK(clk), .RST(rst), .Q(c[338]) );
  DFF \sreg_reg[339]  ( .D(c[339]), .CLK(clk), .RST(rst), .Q(c[337]) );
  DFF \sreg_reg[338]  ( .D(c[338]), .CLK(clk), .RST(rst), .Q(c[336]) );
  DFF \sreg_reg[337]  ( .D(c[337]), .CLK(clk), .RST(rst), .Q(c[335]) );
  DFF \sreg_reg[336]  ( .D(c[336]), .CLK(clk), .RST(rst), .Q(c[334]) );
  DFF \sreg_reg[335]  ( .D(c[335]), .CLK(clk), .RST(rst), .Q(c[333]) );
  DFF \sreg_reg[334]  ( .D(c[334]), .CLK(clk), .RST(rst), .Q(c[332]) );
  DFF \sreg_reg[333]  ( .D(c[333]), .CLK(clk), .RST(rst), .Q(c[331]) );
  DFF \sreg_reg[332]  ( .D(c[332]), .CLK(clk), .RST(rst), .Q(c[330]) );
  DFF \sreg_reg[331]  ( .D(c[331]), .CLK(clk), .RST(rst), .Q(c[329]) );
  DFF \sreg_reg[330]  ( .D(c[330]), .CLK(clk), .RST(rst), .Q(c[328]) );
  DFF \sreg_reg[329]  ( .D(c[329]), .CLK(clk), .RST(rst), .Q(c[327]) );
  DFF \sreg_reg[328]  ( .D(c[328]), .CLK(clk), .RST(rst), .Q(c[326]) );
  DFF \sreg_reg[327]  ( .D(c[327]), .CLK(clk), .RST(rst), .Q(c[325]) );
  DFF \sreg_reg[326]  ( .D(c[326]), .CLK(clk), .RST(rst), .Q(c[324]) );
  DFF \sreg_reg[325]  ( .D(c[325]), .CLK(clk), .RST(rst), .Q(c[323]) );
  DFF \sreg_reg[324]  ( .D(c[324]), .CLK(clk), .RST(rst), .Q(c[322]) );
  DFF \sreg_reg[323]  ( .D(c[323]), .CLK(clk), .RST(rst), .Q(c[321]) );
  DFF \sreg_reg[322]  ( .D(c[322]), .CLK(clk), .RST(rst), .Q(c[320]) );
  DFF \sreg_reg[321]  ( .D(c[321]), .CLK(clk), .RST(rst), .Q(c[319]) );
  DFF \sreg_reg[320]  ( .D(c[320]), .CLK(clk), .RST(rst), .Q(c[318]) );
  DFF \sreg_reg[319]  ( .D(c[319]), .CLK(clk), .RST(rst), .Q(c[317]) );
  DFF \sreg_reg[318]  ( .D(c[318]), .CLK(clk), .RST(rst), .Q(c[316]) );
  DFF \sreg_reg[317]  ( .D(c[317]), .CLK(clk), .RST(rst), .Q(c[315]) );
  DFF \sreg_reg[316]  ( .D(c[316]), .CLK(clk), .RST(rst), .Q(c[314]) );
  DFF \sreg_reg[315]  ( .D(c[315]), .CLK(clk), .RST(rst), .Q(c[313]) );
  DFF \sreg_reg[314]  ( .D(c[314]), .CLK(clk), .RST(rst), .Q(c[312]) );
  DFF \sreg_reg[313]  ( .D(c[313]), .CLK(clk), .RST(rst), .Q(c[311]) );
  DFF \sreg_reg[312]  ( .D(c[312]), .CLK(clk), .RST(rst), .Q(c[310]) );
  DFF \sreg_reg[311]  ( .D(c[311]), .CLK(clk), .RST(rst), .Q(c[309]) );
  DFF \sreg_reg[310]  ( .D(c[310]), .CLK(clk), .RST(rst), .Q(c[308]) );
  DFF \sreg_reg[309]  ( .D(c[309]), .CLK(clk), .RST(rst), .Q(c[307]) );
  DFF \sreg_reg[308]  ( .D(c[308]), .CLK(clk), .RST(rst), .Q(c[306]) );
  DFF \sreg_reg[307]  ( .D(c[307]), .CLK(clk), .RST(rst), .Q(c[305]) );
  DFF \sreg_reg[306]  ( .D(c[306]), .CLK(clk), .RST(rst), .Q(c[304]) );
  DFF \sreg_reg[305]  ( .D(c[305]), .CLK(clk), .RST(rst), .Q(c[303]) );
  DFF \sreg_reg[304]  ( .D(c[304]), .CLK(clk), .RST(rst), .Q(c[302]) );
  DFF \sreg_reg[303]  ( .D(c[303]), .CLK(clk), .RST(rst), .Q(c[301]) );
  DFF \sreg_reg[302]  ( .D(c[302]), .CLK(clk), .RST(rst), .Q(c[300]) );
  DFF \sreg_reg[301]  ( .D(c[301]), .CLK(clk), .RST(rst), .Q(c[299]) );
  DFF \sreg_reg[300]  ( .D(c[300]), .CLK(clk), .RST(rst), .Q(c[298]) );
  DFF \sreg_reg[299]  ( .D(c[299]), .CLK(clk), .RST(rst), .Q(c[297]) );
  DFF \sreg_reg[298]  ( .D(c[298]), .CLK(clk), .RST(rst), .Q(c[296]) );
  DFF \sreg_reg[297]  ( .D(c[297]), .CLK(clk), .RST(rst), .Q(c[295]) );
  DFF \sreg_reg[296]  ( .D(c[296]), .CLK(clk), .RST(rst), .Q(c[294]) );
  DFF \sreg_reg[295]  ( .D(c[295]), .CLK(clk), .RST(rst), .Q(c[293]) );
  DFF \sreg_reg[294]  ( .D(c[294]), .CLK(clk), .RST(rst), .Q(c[292]) );
  DFF \sreg_reg[293]  ( .D(c[293]), .CLK(clk), .RST(rst), .Q(c[291]) );
  DFF \sreg_reg[292]  ( .D(c[292]), .CLK(clk), .RST(rst), .Q(c[290]) );
  DFF \sreg_reg[291]  ( .D(c[291]), .CLK(clk), .RST(rst), .Q(c[289]) );
  DFF \sreg_reg[290]  ( .D(c[290]), .CLK(clk), .RST(rst), .Q(c[288]) );
  DFF \sreg_reg[289]  ( .D(c[289]), .CLK(clk), .RST(rst), .Q(c[287]) );
  DFF \sreg_reg[288]  ( .D(c[288]), .CLK(clk), .RST(rst), .Q(c[286]) );
  DFF \sreg_reg[287]  ( .D(c[287]), .CLK(clk), .RST(rst), .Q(c[285]) );
  DFF \sreg_reg[286]  ( .D(c[286]), .CLK(clk), .RST(rst), .Q(c[284]) );
  DFF \sreg_reg[285]  ( .D(c[285]), .CLK(clk), .RST(rst), .Q(c[283]) );
  DFF \sreg_reg[284]  ( .D(c[284]), .CLK(clk), .RST(rst), .Q(c[282]) );
  DFF \sreg_reg[283]  ( .D(c[283]), .CLK(clk), .RST(rst), .Q(c[281]) );
  DFF \sreg_reg[282]  ( .D(c[282]), .CLK(clk), .RST(rst), .Q(c[280]) );
  DFF \sreg_reg[281]  ( .D(c[281]), .CLK(clk), .RST(rst), .Q(c[279]) );
  DFF \sreg_reg[280]  ( .D(c[280]), .CLK(clk), .RST(rst), .Q(c[278]) );
  DFF \sreg_reg[279]  ( .D(c[279]), .CLK(clk), .RST(rst), .Q(c[277]) );
  DFF \sreg_reg[278]  ( .D(c[278]), .CLK(clk), .RST(rst), .Q(c[276]) );
  DFF \sreg_reg[277]  ( .D(c[277]), .CLK(clk), .RST(rst), .Q(c[275]) );
  DFF \sreg_reg[276]  ( .D(c[276]), .CLK(clk), .RST(rst), .Q(c[274]) );
  DFF \sreg_reg[275]  ( .D(c[275]), .CLK(clk), .RST(rst), .Q(c[273]) );
  DFF \sreg_reg[274]  ( .D(c[274]), .CLK(clk), .RST(rst), .Q(c[272]) );
  DFF \sreg_reg[273]  ( .D(c[273]), .CLK(clk), .RST(rst), .Q(c[271]) );
  DFF \sreg_reg[272]  ( .D(c[272]), .CLK(clk), .RST(rst), .Q(c[270]) );
  DFF \sreg_reg[271]  ( .D(c[271]), .CLK(clk), .RST(rst), .Q(c[269]) );
  DFF \sreg_reg[270]  ( .D(c[270]), .CLK(clk), .RST(rst), .Q(c[268]) );
  DFF \sreg_reg[269]  ( .D(c[269]), .CLK(clk), .RST(rst), .Q(c[267]) );
  DFF \sreg_reg[268]  ( .D(c[268]), .CLK(clk), .RST(rst), .Q(c[266]) );
  DFF \sreg_reg[267]  ( .D(c[267]), .CLK(clk), .RST(rst), .Q(c[265]) );
  DFF \sreg_reg[266]  ( .D(c[266]), .CLK(clk), .RST(rst), .Q(c[264]) );
  DFF \sreg_reg[265]  ( .D(c[265]), .CLK(clk), .RST(rst), .Q(c[263]) );
  DFF \sreg_reg[264]  ( .D(c[264]), .CLK(clk), .RST(rst), .Q(c[262]) );
  DFF \sreg_reg[263]  ( .D(c[263]), .CLK(clk), .RST(rst), .Q(c[261]) );
  DFF \sreg_reg[262]  ( .D(c[262]), .CLK(clk), .RST(rst), .Q(c[260]) );
  DFF \sreg_reg[261]  ( .D(c[261]), .CLK(clk), .RST(rst), .Q(c[259]) );
  DFF \sreg_reg[260]  ( .D(c[260]), .CLK(clk), .RST(rst), .Q(c[258]) );
  DFF \sreg_reg[259]  ( .D(c[259]), .CLK(clk), .RST(rst), .Q(c[257]) );
  DFF \sreg_reg[258]  ( .D(c[258]), .CLK(clk), .RST(rst), .Q(c[256]) );
  DFF \sreg_reg[257]  ( .D(c[257]), .CLK(clk), .RST(rst), .Q(c[255]) );
  DFF \sreg_reg[256]  ( .D(c[256]), .CLK(clk), .RST(rst), .Q(c[254]) );
  DFF \sreg_reg[255]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(c[253]) );
  DFF \sreg_reg[254]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(c[252]) );
  DFF \sreg_reg[253]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(c[251]) );
  DFF \sreg_reg[252]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(c[250]) );
  DFF \sreg_reg[251]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(c[249]) );
  DFF \sreg_reg[250]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(c[248]) );
  DFF \sreg_reg[249]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(c[247]) );
  DFF \sreg_reg[248]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(c[246]) );
  DFF \sreg_reg[247]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(c[245]) );
  DFF \sreg_reg[246]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(c[244]) );
  DFF \sreg_reg[245]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(c[243]) );
  DFF \sreg_reg[244]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(c[242]) );
  DFF \sreg_reg[243]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(c[241]) );
  DFF \sreg_reg[242]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(c[240]) );
  DFF \sreg_reg[241]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(c[239]) );
  DFF \sreg_reg[240]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(c[238]) );
  DFF \sreg_reg[239]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(c[237]) );
  DFF \sreg_reg[238]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(c[236]) );
  DFF \sreg_reg[237]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(c[235]) );
  DFF \sreg_reg[236]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(c[234]) );
  DFF \sreg_reg[235]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(c[233]) );
  DFF \sreg_reg[234]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(c[232]) );
  DFF \sreg_reg[233]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(c[231]) );
  DFF \sreg_reg[232]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(c[230]) );
  DFF \sreg_reg[231]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(c[229]) );
  DFF \sreg_reg[230]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(c[228]) );
  DFF \sreg_reg[229]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(c[227]) );
  DFF \sreg_reg[228]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(c[226]) );
  DFF \sreg_reg[227]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(c[225]) );
  DFF \sreg_reg[226]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(c[224]) );
  DFF \sreg_reg[225]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(c[223]) );
  DFF \sreg_reg[224]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(c[222]) );
  DFF \sreg_reg[223]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(c[221]) );
  DFF \sreg_reg[222]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(c[220]) );
  DFF \sreg_reg[221]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(c[219]) );
  DFF \sreg_reg[220]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(c[218]) );
  DFF \sreg_reg[219]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(c[217]) );
  DFF \sreg_reg[218]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(c[216]) );
  DFF \sreg_reg[217]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(c[215]) );
  DFF \sreg_reg[216]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(c[214]) );
  DFF \sreg_reg[215]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(c[213]) );
  DFF \sreg_reg[214]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(c[212]) );
  DFF \sreg_reg[213]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(c[211]) );
  DFF \sreg_reg[212]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(c[210]) );
  DFF \sreg_reg[211]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(c[209]) );
  DFF \sreg_reg[210]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(c[208]) );
  DFF \sreg_reg[209]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(c[207]) );
  DFF \sreg_reg[208]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(c[206]) );
  DFF \sreg_reg[207]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(c[205]) );
  DFF \sreg_reg[206]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(c[204]) );
  DFF \sreg_reg[205]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(c[203]) );
  DFF \sreg_reg[204]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(c[202]) );
  DFF \sreg_reg[203]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(c[201]) );
  DFF \sreg_reg[202]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(c[200]) );
  DFF \sreg_reg[201]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(c[199]) );
  DFF \sreg_reg[200]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(c[198]) );
  DFF \sreg_reg[199]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(c[197]) );
  DFF \sreg_reg[198]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(c[196]) );
  DFF \sreg_reg[197]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(c[195]) );
  DFF \sreg_reg[196]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(c[194]) );
  DFF \sreg_reg[195]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(c[193]) );
  DFF \sreg_reg[194]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(c[192]) );
  DFF \sreg_reg[193]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(c[191]) );
  DFF \sreg_reg[192]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(c[190]) );
  DFF \sreg_reg[191]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(c[189]) );
  DFF \sreg_reg[190]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(c[188]) );
  DFF \sreg_reg[189]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(c[187]) );
  DFF \sreg_reg[188]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(c[186]) );
  DFF \sreg_reg[187]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(c[185]) );
  DFF \sreg_reg[186]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(c[184]) );
  DFF \sreg_reg[185]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(c[183]) );
  DFF \sreg_reg[184]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(c[182]) );
  DFF \sreg_reg[183]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(c[181]) );
  DFF \sreg_reg[182]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(c[180]) );
  DFF \sreg_reg[181]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(c[179]) );
  DFF \sreg_reg[180]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(c[178]) );
  DFF \sreg_reg[179]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(c[177]) );
  DFF \sreg_reg[178]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(c[176]) );
  DFF \sreg_reg[177]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(c[175]) );
  DFF \sreg_reg[176]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(c[174]) );
  DFF \sreg_reg[175]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(c[173]) );
  DFF \sreg_reg[174]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(c[172]) );
  DFF \sreg_reg[173]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(c[171]) );
  DFF \sreg_reg[172]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(c[170]) );
  DFF \sreg_reg[171]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(c[169]) );
  DFF \sreg_reg[170]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(c[168]) );
  DFF \sreg_reg[169]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(c[167]) );
  DFF \sreg_reg[168]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(c[166]) );
  DFF \sreg_reg[167]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(c[165]) );
  DFF \sreg_reg[166]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(c[164]) );
  DFF \sreg_reg[165]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(c[163]) );
  DFF \sreg_reg[164]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(c[162]) );
  DFF \sreg_reg[163]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(c[161]) );
  DFF \sreg_reg[162]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(c[160]) );
  DFF \sreg_reg[161]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(c[159]) );
  DFF \sreg_reg[160]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(c[158]) );
  DFF \sreg_reg[159]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(c[157]) );
  DFF \sreg_reg[158]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(c[156]) );
  DFF \sreg_reg[157]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(c[155]) );
  DFF \sreg_reg[156]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(c[154]) );
  DFF \sreg_reg[155]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(c[153]) );
  DFF \sreg_reg[154]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(c[152]) );
  DFF \sreg_reg[153]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(c[151]) );
  DFF \sreg_reg[152]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(c[150]) );
  DFF \sreg_reg[151]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(c[149]) );
  DFF \sreg_reg[150]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(c[148]) );
  DFF \sreg_reg[149]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(c[147]) );
  DFF \sreg_reg[148]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(c[146]) );
  DFF \sreg_reg[147]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(c[145]) );
  DFF \sreg_reg[146]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(c[144]) );
  DFF \sreg_reg[145]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(c[143]) );
  DFF \sreg_reg[144]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(c[142]) );
  DFF \sreg_reg[143]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(c[141]) );
  DFF \sreg_reg[142]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(c[140]) );
  DFF \sreg_reg[141]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(c[139]) );
  DFF \sreg_reg[140]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(c[138]) );
  DFF \sreg_reg[139]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(c[137]) );
  DFF \sreg_reg[138]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(c[136]) );
  DFF \sreg_reg[137]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(c[135]) );
  DFF \sreg_reg[136]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(c[134]) );
  DFF \sreg_reg[135]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(c[133]) );
  DFF \sreg_reg[134]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(c[132]) );
  DFF \sreg_reg[133]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(c[131]) );
  DFF \sreg_reg[132]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(c[130]) );
  DFF \sreg_reg[131]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(c[129]) );
  DFF \sreg_reg[130]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(c[128]) );
  DFF \sreg_reg[129]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(c[127]) );
  DFF \sreg_reg[128]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(c[126]) );
  DFF \sreg_reg[127]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[125]) );
  DFF \sreg_reg[126]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[124]) );
  DFF \sreg_reg[125]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[123]) );
  DFF \sreg_reg[124]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[122]) );
  DFF \sreg_reg[123]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[121]) );
  DFF \sreg_reg[122]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[120]) );
  DFF \sreg_reg[121]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[120]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[119]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[118]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[117]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[116]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[115]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[114]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[113]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[112]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[111]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[110]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[109]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[108]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[107]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[106]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[105]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[104]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[103]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[102]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[101]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[100]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[99]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[98]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[97]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[96]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[95]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[94]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[93]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[92]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[91]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[90]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[89]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[88]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[87]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[86]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[85]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[84]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[83]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[82]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[81]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[80]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[79]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[78]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[77]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[76]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[75]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[74]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[73]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[72]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[71]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[70]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[69]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[68]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[67]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[66]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[65]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[64]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[63]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[62]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[61]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[60]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[59]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[58]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[57]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[56]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[55]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[54]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[53]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[52]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[51]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[50]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[49]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[48]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[47]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[46]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[45]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[44]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[43]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[42]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[41]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[40]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[39]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[38]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[37]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[36]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[35]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[34]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[33]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[32]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[31]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[30]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[29]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[28]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[27]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[26]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[25]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[24]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[23]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[22]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[21]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[20]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[19]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[18]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[17]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[16]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[15]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[14]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[13]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[12]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[11]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[10]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[9]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[8]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[7]  ( .D(c[7]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[6]  ( .D(c[6]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[5]  ( .D(c[5]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[4]  ( .D(c[4]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[3]  ( .D(c[3]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[2]  ( .D(c[2]), .CLK(clk), .RST(rst), .Q(c[0]) );
  ADD_N1024_1 ADD_ ( .A({1'b0, 1'b0, sreg[2045:1024]}), .B(clocal), .CI(1'b0), 
        .S({swire, c[1023:1022]}) );
  mult_N1024_CC512_DW02_mult_0 mult_44 ( .A(a), .B(b), .TC(1'b0), .PRODUCT({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, clocal}) );
endmodule

